module b04_reset(clock, RESET_G, nRESET_G, RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_, DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_, DATA_OUT_REG_7_, DATA_OUT_REG_6_, DATA_OUT_REG_5_, DATA_OUT_REG_4_, DATA_OUT_REG_3_, DATA_OUT_REG_2_, DATA_OUT_REG_1_, DATA_OUT_REG_0_);
  input AVERAGE;
  input DATA_IN_0_;
  input DATA_IN_1_;
  input DATA_IN_2_;
  input DATA_IN_3_;
  input DATA_IN_4_;
  input DATA_IN_5_;
  input DATA_IN_6_;
  input DATA_IN_7_;
  output DATA_OUT_REG_0_;
  output DATA_OUT_REG_1_;
  output DATA_OUT_REG_2_;
  output DATA_OUT_REG_3_;
  output DATA_OUT_REG_4_;
  output DATA_OUT_REG_5_;
  output DATA_OUT_REG_6_;
  output DATA_OUT_REG_7_;
  input ENABLE;
  wire REG1_REG_0_;
  wire REG1_REG_1_;
  wire REG1_REG_2_;
  wire REG1_REG_3_;
  wire REG1_REG_4_;
  wire REG1_REG_5_;
  wire REG1_REG_6_;
  wire REG1_REG_7_;
  wire REG2_REG_0_;
  wire REG2_REG_1_;
  wire REG2_REG_2_;
  wire REG2_REG_3_;
  wire REG2_REG_4_;
  wire REG2_REG_5_;
  wire REG2_REG_6_;
  wire REG2_REG_7_;
  wire REG3_REG_0_;
  wire REG3_REG_1_;
  wire REG3_REG_2_;
  wire REG3_REG_3_;
  wire REG3_REG_4_;
  wire REG3_REG_5_;
  wire REG3_REG_6_;
  wire REG3_REG_7_;
  wire REG4_REG_0_;
  wire REG4_REG_1_;
  wire REG4_REG_2_;
  wire REG4_REG_3_;
  wire REG4_REG_4_;
  wire REG4_REG_5_;
  wire REG4_REG_6_;
  wire REG4_REG_7_;
  input RESET_G;
  input RESTART;
  wire RESTART_bF_buf0;
  wire RESTART_bF_buf1;
  wire RESTART_bF_buf2;
  wire RESTART_bF_buf3;
  wire RLAST_REG_0_;
  wire RLAST_REG_1_;
  wire RLAST_REG_2_;
  wire RLAST_REG_3_;
  wire RLAST_REG_4_;
  wire RLAST_REG_5_;
  wire RLAST_REG_6_;
  wire RLAST_REG_7_;
  wire RMAX_REG_0_;
  wire RMAX_REG_1_;
  wire RMAX_REG_2_;
  wire RMAX_REG_3_;
  wire RMAX_REG_4_;
  wire RMAX_REG_5_;
  wire RMAX_REG_6_;
  wire RMAX_REG_7_;
  wire RMIN_REG_0_;
  wire RMIN_REG_1_;
  wire RMIN_REG_2_;
  wire RMIN_REG_3_;
  wire RMIN_REG_4_;
  wire RMIN_REG_5_;
  wire RMIN_REG_6_;
  wire RMIN_REG_7_;
  wire STATO_REG_0_;
  wire STATO_REG_1_;
  wire _abc_3548_n146;
  wire _abc_3548_n147_1;
  wire _abc_3548_n147_1_bF_buf0;
  wire _abc_3548_n147_1_bF_buf1;
  wire _abc_3548_n147_1_bF_buf2;
  wire _abc_3548_n147_1_bF_buf3;
  wire _abc_3548_n147_1_bF_buf4;
  wire _abc_3548_n148;
  wire _abc_3548_n148_bF_buf0;
  wire _abc_3548_n148_bF_buf1;
  wire _abc_3548_n148_bF_buf2;
  wire _abc_3548_n148_bF_buf3;
  wire _abc_3548_n148_bF_buf4;
  wire _abc_3548_n148_bF_buf5;
  wire _abc_3548_n148_bF_buf6;
  wire _abc_3548_n148_bF_buf7;
  wire _abc_3548_n149;
  wire _abc_3548_n150;
  wire _abc_3548_n151;
  wire _abc_3548_n153;
  wire _abc_3548_n154;
  wire _abc_3548_n155;
  wire _abc_3548_n156;
  wire _abc_3548_n157;
  wire _abc_3548_n158;
  wire _abc_3548_n159;
  wire _abc_3548_n160;
  wire _abc_3548_n161;
  wire _abc_3548_n162_1;
  wire _abc_3548_n163;
  wire _abc_3548_n164;
  wire _abc_3548_n165_1;
  wire _abc_3548_n166;
  wire _abc_3548_n167;
  wire _abc_3548_n168;
  wire _abc_3548_n169_1;
  wire _abc_3548_n170;
  wire _abc_3548_n171;
  wire _abc_3548_n172;
  wire _abc_3548_n173;
  wire _abc_3548_n174;
  wire _abc_3548_n175;
  wire _abc_3548_n176;
  wire _abc_3548_n177;
  wire _abc_3548_n178;
  wire _abc_3548_n179_1;
  wire _abc_3548_n180;
  wire _abc_3548_n181;
  wire _abc_3548_n182_1;
  wire _abc_3548_n183;
  wire _abc_3548_n184;
  wire _abc_3548_n185;
  wire _abc_3548_n186;
  wire _abc_3548_n187;
  wire _abc_3548_n188;
  wire _abc_3548_n189;
  wire _abc_3548_n190_1;
  wire _abc_3548_n191;
  wire _abc_3548_n192;
  wire _abc_3548_n193;
  wire _abc_3548_n194;
  wire _abc_3548_n195;
  wire _abc_3548_n196;
  wire _abc_3548_n197;
  wire _abc_3548_n198;
  wire _abc_3548_n199;
  wire _abc_3548_n200;
  wire _abc_3548_n201;
  wire _abc_3548_n202;
  wire _abc_3548_n203;
  wire _abc_3548_n204;
  wire _abc_3548_n205;
  wire _abc_3548_n206;
  wire _abc_3548_n207;
  wire _abc_3548_n208;
  wire _abc_3548_n209_1;
  wire _abc_3548_n210;
  wire _abc_3548_n211_1;
  wire _abc_3548_n212;
  wire _abc_3548_n213;
  wire _abc_3548_n214;
  wire _abc_3548_n215;
  wire _abc_3548_n216;
  wire _abc_3548_n217;
  wire _abc_3548_n218_1;
  wire _abc_3548_n219;
  wire _abc_3548_n220;
  wire _abc_3548_n221;
  wire _abc_3548_n222;
  wire _abc_3548_n223;
  wire _abc_3548_n224;
  wire _abc_3548_n225;
  wire _abc_3548_n226;
  wire _abc_3548_n227;
  wire _abc_3548_n228;
  wire _abc_3548_n229;
  wire _abc_3548_n230;
  wire _abc_3548_n231;
  wire _abc_3548_n232;
  wire _abc_3548_n233;
  wire _abc_3548_n234;
  wire _abc_3548_n235;
  wire _abc_3548_n236;
  wire _abc_3548_n237;
  wire _abc_3548_n238;
  wire _abc_3548_n239_1;
  wire _abc_3548_n240;
  wire _abc_3548_n241_1;
  wire _abc_3548_n242;
  wire _abc_3548_n243;
  wire _abc_3548_n244;
  wire _abc_3548_n245;
  wire _abc_3548_n246;
  wire _abc_3548_n247;
  wire _abc_3548_n248_1;
  wire _abc_3548_n249;
  wire _abc_3548_n250;
  wire _abc_3548_n251;
  wire _abc_3548_n252;
  wire _abc_3548_n253_1;
  wire _abc_3548_n254;
  wire _abc_3548_n255_1;
  wire _abc_3548_n256;
  wire _abc_3548_n257;
  wire _abc_3548_n258;
  wire _abc_3548_n259;
  wire _abc_3548_n260_1;
  wire _abc_3548_n261;
  wire _abc_3548_n262;
  wire _abc_3548_n263_1;
  wire _abc_3548_n264;
  wire _abc_3548_n265_1;
  wire _abc_3548_n266;
  wire _abc_3548_n267;
  wire _abc_3548_n268;
  wire _abc_3548_n269;
  wire _abc_3548_n270_1;
  wire _abc_3548_n271;
  wire _abc_3548_n272_1;
  wire _abc_3548_n273;
  wire _abc_3548_n274;
  wire _abc_3548_n275_1;
  wire _abc_3548_n276;
  wire _abc_3548_n277_1;
  wire _abc_3548_n278;
  wire _abc_3548_n279_1;
  wire _abc_3548_n280_1;
  wire _abc_3548_n281;
  wire _abc_3548_n282_1;
  wire _abc_3548_n283_1;
  wire _abc_3548_n284;
  wire _abc_3548_n285_1;
  wire _abc_3548_n286_1;
  wire _abc_3548_n287;
  wire _abc_3548_n288_1;
  wire _abc_3548_n289;
  wire _abc_3548_n290_1;
  wire _abc_3548_n291;
  wire _abc_3548_n292;
  wire _abc_3548_n293_1;
  wire _abc_3548_n294;
  wire _abc_3548_n295_1;
  wire _abc_3548_n296;
  wire _abc_3548_n297;
  wire _abc_3548_n298_1;
  wire _abc_3548_n299_1;
  wire _abc_3548_n300;
  wire _abc_3548_n301_1;
  wire _abc_3548_n302_1;
  wire _abc_3548_n302_1_bF_buf0;
  wire _abc_3548_n302_1_bF_buf1;
  wire _abc_3548_n302_1_bF_buf2;
  wire _abc_3548_n302_1_bF_buf3;
  wire _abc_3548_n302_1_bF_buf4;
  wire _abc_3548_n302_1_bF_buf5;
  wire _abc_3548_n303;
  wire _abc_3548_n304_1;
  wire _abc_3548_n305;
  wire _abc_3548_n306_1;
  wire _abc_3548_n307;
  wire _abc_3548_n309_1;
  wire _abc_3548_n310;
  wire _abc_3548_n311_1;
  wire _abc_3548_n312;
  wire _abc_3548_n313;
  wire _abc_3548_n314_1;
  wire _abc_3548_n315;
  wire _abc_3548_n316_1;
  wire _abc_3548_n317;
  wire _abc_3548_n318;
  wire _abc_3548_n319_1;
  wire _abc_3548_n320;
  wire _abc_3548_n321_1;
  wire _abc_3548_n322;
  wire _abc_3548_n323;
  wire _abc_3548_n324_1;
  wire _abc_3548_n325_1;
  wire _abc_3548_n326;
  wire _abc_3548_n327_1;
  wire _abc_3548_n328_1;
  wire _abc_3548_n329;
  wire _abc_3548_n330_1;
  wire _abc_3548_n331;
  wire _abc_3548_n332_1;
  wire _abc_3548_n333;
  wire _abc_3548_n334;
  wire _abc_3548_n335_1;
  wire _abc_3548_n336;
  wire _abc_3548_n337_1;
  wire _abc_3548_n338;
  wire _abc_3548_n339;
  wire _abc_3548_n340_1;
  wire _abc_3548_n341_1;
  wire _abc_3548_n342;
  wire _abc_3548_n343_1;
  wire _abc_3548_n345;
  wire _abc_3548_n346_1;
  wire _abc_3548_n347_1;
  wire _abc_3548_n348;
  wire _abc_3548_n349_1;
  wire _abc_3548_n350_1;
  wire _abc_3548_n351;
  wire _abc_3548_n352_1;
  wire _abc_3548_n353;
  wire _abc_3548_n354_1;
  wire _abc_3548_n355;
  wire _abc_3548_n356;
  wire _abc_3548_n357_1;
  wire _abc_3548_n358;
  wire _abc_3548_n359_1;
  wire _abc_3548_n360;
  wire _abc_3548_n361;
  wire _abc_3548_n362_1;
  wire _abc_3548_n363_1;
  wire _abc_3548_n364;
  wire _abc_3548_n365_1;
  wire _abc_3548_n366;
  wire _abc_3548_n367_1;
  wire _abc_3548_n368;
  wire _abc_3548_n369;
  wire _abc_3548_n370_1;
  wire _abc_3548_n371;
  wire _abc_3548_n372;
  wire _abc_3548_n373;
  wire _abc_3548_n374_1;
  wire _abc_3548_n375;
  wire _abc_3548_n376;
  wire _abc_3548_n377_1;
  wire _abc_3548_n378;
  wire _abc_3548_n379;
  wire _abc_3548_n380_1;
  wire _abc_3548_n381;
  wire _abc_3548_n382_1;
  wire _abc_3548_n384_1;
  wire _abc_3548_n385;
  wire _abc_3548_n386;
  wire _abc_3548_n387_1;
  wire _abc_3548_n388;
  wire _abc_3548_n389;
  wire _abc_3548_n390;
  wire _abc_3548_n391;
  wire _abc_3548_n392;
  wire _abc_3548_n393_1;
  wire _abc_3548_n394;
  wire _abc_3548_n395;
  wire _abc_3548_n396_1;
  wire _abc_3548_n397;
  wire _abc_3548_n398;
  wire _abc_3548_n399_1;
  wire _abc_3548_n400;
  wire _abc_3548_n401;
  wire _abc_3548_n402_1;
  wire _abc_3548_n403;
  wire _abc_3548_n404;
  wire _abc_3548_n405_1;
  wire _abc_3548_n406;
  wire _abc_3548_n407;
  wire _abc_3548_n408;
  wire _abc_3548_n409_1;
  wire _abc_3548_n410;
  wire _abc_3548_n411;
  wire _abc_3548_n412;
  wire _abc_3548_n413_1;
  wire _abc_3548_n414;
  wire _abc_3548_n415;
  wire _abc_3548_n416_1;
  wire _abc_3548_n417;
  wire _abc_3548_n418;
  wire _abc_3548_n419;
  wire _abc_3548_n420;
  wire _abc_3548_n421;
  wire _abc_3548_n422;
  wire _abc_3548_n423;
  wire _abc_3548_n424;
  wire _abc_3548_n426;
  wire _abc_3548_n427;
  wire _abc_3548_n428;
  wire _abc_3548_n429;
  wire _abc_3548_n430;
  wire _abc_3548_n431;
  wire _abc_3548_n432;
  wire _abc_3548_n433;
  wire _abc_3548_n434;
  wire _abc_3548_n435;
  wire _abc_3548_n436;
  wire _abc_3548_n437;
  wire _abc_3548_n438;
  wire _abc_3548_n439;
  wire _abc_3548_n440;
  wire _abc_3548_n441;
  wire _abc_3548_n442;
  wire _abc_3548_n443;
  wire _abc_3548_n444;
  wire _abc_3548_n445;
  wire _abc_3548_n446;
  wire _abc_3548_n447;
  wire _abc_3548_n448;
  wire _abc_3548_n449;
  wire _abc_3548_n450;
  wire _abc_3548_n451;
  wire _abc_3548_n452_1;
  wire _abc_3548_n453;
  wire _abc_3548_n454_1;
  wire _abc_3548_n455;
  wire _abc_3548_n456_1;
  wire _abc_3548_n457;
  wire _abc_3548_n458_1;
  wire _abc_3548_n459;
  wire _abc_3548_n460_1;
  wire _abc_3548_n461;
  wire _abc_3548_n462;
  wire _abc_3548_n463_1;
  wire _abc_3548_n464;
  wire _abc_3548_n465_1;
  wire _abc_3548_n466;
  wire _abc_3548_n467_1;
  wire _abc_3548_n468;
  wire _abc_3548_n469;
  wire _abc_3548_n470_1;
  wire _abc_3548_n472_1;
  wire _abc_3548_n473;
  wire _abc_3548_n474_1;
  wire _abc_3548_n475;
  wire _abc_3548_n476_1;
  wire _abc_3548_n477;
  wire _abc_3548_n478_1;
  wire _abc_3548_n479;
  wire _abc_3548_n480_1;
  wire _abc_3548_n481;
  wire _abc_3548_n482_1;
  wire _abc_3548_n483;
  wire _abc_3548_n484_1;
  wire _abc_3548_n485;
  wire _abc_3548_n486_1;
  wire _abc_3548_n487_1;
  wire _abc_3548_n488;
  wire _abc_3548_n489;
  wire _abc_3548_n490;
  wire _abc_3548_n491;
  wire _abc_3548_n492;
  wire _abc_3548_n493;
  wire _abc_3548_n494;
  wire _abc_3548_n495;
  wire _abc_3548_n496;
  wire _abc_3548_n497;
  wire _abc_3548_n498;
  wire _abc_3548_n499;
  wire _abc_3548_n500;
  wire _abc_3548_n501;
  wire _abc_3548_n502;
  wire _abc_3548_n503;
  wire _abc_3548_n504;
  wire _abc_3548_n505;
  wire _abc_3548_n506;
  wire _abc_3548_n507;
  wire _abc_3548_n508;
  wire _abc_3548_n509;
  wire _abc_3548_n510;
  wire _abc_3548_n511;
  wire _abc_3548_n512;
  wire _abc_3548_n513;
  wire _abc_3548_n514;
  wire _abc_3548_n515;
  wire _abc_3548_n516;
  wire _abc_3548_n518;
  wire _abc_3548_n519;
  wire _abc_3548_n520;
  wire _abc_3548_n521;
  wire _abc_3548_n522;
  wire _abc_3548_n523;
  wire _abc_3548_n524;
  wire _abc_3548_n525;
  wire _abc_3548_n526;
  wire _abc_3548_n528;
  wire _abc_3548_n529;
  wire _abc_3548_n530;
  wire _abc_3548_n531;
  wire _abc_3548_n532;
  wire _abc_3548_n534;
  wire _abc_3548_n535;
  wire _abc_3548_n536;
  wire _abc_3548_n538;
  wire _abc_3548_n539;
  wire _abc_3548_n540;
  wire _abc_3548_n542;
  wire _abc_3548_n543;
  wire _abc_3548_n544;
  wire _abc_3548_n546;
  wire _abc_3548_n547;
  wire _abc_3548_n548;
  wire _abc_3548_n550;
  wire _abc_3548_n551;
  wire _abc_3548_n552;
  wire _abc_3548_n554;
  wire _abc_3548_n555;
  wire _abc_3548_n556;
  wire _abc_3548_n558;
  wire _abc_3548_n559;
  wire _abc_3548_n560;
  wire _abc_3548_n562;
  wire _abc_3548_n563;
  wire _abc_3548_n564;
  wire _abc_3548_n566;
  wire _abc_3548_n567;
  wire _abc_3548_n568;
  wire _abc_3548_n570;
  wire _abc_3548_n571;
  wire _abc_3548_n572;
  wire _abc_3548_n574;
  wire _abc_3548_n575;
  wire _abc_3548_n576;
  wire _abc_3548_n578;
  wire _abc_3548_n579;
  wire _abc_3548_n580;
  wire _abc_3548_n582;
  wire _abc_3548_n583;
  wire _abc_3548_n584;
  wire _abc_3548_n586;
  wire _abc_3548_n587;
  wire _abc_3548_n588;
  wire _abc_3548_n590;
  wire _abc_3548_n591;
  wire _abc_3548_n592;
  wire _abc_3548_n594;
  wire _abc_3548_n595;
  wire _abc_3548_n596;
  wire _abc_3548_n598;
  wire _abc_3548_n599;
  wire _abc_3548_n600;
  wire _abc_3548_n602;
  wire _abc_3548_n603;
  wire _abc_3548_n604;
  wire _abc_3548_n606;
  wire _abc_3548_n607;
  wire _abc_3548_n608;
  wire _abc_3548_n610;
  wire _abc_3548_n611;
  wire _abc_3548_n612;
  wire _abc_3548_n614;
  wire _abc_3548_n615;
  wire _abc_3548_n616;
  wire _abc_3548_n618;
  wire _abc_3548_n619;
  wire _abc_3548_n620;
  wire _abc_3548_n622;
  wire _abc_3548_n623;
  wire _abc_3548_n624;
  wire _abc_3548_n626;
  wire _abc_3548_n627;
  wire _abc_3548_n628;
  wire _abc_3548_n630;
  wire _abc_3548_n631;
  wire _abc_3548_n632;
  wire _abc_3548_n634;
  wire _abc_3548_n635;
  wire _abc_3548_n636;
  wire _abc_3548_n638;
  wire _abc_3548_n639;
  wire _abc_3548_n640;
  wire _abc_3548_n642;
  wire _abc_3548_n643;
  wire _abc_3548_n644;
  wire _abc_3548_n646;
  wire _abc_3548_n647;
  wire _abc_3548_n648;
  wire _abc_3548_n650;
  wire _abc_3548_n651;
  wire _abc_3548_n652;
  wire _abc_3548_n654;
  wire _abc_3548_n655;
  wire _abc_3548_n656;
  wire _abc_3548_n658;
  wire _abc_3548_n659;
  wire _abc_3548_n660;
  wire _abc_3548_n662;
  wire _abc_3548_n663;
  wire _abc_3548_n664;
  wire _abc_3548_n665;
  wire _abc_3548_n666;
  wire _abc_3548_n667;
  wire _abc_3548_n668;
  wire _abc_3548_n669;
  wire _abc_3548_n671;
  wire _abc_3548_n672;
  wire _abc_3548_n673;
  wire _abc_3548_n675;
  wire _abc_3548_n676;
  wire _abc_3548_n677;
  wire _abc_3548_n679;
  wire _abc_3548_n680;
  wire _abc_3548_n681;
  wire _abc_3548_n683;
  wire _abc_3548_n684;
  wire _abc_3548_n685;
  wire _abc_3548_n687;
  wire _abc_3548_n688;
  wire _abc_3548_n689;
  wire _abc_3548_n691;
  wire _abc_3548_n692;
  wire _abc_3548_n693;
  wire _abc_3548_n695;
  wire _abc_3548_n696;
  wire _abc_3548_n697;
  wire _abc_3548_n699;
  wire _abc_3548_n700;
  wire _abc_3548_n701;
  wire _abc_3548_n702;
  wire _abc_3548_n703;
  wire _abc_3548_n704;
  wire _abc_3548_n705;
  wire _abc_3548_n706;
  wire _abc_3548_n707;
  wire _abc_3548_n708;
  wire _abc_3548_n709;
  wire _abc_3548_n710;
  wire _abc_3548_n711;
  wire _abc_3548_n712;
  wire _abc_3548_n713;
  wire _abc_3548_n714;
  wire _abc_3548_n715;
  wire _abc_3548_n716;
  wire _abc_3548_n717;
  wire _abc_3548_n718;
  wire _abc_3548_n719;
  wire _abc_3548_n720;
  wire _abc_3548_n721;
  wire _abc_3548_n722;
  wire _abc_3548_n723;
  wire _abc_3548_n724;
  wire _abc_3548_n725;
  wire _abc_3548_n726;
  wire _abc_3548_n727;
  wire _abc_3548_n728;
  wire _abc_3548_n729;
  wire _abc_3548_n730;
  wire _abc_3548_n731;
  wire _abc_3548_n732;
  wire _abc_3548_n733;
  wire _abc_3548_n734;
  wire _abc_3548_n735;
  wire _abc_3548_n736;
  wire _abc_3548_n737;
  wire _abc_3548_n738;
  wire _abc_3548_n739;
  wire _abc_3548_n740;
  wire _abc_3548_n741;
  wire _abc_3548_n742;
  wire _abc_3548_n743;
  wire _abc_3548_n744;
  wire _abc_3548_n745;
  wire _abc_3548_n746;
  wire _abc_3548_n747;
  wire _abc_3548_n748;
  wire _abc_3548_n749;
  wire _abc_3548_n750;
  wire _abc_3548_n751;
  wire _abc_3548_n752;
  wire _abc_3548_n753;
  wire _abc_3548_n754;
  wire _abc_3548_n755;
  wire _abc_3548_n756;
  wire _abc_3548_n757;
  wire _abc_3548_n758;
  wire _abc_3548_n759;
  wire _abc_3548_n760;
  wire _abc_3548_n761;
  wire _abc_3548_n762;
  wire _abc_3548_n763;
  wire _abc_3548_n764;
  wire _abc_3548_n765;
  wire _abc_3548_n766;
  wire _abc_3548_n767;
  wire _abc_3548_n768;
  wire _abc_3548_n769;
  wire _abc_3548_n770;
  wire _abc_3548_n771;
  wire _abc_3548_n772;
  wire _abc_3548_n773;
  wire _abc_3548_n774;
  wire _abc_3548_n775;
  wire _abc_3548_n776;
  wire _abc_3548_n778;
  wire _abc_3548_n779;
  wire _abc_3548_n780;
  wire _abc_3548_n782;
  wire _abc_3548_n783;
  wire _abc_3548_n784;
  wire _abc_3548_n786;
  wire _abc_3548_n787;
  wire _abc_3548_n788;
  wire _abc_3548_n790;
  wire _abc_3548_n791;
  wire _abc_3548_n792;
  wire _abc_3548_n794;
  wire _abc_3548_n795;
  wire _abc_3548_n796;
  wire _abc_3548_n798;
  wire _abc_3548_n799;
  wire _abc_3548_n800;
  wire _abc_3548_n802;
  wire _abc_3548_n803;
  wire _abc_3548_n804;
  wire _abc_3548_n806;
  wire _abc_3548_n807;
  wire _abc_3548_n808;
  wire _abc_3548_n809;
  wire _abc_3548_n810;
  wire _abc_3548_n811;
  wire _abc_3548_n813;
  wire _abc_3548_n814;
  wire _abc_3548_n815;
  wire _abc_3548_n817;
  wire _abc_3548_n818;
  wire _abc_3548_n819;
  wire _abc_3548_n821;
  wire _abc_3548_n822;
  wire _abc_3548_n823;
  wire _abc_3548_n825;
  wire _abc_3548_n826;
  wire _abc_3548_n827;
  wire _abc_3548_n829;
  wire _abc_3548_n830;
  wire _abc_3548_n831;
  wire _abc_3548_n833;
  wire _abc_3548_n834;
  wire _abc_3548_n835;
  wire _abc_3548_n837;
  wire _abc_3548_n838;
  wire _abc_3548_n839;
  wire _abc_3548_n841;
  input clock;
  wire clock_bF_buf0;
  wire clock_bF_buf1;
  wire clock_bF_buf2;
  wire clock_bF_buf3;
  wire clock_bF_buf4;
  wire clock_bF_buf5;
  wire clock_bF_buf6;
  wire clock_bF_buf7;
  wire n104;
  wire n109;
  wire n114;
  wire n119;
  wire n124;
  wire n129;
  wire n134;
  wire n139;
  wire n144;
  wire n149;
  wire n154;
  wire n159;
  wire n164;
  wire n169;
  wire n174;
  wire n179;
  wire n184;
  wire n189;
  wire n194;
  wire n199;
  wire n204;
  wire n209;
  wire n214;
  wire n219;
  wire n224;
  wire n229;
  wire n234;
  wire n239;
  wire n244;
  wire n249;
  wire n254;
  wire n259;
  wire n264;
  wire n269;
  wire n274;
  wire n279;
  wire n284;
  wire n289;
  wire n294;
  wire n299;
  wire n304;
  wire n309;
  wire n314;
  wire n319;
  wire n324;
  wire n328;
  wire n332;
  wire n336;
  wire n340;
  wire n344;
  wire n348;
  wire n352;
  wire n356;
  wire n361;
  wire n44;
  wire n49;
  wire n54;
  wire n59;
  wire n64;
  wire n69;
  wire n74;
  wire n79;
  wire n84;
  wire n89;
  wire n94;
  wire n99;
  input nRESET_G;
  AND2X2 AND2X2_1 ( .A(_abc_3548_n146), .B(STATO_REG_1_), .Y(_abc_3548_n147_1) );
  AND2X2 AND2X2_10 ( .A(_abc_3548_n159), .B(DATA_IN_1_), .Y(_abc_3548_n167) );
  AND2X2 AND2X2_100 ( .A(_abc_3548_n345), .B(_abc_3548_n365_1), .Y(_abc_3548_n368) );
  AND2X2 AND2X2_101 ( .A(_abc_3548_n369), .B(_abc_3548_n347_1), .Y(_abc_3548_n370_1) );
  AND2X2 AND2X2_102 ( .A(_abc_3548_n287), .B(_abc_3548_n372), .Y(_abc_3548_n373) );
  AND2X2 AND2X2_103 ( .A(_abc_3548_n373), .B(_abc_3548_n371), .Y(_abc_3548_n374_1) );
  AND2X2 AND2X2_104 ( .A(_abc_3548_n280_1), .B(_abc_3548_n365_1), .Y(_abc_3548_n375) );
  AND2X2 AND2X2_105 ( .A(_abc_3548_n297), .B(RLAST_REG_2_), .Y(_abc_3548_n376) );
  AND2X2 AND2X2_106 ( .A(_abc_3548_n300), .B(REG4_REG_2_), .Y(_abc_3548_n377_1) );
  AND2X2 AND2X2_107 ( .A(_abc_3548_n302_1), .B(DATA_OUT_REG_2_), .Y(_abc_3548_n378) );
  AND2X2 AND2X2_108 ( .A(_abc_3548_n385), .B(_abc_3548_n357_1), .Y(_abc_3548_n386) );
  AND2X2 AND2X2_109 ( .A(_abc_3548_n388), .B(_abc_3548_n387_1), .Y(_abc_3548_n389) );
  AND2X2 AND2X2_11 ( .A(_abc_3548_n165_1), .B(_abc_3548_n168), .Y(_abc_3548_n169_1) );
  AND2X2 AND2X2_110 ( .A(_abc_3548_n392), .B(_abc_3548_n391), .Y(_abc_3548_n393_1) );
  AND2X2 AND2X2_111 ( .A(_abc_3548_n390), .B(_abc_3548_n394), .Y(_abc_3548_n395) );
  AND2X2 AND2X2_112 ( .A(_abc_3548_n389), .B(_abc_3548_n393_1), .Y(_abc_3548_n397) );
  AND2X2 AND2X2_113 ( .A(_abc_3548_n396_1), .B(_abc_3548_n398), .Y(_abc_3548_n399_1) );
  AND2X2 AND2X2_114 ( .A(_abc_3548_n386), .B(_abc_3548_n399_1), .Y(_abc_3548_n400) );
  AND2X2 AND2X2_115 ( .A(_abc_3548_n401), .B(_abc_3548_n402_1), .Y(_abc_3548_n403) );
  AND2X2 AND2X2_116 ( .A(_abc_3548_n408), .B(_abc_3548_n404), .Y(_abc_3548_n409_1) );
  AND2X2 AND2X2_117 ( .A(_abc_3548_n403), .B(_abc_3548_n367_1), .Y(_abc_3548_n412) );
  AND2X2 AND2X2_118 ( .A(_abc_3548_n414), .B(_abc_3548_n287), .Y(_abc_3548_n415) );
  AND2X2 AND2X2_119 ( .A(_abc_3548_n415), .B(_abc_3548_n410), .Y(_abc_3548_n416_1) );
  AND2X2 AND2X2_12 ( .A(_abc_3548_n159), .B(_abc_3548_n171), .Y(_abc_3548_n172) );
  AND2X2 AND2X2_120 ( .A(_abc_3548_n407), .B(_abc_3548_n280_1), .Y(_abc_3548_n417) );
  AND2X2 AND2X2_121 ( .A(_abc_3548_n297), .B(RLAST_REG_3_), .Y(_abc_3548_n418) );
  AND2X2 AND2X2_122 ( .A(_abc_3548_n300), .B(REG4_REG_3_), .Y(_abc_3548_n419) );
  AND2X2 AND2X2_123 ( .A(_abc_3548_n302_1), .B(DATA_OUT_REG_3_), .Y(_abc_3548_n420) );
  AND2X2 AND2X2_124 ( .A(_abc_3548_n427), .B(_abc_3548_n426), .Y(_abc_3548_n428) );
  AND2X2 AND2X2_125 ( .A(_abc_3548_n431), .B(_abc_3548_n430), .Y(_abc_3548_n432) );
  AND2X2 AND2X2_126 ( .A(_abc_3548_n429), .B(_abc_3548_n433), .Y(_abc_3548_n434) );
  AND2X2 AND2X2_127 ( .A(_abc_3548_n428), .B(_abc_3548_n432), .Y(_abc_3548_n436) );
  AND2X2 AND2X2_128 ( .A(_abc_3548_n435), .B(_abc_3548_n437), .Y(_abc_3548_n438) );
  AND2X2 AND2X2_129 ( .A(_abc_3548_n440), .B(_abc_3548_n398), .Y(_abc_3548_n441) );
  AND2X2 AND2X2_13 ( .A(_abc_3548_n173), .B(RESTART), .Y(_abc_3548_n174) );
  AND2X2 AND2X2_130 ( .A(_abc_3548_n349_1), .B(_abc_3548_n358), .Y(_abc_3548_n443) );
  AND2X2 AND2X2_131 ( .A(_abc_3548_n444), .B(_abc_3548_n396_1), .Y(_abc_3548_n445) );
  AND2X2 AND2X2_132 ( .A(_abc_3548_n442), .B(_abc_3548_n447), .Y(_abc_3548_n448) );
  AND2X2 AND2X2_133 ( .A(_abc_3548_n448), .B(_abc_3548_n280_1), .Y(_abc_3548_n449) );
  AND2X2 AND2X2_134 ( .A(_abc_3548_n297), .B(RLAST_REG_4_), .Y(_abc_3548_n450) );
  AND2X2 AND2X2_135 ( .A(_abc_3548_n300), .B(REG4_REG_4_), .Y(_abc_3548_n451) );
  AND2X2 AND2X2_136 ( .A(_abc_3548_n302_1), .B(DATA_OUT_REG_4_), .Y(_abc_3548_n452_1) );
  AND2X2 AND2X2_137 ( .A(_abc_3548_n413_1), .B(_abc_3548_n370_1), .Y(_abc_3548_n457) );
  AND2X2 AND2X2_138 ( .A(_abc_3548_n446), .B(_abc_3548_n438), .Y(_abc_3548_n458_1) );
  AND2X2 AND2X2_139 ( .A(_abc_3548_n441), .B(_abc_3548_n439), .Y(_abc_3548_n459) );
  AND2X2 AND2X2_14 ( .A(_abc_3548_n177), .B(_abc_3548_n178), .Y(_abc_3548_n179_1) );
  AND2X2 AND2X2_140 ( .A(_abc_3548_n460_1), .B(_abc_3548_n412), .Y(_abc_3548_n461) );
  AND2X2 AND2X2_141 ( .A(_abc_3548_n448), .B(_abc_3548_n408), .Y(_abc_3548_n462) );
  AND2X2 AND2X2_142 ( .A(_abc_3548_n465_1), .B(_abc_3548_n466), .Y(_abc_3548_n467_1) );
  AND2X2 AND2X2_143 ( .A(_abc_3548_n468), .B(_abc_3548_n287), .Y(_abc_3548_n469) );
  AND2X2 AND2X2_144 ( .A(_abc_3548_n469), .B(_abc_3548_n464), .Y(_abc_3548_n470_1) );
  AND2X2 AND2X2_145 ( .A(_abc_3548_n446), .B(_abc_3548_n435), .Y(_abc_3548_n472_1) );
  AND2X2 AND2X2_146 ( .A(_abc_3548_n474_1), .B(_abc_3548_n473), .Y(_abc_3548_n475) );
  AND2X2 AND2X2_147 ( .A(_abc_3548_n478_1), .B(_abc_3548_n477), .Y(_abc_3548_n479) );
  AND2X2 AND2X2_148 ( .A(_abc_3548_n476_1), .B(_abc_3548_n479), .Y(_abc_3548_n480_1) );
  AND2X2 AND2X2_149 ( .A(_abc_3548_n484_1), .B(_abc_3548_n437), .Y(_abc_3548_n485) );
  AND2X2 AND2X2_15 ( .A(_abc_3548_n180), .B(_abc_3548_n181), .Y(_abc_3548_n182_1) );
  AND2X2 AND2X2_150 ( .A(_abc_3548_n441), .B(_abc_3548_n437), .Y(_abc_3548_n488) );
  AND2X2 AND2X2_151 ( .A(_abc_3548_n483), .B(_abc_3548_n435), .Y(_abc_3548_n489) );
  AND2X2 AND2X2_152 ( .A(_abc_3548_n491), .B(_abc_3548_n487_1), .Y(_abc_3548_n492) );
  AND2X2 AND2X2_153 ( .A(_abc_3548_n492), .B(_abc_3548_n280_1), .Y(_abc_3548_n493) );
  AND2X2 AND2X2_154 ( .A(_abc_3548_n297), .B(RLAST_REG_5_), .Y(_abc_3548_n494) );
  AND2X2 AND2X2_155 ( .A(_abc_3548_n300), .B(REG4_REG_5_), .Y(_abc_3548_n495) );
  AND2X2 AND2X2_156 ( .A(_abc_3548_n302_1), .B(DATA_OUT_REG_5_), .Y(_abc_3548_n496) );
  AND2X2 AND2X2_157 ( .A(_abc_3548_n463_1), .B(_abc_3548_n457), .Y(_abc_3548_n501) );
  AND2X2 AND2X2_158 ( .A(_abc_3548_n502), .B(_abc_3548_n485), .Y(_abc_3548_n503) );
  AND2X2 AND2X2_159 ( .A(_abc_3548_n504), .B(_abc_3548_n489), .Y(_abc_3548_n505) );
  AND2X2 AND2X2_16 ( .A(_abc_3548_n183), .B(_abc_3548_n170), .Y(_abc_3548_n184) );
  AND2X2 AND2X2_160 ( .A(_abc_3548_n506), .B(_abc_3548_n461), .Y(_abc_3548_n507) );
  AND2X2 AND2X2_161 ( .A(_abc_3548_n465_1), .B(_abc_3548_n492), .Y(_abc_3548_n508) );
  AND2X2 AND2X2_162 ( .A(_abc_3548_n511), .B(_abc_3548_n512), .Y(_abc_3548_n513) );
  AND2X2 AND2X2_163 ( .A(_abc_3548_n514), .B(_abc_3548_n510), .Y(_abc_3548_n515) );
  AND2X2 AND2X2_164 ( .A(_abc_3548_n515), .B(_abc_3548_n287), .Y(_abc_3548_n516) );
  AND2X2 AND2X2_165 ( .A(_abc_3548_n300), .B(REG4_REG_6_), .Y(_abc_3548_n518) );
  AND2X2 AND2X2_166 ( .A(_abc_3548_n297), .B(RLAST_REG_6_), .Y(_abc_3548_n519) );
  AND2X2 AND2X2_167 ( .A(_abc_3548_n302_1), .B(DATA_OUT_REG_6_), .Y(_abc_3548_n520) );
  AND2X2 AND2X2_168 ( .A(_abc_3548_n511), .B(_abc_3548_n287), .Y(_abc_3548_n525) );
  AND2X2 AND2X2_169 ( .A(_abc_3548_n524), .B(_abc_3548_n525), .Y(_abc_3548_n526) );
  AND2X2 AND2X2_17 ( .A(_abc_3548_n184), .B(_abc_3548_n157), .Y(_abc_3548_n186) );
  AND2X2 AND2X2_170 ( .A(_abc_3548_n300), .B(REG4_REG_7_), .Y(_abc_3548_n528) );
  AND2X2 AND2X2_171 ( .A(_abc_3548_n297), .B(RLAST_REG_7_), .Y(_abc_3548_n529) );
  AND2X2 AND2X2_172 ( .A(_abc_3548_n302_1), .B(DATA_OUT_REG_7_), .Y(_abc_3548_n530) );
  AND2X2 AND2X2_173 ( .A(_abc_3548_n302_1), .B(REG4_REG_0_), .Y(_abc_3548_n534) );
  AND2X2 AND2X2_174 ( .A(_abc_3548_n147_1), .B(REG3_REG_0_), .Y(_abc_3548_n535) );
  AND2X2 AND2X2_175 ( .A(_abc_3548_n302_1), .B(REG4_REG_1_), .Y(_abc_3548_n538) );
  AND2X2 AND2X2_176 ( .A(_abc_3548_n147_1), .B(REG3_REG_1_), .Y(_abc_3548_n539) );
  AND2X2 AND2X2_177 ( .A(_abc_3548_n302_1), .B(REG4_REG_2_), .Y(_abc_3548_n542) );
  AND2X2 AND2X2_178 ( .A(_abc_3548_n147_1), .B(REG3_REG_2_), .Y(_abc_3548_n543) );
  AND2X2 AND2X2_179 ( .A(_abc_3548_n302_1), .B(REG4_REG_3_), .Y(_abc_3548_n546) );
  AND2X2 AND2X2_18 ( .A(_abc_3548_n187), .B(_abc_3548_n185), .Y(_abc_3548_n188) );
  AND2X2 AND2X2_180 ( .A(_abc_3548_n147_1), .B(REG3_REG_3_), .Y(_abc_3548_n547) );
  AND2X2 AND2X2_181 ( .A(_abc_3548_n302_1), .B(REG4_REG_4_), .Y(_abc_3548_n550) );
  AND2X2 AND2X2_182 ( .A(_abc_3548_n147_1), .B(REG3_REG_4_), .Y(_abc_3548_n551) );
  AND2X2 AND2X2_183 ( .A(_abc_3548_n302_1), .B(REG4_REG_5_), .Y(_abc_3548_n554) );
  AND2X2 AND2X2_184 ( .A(_abc_3548_n147_1), .B(REG3_REG_5_), .Y(_abc_3548_n555) );
  AND2X2 AND2X2_185 ( .A(_abc_3548_n302_1), .B(REG4_REG_6_), .Y(_abc_3548_n558) );
  AND2X2 AND2X2_186 ( .A(_abc_3548_n147_1), .B(REG3_REG_6_), .Y(_abc_3548_n559) );
  AND2X2 AND2X2_187 ( .A(_abc_3548_n302_1), .B(REG4_REG_7_), .Y(_abc_3548_n562) );
  AND2X2 AND2X2_188 ( .A(_abc_3548_n147_1), .B(REG3_REG_7_), .Y(_abc_3548_n563) );
  AND2X2 AND2X2_189 ( .A(_abc_3548_n302_1), .B(REG3_REG_0_), .Y(_abc_3548_n566) );
  AND2X2 AND2X2_19 ( .A(DATA_IN_7_), .B(REG4_REG_7_), .Y(_abc_3548_n189) );
  AND2X2 AND2X2_190 ( .A(_abc_3548_n147_1), .B(REG2_REG_0_), .Y(_abc_3548_n567) );
  AND2X2 AND2X2_191 ( .A(_abc_3548_n302_1), .B(REG3_REG_1_), .Y(_abc_3548_n570) );
  AND2X2 AND2X2_192 ( .A(_abc_3548_n147_1), .B(REG2_REG_1_), .Y(_abc_3548_n571) );
  AND2X2 AND2X2_193 ( .A(_abc_3548_n302_1), .B(REG3_REG_2_), .Y(_abc_3548_n574) );
  AND2X2 AND2X2_194 ( .A(_abc_3548_n147_1), .B(REG2_REG_2_), .Y(_abc_3548_n575) );
  AND2X2 AND2X2_195 ( .A(_abc_3548_n302_1), .B(REG3_REG_3_), .Y(_abc_3548_n578) );
  AND2X2 AND2X2_196 ( .A(_abc_3548_n147_1), .B(REG2_REG_3_), .Y(_abc_3548_n579) );
  AND2X2 AND2X2_197 ( .A(_abc_3548_n302_1), .B(REG3_REG_4_), .Y(_abc_3548_n582) );
  AND2X2 AND2X2_198 ( .A(_abc_3548_n147_1), .B(REG2_REG_4_), .Y(_abc_3548_n583) );
  AND2X2 AND2X2_199 ( .A(_abc_3548_n302_1), .B(REG3_REG_5_), .Y(_abc_3548_n586) );
  AND2X2 AND2X2_2 ( .A(_abc_3548_n149), .B(STATO_REG_0_), .Y(_abc_3548_n150) );
  AND2X2 AND2X2_20 ( .A(REG4_REG_1_), .B(DATA_IN_1_), .Y(_abc_3548_n190_1) );
  AND2X2 AND2X2_200 ( .A(_abc_3548_n147_1), .B(REG2_REG_5_), .Y(_abc_3548_n587) );
  AND2X2 AND2X2_201 ( .A(_abc_3548_n302_1), .B(REG3_REG_6_), .Y(_abc_3548_n590) );
  AND2X2 AND2X2_202 ( .A(_abc_3548_n147_1), .B(REG2_REG_6_), .Y(_abc_3548_n591) );
  AND2X2 AND2X2_203 ( .A(_abc_3548_n302_1), .B(REG3_REG_7_), .Y(_abc_3548_n594) );
  AND2X2 AND2X2_204 ( .A(_abc_3548_n147_1), .B(REG2_REG_7_), .Y(_abc_3548_n595) );
  AND2X2 AND2X2_205 ( .A(_abc_3548_n302_1), .B(REG2_REG_0_), .Y(_abc_3548_n598) );
  AND2X2 AND2X2_206 ( .A(_abc_3548_n147_1), .B(REG1_REG_0_), .Y(_abc_3548_n599) );
  AND2X2 AND2X2_207 ( .A(_abc_3548_n302_1), .B(REG2_REG_1_), .Y(_abc_3548_n602) );
  AND2X2 AND2X2_208 ( .A(_abc_3548_n147_1), .B(REG1_REG_1_), .Y(_abc_3548_n603) );
  AND2X2 AND2X2_209 ( .A(_abc_3548_n302_1), .B(REG2_REG_2_), .Y(_abc_3548_n606) );
  AND2X2 AND2X2_21 ( .A(REG4_REG_0_), .B(DATA_IN_0_), .Y(_abc_3548_n191) );
  AND2X2 AND2X2_210 ( .A(_abc_3548_n147_1), .B(REG1_REG_2_), .Y(_abc_3548_n607) );
  AND2X2 AND2X2_211 ( .A(_abc_3548_n302_1), .B(REG2_REG_3_), .Y(_abc_3548_n610) );
  AND2X2 AND2X2_212 ( .A(_abc_3548_n147_1), .B(REG1_REG_3_), .Y(_abc_3548_n611) );
  AND2X2 AND2X2_213 ( .A(_abc_3548_n302_1), .B(REG2_REG_4_), .Y(_abc_3548_n614) );
  AND2X2 AND2X2_214 ( .A(_abc_3548_n147_1), .B(REG1_REG_4_), .Y(_abc_3548_n615) );
  AND2X2 AND2X2_215 ( .A(_abc_3548_n302_1), .B(REG2_REG_5_), .Y(_abc_3548_n618) );
  AND2X2 AND2X2_216 ( .A(_abc_3548_n147_1), .B(REG1_REG_5_), .Y(_abc_3548_n619) );
  AND2X2 AND2X2_217 ( .A(_abc_3548_n302_1), .B(REG2_REG_6_), .Y(_abc_3548_n622) );
  AND2X2 AND2X2_218 ( .A(_abc_3548_n147_1), .B(REG1_REG_6_), .Y(_abc_3548_n623) );
  AND2X2 AND2X2_219 ( .A(_abc_3548_n302_1), .B(REG2_REG_7_), .Y(_abc_3548_n626) );
  AND2X2 AND2X2_22 ( .A(_abc_3548_n193), .B(_abc_3548_n194), .Y(_abc_3548_n195) );
  AND2X2 AND2X2_220 ( .A(_abc_3548_n147_1), .B(REG1_REG_7_), .Y(_abc_3548_n627) );
  AND2X2 AND2X2_221 ( .A(_abc_3548_n302_1), .B(REG1_REG_0_), .Y(_abc_3548_n630) );
  AND2X2 AND2X2_222 ( .A(_abc_3548_n147_1), .B(DATA_IN_0_), .Y(_abc_3548_n631) );
  AND2X2 AND2X2_223 ( .A(_abc_3548_n302_1), .B(REG1_REG_1_), .Y(_abc_3548_n634) );
  AND2X2 AND2X2_224 ( .A(_abc_3548_n147_1), .B(DATA_IN_1_), .Y(_abc_3548_n635) );
  AND2X2 AND2X2_225 ( .A(_abc_3548_n302_1), .B(REG1_REG_2_), .Y(_abc_3548_n638) );
  AND2X2 AND2X2_226 ( .A(_abc_3548_n147_1), .B(DATA_IN_2_), .Y(_abc_3548_n639) );
  AND2X2 AND2X2_227 ( .A(_abc_3548_n302_1), .B(REG1_REG_3_), .Y(_abc_3548_n642) );
  AND2X2 AND2X2_228 ( .A(_abc_3548_n147_1), .B(DATA_IN_3_), .Y(_abc_3548_n643) );
  AND2X2 AND2X2_229 ( .A(_abc_3548_n302_1), .B(REG1_REG_4_), .Y(_abc_3548_n646) );
  AND2X2 AND2X2_23 ( .A(_abc_3548_n192), .B(_abc_3548_n195), .Y(_abc_3548_n196) );
  AND2X2 AND2X2_230 ( .A(_abc_3548_n147_1), .B(DATA_IN_4_), .Y(_abc_3548_n647) );
  AND2X2 AND2X2_231 ( .A(_abc_3548_n302_1), .B(REG1_REG_5_), .Y(_abc_3548_n650) );
  AND2X2 AND2X2_232 ( .A(_abc_3548_n147_1), .B(DATA_IN_5_), .Y(_abc_3548_n651) );
  AND2X2 AND2X2_233 ( .A(_abc_3548_n302_1), .B(REG1_REG_6_), .Y(_abc_3548_n654) );
  AND2X2 AND2X2_234 ( .A(_abc_3548_n147_1), .B(DATA_IN_6_), .Y(_abc_3548_n655) );
  AND2X2 AND2X2_235 ( .A(_abc_3548_n302_1), .B(REG1_REG_7_), .Y(_abc_3548_n658) );
  AND2X2 AND2X2_236 ( .A(_abc_3548_n147_1), .B(DATA_IN_7_), .Y(_abc_3548_n659) );
  AND2X2 AND2X2_237 ( .A(_abc_3548_n146), .B(_abc_3548_n296), .Y(_abc_3548_n662) );
  AND2X2 AND2X2_238 ( .A(_abc_3548_n663), .B(STATO_REG_1_), .Y(_abc_3548_n664) );
  AND2X2 AND2X2_239 ( .A(_abc_3548_n664), .B(DATA_IN_0_), .Y(_abc_3548_n665) );
  AND2X2 AND2X2_24 ( .A(REG4_REG_3_), .B(DATA_IN_3_), .Y(_abc_3548_n197) );
  AND2X2 AND2X2_240 ( .A(_abc_3548_n149), .B(_abc_3548_n146), .Y(_abc_3548_n666) );
  AND2X2 AND2X2_241 ( .A(_abc_3548_n667), .B(RLAST_REG_0_), .Y(_abc_3548_n668) );
  AND2X2 AND2X2_242 ( .A(_abc_3548_n664), .B(DATA_IN_1_), .Y(_abc_3548_n671) );
  AND2X2 AND2X2_243 ( .A(_abc_3548_n667), .B(RLAST_REG_1_), .Y(_abc_3548_n672) );
  AND2X2 AND2X2_244 ( .A(_abc_3548_n664), .B(DATA_IN_2_), .Y(_abc_3548_n675) );
  AND2X2 AND2X2_245 ( .A(_abc_3548_n667), .B(RLAST_REG_2_), .Y(_abc_3548_n676) );
  AND2X2 AND2X2_246 ( .A(_abc_3548_n664), .B(DATA_IN_3_), .Y(_abc_3548_n679) );
  AND2X2 AND2X2_247 ( .A(_abc_3548_n667), .B(RLAST_REG_3_), .Y(_abc_3548_n680) );
  AND2X2 AND2X2_248 ( .A(_abc_3548_n664), .B(DATA_IN_4_), .Y(_abc_3548_n683) );
  AND2X2 AND2X2_249 ( .A(_abc_3548_n667), .B(RLAST_REG_4_), .Y(_abc_3548_n684) );
  AND2X2 AND2X2_25 ( .A(REG4_REG_2_), .B(DATA_IN_2_), .Y(_abc_3548_n198) );
  AND2X2 AND2X2_250 ( .A(_abc_3548_n664), .B(DATA_IN_5_), .Y(_abc_3548_n687) );
  AND2X2 AND2X2_251 ( .A(_abc_3548_n667), .B(RLAST_REG_5_), .Y(_abc_3548_n688) );
  AND2X2 AND2X2_252 ( .A(_abc_3548_n664), .B(DATA_IN_6_), .Y(_abc_3548_n691) );
  AND2X2 AND2X2_253 ( .A(_abc_3548_n667), .B(RLAST_REG_6_), .Y(_abc_3548_n692) );
  AND2X2 AND2X2_254 ( .A(_abc_3548_n664), .B(DATA_IN_7_), .Y(_abc_3548_n695) );
  AND2X2 AND2X2_255 ( .A(_abc_3548_n667), .B(RLAST_REG_7_), .Y(_abc_3548_n696) );
  AND2X2 AND2X2_256 ( .A(_abc_3548_n699), .B(RMAX_REG_7_), .Y(_abc_3548_n700) );
  AND2X2 AND2X2_257 ( .A(_abc_3548_n702), .B(DATA_IN_2_), .Y(_abc_3548_n703) );
  AND2X2 AND2X2_258 ( .A(_abc_3548_n705), .B(RMAX_REG_1_), .Y(_abc_3548_n706) );
  AND2X2 AND2X2_259 ( .A(_abc_3548_n173), .B(DATA_IN_0_), .Y(_abc_3548_n708) );
  AND2X2 AND2X2_26 ( .A(_abc_3548_n201), .B(_abc_3548_n202), .Y(_abc_3548_n203) );
  AND2X2 AND2X2_260 ( .A(_abc_3548_n709), .B(_abc_3548_n707), .Y(_abc_3548_n710) );
  AND2X2 AND2X2_261 ( .A(_abc_3548_n711), .B(_abc_3548_n704), .Y(_abc_3548_n712) );
  AND2X2 AND2X2_262 ( .A(_abc_3548_n202), .B(RMAX_REG_3_), .Y(_abc_3548_n713) );
  AND2X2 AND2X2_263 ( .A(_abc_3548_n714), .B(RMAX_REG_2_), .Y(_abc_3548_n715) );
  AND2X2 AND2X2_264 ( .A(_abc_3548_n253_1), .B(DATA_IN_4_), .Y(_abc_3548_n718) );
  AND2X2 AND2X2_265 ( .A(_abc_3548_n251), .B(DATA_IN_3_), .Y(_abc_3548_n719) );
  AND2X2 AND2X2_266 ( .A(_abc_3548_n717), .B(_abc_3548_n721), .Y(_abc_3548_n722) );
  AND2X2 AND2X2_267 ( .A(_abc_3548_n215), .B(RMAX_REG_5_), .Y(_abc_3548_n723) );
  AND2X2 AND2X2_268 ( .A(_abc_3548_n204), .B(RMAX_REG_4_), .Y(_abc_3548_n724) );
  AND2X2 AND2X2_269 ( .A(_abc_3548_n266), .B(DATA_IN_6_), .Y(_abc_3548_n727) );
  AND2X2 AND2X2_27 ( .A(_abc_3548_n204), .B(_abc_3548_n205), .Y(_abc_3548_n206) );
  AND2X2 AND2X2_270 ( .A(_abc_3548_n264), .B(DATA_IN_5_), .Y(_abc_3548_n728) );
  AND2X2 AND2X2_271 ( .A(_abc_3548_n726), .B(_abc_3548_n730), .Y(_abc_3548_n731) );
  AND2X2 AND2X2_272 ( .A(_abc_3548_n217), .B(RMAX_REG_6_), .Y(_abc_3548_n732) );
  AND2X2 AND2X2_273 ( .A(_abc_3548_n274), .B(DATA_IN_7_), .Y(_abc_3548_n733) );
  AND2X2 AND2X2_274 ( .A(_abc_3548_n735), .B(_abc_3548_n701), .Y(_abc_3548_n736) );
  AND2X2 AND2X2_275 ( .A(_abc_3548_n275_1), .B(DATA_IN_7_), .Y(_abc_3548_n737) );
  AND2X2 AND2X2_276 ( .A(_abc_3548_n714), .B(RMIN_REG_2_), .Y(_abc_3548_n738) );
  AND2X2 AND2X2_277 ( .A(_abc_3548_n705), .B(RMIN_REG_1_), .Y(_abc_3548_n739) );
  AND2X2 AND2X2_278 ( .A(_abc_3548_n154), .B(DATA_IN_1_), .Y(_abc_3548_n741) );
  AND2X2 AND2X2_279 ( .A(_abc_3548_n171), .B(RMIN_REG_0_), .Y(_abc_3548_n743) );
  AND2X2 AND2X2_28 ( .A(_abc_3548_n200), .B(_abc_3548_n208), .Y(_abc_3548_n209_1) );
  AND2X2 AND2X2_280 ( .A(_abc_3548_n742), .B(_abc_3548_n743), .Y(_abc_3548_n744) );
  AND2X2 AND2X2_281 ( .A(_abc_3548_n250), .B(DATA_IN_3_), .Y(_abc_3548_n746) );
  AND2X2 AND2X2_282 ( .A(_abc_3548_n747), .B(_abc_3548_n748), .Y(_abc_3548_n749) );
  AND2X2 AND2X2_283 ( .A(_abc_3548_n745), .B(_abc_3548_n749), .Y(_abc_3548_n750) );
  AND2X2 AND2X2_284 ( .A(_abc_3548_n204), .B(RMIN_REG_4_), .Y(_abc_3548_n751) );
  AND2X2 AND2X2_285 ( .A(_abc_3548_n202), .B(RMIN_REG_3_), .Y(_abc_3548_n752) );
  AND2X2 AND2X2_286 ( .A(_abc_3548_n263_1), .B(DATA_IN_5_), .Y(_abc_3548_n755) );
  AND2X2 AND2X2_287 ( .A(_abc_3548_n254), .B(DATA_IN_4_), .Y(_abc_3548_n756) );
  AND2X2 AND2X2_288 ( .A(_abc_3548_n754), .B(_abc_3548_n758), .Y(_abc_3548_n759) );
  AND2X2 AND2X2_289 ( .A(_abc_3548_n217), .B(RMIN_REG_6_), .Y(_abc_3548_n760) );
  AND2X2 AND2X2_29 ( .A(REG4_REG_5_), .B(DATA_IN_5_), .Y(_abc_3548_n210) );
  AND2X2 AND2X2_290 ( .A(_abc_3548_n215), .B(RMIN_REG_5_), .Y(_abc_3548_n761) );
  AND2X2 AND2X2_291 ( .A(_abc_3548_n267), .B(DATA_IN_6_), .Y(_abc_3548_n764) );
  AND2X2 AND2X2_292 ( .A(_abc_3548_n699), .B(RMIN_REG_7_), .Y(_abc_3548_n765) );
  AND2X2 AND2X2_293 ( .A(_abc_3548_n763), .B(_abc_3548_n767), .Y(_abc_3548_n768) );
  AND2X2 AND2X2_294 ( .A(_abc_3548_n769), .B(STATO_REG_1_), .Y(_abc_3548_n770) );
  AND2X2 AND2X2_295 ( .A(_abc_3548_n770), .B(_abc_3548_n736), .Y(_abc_3548_n771) );
  AND2X2 AND2X2_296 ( .A(_abc_3548_n773), .B(RMIN_REG_0_), .Y(_abc_3548_n774) );
  AND2X2 AND2X2_297 ( .A(_abc_3548_n772), .B(DATA_IN_0_), .Y(_abc_3548_n775) );
  AND2X2 AND2X2_298 ( .A(_abc_3548_n773), .B(RMIN_REG_1_), .Y(_abc_3548_n778) );
  AND2X2 AND2X2_299 ( .A(_abc_3548_n772), .B(DATA_IN_1_), .Y(_abc_3548_n779) );
  AND2X2 AND2X2_3 ( .A(_abc_3548_n154), .B(RESTART), .Y(_abc_3548_n155) );
  AND2X2 AND2X2_30 ( .A(DATA_IN_4_), .B(REG4_REG_4_), .Y(_abc_3548_n211_1) );
  AND2X2 AND2X2_300 ( .A(_abc_3548_n773), .B(RMIN_REG_2_), .Y(_abc_3548_n782) );
  AND2X2 AND2X2_301 ( .A(_abc_3548_n772), .B(DATA_IN_2_), .Y(_abc_3548_n783) );
  AND2X2 AND2X2_302 ( .A(_abc_3548_n773), .B(RMIN_REG_3_), .Y(_abc_3548_n786) );
  AND2X2 AND2X2_303 ( .A(_abc_3548_n772), .B(DATA_IN_3_), .Y(_abc_3548_n787) );
  AND2X2 AND2X2_304 ( .A(_abc_3548_n773), .B(RMIN_REG_4_), .Y(_abc_3548_n790) );
  AND2X2 AND2X2_305 ( .A(_abc_3548_n772), .B(DATA_IN_4_), .Y(_abc_3548_n791) );
  AND2X2 AND2X2_306 ( .A(_abc_3548_n773), .B(RMIN_REG_5_), .Y(_abc_3548_n794) );
  AND2X2 AND2X2_307 ( .A(_abc_3548_n772), .B(DATA_IN_5_), .Y(_abc_3548_n795) );
  AND2X2 AND2X2_308 ( .A(_abc_3548_n773), .B(RMIN_REG_6_), .Y(_abc_3548_n798) );
  AND2X2 AND2X2_309 ( .A(_abc_3548_n772), .B(DATA_IN_6_), .Y(_abc_3548_n799) );
  AND2X2 AND2X2_31 ( .A(_abc_3548_n214), .B(_abc_3548_n215), .Y(_abc_3548_n216) );
  AND2X2 AND2X2_310 ( .A(_abc_3548_n773), .B(RMIN_REG_7_), .Y(_abc_3548_n802) );
  AND2X2 AND2X2_311 ( .A(_abc_3548_n772), .B(DATA_IN_7_), .Y(_abc_3548_n803) );
  AND2X2 AND2X2_312 ( .A(_abc_3548_n806), .B(_abc_3548_n146), .Y(_abc_3548_n807) );
  AND2X2 AND2X2_313 ( .A(_abc_3548_n808), .B(DATA_IN_0_), .Y(_abc_3548_n809) );
  AND2X2 AND2X2_314 ( .A(_abc_3548_n807), .B(RMAX_REG_0_), .Y(_abc_3548_n810) );
  AND2X2 AND2X2_315 ( .A(_abc_3548_n808), .B(DATA_IN_1_), .Y(_abc_3548_n813) );
  AND2X2 AND2X2_316 ( .A(_abc_3548_n807), .B(RMAX_REG_1_), .Y(_abc_3548_n814) );
  AND2X2 AND2X2_317 ( .A(_abc_3548_n808), .B(DATA_IN_2_), .Y(_abc_3548_n817) );
  AND2X2 AND2X2_318 ( .A(_abc_3548_n807), .B(RMAX_REG_2_), .Y(_abc_3548_n818) );
  AND2X2 AND2X2_319 ( .A(_abc_3548_n808), .B(DATA_IN_3_), .Y(_abc_3548_n821) );
  AND2X2 AND2X2_32 ( .A(_abc_3548_n217), .B(_abc_3548_n218_1), .Y(_abc_3548_n219) );
  AND2X2 AND2X2_320 ( .A(_abc_3548_n807), .B(RMAX_REG_3_), .Y(_abc_3548_n822) );
  AND2X2 AND2X2_321 ( .A(_abc_3548_n808), .B(DATA_IN_4_), .Y(_abc_3548_n825) );
  AND2X2 AND2X2_322 ( .A(_abc_3548_n807), .B(RMAX_REG_4_), .Y(_abc_3548_n826) );
  AND2X2 AND2X2_323 ( .A(_abc_3548_n808), .B(DATA_IN_5_), .Y(_abc_3548_n829) );
  AND2X2 AND2X2_324 ( .A(_abc_3548_n807), .B(RMAX_REG_5_), .Y(_abc_3548_n830) );
  AND2X2 AND2X2_325 ( .A(_abc_3548_n808), .B(DATA_IN_6_), .Y(_abc_3548_n833) );
  AND2X2 AND2X2_326 ( .A(_abc_3548_n807), .B(RMAX_REG_6_), .Y(_abc_3548_n834) );
  AND2X2 AND2X2_327 ( .A(_abc_3548_n808), .B(DATA_IN_7_), .Y(_abc_3548_n837) );
  AND2X2 AND2X2_328 ( .A(_abc_3548_n807), .B(RMAX_REG_7_), .Y(_abc_3548_n838) );
  AND2X2 AND2X2_329 ( .A(_abc_3548_n666), .B(_abc_3548_n841), .Y(n361) );
  AND2X2 AND2X2_33 ( .A(_abc_3548_n213), .B(_abc_3548_n221), .Y(_abc_3548_n222) );
  AND2X2 AND2X2_34 ( .A(DATA_IN_6_), .B(REG4_REG_6_), .Y(_abc_3548_n225) );
  AND2X2 AND2X2_35 ( .A(_abc_3548_n226), .B(_abc_3548_n224), .Y(_abc_3548_n227) );
  AND2X2 AND2X2_36 ( .A(_abc_3548_n223), .B(_abc_3548_n227), .Y(_abc_3548_n228) );
  AND2X2 AND2X2_37 ( .A(_abc_3548_n231), .B(ENABLE), .Y(_abc_3548_n232) );
  AND2X2 AND2X2_38 ( .A(_abc_3548_n230), .B(_abc_3548_n232), .Y(_abc_3548_n233) );
  AND2X2 AND2X2_39 ( .A(n356), .B(STATO_REG_1_), .Y(_abc_3548_n235) );
  AND2X2 AND2X2_4 ( .A(_abc_3548_n156), .B(_abc_3548_n153), .Y(_abc_3548_n157) );
  AND2X2 AND2X2_40 ( .A(RMAX_REG_7_), .B(RMIN_REG_7_), .Y(_abc_3548_n236) );
  AND2X2 AND2X2_41 ( .A(RMAX_REG_6_), .B(RMIN_REG_6_), .Y(_abc_3548_n238) );
  AND2X2 AND2X2_42 ( .A(RMIN_REG_1_), .B(RMAX_REG_1_), .Y(_abc_3548_n239_1) );
  AND2X2 AND2X2_43 ( .A(RMIN_REG_0_), .B(RMAX_REG_0_), .Y(_abc_3548_n240) );
  AND2X2 AND2X2_44 ( .A(_abc_3548_n242), .B(_abc_3548_n243), .Y(_abc_3548_n244) );
  AND2X2 AND2X2_45 ( .A(_abc_3548_n241_1), .B(_abc_3548_n244), .Y(_abc_3548_n245) );
  AND2X2 AND2X2_46 ( .A(RMIN_REG_3_), .B(RMAX_REG_3_), .Y(_abc_3548_n246) );
  AND2X2 AND2X2_47 ( .A(RMIN_REG_2_), .B(RMAX_REG_2_), .Y(_abc_3548_n247) );
  AND2X2 AND2X2_48 ( .A(_abc_3548_n250), .B(_abc_3548_n251), .Y(_abc_3548_n252) );
  AND2X2 AND2X2_49 ( .A(_abc_3548_n253_1), .B(_abc_3548_n254), .Y(_abc_3548_n255_1) );
  AND2X2 AND2X2_5 ( .A(_abc_3548_n160), .B(_abc_3548_n158), .Y(_abc_3548_n161) );
  AND2X2 AND2X2_50 ( .A(_abc_3548_n249), .B(_abc_3548_n257), .Y(_abc_3548_n258) );
  AND2X2 AND2X2_51 ( .A(RMIN_REG_5_), .B(RMAX_REG_5_), .Y(_abc_3548_n259) );
  AND2X2 AND2X2_52 ( .A(RMAX_REG_4_), .B(RMIN_REG_4_), .Y(_abc_3548_n260_1) );
  AND2X2 AND2X2_53 ( .A(_abc_3548_n263_1), .B(_abc_3548_n264), .Y(_abc_3548_n265_1) );
  AND2X2 AND2X2_54 ( .A(_abc_3548_n266), .B(_abc_3548_n267), .Y(_abc_3548_n268) );
  AND2X2 AND2X2_55 ( .A(_abc_3548_n262), .B(_abc_3548_n270_1), .Y(_abc_3548_n271) );
  AND2X2 AND2X2_56 ( .A(_abc_3548_n272_1), .B(_abc_3548_n237), .Y(_abc_3548_n273) );
  AND2X2 AND2X2_57 ( .A(_abc_3548_n274), .B(_abc_3548_n275_1), .Y(_abc_3548_n276) );
  AND2X2 AND2X2_58 ( .A(_abc_3548_n278), .B(_abc_3548_n235), .Y(_abc_3548_n279_1) );
  AND2X2 AND2X2_59 ( .A(_abc_3548_n234), .B(_abc_3548_n279_1), .Y(_abc_3548_n280_1) );
  AND2X2 AND2X2_6 ( .A(_abc_3548_n159), .B(REG4_REG_0_), .Y(_abc_3548_n162_1) );
  AND2X2 AND2X2_60 ( .A(_abc_3548_n280_1), .B(_abc_3548_n188), .Y(_abc_3548_n281) );
  AND2X2 AND2X2_61 ( .A(_abc_3548_n282_1), .B(_abc_3548_n235), .Y(_abc_3548_n283_1) );
  AND2X2 AND2X2_62 ( .A(_abc_3548_n235), .B(_abc_3548_n159), .Y(_abc_3548_n284) );
  AND2X2 AND2X2_63 ( .A(_abc_3548_n284), .B(_abc_3548_n232), .Y(_abc_3548_n285_1) );
  AND2X2 AND2X2_64 ( .A(_abc_3548_n229), .B(_abc_3548_n285_1), .Y(_abc_3548_n286_1) );
  AND2X2 AND2X2_65 ( .A(_abc_3548_n175), .B(_abc_3548_n179_1), .Y(_abc_3548_n288_1) );
  AND2X2 AND2X2_66 ( .A(_abc_3548_n188), .B(_abc_3548_n290_1), .Y(_abc_3548_n291) );
  AND2X2 AND2X2_67 ( .A(_abc_3548_n292), .B(_abc_3548_n293_1), .Y(_abc_3548_n294) );
  AND2X2 AND2X2_68 ( .A(_abc_3548_n287), .B(_abc_3548_n294), .Y(_abc_3548_n295_1) );
  AND2X2 AND2X2_69 ( .A(_abc_3548_n284), .B(_abc_3548_n296), .Y(_abc_3548_n297) );
  AND2X2 AND2X2_7 ( .A(RMIN_REG_0_), .B(RESTART), .Y(_abc_3548_n163) );
  AND2X2 AND2X2_70 ( .A(_abc_3548_n297), .B(RLAST_REG_0_), .Y(_abc_3548_n298_1) );
  AND2X2 AND2X2_71 ( .A(ENABLE), .B(AVERAGE), .Y(_abc_3548_n299_1) );
  AND2X2 AND2X2_72 ( .A(_abc_3548_n284), .B(_abc_3548_n299_1), .Y(_abc_3548_n300) );
  AND2X2 AND2X2_73 ( .A(_abc_3548_n300), .B(REG4_REG_0_), .Y(_abc_3548_n301_1) );
  AND2X2 AND2X2_74 ( .A(_abc_3548_n302_1), .B(DATA_OUT_REG_0_), .Y(_abc_3548_n303) );
  AND2X2 AND2X2_75 ( .A(_abc_3548_n310), .B(_abc_3548_n309_1), .Y(_abc_3548_n311_1) );
  AND2X2 AND2X2_76 ( .A(_abc_3548_n314_1), .B(_abc_3548_n313), .Y(_abc_3548_n315) );
  AND2X2 AND2X2_77 ( .A(_abc_3548_n312), .B(_abc_3548_n316_1), .Y(_abc_3548_n317) );
  AND2X2 AND2X2_78 ( .A(_abc_3548_n311_1), .B(_abc_3548_n315), .Y(_abc_3548_n319_1) );
  AND2X2 AND2X2_79 ( .A(_abc_3548_n318), .B(_abc_3548_n320), .Y(_abc_3548_n321_1) );
  AND2X2 AND2X2_8 ( .A(_abc_3548_n161), .B(_abc_3548_n164), .Y(_abc_3548_n165_1) );
  AND2X2 AND2X2_80 ( .A(_abc_3548_n323), .B(_abc_3548_n170), .Y(_abc_3548_n324_1) );
  AND2X2 AND2X2_81 ( .A(_abc_3548_n324_1), .B(_abc_3548_n321_1), .Y(_abc_3548_n325_1) );
  AND2X2 AND2X2_82 ( .A(_abc_3548_n327_1), .B(_abc_3548_n183), .Y(_abc_3548_n328_1) );
  AND2X2 AND2X2_83 ( .A(_abc_3548_n328_1), .B(_abc_3548_n326), .Y(_abc_3548_n329) );
  AND2X2 AND2X2_84 ( .A(_abc_3548_n291), .B(_abc_3548_n330_1), .Y(_abc_3548_n331) );
  AND2X2 AND2X2_85 ( .A(_abc_3548_n332_1), .B(_abc_3548_n333), .Y(_abc_3548_n334) );
  AND2X2 AND2X2_86 ( .A(_abc_3548_n287), .B(_abc_3548_n334), .Y(_abc_3548_n335_1) );
  AND2X2 AND2X2_87 ( .A(_abc_3548_n280_1), .B(_abc_3548_n330_1), .Y(_abc_3548_n336) );
  AND2X2 AND2X2_88 ( .A(_abc_3548_n300), .B(REG4_REG_1_), .Y(_abc_3548_n337_1) );
  AND2X2 AND2X2_89 ( .A(_abc_3548_n297), .B(RLAST_REG_1_), .Y(_abc_3548_n338) );
  AND2X2 AND2X2_9 ( .A(RESTART), .B(RMAX_REG_1_), .Y(_abc_3548_n166) );
  AND2X2 AND2X2_90 ( .A(_abc_3548_n302_1), .B(DATA_OUT_REG_1_), .Y(_abc_3548_n339) );
  AND2X2 AND2X2_91 ( .A(_abc_3548_n328_1), .B(_abc_3548_n318), .Y(_abc_3548_n348) );
  AND2X2 AND2X2_92 ( .A(_abc_3548_n351), .B(_abc_3548_n350_1), .Y(_abc_3548_n352_1) );
  AND2X2 AND2X2_93 ( .A(_abc_3548_n354_1), .B(_abc_3548_n353), .Y(_abc_3548_n355) );
  AND2X2 AND2X2_94 ( .A(_abc_3548_n352_1), .B(_abc_3548_n355), .Y(_abc_3548_n356) );
  AND2X2 AND2X2_95 ( .A(_abc_3548_n357_1), .B(_abc_3548_n358), .Y(_abc_3548_n359_1) );
  AND2X2 AND2X2_96 ( .A(_abc_3548_n349_1), .B(_abc_3548_n360), .Y(_abc_3548_n361) );
  AND2X2 AND2X2_97 ( .A(_abc_3548_n362_1), .B(_abc_3548_n320), .Y(_abc_3548_n363_1) );
  AND2X2 AND2X2_98 ( .A(_abc_3548_n363_1), .B(_abc_3548_n359_1), .Y(_abc_3548_n364) );
  AND2X2 AND2X2_99 ( .A(_abc_3548_n346_1), .B(_abc_3548_n366), .Y(_abc_3548_n367_1) );
  DFFPOSX1 DFFPOSX1_1 ( .CLK(clock), .D(n324), .Q(DATA_OUT_REG_7_) );
  DFFPOSX1 DFFPOSX1_10 ( .CLK(clock), .D(n49), .Q(RMAX_REG_6_) );
  DFFPOSX1 DFFPOSX1_11 ( .CLK(clock), .D(n54), .Q(RMAX_REG_5_) );
  DFFPOSX1 DFFPOSX1_12 ( .CLK(clock), .D(n59), .Q(RMAX_REG_4_) );
  DFFPOSX1 DFFPOSX1_13 ( .CLK(clock), .D(n64), .Q(RMAX_REG_3_) );
  DFFPOSX1 DFFPOSX1_14 ( .CLK(clock), .D(n69), .Q(RMAX_REG_2_) );
  DFFPOSX1 DFFPOSX1_15 ( .CLK(clock), .D(n74), .Q(RMAX_REG_1_) );
  DFFPOSX1 DFFPOSX1_16 ( .CLK(clock), .D(n79), .Q(RMAX_REG_0_) );
  DFFPOSX1 DFFPOSX1_17 ( .CLK(clock), .D(n84), .Q(RMIN_REG_7_) );
  DFFPOSX1 DFFPOSX1_18 ( .CLK(clock), .D(n89), .Q(RMIN_REG_6_) );
  DFFPOSX1 DFFPOSX1_19 ( .CLK(clock), .D(n94), .Q(RMIN_REG_5_) );
  DFFPOSX1 DFFPOSX1_2 ( .CLK(clock), .D(n328), .Q(DATA_OUT_REG_6_) );
  DFFPOSX1 DFFPOSX1_20 ( .CLK(clock), .D(n99), .Q(RMIN_REG_4_) );
  DFFPOSX1 DFFPOSX1_21 ( .CLK(clock), .D(n104), .Q(RMIN_REG_3_) );
  DFFPOSX1 DFFPOSX1_22 ( .CLK(clock), .D(n109), .Q(RMIN_REG_2_) );
  DFFPOSX1 DFFPOSX1_23 ( .CLK(clock), .D(n114), .Q(RMIN_REG_1_) );
  DFFPOSX1 DFFPOSX1_24 ( .CLK(clock), .D(n119), .Q(RMIN_REG_0_) );
  DFFPOSX1 DFFPOSX1_25 ( .CLK(clock), .D(n124), .Q(RLAST_REG_7_) );
  DFFPOSX1 DFFPOSX1_26 ( .CLK(clock), .D(n129), .Q(RLAST_REG_6_) );
  DFFPOSX1 DFFPOSX1_27 ( .CLK(clock), .D(n134), .Q(RLAST_REG_5_) );
  DFFPOSX1 DFFPOSX1_28 ( .CLK(clock), .D(n139), .Q(RLAST_REG_4_) );
  DFFPOSX1 DFFPOSX1_29 ( .CLK(clock), .D(n144), .Q(RLAST_REG_3_) );
  DFFPOSX1 DFFPOSX1_3 ( .CLK(clock), .D(n332), .Q(DATA_OUT_REG_5_) );
  DFFPOSX1 DFFPOSX1_30 ( .CLK(clock), .D(n149), .Q(RLAST_REG_2_) );
  DFFPOSX1 DFFPOSX1_31 ( .CLK(clock), .D(n154), .Q(RLAST_REG_1_) );
  DFFPOSX1 DFFPOSX1_32 ( .CLK(clock), .D(n159), .Q(RLAST_REG_0_) );
  DFFPOSX1 DFFPOSX1_33 ( .CLK(clock), .D(n164), .Q(REG1_REG_7_) );
  DFFPOSX1 DFFPOSX1_34 ( .CLK(clock), .D(n169), .Q(REG1_REG_6_) );
  DFFPOSX1 DFFPOSX1_35 ( .CLK(clock), .D(n174), .Q(REG1_REG_5_) );
  DFFPOSX1 DFFPOSX1_36 ( .CLK(clock), .D(n179), .Q(REG1_REG_4_) );
  DFFPOSX1 DFFPOSX1_37 ( .CLK(clock), .D(n184), .Q(REG1_REG_3_) );
  DFFPOSX1 DFFPOSX1_38 ( .CLK(clock), .D(n189), .Q(REG1_REG_2_) );
  DFFPOSX1 DFFPOSX1_39 ( .CLK(clock), .D(n194), .Q(REG1_REG_1_) );
  DFFPOSX1 DFFPOSX1_4 ( .CLK(clock), .D(n336), .Q(DATA_OUT_REG_4_) );
  DFFPOSX1 DFFPOSX1_40 ( .CLK(clock), .D(n199), .Q(REG1_REG_0_) );
  DFFPOSX1 DFFPOSX1_41 ( .CLK(clock), .D(n204), .Q(REG2_REG_7_) );
  DFFPOSX1 DFFPOSX1_42 ( .CLK(clock), .D(n209), .Q(REG2_REG_6_) );
  DFFPOSX1 DFFPOSX1_43 ( .CLK(clock), .D(n214), .Q(REG2_REG_5_) );
  DFFPOSX1 DFFPOSX1_44 ( .CLK(clock), .D(n219), .Q(REG2_REG_4_) );
  DFFPOSX1 DFFPOSX1_45 ( .CLK(clock), .D(n224), .Q(REG2_REG_3_) );
  DFFPOSX1 DFFPOSX1_46 ( .CLK(clock), .D(n229), .Q(REG2_REG_2_) );
  DFFPOSX1 DFFPOSX1_47 ( .CLK(clock), .D(n234), .Q(REG2_REG_1_) );
  DFFPOSX1 DFFPOSX1_48 ( .CLK(clock), .D(n239), .Q(REG2_REG_0_) );
  DFFPOSX1 DFFPOSX1_49 ( .CLK(clock), .D(n244), .Q(REG3_REG_7_) );
  DFFPOSX1 DFFPOSX1_5 ( .CLK(clock), .D(n340), .Q(DATA_OUT_REG_3_) );
  DFFPOSX1 DFFPOSX1_50 ( .CLK(clock), .D(n249), .Q(REG3_REG_6_) );
  DFFPOSX1 DFFPOSX1_51 ( .CLK(clock), .D(n254), .Q(REG3_REG_5_) );
  DFFPOSX1 DFFPOSX1_52 ( .CLK(clock), .D(n259), .Q(REG3_REG_4_) );
  DFFPOSX1 DFFPOSX1_53 ( .CLK(clock), .D(n264), .Q(REG3_REG_3_) );
  DFFPOSX1 DFFPOSX1_54 ( .CLK(clock), .D(n269), .Q(REG3_REG_2_) );
  DFFPOSX1 DFFPOSX1_55 ( .CLK(clock), .D(n274), .Q(REG3_REG_1_) );
  DFFPOSX1 DFFPOSX1_56 ( .CLK(clock), .D(n279), .Q(REG3_REG_0_) );
  DFFPOSX1 DFFPOSX1_57 ( .CLK(clock), .D(n284), .Q(REG4_REG_7_) );
  DFFPOSX1 DFFPOSX1_58 ( .CLK(clock), .D(n289), .Q(REG4_REG_6_) );
  DFFPOSX1 DFFPOSX1_59 ( .CLK(clock), .D(n294), .Q(REG4_REG_5_) );
  DFFPOSX1 DFFPOSX1_6 ( .CLK(clock), .D(n344), .Q(DATA_OUT_REG_2_) );
  DFFPOSX1 DFFPOSX1_60 ( .CLK(clock), .D(n299), .Q(REG4_REG_4_) );
  DFFPOSX1 DFFPOSX1_61 ( .CLK(clock), .D(n304), .Q(REG4_REG_3_) );
  DFFPOSX1 DFFPOSX1_62 ( .CLK(clock), .D(n309), .Q(REG4_REG_2_) );
  DFFPOSX1 DFFPOSX1_63 ( .CLK(clock), .D(n314), .Q(REG4_REG_1_) );
  DFFPOSX1 DFFPOSX1_64 ( .CLK(clock), .D(n319), .Q(REG4_REG_0_) );
  DFFPOSX1 DFFPOSX1_65 ( .CLK(clock), .D(n356), .Q(STATO_REG_1_) );
  DFFPOSX1 DFFPOSX1_66 ( .CLK(clock), .D(n361), .Q(STATO_REG_0_) );
  DFFPOSX1 DFFPOSX1_7 ( .CLK(clock), .D(n348), .Q(DATA_OUT_REG_1_) );
  DFFPOSX1 DFFPOSX1_8 ( .CLK(clock), .D(n352), .Q(DATA_OUT_REG_0_) );
  DFFPOSX1 DFFPOSX1_9 ( .CLK(clock), .D(n44), .Q(RMAX_REG_7_) );
  INVX1 INVX1_1 ( .A(STATO_REG_0_), .Y(_abc_3548_n146) );
  INVX1 INVX1_10 ( .A(_abc_3548_n168), .Y(_abc_3548_n181) );
  INVX1 INVX1_11 ( .A(_abc_3548_n182_1), .Y(_abc_3548_n183) );
  INVX1 INVX1_12 ( .A(_abc_3548_n186), .Y(_abc_3548_n187) );
  INVX1 INVX1_13 ( .A(REG4_REG_3_), .Y(_abc_3548_n201) );
  INVX1 INVX1_14 ( .A(DATA_IN_3_), .Y(_abc_3548_n202) );
  INVX1 INVX1_15 ( .A(DATA_IN_4_), .Y(_abc_3548_n204) );
  INVX1 INVX1_16 ( .A(REG4_REG_4_), .Y(_abc_3548_n205) );
  INVX1 INVX1_17 ( .A(_abc_3548_n207), .Y(_abc_3548_n208) );
  INVX1 INVX1_18 ( .A(REG4_REG_5_), .Y(_abc_3548_n214) );
  INVX1 INVX1_19 ( .A(DATA_IN_5_), .Y(_abc_3548_n215) );
  INVX1 INVX1_2 ( .A(STATO_REG_1_), .Y(_abc_3548_n149) );
  INVX1 INVX1_20 ( .A(DATA_IN_6_), .Y(_abc_3548_n217) );
  INVX1 INVX1_21 ( .A(REG4_REG_6_), .Y(_abc_3548_n218_1) );
  INVX1 INVX1_22 ( .A(_abc_3548_n220), .Y(_abc_3548_n221) );
  INVX1 INVX1_23 ( .A(_abc_3548_n222), .Y(_abc_3548_n223) );
  INVX1 INVX1_24 ( .A(_abc_3548_n225), .Y(_abc_3548_n226) );
  INVX1 INVX1_25 ( .A(_abc_3548_n229), .Y(_abc_3548_n230) );
  INVX1 INVX1_26 ( .A(AVERAGE), .Y(_abc_3548_n231) );
  INVX1 INVX1_27 ( .A(_abc_3548_n236), .Y(_abc_3548_n237) );
  INVX1 INVX1_28 ( .A(RMIN_REG_3_), .Y(_abc_3548_n250) );
  INVX1 INVX1_29 ( .A(RMAX_REG_3_), .Y(_abc_3548_n251) );
  INVX1 INVX1_3 ( .A(RMIN_REG_1_), .Y(_abc_3548_n154) );
  INVX1 INVX1_30 ( .A(RMAX_REG_4_), .Y(_abc_3548_n253_1) );
  INVX1 INVX1_31 ( .A(RMIN_REG_4_), .Y(_abc_3548_n254) );
  INVX1 INVX1_32 ( .A(_abc_3548_n256), .Y(_abc_3548_n257) );
  INVX1 INVX1_33 ( .A(RMIN_REG_5_), .Y(_abc_3548_n263_1) );
  INVX1 INVX1_34 ( .A(RMAX_REG_5_), .Y(_abc_3548_n264) );
  INVX1 INVX1_35 ( .A(RMAX_REG_6_), .Y(_abc_3548_n266) );
  INVX1 INVX1_36 ( .A(RMIN_REG_6_), .Y(_abc_3548_n267) );
  INVX1 INVX1_37 ( .A(_abc_3548_n269), .Y(_abc_3548_n270_1) );
  INVX1 INVX1_38 ( .A(RMAX_REG_7_), .Y(_abc_3548_n274) );
  INVX1 INVX1_39 ( .A(RMIN_REG_7_), .Y(_abc_3548_n275_1) );
  INVX1 INVX1_4 ( .A(_abc_3548_n155), .Y(_abc_3548_n156) );
  INVX1 INVX1_40 ( .A(_abc_3548_n278), .Y(_abc_3548_n282_1) );
  INVX1 INVX1_41 ( .A(_abc_3548_n289), .Y(_abc_3548_n290_1) );
  INVX1 INVX1_42 ( .A(_abc_3548_n291), .Y(_abc_3548_n292) );
  INVX1 INVX1_43 ( .A(ENABLE), .Y(_abc_3548_n296) );
  INVX1 INVX1_44 ( .A(_abc_3548_n311_1), .Y(_abc_3548_n312) );
  INVX1 INVX1_45 ( .A(_abc_3548_n315), .Y(_abc_3548_n316_1) );
  INVX1 INVX1_46 ( .A(_abc_3548_n317), .Y(_abc_3548_n318) );
  INVX1 INVX1_47 ( .A(_abc_3548_n319_1), .Y(_abc_3548_n320) );
  INVX1 INVX1_48 ( .A(_abc_3548_n157), .Y(_abc_3548_n322) );
  INVX1 INVX1_49 ( .A(_abc_3548_n321_1), .Y(_abc_3548_n326) );
  INVX1 INVX1_5 ( .A(_abc_3548_n169_1), .Y(_abc_3548_n170) );
  INVX1 INVX1_50 ( .A(_abc_3548_n331), .Y(_abc_3548_n332_1) );
  INVX1 INVX1_51 ( .A(_abc_3548_n345), .Y(_abc_3548_n346_1) );
  INVX1 INVX1_52 ( .A(_abc_3548_n356), .Y(_abc_3548_n357_1) );
  INVX1 INVX1_53 ( .A(_abc_3548_n359_1), .Y(_abc_3548_n360) );
  INVX1 INVX1_54 ( .A(_abc_3548_n365_1), .Y(_abc_3548_n366) );
  INVX1 INVX1_55 ( .A(_abc_3548_n370_1), .Y(_abc_3548_n371) );
  INVX1 INVX1_56 ( .A(_abc_3548_n358), .Y(_abc_3548_n384_1) );
  INVX1 INVX1_57 ( .A(_abc_3548_n389), .Y(_abc_3548_n390) );
  INVX1 INVX1_58 ( .A(_abc_3548_n393_1), .Y(_abc_3548_n394) );
  INVX1 INVX1_59 ( .A(_abc_3548_n395), .Y(_abc_3548_n396_1) );
  INVX1 INVX1_6 ( .A(DATA_IN_0_), .Y(_abc_3548_n171) );
  INVX1 INVX1_60 ( .A(_abc_3548_n397), .Y(_abc_3548_n398) );
  INVX1 INVX1_61 ( .A(_abc_3548_n400), .Y(_abc_3548_n401) );
  INVX1 INVX1_62 ( .A(_abc_3548_n367_1), .Y(_abc_3548_n405_1) );
  INVX1 INVX1_63 ( .A(_abc_3548_n402_1), .Y(_abc_3548_n406) );
  INVX1 INVX1_64 ( .A(_abc_3548_n404), .Y(_abc_3548_n411) );
  INVX1 INVX1_65 ( .A(_abc_3548_n428), .Y(_abc_3548_n429) );
  INVX1 INVX1_66 ( .A(_abc_3548_n432), .Y(_abc_3548_n433) );
  INVX1 INVX1_67 ( .A(_abc_3548_n434), .Y(_abc_3548_n435) );
  INVX1 INVX1_68 ( .A(_abc_3548_n436), .Y(_abc_3548_n437) );
  INVX1 INVX1_69 ( .A(_abc_3548_n438), .Y(_abc_3548_n439) );
  INVX1 INVX1_7 ( .A(RMAX_REG_0_), .Y(_abc_3548_n173) );
  INVX1 INVX1_70 ( .A(_abc_3548_n475), .Y(_abc_3548_n476_1) );
  INVX1 INVX1_71 ( .A(_abc_3548_n481), .Y(_abc_3548_n482_1) );
  INVX1 INVX1_72 ( .A(_abc_3548_n483), .Y(_abc_3548_n484_1) );
  INVX1 INVX1_73 ( .A(_abc_3548_n485), .Y(_abc_3548_n486_1) );
  INVX1 INVX1_74 ( .A(_abc_3548_n489), .Y(_abc_3548_n490) );
  INVX1 INVX1_75 ( .A(_abc_3548_n514), .Y(_abc_3548_n524) );
  INVX1 INVX1_76 ( .A(_abc_3548_n662), .Y(_abc_3548_n663) );
  INVX1 INVX1_77 ( .A(DATA_IN_7_), .Y(_abc_3548_n699) );
  INVX1 INVX1_78 ( .A(_abc_3548_n700), .Y(_abc_3548_n701) );
  INVX1 INVX1_79 ( .A(RMAX_REG_2_), .Y(_abc_3548_n702) );
  INVX1 INVX1_8 ( .A(REG4_REG_0_), .Y(_abc_3548_n176) );
  INVX1 INVX1_80 ( .A(_abc_3548_n703), .Y(_abc_3548_n704) );
  INVX1 INVX1_81 ( .A(DATA_IN_1_), .Y(_abc_3548_n705) );
  INVX1 INVX1_82 ( .A(_abc_3548_n708), .Y(_abc_3548_n709) );
  INVX1 INVX1_83 ( .A(DATA_IN_2_), .Y(_abc_3548_n714) );
  INVX1 INVX1_84 ( .A(_abc_3548_n720), .Y(_abc_3548_n721) );
  INVX1 INVX1_85 ( .A(_abc_3548_n729), .Y(_abc_3548_n730) );
  INVX1 INVX1_86 ( .A(_abc_3548_n741), .Y(_abc_3548_n742) );
  INVX1 INVX1_87 ( .A(_abc_3548_n746), .Y(_abc_3548_n747) );
  INVX1 INVX1_88 ( .A(_abc_3548_n757), .Y(_abc_3548_n758) );
  INVX1 INVX1_89 ( .A(_abc_3548_n766), .Y(_abc_3548_n767) );
  INVX1 INVX1_9 ( .A(_abc_3548_n163), .Y(_abc_3548_n178) );
  INVX1 INVX1_90 ( .A(RESET_G), .Y(_abc_3548_n841) );
  INVX2 INVX2_1 ( .A(_abc_3548_n772), .Y(_abc_3548_n773) );
  INVX2 INVX2_2 ( .A(_abc_3548_n807), .Y(_abc_3548_n808) );
  INVX4 INVX4_1 ( .A(RESTART), .Y(_abc_3548_n159) );
  INVX8 INVX8_1 ( .A(nRESET_G), .Y(_abc_3548_n148) );
  INVX8 INVX8_2 ( .A(n356), .Y(_abc_3548_n302_1) );
  OR2X2 OR2X2_1 ( .A(_abc_3548_n150), .B(_abc_3548_n148), .Y(_abc_3548_n151) );
  OR2X2 OR2X2_10 ( .A(_abc_3548_n175), .B(_abc_3548_n179_1), .Y(_abc_3548_n180) );
  OR2X2 OR2X2_100 ( .A(_abc_3548_n452_1), .B(_abc_3548_n148), .Y(_abc_3548_n453) );
  OR2X2 OR2X2_101 ( .A(_abc_3548_n451), .B(_abc_3548_n453), .Y(_abc_3548_n454_1) );
  OR2X2 OR2X2_102 ( .A(_abc_3548_n454_1), .B(_abc_3548_n450), .Y(_abc_3548_n455) );
  OR2X2 OR2X2_103 ( .A(_abc_3548_n449), .B(_abc_3548_n455), .Y(_abc_3548_n456_1) );
  OR2X2 OR2X2_104 ( .A(_abc_3548_n459), .B(_abc_3548_n458_1), .Y(_abc_3548_n460_1) );
  OR2X2 OR2X2_105 ( .A(_abc_3548_n461), .B(_abc_3548_n462), .Y(_abc_3548_n463_1) );
  OR2X2 OR2X2_106 ( .A(_abc_3548_n463_1), .B(_abc_3548_n457), .Y(_abc_3548_n464) );
  OR2X2 OR2X2_107 ( .A(_abc_3548_n448), .B(_abc_3548_n408), .Y(_abc_3548_n465_1) );
  OR2X2 OR2X2_108 ( .A(_abc_3548_n460_1), .B(_abc_3548_n412), .Y(_abc_3548_n466) );
  OR2X2 OR2X2_109 ( .A(_abc_3548_n467_1), .B(_abc_3548_n410), .Y(_abc_3548_n468) );
  OR2X2 OR2X2_11 ( .A(_abc_3548_n184), .B(_abc_3548_n157), .Y(_abc_3548_n185) );
  OR2X2 OR2X2_110 ( .A(_abc_3548_n470_1), .B(_abc_3548_n456_1), .Y(n336) );
  OR2X2 OR2X2_111 ( .A(RESTART), .B(REG4_REG_6_), .Y(_abc_3548_n473) );
  OR2X2 OR2X2_112 ( .A(_abc_3548_n159), .B(RMIN_REG_6_), .Y(_abc_3548_n474_1) );
  OR2X2 OR2X2_113 ( .A(RESTART), .B(DATA_IN_6_), .Y(_abc_3548_n477) );
  OR2X2 OR2X2_114 ( .A(_abc_3548_n159), .B(RMAX_REG_6_), .Y(_abc_3548_n478_1) );
  OR2X2 OR2X2_115 ( .A(_abc_3548_n476_1), .B(_abc_3548_n479), .Y(_abc_3548_n481) );
  OR2X2 OR2X2_116 ( .A(_abc_3548_n482_1), .B(_abc_3548_n480_1), .Y(_abc_3548_n483) );
  OR2X2 OR2X2_117 ( .A(_abc_3548_n472_1), .B(_abc_3548_n486_1), .Y(_abc_3548_n487_1) );
  OR2X2 OR2X2_118 ( .A(_abc_3548_n488), .B(_abc_3548_n490), .Y(_abc_3548_n491) );
  OR2X2 OR2X2_119 ( .A(_abc_3548_n496), .B(_abc_3548_n148), .Y(_abc_3548_n497) );
  OR2X2 OR2X2_12 ( .A(_abc_3548_n190_1), .B(_abc_3548_n191), .Y(_abc_3548_n192) );
  OR2X2 OR2X2_120 ( .A(_abc_3548_n495), .B(_abc_3548_n497), .Y(_abc_3548_n498) );
  OR2X2 OR2X2_121 ( .A(_abc_3548_n498), .B(_abc_3548_n494), .Y(_abc_3548_n499) );
  OR2X2 OR2X2_122 ( .A(_abc_3548_n493), .B(_abc_3548_n499), .Y(_abc_3548_n500) );
  OR2X2 OR2X2_123 ( .A(_abc_3548_n441), .B(_abc_3548_n434), .Y(_abc_3548_n502) );
  OR2X2 OR2X2_124 ( .A(_abc_3548_n446), .B(_abc_3548_n436), .Y(_abc_3548_n504) );
  OR2X2 OR2X2_125 ( .A(_abc_3548_n503), .B(_abc_3548_n505), .Y(_abc_3548_n506) );
  OR2X2 OR2X2_126 ( .A(_abc_3548_n507), .B(_abc_3548_n508), .Y(_abc_3548_n509) );
  OR2X2 OR2X2_127 ( .A(_abc_3548_n509), .B(_abc_3548_n501), .Y(_abc_3548_n510) );
  OR2X2 OR2X2_128 ( .A(_abc_3548_n465_1), .B(_abc_3548_n492), .Y(_abc_3548_n511) );
  OR2X2 OR2X2_129 ( .A(_abc_3548_n506), .B(_abc_3548_n461), .Y(_abc_3548_n512) );
  OR2X2 OR2X2_13 ( .A(REG4_REG_2_), .B(DATA_IN_2_), .Y(_abc_3548_n193) );
  OR2X2 OR2X2_130 ( .A(_abc_3548_n468), .B(_abc_3548_n513), .Y(_abc_3548_n514) );
  OR2X2 OR2X2_131 ( .A(_abc_3548_n516), .B(_abc_3548_n500), .Y(n332) );
  OR2X2 OR2X2_132 ( .A(_abc_3548_n520), .B(_abc_3548_n148), .Y(_abc_3548_n521) );
  OR2X2 OR2X2_133 ( .A(_abc_3548_n519), .B(_abc_3548_n521), .Y(_abc_3548_n522) );
  OR2X2 OR2X2_134 ( .A(_abc_3548_n522), .B(_abc_3548_n518), .Y(_abc_3548_n523) );
  OR2X2 OR2X2_135 ( .A(_abc_3548_n526), .B(_abc_3548_n523), .Y(n328) );
  OR2X2 OR2X2_136 ( .A(_abc_3548_n530), .B(_abc_3548_n148), .Y(_abc_3548_n531) );
  OR2X2 OR2X2_137 ( .A(_abc_3548_n529), .B(_abc_3548_n531), .Y(_abc_3548_n532) );
  OR2X2 OR2X2_138 ( .A(_abc_3548_n532), .B(_abc_3548_n528), .Y(n324) );
  OR2X2 OR2X2_139 ( .A(_abc_3548_n535), .B(_abc_3548_n148), .Y(_abc_3548_n536) );
  OR2X2 OR2X2_14 ( .A(REG4_REG_1_), .B(DATA_IN_1_), .Y(_abc_3548_n194) );
  OR2X2 OR2X2_140 ( .A(_abc_3548_n534), .B(_abc_3548_n536), .Y(n319) );
  OR2X2 OR2X2_141 ( .A(_abc_3548_n539), .B(_abc_3548_n148), .Y(_abc_3548_n540) );
  OR2X2 OR2X2_142 ( .A(_abc_3548_n538), .B(_abc_3548_n540), .Y(n314) );
  OR2X2 OR2X2_143 ( .A(_abc_3548_n543), .B(_abc_3548_n148), .Y(_abc_3548_n544) );
  OR2X2 OR2X2_144 ( .A(_abc_3548_n542), .B(_abc_3548_n544), .Y(n309) );
  OR2X2 OR2X2_145 ( .A(_abc_3548_n547), .B(_abc_3548_n148), .Y(_abc_3548_n548) );
  OR2X2 OR2X2_146 ( .A(_abc_3548_n546), .B(_abc_3548_n548), .Y(n304) );
  OR2X2 OR2X2_147 ( .A(_abc_3548_n551), .B(_abc_3548_n148), .Y(_abc_3548_n552) );
  OR2X2 OR2X2_148 ( .A(_abc_3548_n550), .B(_abc_3548_n552), .Y(n299) );
  OR2X2 OR2X2_149 ( .A(_abc_3548_n555), .B(_abc_3548_n148), .Y(_abc_3548_n556) );
  OR2X2 OR2X2_15 ( .A(_abc_3548_n197), .B(_abc_3548_n198), .Y(_abc_3548_n199) );
  OR2X2 OR2X2_150 ( .A(_abc_3548_n554), .B(_abc_3548_n556), .Y(n294) );
  OR2X2 OR2X2_151 ( .A(_abc_3548_n559), .B(_abc_3548_n148), .Y(_abc_3548_n560) );
  OR2X2 OR2X2_152 ( .A(_abc_3548_n558), .B(_abc_3548_n560), .Y(n289) );
  OR2X2 OR2X2_153 ( .A(_abc_3548_n563), .B(_abc_3548_n148), .Y(_abc_3548_n564) );
  OR2X2 OR2X2_154 ( .A(_abc_3548_n562), .B(_abc_3548_n564), .Y(n284) );
  OR2X2 OR2X2_155 ( .A(_abc_3548_n567), .B(_abc_3548_n148), .Y(_abc_3548_n568) );
  OR2X2 OR2X2_156 ( .A(_abc_3548_n566), .B(_abc_3548_n568), .Y(n279) );
  OR2X2 OR2X2_157 ( .A(_abc_3548_n571), .B(_abc_3548_n148), .Y(_abc_3548_n572) );
  OR2X2 OR2X2_158 ( .A(_abc_3548_n570), .B(_abc_3548_n572), .Y(n274) );
  OR2X2 OR2X2_159 ( .A(_abc_3548_n575), .B(_abc_3548_n148), .Y(_abc_3548_n576) );
  OR2X2 OR2X2_16 ( .A(_abc_3548_n196), .B(_abc_3548_n199), .Y(_abc_3548_n200) );
  OR2X2 OR2X2_160 ( .A(_abc_3548_n574), .B(_abc_3548_n576), .Y(n269) );
  OR2X2 OR2X2_161 ( .A(_abc_3548_n579), .B(_abc_3548_n148), .Y(_abc_3548_n580) );
  OR2X2 OR2X2_162 ( .A(_abc_3548_n578), .B(_abc_3548_n580), .Y(n264) );
  OR2X2 OR2X2_163 ( .A(_abc_3548_n583), .B(_abc_3548_n148), .Y(_abc_3548_n584) );
  OR2X2 OR2X2_164 ( .A(_abc_3548_n582), .B(_abc_3548_n584), .Y(n259) );
  OR2X2 OR2X2_165 ( .A(_abc_3548_n587), .B(_abc_3548_n148), .Y(_abc_3548_n588) );
  OR2X2 OR2X2_166 ( .A(_abc_3548_n586), .B(_abc_3548_n588), .Y(n254) );
  OR2X2 OR2X2_167 ( .A(_abc_3548_n591), .B(_abc_3548_n148), .Y(_abc_3548_n592) );
  OR2X2 OR2X2_168 ( .A(_abc_3548_n590), .B(_abc_3548_n592), .Y(n249) );
  OR2X2 OR2X2_169 ( .A(_abc_3548_n595), .B(_abc_3548_n148), .Y(_abc_3548_n596) );
  OR2X2 OR2X2_17 ( .A(_abc_3548_n203), .B(_abc_3548_n206), .Y(_abc_3548_n207) );
  OR2X2 OR2X2_170 ( .A(_abc_3548_n594), .B(_abc_3548_n596), .Y(n244) );
  OR2X2 OR2X2_171 ( .A(_abc_3548_n599), .B(_abc_3548_n148), .Y(_abc_3548_n600) );
  OR2X2 OR2X2_172 ( .A(_abc_3548_n598), .B(_abc_3548_n600), .Y(n239) );
  OR2X2 OR2X2_173 ( .A(_abc_3548_n603), .B(_abc_3548_n148), .Y(_abc_3548_n604) );
  OR2X2 OR2X2_174 ( .A(_abc_3548_n602), .B(_abc_3548_n604), .Y(n234) );
  OR2X2 OR2X2_175 ( .A(_abc_3548_n607), .B(_abc_3548_n148), .Y(_abc_3548_n608) );
  OR2X2 OR2X2_176 ( .A(_abc_3548_n606), .B(_abc_3548_n608), .Y(n229) );
  OR2X2 OR2X2_177 ( .A(_abc_3548_n611), .B(_abc_3548_n148), .Y(_abc_3548_n612) );
  OR2X2 OR2X2_178 ( .A(_abc_3548_n610), .B(_abc_3548_n612), .Y(n224) );
  OR2X2 OR2X2_179 ( .A(_abc_3548_n615), .B(_abc_3548_n148), .Y(_abc_3548_n616) );
  OR2X2 OR2X2_18 ( .A(_abc_3548_n210), .B(_abc_3548_n211_1), .Y(_abc_3548_n212) );
  OR2X2 OR2X2_180 ( .A(_abc_3548_n614), .B(_abc_3548_n616), .Y(n219) );
  OR2X2 OR2X2_181 ( .A(_abc_3548_n619), .B(_abc_3548_n148), .Y(_abc_3548_n620) );
  OR2X2 OR2X2_182 ( .A(_abc_3548_n618), .B(_abc_3548_n620), .Y(n214) );
  OR2X2 OR2X2_183 ( .A(_abc_3548_n623), .B(_abc_3548_n148), .Y(_abc_3548_n624) );
  OR2X2 OR2X2_184 ( .A(_abc_3548_n622), .B(_abc_3548_n624), .Y(n209) );
  OR2X2 OR2X2_185 ( .A(_abc_3548_n627), .B(_abc_3548_n148), .Y(_abc_3548_n628) );
  OR2X2 OR2X2_186 ( .A(_abc_3548_n626), .B(_abc_3548_n628), .Y(n204) );
  OR2X2 OR2X2_187 ( .A(_abc_3548_n631), .B(_abc_3548_n148), .Y(_abc_3548_n632) );
  OR2X2 OR2X2_188 ( .A(_abc_3548_n630), .B(_abc_3548_n632), .Y(n199) );
  OR2X2 OR2X2_189 ( .A(_abc_3548_n635), .B(_abc_3548_n148), .Y(_abc_3548_n636) );
  OR2X2 OR2X2_19 ( .A(_abc_3548_n209_1), .B(_abc_3548_n212), .Y(_abc_3548_n213) );
  OR2X2 OR2X2_190 ( .A(_abc_3548_n634), .B(_abc_3548_n636), .Y(n194) );
  OR2X2 OR2X2_191 ( .A(_abc_3548_n639), .B(_abc_3548_n148), .Y(_abc_3548_n640) );
  OR2X2 OR2X2_192 ( .A(_abc_3548_n638), .B(_abc_3548_n640), .Y(n189) );
  OR2X2 OR2X2_193 ( .A(_abc_3548_n643), .B(_abc_3548_n148), .Y(_abc_3548_n644) );
  OR2X2 OR2X2_194 ( .A(_abc_3548_n642), .B(_abc_3548_n644), .Y(n184) );
  OR2X2 OR2X2_195 ( .A(_abc_3548_n647), .B(_abc_3548_n148), .Y(_abc_3548_n648) );
  OR2X2 OR2X2_196 ( .A(_abc_3548_n646), .B(_abc_3548_n648), .Y(n179) );
  OR2X2 OR2X2_197 ( .A(_abc_3548_n651), .B(_abc_3548_n148), .Y(_abc_3548_n652) );
  OR2X2 OR2X2_198 ( .A(_abc_3548_n650), .B(_abc_3548_n652), .Y(n174) );
  OR2X2 OR2X2_199 ( .A(_abc_3548_n655), .B(_abc_3548_n148), .Y(_abc_3548_n656) );
  OR2X2 OR2X2_2 ( .A(_abc_3548_n151), .B(_abc_3548_n147_1), .Y(n356) );
  OR2X2 OR2X2_20 ( .A(_abc_3548_n216), .B(_abc_3548_n219), .Y(_abc_3548_n220) );
  OR2X2 OR2X2_200 ( .A(_abc_3548_n654), .B(_abc_3548_n656), .Y(n169) );
  OR2X2 OR2X2_201 ( .A(_abc_3548_n659), .B(_abc_3548_n148), .Y(_abc_3548_n660) );
  OR2X2 OR2X2_202 ( .A(_abc_3548_n658), .B(_abc_3548_n660), .Y(n164) );
  OR2X2 OR2X2_203 ( .A(_abc_3548_n662), .B(_abc_3548_n666), .Y(_abc_3548_n667) );
  OR2X2 OR2X2_204 ( .A(_abc_3548_n668), .B(_abc_3548_n148), .Y(_abc_3548_n669) );
  OR2X2 OR2X2_205 ( .A(_abc_3548_n669), .B(_abc_3548_n665), .Y(n159) );
  OR2X2 OR2X2_206 ( .A(_abc_3548_n672), .B(_abc_3548_n148), .Y(_abc_3548_n673) );
  OR2X2 OR2X2_207 ( .A(_abc_3548_n673), .B(_abc_3548_n671), .Y(n154) );
  OR2X2 OR2X2_208 ( .A(_abc_3548_n676), .B(_abc_3548_n148), .Y(_abc_3548_n677) );
  OR2X2 OR2X2_209 ( .A(_abc_3548_n677), .B(_abc_3548_n675), .Y(n149) );
  OR2X2 OR2X2_21 ( .A(DATA_IN_7_), .B(REG4_REG_7_), .Y(_abc_3548_n224) );
  OR2X2 OR2X2_210 ( .A(_abc_3548_n680), .B(_abc_3548_n148), .Y(_abc_3548_n681) );
  OR2X2 OR2X2_211 ( .A(_abc_3548_n681), .B(_abc_3548_n679), .Y(n144) );
  OR2X2 OR2X2_212 ( .A(_abc_3548_n684), .B(_abc_3548_n148), .Y(_abc_3548_n685) );
  OR2X2 OR2X2_213 ( .A(_abc_3548_n685), .B(_abc_3548_n683), .Y(n139) );
  OR2X2 OR2X2_214 ( .A(_abc_3548_n688), .B(_abc_3548_n148), .Y(_abc_3548_n689) );
  OR2X2 OR2X2_215 ( .A(_abc_3548_n689), .B(_abc_3548_n687), .Y(n134) );
  OR2X2 OR2X2_216 ( .A(_abc_3548_n692), .B(_abc_3548_n148), .Y(_abc_3548_n693) );
  OR2X2 OR2X2_217 ( .A(_abc_3548_n693), .B(_abc_3548_n691), .Y(n129) );
  OR2X2 OR2X2_218 ( .A(_abc_3548_n696), .B(_abc_3548_n148), .Y(_abc_3548_n697) );
  OR2X2 OR2X2_219 ( .A(_abc_3548_n697), .B(_abc_3548_n695), .Y(n124) );
  OR2X2 OR2X2_22 ( .A(_abc_3548_n228), .B(_abc_3548_n189), .Y(_abc_3548_n229) );
  OR2X2 OR2X2_220 ( .A(_abc_3548_n705), .B(RMAX_REG_1_), .Y(_abc_3548_n707) );
  OR2X2 OR2X2_221 ( .A(_abc_3548_n710), .B(_abc_3548_n706), .Y(_abc_3548_n711) );
  OR2X2 OR2X2_222 ( .A(_abc_3548_n713), .B(_abc_3548_n715), .Y(_abc_3548_n716) );
  OR2X2 OR2X2_223 ( .A(_abc_3548_n712), .B(_abc_3548_n716), .Y(_abc_3548_n717) );
  OR2X2 OR2X2_224 ( .A(_abc_3548_n718), .B(_abc_3548_n719), .Y(_abc_3548_n720) );
  OR2X2 OR2X2_225 ( .A(_abc_3548_n723), .B(_abc_3548_n724), .Y(_abc_3548_n725) );
  OR2X2 OR2X2_226 ( .A(_abc_3548_n722), .B(_abc_3548_n725), .Y(_abc_3548_n726) );
  OR2X2 OR2X2_227 ( .A(_abc_3548_n727), .B(_abc_3548_n728), .Y(_abc_3548_n729) );
  OR2X2 OR2X2_228 ( .A(_abc_3548_n732), .B(_abc_3548_n733), .Y(_abc_3548_n734) );
  OR2X2 OR2X2_229 ( .A(_abc_3548_n731), .B(_abc_3548_n734), .Y(_abc_3548_n735) );
  OR2X2 OR2X2_23 ( .A(_abc_3548_n233), .B(RESTART), .Y(_abc_3548_n234) );
  OR2X2 OR2X2_230 ( .A(_abc_3548_n738), .B(_abc_3548_n739), .Y(_abc_3548_n740) );
  OR2X2 OR2X2_231 ( .A(_abc_3548_n744), .B(_abc_3548_n740), .Y(_abc_3548_n745) );
  OR2X2 OR2X2_232 ( .A(_abc_3548_n714), .B(RMIN_REG_2_), .Y(_abc_3548_n748) );
  OR2X2 OR2X2_233 ( .A(_abc_3548_n751), .B(_abc_3548_n752), .Y(_abc_3548_n753) );
  OR2X2 OR2X2_234 ( .A(_abc_3548_n750), .B(_abc_3548_n753), .Y(_abc_3548_n754) );
  OR2X2 OR2X2_235 ( .A(_abc_3548_n755), .B(_abc_3548_n756), .Y(_abc_3548_n757) );
  OR2X2 OR2X2_236 ( .A(_abc_3548_n760), .B(_abc_3548_n761), .Y(_abc_3548_n762) );
  OR2X2 OR2X2_237 ( .A(_abc_3548_n759), .B(_abc_3548_n762), .Y(_abc_3548_n763) );
  OR2X2 OR2X2_238 ( .A(_abc_3548_n764), .B(_abc_3548_n765), .Y(_abc_3548_n766) );
  OR2X2 OR2X2_239 ( .A(_abc_3548_n768), .B(_abc_3548_n737), .Y(_abc_3548_n769) );
  OR2X2 OR2X2_24 ( .A(_abc_3548_n239_1), .B(_abc_3548_n240), .Y(_abc_3548_n241_1) );
  OR2X2 OR2X2_240 ( .A(_abc_3548_n771), .B(STATO_REG_0_), .Y(_abc_3548_n772) );
  OR2X2 OR2X2_241 ( .A(_abc_3548_n775), .B(_abc_3548_n148), .Y(_abc_3548_n776) );
  OR2X2 OR2X2_242 ( .A(_abc_3548_n776), .B(_abc_3548_n774), .Y(n119) );
  OR2X2 OR2X2_243 ( .A(_abc_3548_n779), .B(_abc_3548_n148), .Y(_abc_3548_n780) );
  OR2X2 OR2X2_244 ( .A(_abc_3548_n780), .B(_abc_3548_n778), .Y(n114) );
  OR2X2 OR2X2_245 ( .A(_abc_3548_n783), .B(_abc_3548_n148), .Y(_abc_3548_n784) );
  OR2X2 OR2X2_246 ( .A(_abc_3548_n784), .B(_abc_3548_n782), .Y(n109) );
  OR2X2 OR2X2_247 ( .A(_abc_3548_n787), .B(_abc_3548_n148), .Y(_abc_3548_n788) );
  OR2X2 OR2X2_248 ( .A(_abc_3548_n788), .B(_abc_3548_n786), .Y(n104) );
  OR2X2 OR2X2_249 ( .A(_abc_3548_n791), .B(_abc_3548_n148), .Y(_abc_3548_n792) );
  OR2X2 OR2X2_25 ( .A(RMIN_REG_2_), .B(RMAX_REG_2_), .Y(_abc_3548_n242) );
  OR2X2 OR2X2_250 ( .A(_abc_3548_n792), .B(_abc_3548_n790), .Y(n99) );
  OR2X2 OR2X2_251 ( .A(_abc_3548_n795), .B(_abc_3548_n148), .Y(_abc_3548_n796) );
  OR2X2 OR2X2_252 ( .A(_abc_3548_n796), .B(_abc_3548_n794), .Y(n94) );
  OR2X2 OR2X2_253 ( .A(_abc_3548_n799), .B(_abc_3548_n148), .Y(_abc_3548_n800) );
  OR2X2 OR2X2_254 ( .A(_abc_3548_n800), .B(_abc_3548_n798), .Y(n89) );
  OR2X2 OR2X2_255 ( .A(_abc_3548_n803), .B(_abc_3548_n148), .Y(_abc_3548_n804) );
  OR2X2 OR2X2_256 ( .A(_abc_3548_n804), .B(_abc_3548_n802), .Y(n84) );
  OR2X2 OR2X2_257 ( .A(_abc_3548_n736), .B(_abc_3548_n149), .Y(_abc_3548_n806) );
  OR2X2 OR2X2_258 ( .A(_abc_3548_n810), .B(_abc_3548_n148), .Y(_abc_3548_n811) );
  OR2X2 OR2X2_259 ( .A(_abc_3548_n811), .B(_abc_3548_n809), .Y(n79) );
  OR2X2 OR2X2_26 ( .A(RMIN_REG_1_), .B(RMAX_REG_1_), .Y(_abc_3548_n243) );
  OR2X2 OR2X2_260 ( .A(_abc_3548_n814), .B(_abc_3548_n148), .Y(_abc_3548_n815) );
  OR2X2 OR2X2_261 ( .A(_abc_3548_n815), .B(_abc_3548_n813), .Y(n74) );
  OR2X2 OR2X2_262 ( .A(_abc_3548_n818), .B(_abc_3548_n148), .Y(_abc_3548_n819) );
  OR2X2 OR2X2_263 ( .A(_abc_3548_n819), .B(_abc_3548_n817), .Y(n69) );
  OR2X2 OR2X2_264 ( .A(_abc_3548_n822), .B(_abc_3548_n148), .Y(_abc_3548_n823) );
  OR2X2 OR2X2_265 ( .A(_abc_3548_n823), .B(_abc_3548_n821), .Y(n64) );
  OR2X2 OR2X2_266 ( .A(_abc_3548_n826), .B(_abc_3548_n148), .Y(_abc_3548_n827) );
  OR2X2 OR2X2_267 ( .A(_abc_3548_n827), .B(_abc_3548_n825), .Y(n59) );
  OR2X2 OR2X2_268 ( .A(_abc_3548_n830), .B(_abc_3548_n148), .Y(_abc_3548_n831) );
  OR2X2 OR2X2_269 ( .A(_abc_3548_n831), .B(_abc_3548_n829), .Y(n54) );
  OR2X2 OR2X2_27 ( .A(_abc_3548_n246), .B(_abc_3548_n247), .Y(_abc_3548_n248_1) );
  OR2X2 OR2X2_270 ( .A(_abc_3548_n834), .B(_abc_3548_n148), .Y(_abc_3548_n835) );
  OR2X2 OR2X2_271 ( .A(_abc_3548_n835), .B(_abc_3548_n833), .Y(n49) );
  OR2X2 OR2X2_272 ( .A(_abc_3548_n838), .B(_abc_3548_n148), .Y(_abc_3548_n839) );
  OR2X2 OR2X2_273 ( .A(_abc_3548_n839), .B(_abc_3548_n837), .Y(n44) );
  OR2X2 OR2X2_28 ( .A(_abc_3548_n245), .B(_abc_3548_n248_1), .Y(_abc_3548_n249) );
  OR2X2 OR2X2_29 ( .A(_abc_3548_n252), .B(_abc_3548_n255_1), .Y(_abc_3548_n256) );
  OR2X2 OR2X2_3 ( .A(RESTART), .B(REG4_REG_1_), .Y(_abc_3548_n153) );
  OR2X2 OR2X2_30 ( .A(_abc_3548_n259), .B(_abc_3548_n260_1), .Y(_abc_3548_n261) );
  OR2X2 OR2X2_31 ( .A(_abc_3548_n258), .B(_abc_3548_n261), .Y(_abc_3548_n262) );
  OR2X2 OR2X2_32 ( .A(_abc_3548_n265_1), .B(_abc_3548_n268), .Y(_abc_3548_n269) );
  OR2X2 OR2X2_33 ( .A(_abc_3548_n271), .B(_abc_3548_n238), .Y(_abc_3548_n272_1) );
  OR2X2 OR2X2_34 ( .A(_abc_3548_n273), .B(_abc_3548_n276), .Y(_abc_3548_n277_1) );
  OR2X2 OR2X2_35 ( .A(_abc_3548_n277_1), .B(_abc_3548_n159), .Y(_abc_3548_n278) );
  OR2X2 OR2X2_36 ( .A(_abc_3548_n283_1), .B(_abc_3548_n286_1), .Y(_abc_3548_n287) );
  OR2X2 OR2X2_37 ( .A(_abc_3548_n288_1), .B(_abc_3548_n165_1), .Y(_abc_3548_n289) );
  OR2X2 OR2X2_38 ( .A(_abc_3548_n188), .B(_abc_3548_n290_1), .Y(_abc_3548_n293_1) );
  OR2X2 OR2X2_39 ( .A(_abc_3548_n303), .B(_abc_3548_n148), .Y(_abc_3548_n304_1) );
  OR2X2 OR2X2_4 ( .A(RESTART), .B(DATA_IN_0_), .Y(_abc_3548_n158) );
  OR2X2 OR2X2_40 ( .A(_abc_3548_n301_1), .B(_abc_3548_n304_1), .Y(_abc_3548_n305) );
  OR2X2 OR2X2_41 ( .A(_abc_3548_n305), .B(_abc_3548_n298_1), .Y(_abc_3548_n306_1) );
  OR2X2 OR2X2_42 ( .A(_abc_3548_n295_1), .B(_abc_3548_n306_1), .Y(_abc_3548_n307) );
  OR2X2 OR2X2_43 ( .A(_abc_3548_n307), .B(_abc_3548_n281), .Y(n352) );
  OR2X2 OR2X2_44 ( .A(RESTART), .B(REG4_REG_2_), .Y(_abc_3548_n309_1) );
  OR2X2 OR2X2_45 ( .A(_abc_3548_n159), .B(RMIN_REG_2_), .Y(_abc_3548_n310) );
  OR2X2 OR2X2_46 ( .A(RESTART), .B(DATA_IN_2_), .Y(_abc_3548_n313) );
  OR2X2 OR2X2_47 ( .A(_abc_3548_n159), .B(RMAX_REG_2_), .Y(_abc_3548_n314_1) );
  OR2X2 OR2X2_48 ( .A(_abc_3548_n182_1), .B(_abc_3548_n322), .Y(_abc_3548_n323) );
  OR2X2 OR2X2_49 ( .A(_abc_3548_n169_1), .B(_abc_3548_n157), .Y(_abc_3548_n327_1) );
  OR2X2 OR2X2_5 ( .A(_abc_3548_n159), .B(RMAX_REG_0_), .Y(_abc_3548_n160) );
  OR2X2 OR2X2_50 ( .A(_abc_3548_n325_1), .B(_abc_3548_n329), .Y(_abc_3548_n330_1) );
  OR2X2 OR2X2_51 ( .A(_abc_3548_n291), .B(_abc_3548_n330_1), .Y(_abc_3548_n333) );
  OR2X2 OR2X2_52 ( .A(_abc_3548_n339), .B(_abc_3548_n148), .Y(_abc_3548_n340_1) );
  OR2X2 OR2X2_53 ( .A(_abc_3548_n338), .B(_abc_3548_n340_1), .Y(_abc_3548_n341_1) );
  OR2X2 OR2X2_54 ( .A(_abc_3548_n341_1), .B(_abc_3548_n337_1), .Y(_abc_3548_n342) );
  OR2X2 OR2X2_55 ( .A(_abc_3548_n336), .B(_abc_3548_n342), .Y(_abc_3548_n343_1) );
  OR2X2 OR2X2_56 ( .A(_abc_3548_n343_1), .B(_abc_3548_n335_1), .Y(n348) );
  OR2X2 OR2X2_57 ( .A(_abc_3548_n293_1), .B(_abc_3548_n330_1), .Y(_abc_3548_n345) );
  OR2X2 OR2X2_58 ( .A(_abc_3548_n346_1), .B(_abc_3548_n331), .Y(_abc_3548_n347_1) );
  OR2X2 OR2X2_59 ( .A(_abc_3548_n348), .B(_abc_3548_n319_1), .Y(_abc_3548_n349_1) );
  OR2X2 OR2X2_6 ( .A(_abc_3548_n162_1), .B(_abc_3548_n163), .Y(_abc_3548_n164) );
  OR2X2 OR2X2_60 ( .A(RESTART), .B(REG4_REG_3_), .Y(_abc_3548_n350_1) );
  OR2X2 OR2X2_61 ( .A(_abc_3548_n159), .B(RMIN_REG_3_), .Y(_abc_3548_n351) );
  OR2X2 OR2X2_62 ( .A(RESTART), .B(DATA_IN_3_), .Y(_abc_3548_n353) );
  OR2X2 OR2X2_63 ( .A(_abc_3548_n159), .B(RMAX_REG_3_), .Y(_abc_3548_n354_1) );
  OR2X2 OR2X2_64 ( .A(_abc_3548_n352_1), .B(_abc_3548_n355), .Y(_abc_3548_n358) );
  OR2X2 OR2X2_65 ( .A(_abc_3548_n324_1), .B(_abc_3548_n317), .Y(_abc_3548_n362_1) );
  OR2X2 OR2X2_66 ( .A(_abc_3548_n364), .B(_abc_3548_n361), .Y(_abc_3548_n365_1) );
  OR2X2 OR2X2_67 ( .A(_abc_3548_n367_1), .B(_abc_3548_n368), .Y(_abc_3548_n369) );
  OR2X2 OR2X2_68 ( .A(_abc_3548_n347_1), .B(_abc_3548_n365_1), .Y(_abc_3548_n372) );
  OR2X2 OR2X2_69 ( .A(_abc_3548_n378), .B(_abc_3548_n148), .Y(_abc_3548_n379) );
  OR2X2 OR2X2_7 ( .A(_abc_3548_n167), .B(_abc_3548_n166), .Y(_abc_3548_n168) );
  OR2X2 OR2X2_70 ( .A(_abc_3548_n377_1), .B(_abc_3548_n379), .Y(_abc_3548_n380_1) );
  OR2X2 OR2X2_71 ( .A(_abc_3548_n380_1), .B(_abc_3548_n376), .Y(_abc_3548_n381) );
  OR2X2 OR2X2_72 ( .A(_abc_3548_n375), .B(_abc_3548_n381), .Y(_abc_3548_n382_1) );
  OR2X2 OR2X2_73 ( .A(_abc_3548_n374_1), .B(_abc_3548_n382_1), .Y(n344) );
  OR2X2 OR2X2_74 ( .A(_abc_3548_n363_1), .B(_abc_3548_n384_1), .Y(_abc_3548_n385) );
  OR2X2 OR2X2_75 ( .A(RESTART), .B(REG4_REG_4_), .Y(_abc_3548_n387_1) );
  OR2X2 OR2X2_76 ( .A(_abc_3548_n159), .B(RMIN_REG_4_), .Y(_abc_3548_n388) );
  OR2X2 OR2X2_77 ( .A(RESTART), .B(DATA_IN_4_), .Y(_abc_3548_n391) );
  OR2X2 OR2X2_78 ( .A(_abc_3548_n159), .B(RMAX_REG_4_), .Y(_abc_3548_n392) );
  OR2X2 OR2X2_79 ( .A(_abc_3548_n386), .B(_abc_3548_n399_1), .Y(_abc_3548_n402_1) );
  OR2X2 OR2X2_8 ( .A(_abc_3548_n172), .B(_abc_3548_n174), .Y(_abc_3548_n175) );
  OR2X2 OR2X2_80 ( .A(_abc_3548_n403), .B(_abc_3548_n367_1), .Y(_abc_3548_n404) );
  OR2X2 OR2X2_81 ( .A(_abc_3548_n406), .B(_abc_3548_n400), .Y(_abc_3548_n407) );
  OR2X2 OR2X2_82 ( .A(_abc_3548_n407), .B(_abc_3548_n405_1), .Y(_abc_3548_n408) );
  OR2X2 OR2X2_83 ( .A(_abc_3548_n409_1), .B(_abc_3548_n371), .Y(_abc_3548_n410) );
  OR2X2 OR2X2_84 ( .A(_abc_3548_n411), .B(_abc_3548_n412), .Y(_abc_3548_n413_1) );
  OR2X2 OR2X2_85 ( .A(_abc_3548_n413_1), .B(_abc_3548_n370_1), .Y(_abc_3548_n414) );
  OR2X2 OR2X2_86 ( .A(_abc_3548_n420), .B(_abc_3548_n148), .Y(_abc_3548_n421) );
  OR2X2 OR2X2_87 ( .A(_abc_3548_n419), .B(_abc_3548_n421), .Y(_abc_3548_n422) );
  OR2X2 OR2X2_88 ( .A(_abc_3548_n422), .B(_abc_3548_n418), .Y(_abc_3548_n423) );
  OR2X2 OR2X2_89 ( .A(_abc_3548_n417), .B(_abc_3548_n423), .Y(_abc_3548_n424) );
  OR2X2 OR2X2_9 ( .A(_abc_3548_n176), .B(RESTART), .Y(_abc_3548_n177) );
  OR2X2 OR2X2_90 ( .A(_abc_3548_n416_1), .B(_abc_3548_n424), .Y(n340) );
  OR2X2 OR2X2_91 ( .A(RESTART), .B(REG4_REG_5_), .Y(_abc_3548_n426) );
  OR2X2 OR2X2_92 ( .A(_abc_3548_n159), .B(RMIN_REG_5_), .Y(_abc_3548_n427) );
  OR2X2 OR2X2_93 ( .A(RESTART), .B(DATA_IN_5_), .Y(_abc_3548_n430) );
  OR2X2 OR2X2_94 ( .A(_abc_3548_n159), .B(RMAX_REG_5_), .Y(_abc_3548_n431) );
  OR2X2 OR2X2_95 ( .A(_abc_3548_n386), .B(_abc_3548_n395), .Y(_abc_3548_n440) );
  OR2X2 OR2X2_96 ( .A(_abc_3548_n441), .B(_abc_3548_n439), .Y(_abc_3548_n442) );
  OR2X2 OR2X2_97 ( .A(_abc_3548_n443), .B(_abc_3548_n356), .Y(_abc_3548_n444) );
  OR2X2 OR2X2_98 ( .A(_abc_3548_n445), .B(_abc_3548_n397), .Y(_abc_3548_n446) );
  OR2X2 OR2X2_99 ( .A(_abc_3548_n446), .B(_abc_3548_n438), .Y(_abc_3548_n447) );
endmodule