module b04_reset(clock, RESET_G, nRESET_G, RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_, DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_, DATA_OUT_REG_7_, DATA_OUT_REG_6_, DATA_OUT_REG_5_, DATA_OUT_REG_4_, DATA_OUT_REG_3_, DATA_OUT_REG_2_, DATA_OUT_REG_1_, DATA_OUT_REG_0_);

input AVERAGE;
input DATA_IN_0_;
input DATA_IN_1_;
input DATA_IN_2_;
input DATA_IN_3_;
input DATA_IN_4_;
input DATA_IN_5_;
input DATA_IN_6_;
input DATA_IN_7_;
output DATA_OUT_REG_0_;
output DATA_OUT_REG_1_;
output DATA_OUT_REG_2_;
output DATA_OUT_REG_3_;
output DATA_OUT_REG_4_;
output DATA_OUT_REG_5_;
output DATA_OUT_REG_6_;
output DATA_OUT_REG_7_;
input ENABLE;
wire REG1_REG_0_; 
wire REG1_REG_1_; 
wire REG1_REG_2_; 
wire REG1_REG_3_; 
wire REG1_REG_4_; 
wire REG1_REG_5_; 
wire REG1_REG_6_; 
wire REG1_REG_7_; 
wire REG2_REG_0_; 
wire REG2_REG_1_; 
wire REG2_REG_2_; 
wire REG2_REG_3_; 
wire REG2_REG_4_; 
wire REG2_REG_5_; 
wire REG2_REG_6_; 
wire REG2_REG_7_; 
wire REG3_REG_0_; 
wire REG3_REG_1_; 
wire REG3_REG_2_; 
wire REG3_REG_3_; 
wire REG3_REG_4_; 
wire REG3_REG_5_; 
wire REG3_REG_6_; 
wire REG3_REG_7_; 
wire REG4_REG_0_; 
wire REG4_REG_1_; 
wire REG4_REG_2_; 
wire REG4_REG_3_; 
wire REG4_REG_4_; 
wire REG4_REG_5_; 
wire REG4_REG_6_; 
wire REG4_REG_7_; 
input RESET_G;
input RESTART;
wire RESTART_bF_buf0; 
wire RESTART_bF_buf1; 
wire RESTART_bF_buf2; 
wire RESTART_bF_buf3; 
wire RESTART_bF_buf4; 
wire RESTART_bF_buf5; 
wire RLAST_REG_0_; 
wire RLAST_REG_1_; 
wire RLAST_REG_2_; 
wire RLAST_REG_3_; 
wire RLAST_REG_4_; 
wire RLAST_REG_5_; 
wire RLAST_REG_6_; 
wire RLAST_REG_7_; 
wire RMAX_REG_0_; 
wire RMAX_REG_1_; 
wire RMAX_REG_2_; 
wire RMAX_REG_3_; 
wire RMAX_REG_4_; 
wire RMAX_REG_5_; 
wire RMAX_REG_6_; 
wire RMAX_REG_7_; 
wire RMIN_REG_0_; 
wire RMIN_REG_1_; 
wire RMIN_REG_2_; 
wire RMIN_REG_3_; 
wire RMIN_REG_4_; 
wire RMIN_REG_5_; 
wire RMIN_REG_6_; 
wire RMIN_REG_7_; 
wire STATO_REG_0_; 
wire STATO_REG_1_; 
wire _abc_3576_new_n146_; 
wire _abc_3576_new_n147_; 
wire _abc_3576_new_n147__bF_buf0; 
wire _abc_3576_new_n147__bF_buf1; 
wire _abc_3576_new_n147__bF_buf2; 
wire _abc_3576_new_n147__bF_buf3; 
wire _abc_3576_new_n147__bF_buf4; 
wire _abc_3576_new_n147__bF_buf5; 
wire _abc_3576_new_n148_; 
wire _abc_3576_new_n150_; 
wire _abc_3576_new_n151_; 
wire _abc_3576_new_n152_; 
wire _abc_3576_new_n153_; 
wire _abc_3576_new_n154_; 
wire _abc_3576_new_n155_; 
wire _abc_3576_new_n156_; 
wire _abc_3576_new_n157_; 
wire _abc_3576_new_n158_; 
wire _abc_3576_new_n159_; 
wire _abc_3576_new_n160_; 
wire _abc_3576_new_n161_; 
wire _abc_3576_new_n162_; 
wire _abc_3576_new_n163_; 
wire _abc_3576_new_n164_; 
wire _abc_3576_new_n165_; 
wire _abc_3576_new_n166_; 
wire _abc_3576_new_n167_; 
wire _abc_3576_new_n168_; 
wire _abc_3576_new_n169_; 
wire _abc_3576_new_n170_; 
wire _abc_3576_new_n171_; 
wire _abc_3576_new_n172_; 
wire _abc_3576_new_n173_; 
wire _abc_3576_new_n174_; 
wire _abc_3576_new_n175_; 
wire _abc_3576_new_n176_; 
wire _abc_3576_new_n177_; 
wire _abc_3576_new_n178_; 
wire _abc_3576_new_n179_; 
wire _abc_3576_new_n180_; 
wire _abc_3576_new_n181_; 
wire _abc_3576_new_n182_; 
wire _abc_3576_new_n183_; 
wire _abc_3576_new_n184_; 
wire _abc_3576_new_n185_; 
wire _abc_3576_new_n186_; 
wire _abc_3576_new_n187_; 
wire _abc_3576_new_n188_; 
wire _abc_3576_new_n189_; 
wire _abc_3576_new_n190_; 
wire _abc_3576_new_n191_; 
wire _abc_3576_new_n192_; 
wire _abc_3576_new_n193_; 
wire _abc_3576_new_n194_; 
wire _abc_3576_new_n195_; 
wire _abc_3576_new_n196_; 
wire _abc_3576_new_n197_; 
wire _abc_3576_new_n198_; 
wire _abc_3576_new_n199_; 
wire _abc_3576_new_n200_; 
wire _abc_3576_new_n201_; 
wire _abc_3576_new_n202_; 
wire _abc_3576_new_n203_; 
wire _abc_3576_new_n204_; 
wire _abc_3576_new_n205_; 
wire _abc_3576_new_n206_; 
wire _abc_3576_new_n207_; 
wire _abc_3576_new_n208_; 
wire _abc_3576_new_n209_; 
wire _abc_3576_new_n210_; 
wire _abc_3576_new_n211_; 
wire _abc_3576_new_n212_; 
wire _abc_3576_new_n213_; 
wire _abc_3576_new_n214_; 
wire _abc_3576_new_n215_; 
wire _abc_3576_new_n216_; 
wire _abc_3576_new_n217_; 
wire _abc_3576_new_n218_; 
wire _abc_3576_new_n219_; 
wire _abc_3576_new_n220_; 
wire _abc_3576_new_n221_; 
wire _abc_3576_new_n222_; 
wire _abc_3576_new_n223_; 
wire _abc_3576_new_n224_; 
wire _abc_3576_new_n225_; 
wire _abc_3576_new_n226_; 
wire _abc_3576_new_n227_; 
wire _abc_3576_new_n228_; 
wire _abc_3576_new_n229_; 
wire _abc_3576_new_n230_; 
wire _abc_3576_new_n231_; 
wire _abc_3576_new_n232_; 
wire _abc_3576_new_n233_; 
wire _abc_3576_new_n234_; 
wire _abc_3576_new_n235_; 
wire _abc_3576_new_n236_; 
wire _abc_3576_new_n237_; 
wire _abc_3576_new_n238_; 
wire _abc_3576_new_n239_; 
wire _abc_3576_new_n240_; 
wire _abc_3576_new_n241_; 
wire _abc_3576_new_n242_; 
wire _abc_3576_new_n243_; 
wire _abc_3576_new_n244_; 
wire _abc_3576_new_n245_; 
wire _abc_3576_new_n246_; 
wire _abc_3576_new_n247_; 
wire _abc_3576_new_n248_; 
wire _abc_3576_new_n249_; 
wire _abc_3576_new_n250_; 
wire _abc_3576_new_n251_; 
wire _abc_3576_new_n252_; 
wire _abc_3576_new_n253_; 
wire _abc_3576_new_n254_; 
wire _abc_3576_new_n256_; 
wire _abc_3576_new_n257_; 
wire _abc_3576_new_n258_; 
wire _abc_3576_new_n259_; 
wire _abc_3576_new_n260_; 
wire _abc_3576_new_n261_; 
wire _abc_3576_new_n262_; 
wire _abc_3576_new_n263_; 
wire _abc_3576_new_n264_; 
wire _abc_3576_new_n265_; 
wire _abc_3576_new_n266_; 
wire _abc_3576_new_n267_; 
wire _abc_3576_new_n268_; 
wire _abc_3576_new_n269_; 
wire _abc_3576_new_n270_; 
wire _abc_3576_new_n271_; 
wire _abc_3576_new_n272_; 
wire _abc_3576_new_n273_; 
wire _abc_3576_new_n274_; 
wire _abc_3576_new_n275_; 
wire _abc_3576_new_n276_; 
wire _abc_3576_new_n277_; 
wire _abc_3576_new_n278_; 
wire _abc_3576_new_n279_; 
wire _abc_3576_new_n281_; 
wire _abc_3576_new_n282_; 
wire _abc_3576_new_n283_; 
wire _abc_3576_new_n284_; 
wire _abc_3576_new_n285_; 
wire _abc_3576_new_n286_; 
wire _abc_3576_new_n287_; 
wire _abc_3576_new_n288_; 
wire _abc_3576_new_n289_; 
wire _abc_3576_new_n290_; 
wire _abc_3576_new_n291_; 
wire _abc_3576_new_n292_; 
wire _abc_3576_new_n293_; 
wire _abc_3576_new_n294_; 
wire _abc_3576_new_n295_; 
wire _abc_3576_new_n296_; 
wire _abc_3576_new_n297_; 
wire _abc_3576_new_n298_; 
wire _abc_3576_new_n299_; 
wire _abc_3576_new_n300_; 
wire _abc_3576_new_n301_; 
wire _abc_3576_new_n302_; 
wire _abc_3576_new_n303_; 
wire _abc_3576_new_n304_; 
wire _abc_3576_new_n305_; 
wire _abc_3576_new_n306_; 
wire _abc_3576_new_n307_; 
wire _abc_3576_new_n308_; 
wire _abc_3576_new_n309_; 
wire _abc_3576_new_n311_; 
wire _abc_3576_new_n312_; 
wire _abc_3576_new_n313_; 
wire _abc_3576_new_n314_; 
wire _abc_3576_new_n315_; 
wire _abc_3576_new_n316_; 
wire _abc_3576_new_n317_; 
wire _abc_3576_new_n318_; 
wire _abc_3576_new_n319_; 
wire _abc_3576_new_n320_; 
wire _abc_3576_new_n321_; 
wire _abc_3576_new_n322_; 
wire _abc_3576_new_n323_; 
wire _abc_3576_new_n324_; 
wire _abc_3576_new_n325_; 
wire _abc_3576_new_n326_; 
wire _abc_3576_new_n327_; 
wire _abc_3576_new_n328_; 
wire _abc_3576_new_n329_; 
wire _abc_3576_new_n330_; 
wire _abc_3576_new_n331_; 
wire _abc_3576_new_n332_; 
wire _abc_3576_new_n333_; 
wire _abc_3576_new_n334_; 
wire _abc_3576_new_n335_; 
wire _abc_3576_new_n336_; 
wire _abc_3576_new_n337_; 
wire _abc_3576_new_n338_; 
wire _abc_3576_new_n339_; 
wire _abc_3576_new_n340_; 
wire _abc_3576_new_n341_; 
wire _abc_3576_new_n342_; 
wire _abc_3576_new_n343_; 
wire _abc_3576_new_n344_; 
wire _abc_3576_new_n345_; 
wire _abc_3576_new_n346_; 
wire _abc_3576_new_n347_; 
wire _abc_3576_new_n348_; 
wire _abc_3576_new_n349_; 
wire _abc_3576_new_n350_; 
wire _abc_3576_new_n351_; 
wire _abc_3576_new_n352_; 
wire _abc_3576_new_n354_; 
wire _abc_3576_new_n355_; 
wire _abc_3576_new_n356_; 
wire _abc_3576_new_n357_; 
wire _abc_3576_new_n358_; 
wire _abc_3576_new_n359_; 
wire _abc_3576_new_n360_; 
wire _abc_3576_new_n361_; 
wire _abc_3576_new_n362_; 
wire _abc_3576_new_n363_; 
wire _abc_3576_new_n364_; 
wire _abc_3576_new_n365_; 
wire _abc_3576_new_n366_; 
wire _abc_3576_new_n367_; 
wire _abc_3576_new_n368_; 
wire _abc_3576_new_n369_; 
wire _abc_3576_new_n370_; 
wire _abc_3576_new_n371_; 
wire _abc_3576_new_n372_; 
wire _abc_3576_new_n373_; 
wire _abc_3576_new_n374_; 
wire _abc_3576_new_n375_; 
wire _abc_3576_new_n376_; 
wire _abc_3576_new_n377_; 
wire _abc_3576_new_n378_; 
wire _abc_3576_new_n380_; 
wire _abc_3576_new_n381_; 
wire _abc_3576_new_n382_; 
wire _abc_3576_new_n383_; 
wire _abc_3576_new_n384_; 
wire _abc_3576_new_n385_; 
wire _abc_3576_new_n386_; 
wire _abc_3576_new_n387_; 
wire _abc_3576_new_n388_; 
wire _abc_3576_new_n389_; 
wire _abc_3576_new_n390_; 
wire _abc_3576_new_n391_; 
wire _abc_3576_new_n392_; 
wire _abc_3576_new_n393_; 
wire _abc_3576_new_n394_; 
wire _abc_3576_new_n395_; 
wire _abc_3576_new_n396_; 
wire _abc_3576_new_n397_; 
wire _abc_3576_new_n398_; 
wire _abc_3576_new_n399_; 
wire _abc_3576_new_n400_; 
wire _abc_3576_new_n401_; 
wire _abc_3576_new_n402_; 
wire _abc_3576_new_n403_; 
wire _abc_3576_new_n404_; 
wire _abc_3576_new_n405_; 
wire _abc_3576_new_n406_; 
wire _abc_3576_new_n407_; 
wire _abc_3576_new_n408_; 
wire _abc_3576_new_n410_; 
wire _abc_3576_new_n411_; 
wire _abc_3576_new_n412_; 
wire _abc_3576_new_n413_; 
wire _abc_3576_new_n414_; 
wire _abc_3576_new_n416_; 
wire _abc_3576_new_n417_; 
wire _abc_3576_new_n419_; 
wire _abc_3576_new_n419__bF_buf0; 
wire _abc_3576_new_n419__bF_buf1; 
wire _abc_3576_new_n419__bF_buf2; 
wire _abc_3576_new_n419__bF_buf3; 
wire _abc_3576_new_n419__bF_buf4; 
wire _abc_3576_new_n420_; 
wire _abc_3576_new_n422_; 
wire _abc_3576_new_n424_; 
wire _abc_3576_new_n426_; 
wire _abc_3576_new_n428_; 
wire _abc_3576_new_n430_; 
wire _abc_3576_new_n432_; 
wire _abc_3576_new_n434_; 
wire _abc_3576_new_n436_; 
wire _abc_3576_new_n437_; 
wire _abc_3576_new_n439_; 
wire _abc_3576_new_n440_; 
wire _abc_3576_new_n442_; 
wire _abc_3576_new_n443_; 
wire _abc_3576_new_n445_; 
wire _abc_3576_new_n446_; 
wire _abc_3576_new_n448_; 
wire _abc_3576_new_n449_; 
wire _abc_3576_new_n451_; 
wire _abc_3576_new_n452_; 
wire _abc_3576_new_n454_; 
wire _abc_3576_new_n455_; 
wire _abc_3576_new_n457_; 
wire _abc_3576_new_n458_; 
wire _abc_3576_new_n460_; 
wire _abc_3576_new_n461_; 
wire _abc_3576_new_n463_; 
wire _abc_3576_new_n464_; 
wire _abc_3576_new_n466_; 
wire _abc_3576_new_n467_; 
wire _abc_3576_new_n469_; 
wire _abc_3576_new_n470_; 
wire _abc_3576_new_n472_; 
wire _abc_3576_new_n473_; 
wire _abc_3576_new_n475_; 
wire _abc_3576_new_n476_; 
wire _abc_3576_new_n478_; 
wire _abc_3576_new_n479_; 
wire _abc_3576_new_n481_; 
wire _abc_3576_new_n482_; 
wire _abc_3576_new_n484_; 
wire _abc_3576_new_n485_; 
wire _abc_3576_new_n487_; 
wire _abc_3576_new_n488_; 
wire _abc_3576_new_n490_; 
wire _abc_3576_new_n491_; 
wire _abc_3576_new_n493_; 
wire _abc_3576_new_n494_; 
wire _abc_3576_new_n496_; 
wire _abc_3576_new_n497_; 
wire _abc_3576_new_n499_; 
wire _abc_3576_new_n500_; 
wire _abc_3576_new_n502_; 
wire _abc_3576_new_n503_; 
wire _abc_3576_new_n505_; 
wire _abc_3576_new_n506_; 
wire _abc_3576_new_n508_; 
wire _abc_3576_new_n509_; 
wire _abc_3576_new_n510_; 
wire _abc_3576_new_n511_; 
wire _abc_3576_new_n513_; 
wire _abc_3576_new_n514_; 
wire _abc_3576_new_n516_; 
wire _abc_3576_new_n517_; 
wire _abc_3576_new_n518_; 
wire _abc_3576_new_n520_; 
wire _abc_3576_new_n521_; 
wire _abc_3576_new_n523_; 
wire _abc_3576_new_n524_; 
wire _abc_3576_new_n525_; 
wire _abc_3576_new_n527_; 
wire _abc_3576_new_n528_; 
wire _abc_3576_new_n530_; 
wire _abc_3576_new_n531_; 
wire _abc_3576_new_n533_; 
wire _abc_3576_new_n534_; 
wire _abc_3576_new_n535_; 
wire _abc_3576_new_n537_; 
wire _abc_3576_new_n538_; 
wire _abc_3576_new_n539_; 
wire _abc_3576_new_n540_; 
wire _abc_3576_new_n541_; 
wire _abc_3576_new_n542_; 
wire _abc_3576_new_n543_; 
wire _abc_3576_new_n544_; 
wire _abc_3576_new_n545_; 
wire _abc_3576_new_n546_; 
wire _abc_3576_new_n547_; 
wire _abc_3576_new_n548_; 
wire _abc_3576_new_n549_; 
wire _abc_3576_new_n550_; 
wire _abc_3576_new_n551_; 
wire _abc_3576_new_n552_; 
wire _abc_3576_new_n553_; 
wire _abc_3576_new_n554_; 
wire _abc_3576_new_n555_; 
wire _abc_3576_new_n556_; 
wire _abc_3576_new_n557_; 
wire _abc_3576_new_n558_; 
wire _abc_3576_new_n559_; 
wire _abc_3576_new_n560_; 
wire _abc_3576_new_n561_; 
wire _abc_3576_new_n562_; 
wire _abc_3576_new_n563_; 
wire _abc_3576_new_n564_; 
wire _abc_3576_new_n565_; 
wire _abc_3576_new_n566_; 
wire _abc_3576_new_n567_; 
wire _abc_3576_new_n568_; 
wire _abc_3576_new_n569_; 
wire _abc_3576_new_n570_; 
wire _abc_3576_new_n572_; 
wire _abc_3576_new_n573_; 
wire _abc_3576_new_n575_; 
wire _abc_3576_new_n576_; 
wire _abc_3576_new_n578_; 
wire _abc_3576_new_n579_; 
wire _abc_3576_new_n581_; 
wire _abc_3576_new_n582_; 
wire _abc_3576_new_n584_; 
wire _abc_3576_new_n585_; 
wire _abc_3576_new_n587_; 
wire _abc_3576_new_n588_; 
wire _abc_3576_new_n590_; 
wire _abc_3576_new_n591_; 
wire _abc_3576_new_n593_; 
wire _abc_3576_new_n594_; 
wire _abc_3576_new_n595_; 
wire _abc_3576_new_n596_; 
wire _abc_3576_new_n598_; 
wire _abc_3576_new_n600_; 
wire _abc_3576_new_n602_; 
wire _abc_3576_new_n604_; 
wire _abc_3576_new_n606_; 
wire _abc_3576_new_n608_; 
wire _abc_3576_new_n610_; 
wire _auto_iopadmap_cc_368_execute_4044; 
wire _auto_iopadmap_cc_368_execute_4046; 
wire _auto_iopadmap_cc_368_execute_4048; 
wire _auto_iopadmap_cc_368_execute_4050; 
wire _auto_iopadmap_cc_368_execute_4052; 
wire _auto_iopadmap_cc_368_execute_4054; 
wire _auto_iopadmap_cc_368_execute_4056; 
wire _auto_iopadmap_cc_368_execute_4058; 
input clock;
wire clock_bF_buf0; 
wire clock_bF_buf1; 
wire clock_bF_buf2; 
wire clock_bF_buf3; 
wire clock_bF_buf4; 
wire clock_bF_buf5; 
wire clock_bF_buf6; 
wire clock_bF_buf7; 
wire n104; 
wire n109; 
wire n114; 
wire n119; 
wire n124; 
wire n129; 
wire n134; 
wire n139; 
wire n144; 
wire n149; 
wire n154; 
wire n159; 
wire n164; 
wire n169; 
wire n174; 
wire n179; 
wire n184; 
wire n189; 
wire n194; 
wire n199; 
wire n204; 
wire n209; 
wire n214; 
wire n219; 
wire n224; 
wire n229; 
wire n234; 
wire n239; 
wire n244; 
wire n249; 
wire n254; 
wire n259; 
wire n264; 
wire n269; 
wire n274; 
wire n279; 
wire n284; 
wire n289; 
wire n294; 
wire n299; 
wire n304; 
wire n309; 
wire n314; 
wire n319; 
wire n324; 
wire n328; 
wire n332; 
wire n336; 
wire n340; 
wire n344; 
wire n348; 
wire n352; 
wire n356; 
wire n356_bF_buf0; 
wire n356_bF_buf1; 
wire n356_bF_buf2; 
wire n356_bF_buf3; 
wire n356_bF_buf4; 
wire n356_bF_buf5; 
wire n361; 
wire n44; 
wire n49; 
wire n54; 
wire n59; 
wire n64; 
wire n69; 
wire n74; 
wire n79; 
wire n84; 
wire n89; 
wire n94; 
wire n99; 
input nRESET_G;
wire nRESET_G_bF_buf0; 
wire nRESET_G_bF_buf1; 
wire nRESET_G_bF_buf2; 
wire nRESET_G_bF_buf3; 
AND2X2 AND2X2_1 ( .A(_abc_3576_new_n211_), .B(_abc_3576_new_n241_), .Y(_abc_3576_new_n242_));
AND2X2 AND2X2_2 ( .A(_abc_3576_new_n242_), .B(_abc_3576_new_n240_), .Y(_abc_3576_new_n243_));
AND2X2 AND2X2_3 ( .A(AVERAGE), .B(ENABLE), .Y(_abc_3576_new_n246_));
AND2X2 AND2X2_4 ( .A(_abc_3576_new_n289_), .B(_abc_3576_new_n292_), .Y(_abc_3576_new_n293_));
AND2X2 AND2X2_5 ( .A(_abc_3576_new_n272_), .B(_abc_3576_new_n301_), .Y(_abc_3576_new_n302_));
AND2X2 AND2X2_6 ( .A(_abc_3576_new_n416_), .B(nRESET_G_bF_buf0), .Y(_abc_3576_new_n417_));
AND2X2 AND2X2_7 ( .A(_abc_3576_new_n551_), .B(_abc_3576_new_n537_), .Y(_abc_3576_new_n552_));
AOI21X1 AOI21X1_1 ( .A(_abc_3576_new_n146_), .B(STATO_REG_0_), .C(_abc_3576_new_n147__bF_buf5), .Y(_abc_3576_new_n148_));
AOI21X1 AOI21X1_10 ( .A(REG4_REG_1_), .B(_abc_3576_new_n248_), .C(_abc_3576_new_n278_), .Y(_abc_3576_new_n279_));
AOI21X1 AOI21X1_11 ( .A(_abc_3576_new_n296_), .B(_abc_3576_new_n281_), .C(_abc_3576_new_n293_), .Y(_abc_3576_new_n297_));
AOI21X1 AOI21X1_12 ( .A(_abc_3576_new_n299_), .B(_abc_3576_new_n294_), .C(_abc_3576_new_n298_), .Y(_abc_3576_new_n300_));
AOI21X1 AOI21X1_13 ( .A(_abc_3576_new_n305_), .B(RLAST_REG_2_), .C(_abc_3576_new_n307_), .Y(_abc_3576_new_n308_));
AOI21X1 AOI21X1_14 ( .A(_abc_3576_new_n251_), .B(_auto_iopadmap_cc_368_execute_4050), .C(_abc_3576_new_n147__bF_buf1), .Y(_abc_3576_new_n313_));
AOI21X1 AOI21X1_15 ( .A(_abc_3576_new_n338_), .B(_abc_3576_new_n339_), .C(_abc_3576_new_n187_), .Y(_abc_3576_new_n340_));
AOI21X1 AOI21X1_16 ( .A(_abc_3576_new_n342_), .B(_abc_3576_new_n343_), .C(_abc_3576_new_n317_), .Y(_abc_3576_new_n344_));
AOI21X1 AOI21X1_17 ( .A(_abc_3576_new_n326_), .B(_abc_3576_new_n289_), .C(_abc_3576_new_n330_), .Y(_abc_3576_new_n345_));
AOI21X1 AOI21X1_18 ( .A(_abc_3576_new_n332_), .B(_abc_3576_new_n346_), .C(_abc_3576_new_n341_), .Y(_abc_3576_new_n354_));
AOI21X1 AOI21X1_19 ( .A(_abc_3576_new_n365_), .B(_abc_3576_new_n328_), .C(_abc_3576_new_n363_), .Y(_abc_3576_new_n368_));
AOI21X1 AOI21X1_2 ( .A(_abc_3576_new_n154_), .B(_abc_3576_new_n177_), .C(_abc_3576_new_n157_), .Y(_abc_3576_new_n178_));
AOI21X1 AOI21X1_20 ( .A(_abc_3576_new_n333_), .B(_abc_3576_new_n324_), .C(_abc_3576_new_n361_), .Y(_abc_3576_new_n369_));
AOI21X1 AOI21X1_21 ( .A(_abc_3576_new_n251_), .B(_auto_iopadmap_cc_368_execute_4052), .C(_abc_3576_new_n147__bF_buf0), .Y(_abc_3576_new_n376_));
AOI21X1 AOI21X1_22 ( .A(RLAST_REG_4_), .B(_abc_3576_new_n305_), .C(_abc_3576_new_n377_), .Y(_abc_3576_new_n378_));
AOI21X1 AOI21X1_23 ( .A(_abc_3576_new_n391_), .B(_abc_3576_new_n393_), .C(_abc_3576_new_n380_), .Y(_abc_3576_new_n394_));
AOI21X1 AOI21X1_24 ( .A(_abc_3576_new_n248_), .B(REG4_REG_5_), .C(_abc_3576_new_n405_), .Y(_abc_3576_new_n406_));
AOI21X1 AOI21X1_25 ( .A(_abc_3576_new_n243_), .B(_abc_3576_new_n402_), .C(_abc_3576_new_n407_), .Y(_abc_3576_new_n408_));
AOI21X1 AOI21X1_26 ( .A(_abc_3576_new_n251_), .B(_auto_iopadmap_cc_368_execute_4056), .C(_abc_3576_new_n147__bF_buf5), .Y(_abc_3576_new_n411_));
AOI21X1 AOI21X1_27 ( .A(REG4_REG_6_), .B(_abc_3576_new_n248_), .C(_abc_3576_new_n412_), .Y(_abc_3576_new_n413_));
AOI21X1 AOI21X1_28 ( .A(_abc_3576_new_n419__bF_buf4), .B(REG3_REG_0_), .C(_abc_3576_new_n147__bF_buf4), .Y(_abc_3576_new_n420_));
AOI21X1 AOI21X1_29 ( .A(_abc_3576_new_n419__bF_buf3), .B(REG3_REG_1_), .C(_abc_3576_new_n147__bF_buf3), .Y(_abc_3576_new_n422_));
AOI21X1 AOI21X1_3 ( .A(_abc_3576_new_n194_), .B(_abc_3576_new_n195_), .C(_abc_3576_new_n200_), .Y(_abc_3576_new_n201_));
AOI21X1 AOI21X1_30 ( .A(_abc_3576_new_n419__bF_buf2), .B(REG3_REG_2_), .C(_abc_3576_new_n147__bF_buf2), .Y(_abc_3576_new_n424_));
AOI21X1 AOI21X1_31 ( .A(_abc_3576_new_n419__bF_buf1), .B(REG3_REG_3_), .C(_abc_3576_new_n147__bF_buf1), .Y(_abc_3576_new_n426_));
AOI21X1 AOI21X1_32 ( .A(_abc_3576_new_n419__bF_buf0), .B(REG3_REG_4_), .C(_abc_3576_new_n147__bF_buf0), .Y(_abc_3576_new_n428_));
AOI21X1 AOI21X1_33 ( .A(_abc_3576_new_n419__bF_buf4), .B(REG3_REG_5_), .C(_abc_3576_new_n147__bF_buf5), .Y(_abc_3576_new_n430_));
AOI21X1 AOI21X1_34 ( .A(_abc_3576_new_n419__bF_buf3), .B(REG3_REG_6_), .C(_abc_3576_new_n147__bF_buf4), .Y(_abc_3576_new_n432_));
AOI21X1 AOI21X1_35 ( .A(_abc_3576_new_n419__bF_buf2), .B(REG3_REG_7_), .C(_abc_3576_new_n147__bF_buf3), .Y(_abc_3576_new_n434_));
AOI21X1 AOI21X1_36 ( .A(_abc_3576_new_n419__bF_buf1), .B(REG2_REG_0_), .C(_abc_3576_new_n147__bF_buf2), .Y(_abc_3576_new_n437_));
AOI21X1 AOI21X1_37 ( .A(_abc_3576_new_n419__bF_buf0), .B(REG2_REG_1_), .C(_abc_3576_new_n147__bF_buf1), .Y(_abc_3576_new_n440_));
AOI21X1 AOI21X1_38 ( .A(_abc_3576_new_n419__bF_buf4), .B(REG2_REG_2_), .C(_abc_3576_new_n147__bF_buf0), .Y(_abc_3576_new_n443_));
AOI21X1 AOI21X1_39 ( .A(_abc_3576_new_n419__bF_buf3), .B(REG2_REG_3_), .C(_abc_3576_new_n147__bF_buf5), .Y(_abc_3576_new_n446_));
AOI21X1 AOI21X1_4 ( .A(_abc_3576_new_n214_), .B(_abc_3576_new_n215_), .C(_abc_3576_new_n220_), .Y(_abc_3576_new_n221_));
AOI21X1 AOI21X1_40 ( .A(_abc_3576_new_n419__bF_buf2), .B(REG2_REG_4_), .C(_abc_3576_new_n147__bF_buf4), .Y(_abc_3576_new_n449_));
AOI21X1 AOI21X1_41 ( .A(_abc_3576_new_n419__bF_buf1), .B(REG2_REG_5_), .C(_abc_3576_new_n147__bF_buf3), .Y(_abc_3576_new_n452_));
AOI21X1 AOI21X1_42 ( .A(_abc_3576_new_n419__bF_buf0), .B(REG2_REG_6_), .C(_abc_3576_new_n147__bF_buf2), .Y(_abc_3576_new_n455_));
AOI21X1 AOI21X1_43 ( .A(_abc_3576_new_n419__bF_buf4), .B(REG2_REG_7_), .C(_abc_3576_new_n147__bF_buf1), .Y(_abc_3576_new_n458_));
AOI21X1 AOI21X1_44 ( .A(_abc_3576_new_n419__bF_buf3), .B(REG1_REG_0_), .C(_abc_3576_new_n147__bF_buf0), .Y(_abc_3576_new_n461_));
AOI21X1 AOI21X1_45 ( .A(_abc_3576_new_n419__bF_buf2), .B(REG1_REG_1_), .C(_abc_3576_new_n147__bF_buf5), .Y(_abc_3576_new_n464_));
AOI21X1 AOI21X1_46 ( .A(_abc_3576_new_n419__bF_buf1), .B(REG1_REG_2_), .C(_abc_3576_new_n147__bF_buf4), .Y(_abc_3576_new_n467_));
AOI21X1 AOI21X1_47 ( .A(_abc_3576_new_n419__bF_buf0), .B(REG1_REG_3_), .C(_abc_3576_new_n147__bF_buf3), .Y(_abc_3576_new_n470_));
AOI21X1 AOI21X1_48 ( .A(_abc_3576_new_n419__bF_buf4), .B(REG1_REG_4_), .C(_abc_3576_new_n147__bF_buf2), .Y(_abc_3576_new_n473_));
AOI21X1 AOI21X1_49 ( .A(_abc_3576_new_n419__bF_buf3), .B(REG1_REG_5_), .C(_abc_3576_new_n147__bF_buf1), .Y(_abc_3576_new_n476_));
AOI21X1 AOI21X1_5 ( .A(_abc_3576_new_n234_), .B(_abc_3576_new_n211_), .C(_abc_3576_new_n189_), .Y(_abc_3576_new_n235_));
AOI21X1 AOI21X1_50 ( .A(_abc_3576_new_n419__bF_buf2), .B(REG1_REG_6_), .C(_abc_3576_new_n147__bF_buf0), .Y(_abc_3576_new_n479_));
AOI21X1 AOI21X1_51 ( .A(_abc_3576_new_n419__bF_buf1), .B(REG1_REG_7_), .C(_abc_3576_new_n147__bF_buf5), .Y(_abc_3576_new_n482_));
AOI21X1 AOI21X1_52 ( .A(_abc_3576_new_n419__bF_buf0), .B(DATA_IN_0_), .C(_abc_3576_new_n147__bF_buf4), .Y(_abc_3576_new_n485_));
AOI21X1 AOI21X1_53 ( .A(_abc_3576_new_n419__bF_buf4), .B(DATA_IN_1_), .C(_abc_3576_new_n147__bF_buf3), .Y(_abc_3576_new_n488_));
AOI21X1 AOI21X1_54 ( .A(_abc_3576_new_n419__bF_buf3), .B(DATA_IN_2_), .C(_abc_3576_new_n147__bF_buf2), .Y(_abc_3576_new_n491_));
AOI21X1 AOI21X1_55 ( .A(_abc_3576_new_n419__bF_buf2), .B(DATA_IN_3_), .C(_abc_3576_new_n147__bF_buf1), .Y(_abc_3576_new_n494_));
AOI21X1 AOI21X1_56 ( .A(_abc_3576_new_n419__bF_buf1), .B(DATA_IN_4_), .C(_abc_3576_new_n147__bF_buf0), .Y(_abc_3576_new_n497_));
AOI21X1 AOI21X1_57 ( .A(_abc_3576_new_n419__bF_buf0), .B(DATA_IN_5_), .C(_abc_3576_new_n147__bF_buf5), .Y(_abc_3576_new_n500_));
AOI21X1 AOI21X1_58 ( .A(_abc_3576_new_n419__bF_buf4), .B(DATA_IN_6_), .C(_abc_3576_new_n147__bF_buf4), .Y(_abc_3576_new_n503_));
AOI21X1 AOI21X1_59 ( .A(_abc_3576_new_n419__bF_buf3), .B(DATA_IN_7_), .C(_abc_3576_new_n147__bF_buf3), .Y(_abc_3576_new_n506_));
AOI21X1 AOI21X1_6 ( .A(_abc_3576_new_n251_), .B(_auto_iopadmap_cc_368_execute_4044), .C(_abc_3576_new_n147__bF_buf3), .Y(_abc_3576_new_n252_));
AOI21X1 AOI21X1_60 ( .A(_abc_3576_new_n223_), .B(RMAX_REG_5_), .C(_abc_3576_new_n546_), .Y(_abc_3576_new_n547_));
AOI21X1 AOI21X1_61 ( .A(_abc_3576_new_n563_), .B(_abc_3576_new_n564_), .C(_abc_3576_new_n565_), .Y(_abc_3576_new_n566_));
AOI21X1 AOI21X1_62 ( .A(_abc_3576_new_n595_), .B(RMAX_REG_0_), .C(_abc_3576_new_n147__bF_buf2), .Y(_abc_3576_new_n596_));
AOI21X1 AOI21X1_63 ( .A(_abc_3576_new_n595_), .B(RMAX_REG_1_), .C(_abc_3576_new_n147__bF_buf1), .Y(_abc_3576_new_n598_));
AOI21X1 AOI21X1_64 ( .A(_abc_3576_new_n595_), .B(RMAX_REG_2_), .C(_abc_3576_new_n147__bF_buf0), .Y(_abc_3576_new_n600_));
AOI21X1 AOI21X1_65 ( .A(_abc_3576_new_n595_), .B(RMAX_REG_3_), .C(_abc_3576_new_n147__bF_buf5), .Y(_abc_3576_new_n602_));
AOI21X1 AOI21X1_66 ( .A(_abc_3576_new_n595_), .B(RMAX_REG_4_), .C(_abc_3576_new_n147__bF_buf4), .Y(_abc_3576_new_n604_));
AOI21X1 AOI21X1_67 ( .A(_abc_3576_new_n595_), .B(RMAX_REG_5_), .C(_abc_3576_new_n147__bF_buf3), .Y(_abc_3576_new_n606_));
AOI21X1 AOI21X1_68 ( .A(_abc_3576_new_n595_), .B(RMAX_REG_6_), .C(_abc_3576_new_n147__bF_buf2), .Y(_abc_3576_new_n608_));
AOI21X1 AOI21X1_69 ( .A(_abc_3576_new_n595_), .B(RMAX_REG_7_), .C(_abc_3576_new_n147__bF_buf1), .Y(_abc_3576_new_n610_));
AOI21X1 AOI21X1_7 ( .A(REG4_REG_0_), .B(_abc_3576_new_n248_), .C(_abc_3576_new_n253_), .Y(_abc_3576_new_n254_));
AOI21X1 AOI21X1_8 ( .A(_abc_3576_new_n159_), .B(_abc_3576_new_n267_), .C(_abc_3576_new_n266_), .Y(_abc_3576_new_n268_));
AOI21X1 AOI21X1_9 ( .A(_abc_3576_new_n251_), .B(_auto_iopadmap_cc_368_execute_4046), .C(_abc_3576_new_n147__bF_buf2), .Y(_abc_3576_new_n277_));
AOI22X1 AOI22X1_1 ( .A(_abc_3576_new_n181_), .B(_abc_3576_new_n179_), .C(_abc_3576_new_n182_), .D(_abc_3576_new_n184_), .Y(_abc_3576_new_n185_));
AOI22X1 AOI22X1_10 ( .A(_abc_3576_new_n341_), .B(_abc_3576_new_n318_), .C(_abc_3576_new_n349_), .D(_abc_3576_new_n348_), .Y(_abc_3576_new_n350_));
AOI22X1 AOI22X1_11 ( .A(_abc_3576_new_n235_), .B(_abc_3576_new_n351_), .C(_abc_3576_new_n335_), .D(_abc_3576_new_n243_), .Y(_abc_3576_new_n352_));
AOI22X1 AOI22X1_12 ( .A(_abc_3576_new_n395_), .B(_abc_3576_new_n354_), .C(_abc_3576_new_n397_), .D(_abc_3576_new_n396_), .Y(_abc_3576_new_n398_));
AOI22X1 AOI22X1_13 ( .A(_auto_iopadmap_cc_368_execute_4058), .B(_abc_3576_new_n251_), .C(RLAST_REG_7_), .D(_abc_3576_new_n305_), .Y(_abc_3576_new_n416_));
AOI22X1 AOI22X1_14 ( .A(_abc_3576_new_n286_), .B(DATA_IN_3_), .C(DATA_IN_4_), .D(_abc_3576_new_n195_), .Y(_abc_3576_new_n544_));
AOI22X1 AOI22X1_15 ( .A(_abc_3576_new_n203_), .B(DATA_IN_5_), .C(DATA_IN_6_), .D(_abc_3576_new_n192_), .Y(_abc_3576_new_n548_));
AOI22X1 AOI22X1_16 ( .A(_abc_3576_new_n228_), .B(RMAX_REG_6_), .C(DATA_IN_7_), .D(_abc_3576_new_n191_), .Y(_abc_3576_new_n550_));
AOI22X1 AOI22X1_17 ( .A(_abc_3576_new_n153_), .B(RMIN_REG_1_), .C(_abc_3576_new_n257_), .D(RMIN_REG_2_), .Y(_abc_3576_new_n555_));
AOI22X1 AOI22X1_18 ( .A(_abc_3576_new_n290_), .B(RMIN_REG_3_), .C(_abc_3576_new_n215_), .D(RMIN_REG_4_), .Y(_abc_3576_new_n558_));
AOI22X1 AOI22X1_19 ( .A(_abc_3576_new_n202_), .B(DATA_IN_5_), .C(DATA_IN_4_), .D(_abc_3576_new_n194_), .Y(_abc_3576_new_n560_));
AOI22X1 AOI22X1_2 ( .A(RMIN_REG_0_), .B(RMAX_REG_0_), .C(RMIN_REG_1_), .D(RMAX_REG_1_), .Y(_abc_3576_new_n196_));
AOI22X1 AOI22X1_20 ( .A(_abc_3576_new_n228_), .B(RMIN_REG_6_), .C(DATA_IN_7_), .D(_abc_3576_new_n190_), .Y(_abc_3576_new_n564_));
AOI22X1 AOI22X1_3 ( .A(RMIN_REG_2_), .B(RMAX_REG_2_), .C(RMIN_REG_3_), .D(RMAX_REG_3_), .Y(_abc_3576_new_n198_));
AOI22X1 AOI22X1_4 ( .A(REG4_REG_0_), .B(DATA_IN_0_), .C(REG4_REG_1_), .D(DATA_IN_1_), .Y(_abc_3576_new_n216_));
AOI22X1 AOI22X1_5 ( .A(DATA_IN_3_), .B(REG4_REG_3_), .C(REG4_REG_2_), .D(DATA_IN_2_), .Y(_abc_3576_new_n218_));
AOI22X1 AOI22X1_6 ( .A(_abc_3576_new_n260_), .B(_abc_3576_new_n265_), .C(_abc_3576_new_n156_), .D(_abc_3576_new_n269_), .Y(_abc_3576_new_n270_));
AOI22X1 AOI22X1_7 ( .A(_abc_3576_new_n163_), .B(_abc_3576_new_n166_), .C(_abc_3576_new_n152_), .D(_abc_3576_new_n155_), .Y(_abc_3576_new_n295_));
AOI22X1 AOI22X1_8 ( .A(REG4_REG_2_), .B(_abc_3576_new_n248_), .C(_abc_3576_new_n301_), .D(_abc_3576_new_n243_), .Y(_abc_3576_new_n309_));
AOI22X1 AOI22X1_9 ( .A(_abc_3576_new_n167_), .B(_abc_3576_new_n170_), .C(_abc_3576_new_n238_), .D(_abc_3576_new_n237_), .Y(_abc_3576_new_n316_));
BUFX2 BUFX2_1 ( .A(nRESET_G), .Y(nRESET_G_bF_buf2));
BUFX2 BUFX2_10 ( .A(_auto_iopadmap_cc_368_execute_4056), .Y(DATA_OUT_REG_6_));
BUFX2 BUFX2_11 ( .A(_auto_iopadmap_cc_368_execute_4058), .Y(DATA_OUT_REG_7_));
BUFX2 BUFX2_2 ( .A(nRESET_G), .Y(nRESET_G_bF_buf1));
BUFX2 BUFX2_3 ( .A(nRESET_G), .Y(nRESET_G_bF_buf0));
BUFX2 BUFX2_4 ( .A(_auto_iopadmap_cc_368_execute_4044), .Y(DATA_OUT_REG_0_));
BUFX2 BUFX2_5 ( .A(_auto_iopadmap_cc_368_execute_4046), .Y(DATA_OUT_REG_1_));
BUFX2 BUFX2_6 ( .A(_auto_iopadmap_cc_368_execute_4048), .Y(DATA_OUT_REG_2_));
BUFX2 BUFX2_7 ( .A(_auto_iopadmap_cc_368_execute_4050), .Y(DATA_OUT_REG_3_));
BUFX2 BUFX2_8 ( .A(_auto_iopadmap_cc_368_execute_4052), .Y(DATA_OUT_REG_4_));
BUFX2 BUFX2_9 ( .A(_auto_iopadmap_cc_368_execute_4054), .Y(DATA_OUT_REG_5_));
BUFX4 BUFX4_1 ( .A(clock), .Y(clock_bF_buf7));
BUFX4 BUFX4_10 ( .A(_abc_3576_new_n147_), .Y(_abc_3576_new_n147__bF_buf4));
BUFX4 BUFX4_11 ( .A(_abc_3576_new_n147_), .Y(_abc_3576_new_n147__bF_buf3));
BUFX4 BUFX4_12 ( .A(_abc_3576_new_n147_), .Y(_abc_3576_new_n147__bF_buf2));
BUFX4 BUFX4_13 ( .A(_abc_3576_new_n147_), .Y(_abc_3576_new_n147__bF_buf1));
BUFX4 BUFX4_14 ( .A(_abc_3576_new_n147_), .Y(_abc_3576_new_n147__bF_buf0));
BUFX4 BUFX4_15 ( .A(nRESET_G), .Y(nRESET_G_bF_buf3));
BUFX4 BUFX4_16 ( .A(RESTART), .Y(RESTART_bF_buf5));
BUFX4 BUFX4_17 ( .A(RESTART), .Y(RESTART_bF_buf4));
BUFX4 BUFX4_18 ( .A(RESTART), .Y(RESTART_bF_buf3));
BUFX4 BUFX4_19 ( .A(RESTART), .Y(RESTART_bF_buf2));
BUFX4 BUFX4_2 ( .A(clock), .Y(clock_bF_buf6));
BUFX4 BUFX4_20 ( .A(RESTART), .Y(RESTART_bF_buf1));
BUFX4 BUFX4_21 ( .A(RESTART), .Y(RESTART_bF_buf0));
BUFX4 BUFX4_22 ( .A(_abc_3576_new_n419_), .Y(_abc_3576_new_n419__bF_buf4));
BUFX4 BUFX4_23 ( .A(_abc_3576_new_n419_), .Y(_abc_3576_new_n419__bF_buf3));
BUFX4 BUFX4_24 ( .A(_abc_3576_new_n419_), .Y(_abc_3576_new_n419__bF_buf2));
BUFX4 BUFX4_25 ( .A(_abc_3576_new_n419_), .Y(_abc_3576_new_n419__bF_buf1));
BUFX4 BUFX4_26 ( .A(_abc_3576_new_n419_), .Y(_abc_3576_new_n419__bF_buf0));
BUFX4 BUFX4_27 ( .A(n356), .Y(n356_bF_buf5));
BUFX4 BUFX4_28 ( .A(n356), .Y(n356_bF_buf4));
BUFX4 BUFX4_29 ( .A(n356), .Y(n356_bF_buf3));
BUFX4 BUFX4_3 ( .A(clock), .Y(clock_bF_buf5));
BUFX4 BUFX4_30 ( .A(n356), .Y(n356_bF_buf2));
BUFX4 BUFX4_31 ( .A(n356), .Y(n356_bF_buf1));
BUFX4 BUFX4_32 ( .A(n356), .Y(n356_bF_buf0));
BUFX4 BUFX4_4 ( .A(clock), .Y(clock_bF_buf4));
BUFX4 BUFX4_5 ( .A(clock), .Y(clock_bF_buf3));
BUFX4 BUFX4_6 ( .A(clock), .Y(clock_bF_buf2));
BUFX4 BUFX4_7 ( .A(clock), .Y(clock_bF_buf1));
BUFX4 BUFX4_8 ( .A(clock), .Y(clock_bF_buf0));
BUFX4 BUFX4_9 ( .A(_abc_3576_new_n147_), .Y(_abc_3576_new_n147__bF_buf5));
DFFPOSX1 DFFPOSX1_1 ( .CLK(clock_bF_buf7), .D(n324), .Q(_auto_iopadmap_cc_368_execute_4058));
DFFPOSX1 DFFPOSX1_10 ( .CLK(clock_bF_buf6), .D(n49), .Q(RMAX_REG_6_));
DFFPOSX1 DFFPOSX1_11 ( .CLK(clock_bF_buf5), .D(n54), .Q(RMAX_REG_5_));
DFFPOSX1 DFFPOSX1_12 ( .CLK(clock_bF_buf4), .D(n59), .Q(RMAX_REG_4_));
DFFPOSX1 DFFPOSX1_13 ( .CLK(clock_bF_buf3), .D(n64), .Q(RMAX_REG_3_));
DFFPOSX1 DFFPOSX1_14 ( .CLK(clock_bF_buf2), .D(n69), .Q(RMAX_REG_2_));
DFFPOSX1 DFFPOSX1_15 ( .CLK(clock_bF_buf1), .D(n74), .Q(RMAX_REG_1_));
DFFPOSX1 DFFPOSX1_16 ( .CLK(clock_bF_buf0), .D(n79), .Q(RMAX_REG_0_));
DFFPOSX1 DFFPOSX1_17 ( .CLK(clock_bF_buf7), .D(n84), .Q(RMIN_REG_7_));
DFFPOSX1 DFFPOSX1_18 ( .CLK(clock_bF_buf6), .D(n89), .Q(RMIN_REG_6_));
DFFPOSX1 DFFPOSX1_19 ( .CLK(clock_bF_buf5), .D(n94), .Q(RMIN_REG_5_));
DFFPOSX1 DFFPOSX1_2 ( .CLK(clock_bF_buf6), .D(n332), .Q(_auto_iopadmap_cc_368_execute_4054));
DFFPOSX1 DFFPOSX1_20 ( .CLK(clock_bF_buf4), .D(n99), .Q(RMIN_REG_4_));
DFFPOSX1 DFFPOSX1_21 ( .CLK(clock_bF_buf3), .D(n104), .Q(RMIN_REG_3_));
DFFPOSX1 DFFPOSX1_22 ( .CLK(clock_bF_buf2), .D(n109), .Q(RMIN_REG_2_));
DFFPOSX1 DFFPOSX1_23 ( .CLK(clock_bF_buf1), .D(n114), .Q(RMIN_REG_1_));
DFFPOSX1 DFFPOSX1_24 ( .CLK(clock_bF_buf0), .D(n119), .Q(RMIN_REG_0_));
DFFPOSX1 DFFPOSX1_25 ( .CLK(clock_bF_buf7), .D(n124), .Q(RLAST_REG_7_));
DFFPOSX1 DFFPOSX1_26 ( .CLK(clock_bF_buf6), .D(n129), .Q(RLAST_REG_6_));
DFFPOSX1 DFFPOSX1_27 ( .CLK(clock_bF_buf5), .D(n134), .Q(RLAST_REG_5_));
DFFPOSX1 DFFPOSX1_28 ( .CLK(clock_bF_buf4), .D(n139), .Q(RLAST_REG_4_));
DFFPOSX1 DFFPOSX1_29 ( .CLK(clock_bF_buf3), .D(n144), .Q(RLAST_REG_3_));
DFFPOSX1 DFFPOSX1_3 ( .CLK(clock_bF_buf5), .D(n344), .Q(_auto_iopadmap_cc_368_execute_4048));
DFFPOSX1 DFFPOSX1_30 ( .CLK(clock_bF_buf2), .D(n149), .Q(RLAST_REG_2_));
DFFPOSX1 DFFPOSX1_31 ( .CLK(clock_bF_buf1), .D(n154), .Q(RLAST_REG_1_));
DFFPOSX1 DFFPOSX1_32 ( .CLK(clock_bF_buf0), .D(n159), .Q(RLAST_REG_0_));
DFFPOSX1 DFFPOSX1_33 ( .CLK(clock_bF_buf7), .D(n164), .Q(REG1_REG_7_));
DFFPOSX1 DFFPOSX1_34 ( .CLK(clock_bF_buf6), .D(n169), .Q(REG1_REG_6_));
DFFPOSX1 DFFPOSX1_35 ( .CLK(clock_bF_buf5), .D(n174), .Q(REG1_REG_5_));
DFFPOSX1 DFFPOSX1_36 ( .CLK(clock_bF_buf4), .D(n179), .Q(REG1_REG_4_));
DFFPOSX1 DFFPOSX1_37 ( .CLK(clock_bF_buf3), .D(n184), .Q(REG1_REG_3_));
DFFPOSX1 DFFPOSX1_38 ( .CLK(clock_bF_buf2), .D(n189), .Q(REG1_REG_2_));
DFFPOSX1 DFFPOSX1_39 ( .CLK(clock_bF_buf1), .D(n194), .Q(REG1_REG_1_));
DFFPOSX1 DFFPOSX1_4 ( .CLK(clock_bF_buf4), .D(n336), .Q(_auto_iopadmap_cc_368_execute_4052));
DFFPOSX1 DFFPOSX1_40 ( .CLK(clock_bF_buf0), .D(n199), .Q(REG1_REG_0_));
DFFPOSX1 DFFPOSX1_41 ( .CLK(clock_bF_buf7), .D(n204), .Q(REG2_REG_7_));
DFFPOSX1 DFFPOSX1_42 ( .CLK(clock_bF_buf6), .D(n209), .Q(REG2_REG_6_));
DFFPOSX1 DFFPOSX1_43 ( .CLK(clock_bF_buf5), .D(n214), .Q(REG2_REG_5_));
DFFPOSX1 DFFPOSX1_44 ( .CLK(clock_bF_buf4), .D(n219), .Q(REG2_REG_4_));
DFFPOSX1 DFFPOSX1_45 ( .CLK(clock_bF_buf3), .D(n224), .Q(REG2_REG_3_));
DFFPOSX1 DFFPOSX1_46 ( .CLK(clock_bF_buf2), .D(n229), .Q(REG2_REG_2_));
DFFPOSX1 DFFPOSX1_47 ( .CLK(clock_bF_buf1), .D(n234), .Q(REG2_REG_1_));
DFFPOSX1 DFFPOSX1_48 ( .CLK(clock_bF_buf0), .D(n239), .Q(REG2_REG_0_));
DFFPOSX1 DFFPOSX1_49 ( .CLK(clock_bF_buf7), .D(n244), .Q(REG3_REG_7_));
DFFPOSX1 DFFPOSX1_5 ( .CLK(clock_bF_buf3), .D(n340), .Q(_auto_iopadmap_cc_368_execute_4050));
DFFPOSX1 DFFPOSX1_50 ( .CLK(clock_bF_buf6), .D(n249), .Q(REG3_REG_6_));
DFFPOSX1 DFFPOSX1_51 ( .CLK(clock_bF_buf5), .D(n254), .Q(REG3_REG_5_));
DFFPOSX1 DFFPOSX1_52 ( .CLK(clock_bF_buf4), .D(n259), .Q(REG3_REG_4_));
DFFPOSX1 DFFPOSX1_53 ( .CLK(clock_bF_buf3), .D(n264), .Q(REG3_REG_3_));
DFFPOSX1 DFFPOSX1_54 ( .CLK(clock_bF_buf2), .D(n269), .Q(REG3_REG_2_));
DFFPOSX1 DFFPOSX1_55 ( .CLK(clock_bF_buf1), .D(n274), .Q(REG3_REG_1_));
DFFPOSX1 DFFPOSX1_56 ( .CLK(clock_bF_buf0), .D(n279), .Q(REG3_REG_0_));
DFFPOSX1 DFFPOSX1_57 ( .CLK(clock_bF_buf7), .D(n284), .Q(REG4_REG_7_));
DFFPOSX1 DFFPOSX1_58 ( .CLK(clock_bF_buf6), .D(n289), .Q(REG4_REG_6_));
DFFPOSX1 DFFPOSX1_59 ( .CLK(clock_bF_buf5), .D(n294), .Q(REG4_REG_5_));
DFFPOSX1 DFFPOSX1_6 ( .CLK(clock_bF_buf2), .D(n328), .Q(_auto_iopadmap_cc_368_execute_4056));
DFFPOSX1 DFFPOSX1_60 ( .CLK(clock_bF_buf4), .D(n299), .Q(REG4_REG_4_));
DFFPOSX1 DFFPOSX1_61 ( .CLK(clock_bF_buf3), .D(n304), .Q(REG4_REG_3_));
DFFPOSX1 DFFPOSX1_62 ( .CLK(clock_bF_buf2), .D(n309), .Q(REG4_REG_2_));
DFFPOSX1 DFFPOSX1_63 ( .CLK(clock_bF_buf1), .D(n314), .Q(REG4_REG_1_));
DFFPOSX1 DFFPOSX1_64 ( .CLK(clock_bF_buf0), .D(n319), .Q(REG4_REG_0_));
DFFPOSX1 DFFPOSX1_65 ( .CLK(clock_bF_buf7), .D(n356_bF_buf0), .Q(STATO_REG_1_));
DFFPOSX1 DFFPOSX1_66 ( .CLK(clock_bF_buf6), .D(n361), .Q(STATO_REG_0_));
DFFPOSX1 DFFPOSX1_7 ( .CLK(clock_bF_buf1), .D(n348), .Q(_auto_iopadmap_cc_368_execute_4046));
DFFPOSX1 DFFPOSX1_8 ( .CLK(clock_bF_buf0), .D(n352), .Q(_auto_iopadmap_cc_368_execute_4044));
DFFPOSX1 DFFPOSX1_9 ( .CLK(clock_bF_buf7), .D(n44), .Q(RMAX_REG_7_));
INVX1 INVX1_1 ( .A(REG4_REG_1_), .Y(_abc_3576_new_n150_));
INVX1 INVX1_10 ( .A(RMAX_REG_5_), .Y(_abc_3576_new_n203_));
INVX1 INVX1_11 ( .A(_abc_3576_new_n205_), .Y(_abc_3576_new_n206_));
INVX1 INVX1_12 ( .A(REG4_REG_7_), .Y(_abc_3576_new_n213_));
INVX1 INVX1_13 ( .A(REG4_REG_5_), .Y(_abc_3576_new_n222_));
INVX1 INVX1_14 ( .A(REG4_REG_6_), .Y(_abc_3576_new_n229_));
INVX1 INVX1_15 ( .A(ENABLE), .Y(_abc_3576_new_n232_));
INVX1 INVX1_16 ( .A(_abc_3576_new_n233_), .Y(_abc_3576_new_n239_));
INVX1 INVX1_17 ( .A(_abc_3576_new_n189_), .Y(_abc_3576_new_n241_));
INVX1 INVX1_18 ( .A(RLAST_REG_0_), .Y(_abc_3576_new_n249_));
INVX1 INVX1_19 ( .A(REG4_REG_2_), .Y(_abc_3576_new_n261_));
INVX1 INVX1_2 ( .A(DATA_IN_0_), .Y(_abc_3576_new_n161_));
INVX1 INVX1_20 ( .A(RLAST_REG_1_), .Y(_abc_3576_new_n276_));
INVX1 INVX1_21 ( .A(REG4_REG_3_), .Y(_abc_3576_new_n282_));
INVX1 INVX1_22 ( .A(_abc_3576_new_n284_), .Y(_abc_3576_new_n285_));
INVX1 INVX1_23 ( .A(RMAX_REG_3_), .Y(_abc_3576_new_n286_));
INVX1 INVX1_24 ( .A(_abc_3576_new_n250_), .Y(_abc_3576_new_n305_));
INVX1 INVX1_25 ( .A(_auto_iopadmap_cc_368_execute_4048), .Y(_abc_3576_new_n306_));
INVX1 INVX1_26 ( .A(RLAST_REG_3_), .Y(_abc_3576_new_n312_));
INVX1 INVX1_27 ( .A(_abc_3576_new_n324_), .Y(_abc_3576_new_n325_));
INVX1 INVX1_28 ( .A(_abc_3576_new_n328_), .Y(_abc_3576_new_n329_));
INVX1 INVX1_29 ( .A(_abc_3576_new_n330_), .Y(_abc_3576_new_n331_));
INVX1 INVX1_3 ( .A(REG4_REG_0_), .Y(_abc_3576_new_n164_));
INVX1 INVX1_30 ( .A(_abc_3576_new_n334_), .Y(_abc_3576_new_n335_));
INVX1 INVX1_31 ( .A(_abc_3576_new_n346_), .Y(_abc_3576_new_n347_));
INVX1 INVX1_32 ( .A(_abc_3576_new_n350_), .Y(_abc_3576_new_n351_));
INVX1 INVX1_33 ( .A(_abc_3576_new_n361_), .Y(_abc_3576_new_n363_));
INVX1 INVX1_34 ( .A(_abc_3576_new_n385_), .Y(_abc_3576_new_n386_));
INVX1 INVX1_35 ( .A(_abc_3576_new_n389_), .Y(_abc_3576_new_n390_));
INVX1 INVX1_36 ( .A(RLAST_REG_5_), .Y(_abc_3576_new_n403_));
INVX1 INVX1_37 ( .A(_auto_iopadmap_cc_368_execute_4054), .Y(_abc_3576_new_n404_));
INVX1 INVX1_38 ( .A(RLAST_REG_6_), .Y(_abc_3576_new_n410_));
INVX1 INVX1_39 ( .A(REG3_REG_0_), .Y(_abc_3576_new_n436_));
INVX1 INVX1_4 ( .A(_abc_3576_new_n172_), .Y(_abc_3576_new_n173_));
INVX1 INVX1_40 ( .A(REG3_REG_1_), .Y(_abc_3576_new_n439_));
INVX1 INVX1_41 ( .A(REG3_REG_2_), .Y(_abc_3576_new_n442_));
INVX1 INVX1_42 ( .A(REG3_REG_3_), .Y(_abc_3576_new_n445_));
INVX1 INVX1_43 ( .A(REG3_REG_4_), .Y(_abc_3576_new_n448_));
INVX1 INVX1_44 ( .A(REG3_REG_5_), .Y(_abc_3576_new_n451_));
INVX1 INVX1_45 ( .A(REG3_REG_6_), .Y(_abc_3576_new_n454_));
INVX1 INVX1_46 ( .A(REG3_REG_7_), .Y(_abc_3576_new_n457_));
INVX1 INVX1_47 ( .A(REG2_REG_0_), .Y(_abc_3576_new_n460_));
INVX1 INVX1_48 ( .A(REG2_REG_1_), .Y(_abc_3576_new_n463_));
INVX1 INVX1_49 ( .A(REG2_REG_2_), .Y(_abc_3576_new_n466_));
INVX1 INVX1_5 ( .A(RMIN_REG_1_), .Y(_abc_3576_new_n180_));
INVX1 INVX1_50 ( .A(REG2_REG_3_), .Y(_abc_3576_new_n469_));
INVX1 INVX1_51 ( .A(REG2_REG_4_), .Y(_abc_3576_new_n472_));
INVX1 INVX1_52 ( .A(REG2_REG_5_), .Y(_abc_3576_new_n475_));
INVX1 INVX1_53 ( .A(REG2_REG_6_), .Y(_abc_3576_new_n478_));
INVX1 INVX1_54 ( .A(REG2_REG_7_), .Y(_abc_3576_new_n481_));
INVX1 INVX1_55 ( .A(REG1_REG_0_), .Y(_abc_3576_new_n484_));
INVX1 INVX1_56 ( .A(REG1_REG_1_), .Y(_abc_3576_new_n487_));
INVX1 INVX1_57 ( .A(REG1_REG_2_), .Y(_abc_3576_new_n490_));
INVX1 INVX1_58 ( .A(REG1_REG_3_), .Y(_abc_3576_new_n493_));
INVX1 INVX1_59 ( .A(REG1_REG_4_), .Y(_abc_3576_new_n496_));
INVX1 INVX1_6 ( .A(RMAX_REG_1_), .Y(_abc_3576_new_n183_));
INVX1 INVX1_60 ( .A(REG1_REG_5_), .Y(_abc_3576_new_n499_));
INVX1 INVX1_61 ( .A(REG1_REG_6_), .Y(_abc_3576_new_n502_));
INVX1 INVX1_62 ( .A(REG1_REG_7_), .Y(_abc_3576_new_n505_));
INVX1 INVX1_63 ( .A(_abc_3576_new_n510_), .Y(_abc_3576_new_n511_));
INVX1 INVX1_64 ( .A(_abc_3576_new_n513_), .Y(_abc_3576_new_n514_));
INVX1 INVX1_65 ( .A(RLAST_REG_2_), .Y(_abc_3576_new_n516_));
INVX1 INVX1_66 ( .A(_abc_3576_new_n517_), .Y(_abc_3576_new_n518_));
INVX1 INVX1_67 ( .A(_abc_3576_new_n520_), .Y(_abc_3576_new_n521_));
INVX1 INVX1_68 ( .A(RLAST_REG_4_), .Y(_abc_3576_new_n523_));
INVX1 INVX1_69 ( .A(_abc_3576_new_n524_), .Y(_abc_3576_new_n525_));
INVX1 INVX1_7 ( .A(RMAX_REG_6_), .Y(_abc_3576_new_n192_));
INVX1 INVX1_70 ( .A(_abc_3576_new_n527_), .Y(_abc_3576_new_n528_));
INVX1 INVX1_71 ( .A(_abc_3576_new_n530_), .Y(_abc_3576_new_n531_));
INVX1 INVX1_72 ( .A(RLAST_REG_7_), .Y(_abc_3576_new_n533_));
INVX1 INVX1_73 ( .A(_abc_3576_new_n534_), .Y(_abc_3576_new_n535_));
INVX1 INVX1_74 ( .A(_abc_3576_new_n548_), .Y(_abc_3576_new_n549_));
INVX1 INVX1_8 ( .A(RMIN_REG_6_), .Y(_abc_3576_new_n193_));
INVX1 INVX1_9 ( .A(RMIN_REG_4_), .Y(_abc_3576_new_n194_));
INVX2 INVX2_1 ( .A(STATO_REG_1_), .Y(_abc_3576_new_n146_));
INVX2 INVX2_10 ( .A(DATA_IN_5_), .Y(_abc_3576_new_n223_));
INVX2 INVX2_11 ( .A(_abc_3576_new_n247_), .Y(_abc_3576_new_n248_));
INVX2 INVX2_12 ( .A(n356_bF_buf5), .Y(_abc_3576_new_n251_));
INVX2 INVX2_13 ( .A(DATA_IN_2_), .Y(_abc_3576_new_n257_));
INVX2 INVX2_14 ( .A(DATA_IN_3_), .Y(_abc_3576_new_n290_));
INVX2 INVX2_2 ( .A(RESTART_bF_buf5), .Y(_abc_3576_new_n176_));
INVX2 INVX2_3 ( .A(RMIN_REG_7_), .Y(_abc_3576_new_n190_));
INVX2 INVX2_4 ( .A(RMAX_REG_7_), .Y(_abc_3576_new_n191_));
INVX2 INVX2_5 ( .A(RMAX_REG_4_), .Y(_abc_3576_new_n195_));
INVX2 INVX2_6 ( .A(RMIN_REG_5_), .Y(_abc_3576_new_n202_));
INVX2 INVX2_7 ( .A(DATA_IN_7_), .Y(_abc_3576_new_n212_));
INVX2 INVX2_8 ( .A(REG4_REG_4_), .Y(_abc_3576_new_n214_));
INVX2 INVX2_9 ( .A(DATA_IN_4_), .Y(_abc_3576_new_n215_));
INVX4 INVX4_1 ( .A(DATA_IN_1_), .Y(_abc_3576_new_n153_));
INVX4 INVX4_2 ( .A(STATO_REG_0_), .Y(_abc_3576_new_n188_));
INVX4 INVX4_3 ( .A(DATA_IN_6_), .Y(_abc_3576_new_n228_));
INVX4 INVX4_4 ( .A(_abc_3576_new_n567_), .Y(_abc_3576_new_n568_));
INVX8 INVX8_1 ( .A(nRESET_G_bF_buf3), .Y(_abc_3576_new_n147_));
MUX2X1 MUX2X1_1 ( .A(RMIN_REG_1_), .B(REG4_REG_1_), .S(RESTART_bF_buf1), .Y(_abc_3576_new_n157_));
MUX2X1 MUX2X1_2 ( .A(RMAX_REG_1_), .B(DATA_IN_1_), .S(RESTART_bF_buf0), .Y(_abc_3576_new_n158_));
MUX2X1 MUX2X1_3 ( .A(RMAX_REG_0_), .B(DATA_IN_0_), .S(RESTART_bF_buf1), .Y(_abc_3576_new_n168_));
MUX2X1 MUX2X1_4 ( .A(RMIN_REG_0_), .B(REG4_REG_0_), .S(RESTART_bF_buf0), .Y(_abc_3576_new_n169_));
MUX2X1 MUX2X1_5 ( .A(RMIN_REG_2_), .B(REG4_REG_2_), .S(RESTART_bF_buf5), .Y(_abc_3576_new_n256_));
MUX2X1 MUX2X1_6 ( .A(RMAX_REG_2_), .B(DATA_IN_2_), .S(RESTART_bF_buf0), .Y(_abc_3576_new_n264_));
NAND2X1 NAND2X1_1 ( .A(RESTART_bF_buf5), .B(RMIN_REG_1_), .Y(_abc_3576_new_n151_));
NAND2X1 NAND2X1_10 ( .A(_abc_3576_new_n170_), .B(_abc_3576_new_n167_), .Y(_abc_3576_new_n171_));
NAND2X1 NAND2X1_11 ( .A(DATA_IN_1_), .B(_abc_3576_new_n176_), .Y(_abc_3576_new_n177_));
NAND2X1 NAND2X1_12 ( .A(RESTART_bF_buf3), .B(_abc_3576_new_n180_), .Y(_abc_3576_new_n181_));
NAND2X1 NAND2X1_13 ( .A(_abc_3576_new_n176_), .B(_abc_3576_new_n153_), .Y(_abc_3576_new_n182_));
NAND2X1 NAND2X1_14 ( .A(RESTART_bF_buf2), .B(_abc_3576_new_n183_), .Y(_abc_3576_new_n184_));
NAND2X1 NAND2X1_15 ( .A(_abc_3576_new_n190_), .B(_abc_3576_new_n191_), .Y(_abc_3576_new_n210_));
NAND2X1 NAND2X1_16 ( .A(_abc_3576_new_n246_), .B(_abc_3576_new_n245_), .Y(_abc_3576_new_n247_));
NAND2X1 NAND2X1_17 ( .A(_abc_3576_new_n232_), .B(_abc_3576_new_n245_), .Y(_abc_3576_new_n250_));
NAND2X1 NAND2X1_18 ( .A(RESTART_bF_buf4), .B(RMAX_REG_2_), .Y(_abc_3576_new_n258_));
NAND2X1 NAND2X1_19 ( .A(_abc_3576_new_n256_), .B(_abc_3576_new_n259_), .Y(_abc_3576_new_n260_));
NAND2X1 NAND2X1_2 ( .A(RESTART_bF_buf3), .B(RMAX_REG_1_), .Y(_abc_3576_new_n154_));
NAND2X1 NAND2X1_20 ( .A(RESTART_bF_buf2), .B(RMIN_REG_2_), .Y(_abc_3576_new_n262_));
NAND2X1 NAND2X1_21 ( .A(_abc_3576_new_n264_), .B(_abc_3576_new_n263_), .Y(_abc_3576_new_n265_));
NAND2X1 NAND2X1_22 ( .A(_abc_3576_new_n260_), .B(_abc_3576_new_n265_), .Y(_abc_3576_new_n266_));
NAND2X1 NAND2X1_23 ( .A(_abc_3576_new_n172_), .B(_abc_3576_new_n271_), .Y(_abc_3576_new_n272_));
NAND2X1 NAND2X1_24 ( .A(_abc_3576_new_n271_), .B(_abc_3576_new_n243_), .Y(_abc_3576_new_n275_));
NAND2X1 NAND2X1_25 ( .A(_abc_3576_new_n256_), .B(_abc_3576_new_n264_), .Y(_abc_3576_new_n281_));
NAND2X1 NAND2X1_26 ( .A(RESTART_bF_buf5), .B(RMIN_REG_3_), .Y(_abc_3576_new_n283_));
NAND2X1 NAND2X1_27 ( .A(RESTART_bF_buf3), .B(_abc_3576_new_n286_), .Y(_abc_3576_new_n287_));
NAND2X1 NAND2X1_28 ( .A(_abc_3576_new_n288_), .B(_abc_3576_new_n285_), .Y(_abc_3576_new_n289_));
NAND2X1 NAND2X1_29 ( .A(_abc_3576_new_n176_), .B(_abc_3576_new_n290_), .Y(_abc_3576_new_n291_));
NAND2X1 NAND2X1_3 ( .A(_abc_3576_new_n152_), .B(_abc_3576_new_n155_), .Y(_abc_3576_new_n156_));
NAND2X1 NAND2X1_30 ( .A(_abc_3576_new_n263_), .B(_abc_3576_new_n259_), .Y(_abc_3576_new_n294_));
NAND2X1 NAND2X1_31 ( .A(_abc_3576_new_n292_), .B(_abc_3576_new_n289_), .Y(_abc_3576_new_n298_));
NAND2X1 NAND2X1_32 ( .A(RESTART_bF_buf1), .B(RMIN_REG_4_), .Y(_abc_3576_new_n320_));
NAND2X1 NAND2X1_33 ( .A(RESTART_bF_buf5), .B(RMAX_REG_4_), .Y(_abc_3576_new_n322_));
NAND2X1 NAND2X1_34 ( .A(_abc_3576_new_n321_), .B(_abc_3576_new_n323_), .Y(_abc_3576_new_n324_));
NAND2X1 NAND2X1_35 ( .A(_abc_3576_new_n289_), .B(_abc_3576_new_n326_), .Y(_abc_3576_new_n327_));
NAND2X1 NAND2X1_36 ( .A(_abc_3576_new_n331_), .B(_abc_3576_new_n327_), .Y(_abc_3576_new_n332_));
NAND2X1 NAND2X1_37 ( .A(_abc_3576_new_n281_), .B(_abc_3576_new_n294_), .Y(_abc_3576_new_n337_));
NAND2X1 NAND2X1_38 ( .A(RESTART_bF_buf3), .B(_abc_3576_new_n203_), .Y(_abc_3576_new_n355_));
NAND2X1 NAND2X1_39 ( .A(RESTART_bF_buf1), .B(_abc_3576_new_n202_), .Y(_abc_3576_new_n357_));
NAND2X1 NAND2X1_4 ( .A(_abc_3576_new_n157_), .B(_abc_3576_new_n158_), .Y(_abc_3576_new_n159_));
NAND2X1 NAND2X1_40 ( .A(_abc_3576_new_n356_), .B(_abc_3576_new_n358_), .Y(_abc_3576_new_n360_));
NAND2X1 NAND2X1_41 ( .A(_abc_3576_new_n360_), .B(_abc_3576_new_n359_), .Y(_abc_3576_new_n361_));
NAND2X1 NAND2X1_42 ( .A(_abc_3576_new_n370_), .B(_abc_3576_new_n367_), .Y(_abc_3576_new_n371_));
NAND2X1 NAND2X1_43 ( .A(_abc_3576_new_n371_), .B(_abc_3576_new_n351_), .Y(_abc_3576_new_n372_));
NAND2X1 NAND2X1_44 ( .A(RESTART_bF_buf5), .B(RMIN_REG_6_), .Y(_abc_3576_new_n382_));
NAND2X1 NAND2X1_45 ( .A(RESTART_bF_buf3), .B(RMAX_REG_6_), .Y(_abc_3576_new_n384_));
NAND2X1 NAND2X1_46 ( .A(_abc_3576_new_n383_), .B(_abc_3576_new_n386_), .Y(_abc_3576_new_n388_));
NAND2X1 NAND2X1_47 ( .A(_abc_3576_new_n388_), .B(_abc_3576_new_n387_), .Y(_abc_3576_new_n389_));
NAND2X1 NAND2X1_48 ( .A(_abc_3576_new_n362_), .B(_abc_3576_new_n366_), .Y(_abc_3576_new_n395_));
NAND2X1 NAND2X1_49 ( .A(_abc_3576_new_n235_), .B(_abc_3576_new_n400_), .Y(_abc_3576_new_n401_));
NAND2X1 NAND2X1_5 ( .A(_abc_3576_new_n159_), .B(_abc_3576_new_n156_), .Y(_abc_3576_new_n160_));
NAND2X1 NAND2X1_50 ( .A(_abc_3576_new_n391_), .B(_abc_3576_new_n393_), .Y(_abc_3576_new_n402_));
NAND2X1 NAND2X1_51 ( .A(RMAX_REG_7_), .B(_abc_3576_new_n212_), .Y(_abc_3576_new_n537_));
NAND2X1 NAND2X1_52 ( .A(RMAX_REG_2_), .B(_abc_3576_new_n257_), .Y(_abc_3576_new_n542_));
NAND2X1 NAND2X1_53 ( .A(_abc_3576_new_n560_), .B(_abc_3576_new_n559_), .Y(_abc_3576_new_n561_));
NAND2X1 NAND2X1_54 ( .A(_abc_3576_new_n566_), .B(_abc_3576_new_n552_), .Y(_abc_3576_new_n567_));
NAND2X1 NAND2X1_55 ( .A(_abc_3576_new_n146_), .B(_abc_3576_new_n188_), .Y(_abc_3576_new_n593_));
NAND2X1 NAND2X1_6 ( .A(RESTART_bF_buf5), .B(RMAX_REG_0_), .Y(_abc_3576_new_n162_));
NAND2X1 NAND2X1_7 ( .A(RMIN_REG_0_), .B(RESTART_bF_buf3), .Y(_abc_3576_new_n165_));
NAND2X1 NAND2X1_8 ( .A(_abc_3576_new_n163_), .B(_abc_3576_new_n166_), .Y(_abc_3576_new_n167_));
NAND2X1 NAND2X1_9 ( .A(_abc_3576_new_n168_), .B(_abc_3576_new_n169_), .Y(_abc_3576_new_n170_));
NAND3X1 NAND3X1_1 ( .A(_abc_3576_new_n159_), .B(_abc_3576_new_n167_), .C(_abc_3576_new_n156_), .Y(_abc_3576_new_n174_));
NAND3X1 NAND3X1_10 ( .A(_abc_3576_new_n274_), .B(_abc_3576_new_n279_), .C(_abc_3576_new_n275_), .Y(n348));
NAND3X1 NAND3X1_11 ( .A(_abc_3576_new_n291_), .B(_abc_3576_new_n287_), .C(_abc_3576_new_n284_), .Y(_abc_3576_new_n292_));
NAND3X1 NAND3X1_12 ( .A(_abc_3576_new_n159_), .B(_abc_3576_new_n281_), .C(_abc_3576_new_n267_), .Y(_abc_3576_new_n299_));
NAND3X1 NAND3X1_13 ( .A(_abc_3576_new_n304_), .B(_abc_3576_new_n308_), .C(_abc_3576_new_n309_), .Y(n344));
NAND3X1 NAND3X1_14 ( .A(_abc_3576_new_n172_), .B(_abc_3576_new_n271_), .C(_abc_3576_new_n301_), .Y(_abc_3576_new_n318_));
NAND3X1 NAND3X1_15 ( .A(_abc_3576_new_n294_), .B(_abc_3576_new_n292_), .C(_abc_3576_new_n299_), .Y(_abc_3576_new_n326_));
NAND3X1 NAND3X1_16 ( .A(_abc_3576_new_n289_), .B(_abc_3576_new_n328_), .C(_abc_3576_new_n326_), .Y(_abc_3576_new_n333_));
NAND3X1 NAND3X1_17 ( .A(_abc_3576_new_n159_), .B(_abc_3576_new_n267_), .C(_abc_3576_new_n266_), .Y(_abc_3576_new_n339_));
NAND3X1 NAND3X1_18 ( .A(_abc_3576_new_n294_), .B(_abc_3576_new_n299_), .C(_abc_3576_new_n298_), .Y(_abc_3576_new_n342_));
NAND3X1 NAND3X1_19 ( .A(_abc_3576_new_n281_), .B(_abc_3576_new_n296_), .C(_abc_3576_new_n293_), .Y(_abc_3576_new_n343_));
NAND3X1 NAND3X1_2 ( .A(_abc_3576_new_n174_), .B(_abc_3576_new_n171_), .C(_abc_3576_new_n186_), .Y(_abc_3576_new_n187_));
NAND3X1 NAND3X1_20 ( .A(_abc_3576_new_n289_), .B(_abc_3576_new_n326_), .C(_abc_3576_new_n330_), .Y(_abc_3576_new_n346_));
NAND3X1 NAND3X1_21 ( .A(_abc_3576_new_n332_), .B(_abc_3576_new_n346_), .C(_abc_3576_new_n341_), .Y(_abc_3576_new_n349_));
NAND3X1 NAND3X1_22 ( .A(_abc_3576_new_n324_), .B(_abc_3576_new_n361_), .C(_abc_3576_new_n333_), .Y(_abc_3576_new_n362_));
NAND3X1 NAND3X1_23 ( .A(_abc_3576_new_n281_), .B(_abc_3576_new_n289_), .C(_abc_3576_new_n296_), .Y(_abc_3576_new_n364_));
NAND3X1 NAND3X1_24 ( .A(_abc_3576_new_n292_), .B(_abc_3576_new_n324_), .C(_abc_3576_new_n364_), .Y(_abc_3576_new_n365_));
NAND3X1 NAND3X1_25 ( .A(_abc_3576_new_n328_), .B(_abc_3576_new_n363_), .C(_abc_3576_new_n365_), .Y(_abc_3576_new_n366_));
NAND3X1 NAND3X1_26 ( .A(_abc_3576_new_n362_), .B(_abc_3576_new_n366_), .C(_abc_3576_new_n354_), .Y(_abc_3576_new_n367_));
NAND3X1 NAND3X1_27 ( .A(_abc_3576_new_n367_), .B(_abc_3576_new_n370_), .C(_abc_3576_new_n350_), .Y(_abc_3576_new_n373_));
NAND3X1 NAND3X1_28 ( .A(_abc_3576_new_n235_), .B(_abc_3576_new_n373_), .C(_abc_3576_new_n372_), .Y(_abc_3576_new_n374_));
NAND3X1 NAND3X1_29 ( .A(_abc_3576_new_n362_), .B(_abc_3576_new_n366_), .C(_abc_3576_new_n243_), .Y(_abc_3576_new_n375_));
NAND3X1 NAND3X1_3 ( .A(RESTART_bF_buf1), .B(_abc_3576_new_n210_), .C(_abc_3576_new_n209_), .Y(_abc_3576_new_n211_));
NAND3X1 NAND3X1_30 ( .A(_abc_3576_new_n378_), .B(_abc_3576_new_n374_), .C(_abc_3576_new_n375_), .Y(n336));
NAND3X1 NAND3X1_31 ( .A(_abc_3576_new_n324_), .B(_abc_3576_new_n359_), .C(_abc_3576_new_n333_), .Y(_abc_3576_new_n381_));
NAND3X1 NAND3X1_32 ( .A(_abc_3576_new_n360_), .B(_abc_3576_new_n390_), .C(_abc_3576_new_n381_), .Y(_abc_3576_new_n391_));
NAND3X1 NAND3X1_33 ( .A(_abc_3576_new_n328_), .B(_abc_3576_new_n360_), .C(_abc_3576_new_n365_), .Y(_abc_3576_new_n392_));
NAND3X1 NAND3X1_34 ( .A(_abc_3576_new_n359_), .B(_abc_3576_new_n389_), .C(_abc_3576_new_n392_), .Y(_abc_3576_new_n393_));
NAND3X1 NAND3X1_35 ( .A(_abc_3576_new_n359_), .B(_abc_3576_new_n390_), .C(_abc_3576_new_n392_), .Y(_abc_3576_new_n396_));
NAND3X1 NAND3X1_36 ( .A(_abc_3576_new_n360_), .B(_abc_3576_new_n389_), .C(_abc_3576_new_n381_), .Y(_abc_3576_new_n397_));
NAND3X1 NAND3X1_37 ( .A(_abc_3576_new_n380_), .B(_abc_3576_new_n402_), .C(_abc_3576_new_n235_), .Y(_abc_3576_new_n414_));
NAND3X1 NAND3X1_38 ( .A(_abc_3576_new_n188_), .B(RMIN_REG_0_), .C(_abc_3576_new_n567_), .Y(_abc_3576_new_n570_));
NAND3X1 NAND3X1_39 ( .A(nRESET_G_bF_buf3), .B(_abc_3576_new_n570_), .C(_abc_3576_new_n569_), .Y(n119));
NAND3X1 NAND3X1_4 ( .A(_abc_3576_new_n176_), .B(_abc_3576_new_n233_), .C(_abc_3576_new_n231_), .Y(_abc_3576_new_n234_));
NAND3X1 NAND3X1_40 ( .A(_abc_3576_new_n188_), .B(RMIN_REG_1_), .C(_abc_3576_new_n567_), .Y(_abc_3576_new_n573_));
NAND3X1 NAND3X1_41 ( .A(nRESET_G_bF_buf2), .B(_abc_3576_new_n573_), .C(_abc_3576_new_n572_), .Y(n114));
NAND3X1 NAND3X1_42 ( .A(_abc_3576_new_n188_), .B(RMIN_REG_2_), .C(_abc_3576_new_n567_), .Y(_abc_3576_new_n575_));
NAND3X1 NAND3X1_43 ( .A(nRESET_G_bF_buf1), .B(_abc_3576_new_n575_), .C(_abc_3576_new_n576_), .Y(n109));
NAND3X1 NAND3X1_44 ( .A(_abc_3576_new_n188_), .B(RMIN_REG_3_), .C(_abc_3576_new_n567_), .Y(_abc_3576_new_n579_));
NAND3X1 NAND3X1_45 ( .A(nRESET_G_bF_buf0), .B(_abc_3576_new_n579_), .C(_abc_3576_new_n578_), .Y(n104));
NAND3X1 NAND3X1_46 ( .A(_abc_3576_new_n188_), .B(RMIN_REG_4_), .C(_abc_3576_new_n567_), .Y(_abc_3576_new_n581_));
NAND3X1 NAND3X1_47 ( .A(nRESET_G_bF_buf3), .B(_abc_3576_new_n581_), .C(_abc_3576_new_n582_), .Y(n99));
NAND3X1 NAND3X1_48 ( .A(_abc_3576_new_n188_), .B(RMIN_REG_5_), .C(_abc_3576_new_n567_), .Y(_abc_3576_new_n584_));
NAND3X1 NAND3X1_49 ( .A(nRESET_G_bF_buf2), .B(_abc_3576_new_n584_), .C(_abc_3576_new_n585_), .Y(n94));
NAND3X1 NAND3X1_5 ( .A(_abc_3576_new_n173_), .B(_abc_3576_new_n187_), .C(_abc_3576_new_n235_), .Y(_abc_3576_new_n236_));
NAND3X1 NAND3X1_50 ( .A(_abc_3576_new_n188_), .B(RMIN_REG_6_), .C(_abc_3576_new_n567_), .Y(_abc_3576_new_n587_));
NAND3X1 NAND3X1_51 ( .A(nRESET_G_bF_buf1), .B(_abc_3576_new_n587_), .C(_abc_3576_new_n588_), .Y(n89));
NAND3X1 NAND3X1_52 ( .A(_abc_3576_new_n188_), .B(RMIN_REG_7_), .C(_abc_3576_new_n567_), .Y(_abc_3576_new_n590_));
NAND3X1 NAND3X1_53 ( .A(nRESET_G_bF_buf0), .B(_abc_3576_new_n590_), .C(_abc_3576_new_n591_), .Y(n84));
NAND3X1 NAND3X1_6 ( .A(_abc_3576_new_n159_), .B(_abc_3576_new_n156_), .C(_abc_3576_new_n175_), .Y(_abc_3576_new_n238_));
NAND3X1 NAND3X1_7 ( .A(_abc_3576_new_n237_), .B(_abc_3576_new_n238_), .C(_abc_3576_new_n243_), .Y(_abc_3576_new_n244_));
NAND3X1 NAND3X1_8 ( .A(_abc_3576_new_n236_), .B(_abc_3576_new_n254_), .C(_abc_3576_new_n244_), .Y(n352));
NAND3X1 NAND3X1_9 ( .A(_abc_3576_new_n272_), .B(_abc_3576_new_n273_), .C(_abc_3576_new_n235_), .Y(_abc_3576_new_n274_));
NOR2X1 NOR2X1_1 ( .A(_abc_3576_new_n160_), .B(_abc_3576_new_n171_), .Y(_abc_3576_new_n172_));
NOR2X1 NOR2X1_10 ( .A(_abc_3576_new_n282_), .B(_abc_3576_new_n247_), .Y(_abc_3576_new_n311_));
NOR2X1 NOR2X1_11 ( .A(_abc_3576_new_n311_), .B(_abc_3576_new_n314_), .Y(_abc_3576_new_n315_));
NOR2X1 NOR2X1_12 ( .A(_abc_3576_new_n325_), .B(_abc_3576_new_n329_), .Y(_abc_3576_new_n330_));
NOR2X1 NOR2X1_13 ( .A(_abc_3576_new_n335_), .B(_abc_3576_new_n319_), .Y(_abc_3576_new_n336_));
NOR2X1 NOR2X1_14 ( .A(STATO_REG_0_), .B(_abc_3576_new_n146_), .Y(_abc_3576_new_n419_));
NOR2X1 NOR2X1_15 ( .A(RMAX_REG_0_), .B(_abc_3576_new_n538_), .Y(_abc_3576_new_n539_));
NOR2X1 NOR2X1_16 ( .A(_abc_3576_new_n540_), .B(_abc_3576_new_n539_), .Y(_abc_3576_new_n541_));
NOR2X1 NOR2X1_17 ( .A(RMIN_REG_3_), .B(_abc_3576_new_n290_), .Y(_abc_3576_new_n553_));
NOR2X1 NOR2X1_18 ( .A(RESET_G), .B(_abc_3576_new_n593_), .Y(n361));
NOR2X1 NOR2X1_2 ( .A(_abc_3576_new_n168_), .B(_abc_3576_new_n169_), .Y(_abc_3576_new_n175_));
NOR2X1 NOR2X1_3 ( .A(_abc_3576_new_n224_), .B(_abc_3576_new_n221_), .Y(_abc_3576_new_n225_));
NOR2X1 NOR2X1_4 ( .A(_abc_3576_new_n226_), .B(_abc_3576_new_n225_), .Y(_abc_3576_new_n227_));
NOR2X1 NOR2X1_5 ( .A(AVERAGE), .B(_abc_3576_new_n232_), .Y(_abc_3576_new_n233_));
NOR2X1 NOR2X1_6 ( .A(RESTART_bF_buf0), .B(_abc_3576_new_n189_), .Y(_abc_3576_new_n245_));
NOR2X1 NOR2X1_7 ( .A(_abc_3576_new_n268_), .B(_abc_3576_new_n270_), .Y(_abc_3576_new_n271_));
NOR2X1 NOR2X1_8 ( .A(_abc_3576_new_n300_), .B(_abc_3576_new_n297_), .Y(_abc_3576_new_n301_));
NOR2X1 NOR2X1_9 ( .A(_abc_3576_new_n301_), .B(_abc_3576_new_n272_), .Y(_abc_3576_new_n303_));
NOR3X1 NOR3X1_1 ( .A(_abc_3576_new_n398_), .B(_abc_3576_new_n394_), .C(_abc_3576_new_n373_), .Y(_abc_3576_new_n399_));
OAI21X1 OAI21X1_1 ( .A(_abc_3576_new_n146_), .B(STATO_REG_0_), .C(_abc_3576_new_n148_), .Y(n356));
OAI21X1 OAI21X1_10 ( .A(_abc_3576_new_n204_), .B(_abc_3576_new_n201_), .C(_abc_3576_new_n206_), .Y(_abc_3576_new_n207_));
OAI21X1 OAI21X1_100 ( .A(_abc_3576_new_n212_), .B(_abc_3576_new_n509_), .C(nRESET_G_bF_buf0), .Y(_abc_3576_new_n534_));
OAI21X1 OAI21X1_101 ( .A(_abc_3576_new_n533_), .B(_abc_3576_new_n508_), .C(_abc_3576_new_n535_), .Y(n124));
OAI21X1 OAI21X1_102 ( .A(DATA_IN_1_), .B(_abc_3576_new_n183_), .C(DATA_IN_0_), .Y(_abc_3576_new_n538_));
OAI21X1 OAI21X1_103 ( .A(DATA_IN_3_), .B(_abc_3576_new_n286_), .C(_abc_3576_new_n542_), .Y(_abc_3576_new_n543_));
OAI21X1 OAI21X1_104 ( .A(_abc_3576_new_n543_), .B(_abc_3576_new_n541_), .C(_abc_3576_new_n544_), .Y(_abc_3576_new_n545_));
OAI21X1 OAI21X1_105 ( .A(DATA_IN_4_), .B(_abc_3576_new_n195_), .C(_abc_3576_new_n545_), .Y(_abc_3576_new_n546_));
OAI21X1 OAI21X1_106 ( .A(_abc_3576_new_n549_), .B(_abc_3576_new_n547_), .C(_abc_3576_new_n550_), .Y(_abc_3576_new_n551_));
OAI21X1 OAI21X1_107 ( .A(RMIN_REG_1_), .B(_abc_3576_new_n153_), .C(RMIN_REG_0_), .Y(_abc_3576_new_n554_));
OAI21X1 OAI21X1_108 ( .A(DATA_IN_0_), .B(_abc_3576_new_n554_), .C(_abc_3576_new_n555_), .Y(_abc_3576_new_n556_));
OAI21X1 OAI21X1_109 ( .A(_abc_3576_new_n257_), .B(RMIN_REG_2_), .C(_abc_3576_new_n556_), .Y(_abc_3576_new_n557_));
OAI21X1 OAI21X1_11 ( .A(_abc_3576_new_n192_), .B(_abc_3576_new_n193_), .C(_abc_3576_new_n207_), .Y(_abc_3576_new_n208_));
OAI21X1 OAI21X1_110 ( .A(_abc_3576_new_n553_), .B(_abc_3576_new_n557_), .C(_abc_3576_new_n558_), .Y(_abc_3576_new_n559_));
OAI21X1 OAI21X1_111 ( .A(DATA_IN_5_), .B(_abc_3576_new_n202_), .C(_abc_3576_new_n561_), .Y(_abc_3576_new_n562_));
OAI21X1 OAI21X1_112 ( .A(_abc_3576_new_n228_), .B(RMIN_REG_6_), .C(_abc_3576_new_n562_), .Y(_abc_3576_new_n563_));
OAI21X1 OAI21X1_113 ( .A(DATA_IN_7_), .B(_abc_3576_new_n190_), .C(STATO_REG_1_), .Y(_abc_3576_new_n565_));
OAI21X1 OAI21X1_114 ( .A(STATO_REG_0_), .B(_abc_3576_new_n568_), .C(DATA_IN_0_), .Y(_abc_3576_new_n569_));
OAI21X1 OAI21X1_115 ( .A(STATO_REG_0_), .B(_abc_3576_new_n568_), .C(DATA_IN_1_), .Y(_abc_3576_new_n572_));
OAI21X1 OAI21X1_116 ( .A(STATO_REG_0_), .B(_abc_3576_new_n568_), .C(DATA_IN_2_), .Y(_abc_3576_new_n576_));
OAI21X1 OAI21X1_117 ( .A(STATO_REG_0_), .B(_abc_3576_new_n568_), .C(DATA_IN_3_), .Y(_abc_3576_new_n578_));
OAI21X1 OAI21X1_118 ( .A(STATO_REG_0_), .B(_abc_3576_new_n568_), .C(DATA_IN_4_), .Y(_abc_3576_new_n582_));
OAI21X1 OAI21X1_119 ( .A(STATO_REG_0_), .B(_abc_3576_new_n568_), .C(DATA_IN_5_), .Y(_abc_3576_new_n585_));
OAI21X1 OAI21X1_12 ( .A(_abc_3576_new_n190_), .B(_abc_3576_new_n191_), .C(_abc_3576_new_n208_), .Y(_abc_3576_new_n209_));
OAI21X1 OAI21X1_120 ( .A(STATO_REG_0_), .B(_abc_3576_new_n568_), .C(DATA_IN_6_), .Y(_abc_3576_new_n588_));
OAI21X1 OAI21X1_121 ( .A(STATO_REG_0_), .B(_abc_3576_new_n568_), .C(DATA_IN_7_), .Y(_abc_3576_new_n591_));
OAI21X1 OAI21X1_122 ( .A(DATA_IN_7_), .B(_abc_3576_new_n191_), .C(_abc_3576_new_n551_), .Y(_abc_3576_new_n594_));
OAI21X1 OAI21X1_123 ( .A(STATO_REG_0_), .B(_abc_3576_new_n594_), .C(_abc_3576_new_n593_), .Y(_abc_3576_new_n595_));
OAI21X1 OAI21X1_124 ( .A(_abc_3576_new_n161_), .B(_abc_3576_new_n595_), .C(_abc_3576_new_n596_), .Y(n79));
OAI21X1 OAI21X1_125 ( .A(_abc_3576_new_n153_), .B(_abc_3576_new_n595_), .C(_abc_3576_new_n598_), .Y(n74));
OAI21X1 OAI21X1_126 ( .A(_abc_3576_new_n257_), .B(_abc_3576_new_n595_), .C(_abc_3576_new_n600_), .Y(n69));
OAI21X1 OAI21X1_127 ( .A(_abc_3576_new_n290_), .B(_abc_3576_new_n595_), .C(_abc_3576_new_n602_), .Y(n64));
OAI21X1 OAI21X1_128 ( .A(_abc_3576_new_n215_), .B(_abc_3576_new_n595_), .C(_abc_3576_new_n604_), .Y(n59));
OAI21X1 OAI21X1_129 ( .A(_abc_3576_new_n223_), .B(_abc_3576_new_n595_), .C(_abc_3576_new_n606_), .Y(n54));
OAI21X1 OAI21X1_13 ( .A(_abc_3576_new_n217_), .B(_abc_3576_new_n216_), .C(_abc_3576_new_n218_), .Y(_abc_3576_new_n219_));
OAI21X1 OAI21X1_130 ( .A(_abc_3576_new_n228_), .B(_abc_3576_new_n595_), .C(_abc_3576_new_n608_), .Y(n49));
OAI21X1 OAI21X1_131 ( .A(_abc_3576_new_n212_), .B(_abc_3576_new_n595_), .C(_abc_3576_new_n610_), .Y(n44));
OAI21X1 OAI21X1_14 ( .A(DATA_IN_3_), .B(REG4_REG_3_), .C(_abc_3576_new_n219_), .Y(_abc_3576_new_n220_));
OAI21X1 OAI21X1_15 ( .A(_abc_3576_new_n178_), .B(_abc_3576_new_n185_), .C(_abc_3576_new_n167_), .Y(_abc_3576_new_n237_));
OAI21X1 OAI21X1_16 ( .A(_abc_3576_new_n239_), .B(_abc_3576_new_n231_), .C(_abc_3576_new_n176_), .Y(_abc_3576_new_n240_));
OAI21X1 OAI21X1_17 ( .A(_abc_3576_new_n249_), .B(_abc_3576_new_n250_), .C(_abc_3576_new_n252_), .Y(_abc_3576_new_n253_));
OAI21X1 OAI21X1_18 ( .A(RESTART_bF_buf3), .B(_abc_3576_new_n257_), .C(_abc_3576_new_n258_), .Y(_abc_3576_new_n259_));
OAI21X1 OAI21X1_19 ( .A(RESTART_bF_buf1), .B(_abc_3576_new_n261_), .C(_abc_3576_new_n262_), .Y(_abc_3576_new_n263_));
OAI21X1 OAI21X1_2 ( .A(RESTART_bF_buf4), .B(_abc_3576_new_n150_), .C(_abc_3576_new_n151_), .Y(_abc_3576_new_n152_));
OAI21X1 OAI21X1_20 ( .A(_abc_3576_new_n152_), .B(_abc_3576_new_n155_), .C(_abc_3576_new_n175_), .Y(_abc_3576_new_n269_));
OAI21X1 OAI21X1_21 ( .A(_abc_3576_new_n268_), .B(_abc_3576_new_n270_), .C(_abc_3576_new_n173_), .Y(_abc_3576_new_n273_));
OAI21X1 OAI21X1_22 ( .A(_abc_3576_new_n276_), .B(_abc_3576_new_n250_), .C(_abc_3576_new_n277_), .Y(_abc_3576_new_n278_));
OAI21X1 OAI21X1_23 ( .A(RESTART_bF_buf4), .B(_abc_3576_new_n282_), .C(_abc_3576_new_n283_), .Y(_abc_3576_new_n284_));
OAI21X1 OAI21X1_24 ( .A(RESTART_bF_buf2), .B(DATA_IN_3_), .C(_abc_3576_new_n287_), .Y(_abc_3576_new_n288_));
OAI21X1 OAI21X1_25 ( .A(_abc_3576_new_n185_), .B(_abc_3576_new_n295_), .C(_abc_3576_new_n294_), .Y(_abc_3576_new_n296_));
OAI21X1 OAI21X1_26 ( .A(_abc_3576_new_n302_), .B(_abc_3576_new_n303_), .C(_abc_3576_new_n235_), .Y(_abc_3576_new_n304_));
OAI21X1 OAI21X1_27 ( .A(_abc_3576_new_n306_), .B(n356_bF_buf4), .C(nRESET_G_bF_buf2), .Y(_abc_3576_new_n307_));
OAI21X1 OAI21X1_28 ( .A(_abc_3576_new_n312_), .B(_abc_3576_new_n250_), .C(_abc_3576_new_n313_), .Y(_abc_3576_new_n314_));
OAI21X1 OAI21X1_29 ( .A(_abc_3576_new_n268_), .B(_abc_3576_new_n270_), .C(_abc_3576_new_n316_), .Y(_abc_3576_new_n317_));
OAI21X1 OAI21X1_3 ( .A(RESTART_bF_buf2), .B(_abc_3576_new_n153_), .C(_abc_3576_new_n154_), .Y(_abc_3576_new_n155_));
OAI21X1 OAI21X1_30 ( .A(_abc_3576_new_n317_), .B(_abc_3576_new_n301_), .C(_abc_3576_new_n318_), .Y(_abc_3576_new_n319_));
OAI21X1 OAI21X1_31 ( .A(RESTART_bF_buf0), .B(_abc_3576_new_n214_), .C(_abc_3576_new_n320_), .Y(_abc_3576_new_n321_));
OAI21X1 OAI21X1_32 ( .A(RESTART_bF_buf4), .B(_abc_3576_new_n215_), .C(_abc_3576_new_n322_), .Y(_abc_3576_new_n323_));
OAI21X1 OAI21X1_33 ( .A(_abc_3576_new_n325_), .B(_abc_3576_new_n333_), .C(_abc_3576_new_n332_), .Y(_abc_3576_new_n334_));
OAI21X1 OAI21X1_34 ( .A(_abc_3576_new_n185_), .B(_abc_3576_new_n295_), .C(_abc_3576_new_n337_), .Y(_abc_3576_new_n338_));
OAI21X1 OAI21X1_35 ( .A(_abc_3576_new_n297_), .B(_abc_3576_new_n300_), .C(_abc_3576_new_n340_), .Y(_abc_3576_new_n341_));
OAI21X1 OAI21X1_36 ( .A(_abc_3576_new_n345_), .B(_abc_3576_new_n347_), .C(_abc_3576_new_n344_), .Y(_abc_3576_new_n348_));
OAI21X1 OAI21X1_37 ( .A(_abc_3576_new_n336_), .B(_abc_3576_new_n352_), .C(_abc_3576_new_n315_), .Y(n340));
OAI21X1 OAI21X1_38 ( .A(RESTART_bF_buf2), .B(DATA_IN_5_), .C(_abc_3576_new_n355_), .Y(_abc_3576_new_n356_));
OAI21X1 OAI21X1_39 ( .A(RESTART_bF_buf0), .B(REG4_REG_5_), .C(_abc_3576_new_n357_), .Y(_abc_3576_new_n358_));
OAI21X1 OAI21X1_4 ( .A(RESTART_bF_buf4), .B(_abc_3576_new_n161_), .C(_abc_3576_new_n162_), .Y(_abc_3576_new_n163_));
OAI21X1 OAI21X1_40 ( .A(_abc_3576_new_n368_), .B(_abc_3576_new_n369_), .C(_abc_3576_new_n348_), .Y(_abc_3576_new_n370_));
OAI21X1 OAI21X1_41 ( .A(_abc_3576_new_n214_), .B(_abc_3576_new_n247_), .C(_abc_3576_new_n376_), .Y(_abc_3576_new_n377_));
OAI21X1 OAI21X1_42 ( .A(_abc_3576_new_n368_), .B(_abc_3576_new_n369_), .C(_abc_3576_new_n354_), .Y(_abc_3576_new_n380_));
OAI21X1 OAI21X1_43 ( .A(RESTART_bF_buf4), .B(_abc_3576_new_n229_), .C(_abc_3576_new_n382_), .Y(_abc_3576_new_n383_));
OAI21X1 OAI21X1_44 ( .A(RESTART_bF_buf2), .B(_abc_3576_new_n228_), .C(_abc_3576_new_n384_), .Y(_abc_3576_new_n385_));
OAI21X1 OAI21X1_45 ( .A(_abc_3576_new_n398_), .B(_abc_3576_new_n394_), .C(_abc_3576_new_n373_), .Y(_abc_3576_new_n400_));
OAI21X1 OAI21X1_46 ( .A(_abc_3576_new_n404_), .B(n356_bF_buf3), .C(nRESET_G_bF_buf1), .Y(_abc_3576_new_n405_));
OAI21X1 OAI21X1_47 ( .A(_abc_3576_new_n403_), .B(_abc_3576_new_n250_), .C(_abc_3576_new_n406_), .Y(_abc_3576_new_n407_));
OAI21X1 OAI21X1_48 ( .A(_abc_3576_new_n399_), .B(_abc_3576_new_n401_), .C(_abc_3576_new_n408_), .Y(n332));
OAI21X1 OAI21X1_49 ( .A(_abc_3576_new_n410_), .B(_abc_3576_new_n250_), .C(_abc_3576_new_n411_), .Y(_abc_3576_new_n412_));
OAI21X1 OAI21X1_5 ( .A(RESTART_bF_buf2), .B(_abc_3576_new_n164_), .C(_abc_3576_new_n165_), .Y(_abc_3576_new_n166_));
OAI21X1 OAI21X1_50 ( .A(_abc_3576_new_n373_), .B(_abc_3576_new_n414_), .C(_abc_3576_new_n413_), .Y(n328));
OAI21X1 OAI21X1_51 ( .A(_abc_3576_new_n213_), .B(_abc_3576_new_n247_), .C(_abc_3576_new_n417_), .Y(n324));
OAI21X1 OAI21X1_52 ( .A(_abc_3576_new_n164_), .B(n356_bF_buf2), .C(_abc_3576_new_n420_), .Y(n319));
OAI21X1 OAI21X1_53 ( .A(_abc_3576_new_n150_), .B(n356_bF_buf1), .C(_abc_3576_new_n422_), .Y(n314));
OAI21X1 OAI21X1_54 ( .A(_abc_3576_new_n261_), .B(n356_bF_buf0), .C(_abc_3576_new_n424_), .Y(n309));
OAI21X1 OAI21X1_55 ( .A(_abc_3576_new_n282_), .B(n356_bF_buf5), .C(_abc_3576_new_n426_), .Y(n304));
OAI21X1 OAI21X1_56 ( .A(_abc_3576_new_n214_), .B(n356_bF_buf4), .C(_abc_3576_new_n428_), .Y(n299));
OAI21X1 OAI21X1_57 ( .A(_abc_3576_new_n222_), .B(n356_bF_buf3), .C(_abc_3576_new_n430_), .Y(n294));
OAI21X1 OAI21X1_58 ( .A(_abc_3576_new_n229_), .B(n356_bF_buf2), .C(_abc_3576_new_n432_), .Y(n289));
OAI21X1 OAI21X1_59 ( .A(_abc_3576_new_n213_), .B(n356_bF_buf1), .C(_abc_3576_new_n434_), .Y(n284));
OAI21X1 OAI21X1_6 ( .A(_abc_3576_new_n178_), .B(_abc_3576_new_n185_), .C(_abc_3576_new_n175_), .Y(_abc_3576_new_n186_));
OAI21X1 OAI21X1_60 ( .A(_abc_3576_new_n436_), .B(n356_bF_buf0), .C(_abc_3576_new_n437_), .Y(n279));
OAI21X1 OAI21X1_61 ( .A(_abc_3576_new_n439_), .B(n356_bF_buf5), .C(_abc_3576_new_n440_), .Y(n274));
OAI21X1 OAI21X1_62 ( .A(_abc_3576_new_n442_), .B(n356_bF_buf4), .C(_abc_3576_new_n443_), .Y(n269));
OAI21X1 OAI21X1_63 ( .A(_abc_3576_new_n445_), .B(n356_bF_buf3), .C(_abc_3576_new_n446_), .Y(n264));
OAI21X1 OAI21X1_64 ( .A(_abc_3576_new_n448_), .B(n356_bF_buf2), .C(_abc_3576_new_n449_), .Y(n259));
OAI21X1 OAI21X1_65 ( .A(_abc_3576_new_n451_), .B(n356_bF_buf1), .C(_abc_3576_new_n452_), .Y(n254));
OAI21X1 OAI21X1_66 ( .A(_abc_3576_new_n454_), .B(n356_bF_buf0), .C(_abc_3576_new_n455_), .Y(n249));
OAI21X1 OAI21X1_67 ( .A(_abc_3576_new_n457_), .B(n356_bF_buf5), .C(_abc_3576_new_n458_), .Y(n244));
OAI21X1 OAI21X1_68 ( .A(_abc_3576_new_n460_), .B(n356_bF_buf4), .C(_abc_3576_new_n461_), .Y(n239));
OAI21X1 OAI21X1_69 ( .A(_abc_3576_new_n463_), .B(n356_bF_buf3), .C(_abc_3576_new_n464_), .Y(n234));
OAI21X1 OAI21X1_7 ( .A(_abc_3576_new_n147__bF_buf4), .B(_abc_3576_new_n188_), .C(STATO_REG_1_), .Y(_abc_3576_new_n189_));
OAI21X1 OAI21X1_70 ( .A(_abc_3576_new_n466_), .B(n356_bF_buf2), .C(_abc_3576_new_n467_), .Y(n229));
OAI21X1 OAI21X1_71 ( .A(_abc_3576_new_n469_), .B(n356_bF_buf1), .C(_abc_3576_new_n470_), .Y(n224));
OAI21X1 OAI21X1_72 ( .A(_abc_3576_new_n472_), .B(n356_bF_buf0), .C(_abc_3576_new_n473_), .Y(n219));
OAI21X1 OAI21X1_73 ( .A(_abc_3576_new_n475_), .B(n356_bF_buf5), .C(_abc_3576_new_n476_), .Y(n214));
OAI21X1 OAI21X1_74 ( .A(_abc_3576_new_n478_), .B(n356_bF_buf4), .C(_abc_3576_new_n479_), .Y(n209));
OAI21X1 OAI21X1_75 ( .A(_abc_3576_new_n481_), .B(n356_bF_buf3), .C(_abc_3576_new_n482_), .Y(n204));
OAI21X1 OAI21X1_76 ( .A(_abc_3576_new_n484_), .B(n356_bF_buf2), .C(_abc_3576_new_n485_), .Y(n199));
OAI21X1 OAI21X1_77 ( .A(_abc_3576_new_n487_), .B(n356_bF_buf1), .C(_abc_3576_new_n488_), .Y(n194));
OAI21X1 OAI21X1_78 ( .A(_abc_3576_new_n490_), .B(n356_bF_buf0), .C(_abc_3576_new_n491_), .Y(n189));
OAI21X1 OAI21X1_79 ( .A(_abc_3576_new_n493_), .B(n356_bF_buf5), .C(_abc_3576_new_n494_), .Y(n184));
OAI21X1 OAI21X1_8 ( .A(_abc_3576_new_n197_), .B(_abc_3576_new_n196_), .C(_abc_3576_new_n198_), .Y(_abc_3576_new_n199_));
OAI21X1 OAI21X1_80 ( .A(_abc_3576_new_n496_), .B(n356_bF_buf4), .C(_abc_3576_new_n497_), .Y(n179));
OAI21X1 OAI21X1_81 ( .A(_abc_3576_new_n499_), .B(n356_bF_buf3), .C(_abc_3576_new_n500_), .Y(n174));
OAI21X1 OAI21X1_82 ( .A(_abc_3576_new_n502_), .B(n356_bF_buf2), .C(_abc_3576_new_n503_), .Y(n169));
OAI21X1 OAI21X1_83 ( .A(_abc_3576_new_n505_), .B(n356_bF_buf1), .C(_abc_3576_new_n506_), .Y(n164));
OAI21X1 OAI21X1_84 ( .A(_abc_3576_new_n146_), .B(_abc_3576_new_n232_), .C(_abc_3576_new_n188_), .Y(_abc_3576_new_n508_));
OAI21X1 OAI21X1_85 ( .A(STATO_REG_0_), .B(ENABLE), .C(STATO_REG_1_), .Y(_abc_3576_new_n509_));
OAI21X1 OAI21X1_86 ( .A(_abc_3576_new_n161_), .B(_abc_3576_new_n509_), .C(nRESET_G_bF_buf3), .Y(_abc_3576_new_n510_));
OAI21X1 OAI21X1_87 ( .A(_abc_3576_new_n249_), .B(_abc_3576_new_n508_), .C(_abc_3576_new_n511_), .Y(n159));
OAI21X1 OAI21X1_88 ( .A(_abc_3576_new_n153_), .B(_abc_3576_new_n509_), .C(nRESET_G_bF_buf2), .Y(_abc_3576_new_n513_));
OAI21X1 OAI21X1_89 ( .A(_abc_3576_new_n276_), .B(_abc_3576_new_n508_), .C(_abc_3576_new_n514_), .Y(n154));
OAI21X1 OAI21X1_9 ( .A(RMIN_REG_3_), .B(RMAX_REG_3_), .C(_abc_3576_new_n199_), .Y(_abc_3576_new_n200_));
OAI21X1 OAI21X1_90 ( .A(_abc_3576_new_n257_), .B(_abc_3576_new_n509_), .C(nRESET_G_bF_buf1), .Y(_abc_3576_new_n517_));
OAI21X1 OAI21X1_91 ( .A(_abc_3576_new_n516_), .B(_abc_3576_new_n508_), .C(_abc_3576_new_n518_), .Y(n149));
OAI21X1 OAI21X1_92 ( .A(_abc_3576_new_n290_), .B(_abc_3576_new_n509_), .C(nRESET_G_bF_buf0), .Y(_abc_3576_new_n520_));
OAI21X1 OAI21X1_93 ( .A(_abc_3576_new_n312_), .B(_abc_3576_new_n508_), .C(_abc_3576_new_n521_), .Y(n144));
OAI21X1 OAI21X1_94 ( .A(_abc_3576_new_n215_), .B(_abc_3576_new_n509_), .C(nRESET_G_bF_buf3), .Y(_abc_3576_new_n524_));
OAI21X1 OAI21X1_95 ( .A(_abc_3576_new_n523_), .B(_abc_3576_new_n508_), .C(_abc_3576_new_n525_), .Y(n139));
OAI21X1 OAI21X1_96 ( .A(_abc_3576_new_n223_), .B(_abc_3576_new_n509_), .C(nRESET_G_bF_buf2), .Y(_abc_3576_new_n527_));
OAI21X1 OAI21X1_97 ( .A(_abc_3576_new_n403_), .B(_abc_3576_new_n508_), .C(_abc_3576_new_n528_), .Y(n134));
OAI21X1 OAI21X1_98 ( .A(_abc_3576_new_n228_), .B(_abc_3576_new_n509_), .C(nRESET_G_bF_buf1), .Y(_abc_3576_new_n530_));
OAI21X1 OAI21X1_99 ( .A(_abc_3576_new_n410_), .B(_abc_3576_new_n508_), .C(_abc_3576_new_n531_), .Y(n129));
OAI22X1 OAI22X1_1 ( .A(RMIN_REG_1_), .B(RMAX_REG_1_), .C(RMIN_REG_2_), .D(RMAX_REG_2_), .Y(_abc_3576_new_n197_));
OAI22X1 OAI22X1_10 ( .A(RMAX_REG_1_), .B(_abc_3576_new_n153_), .C(_abc_3576_new_n257_), .D(RMAX_REG_2_), .Y(_abc_3576_new_n540_));
OAI22X1 OAI22X1_2 ( .A(_abc_3576_new_n202_), .B(_abc_3576_new_n203_), .C(_abc_3576_new_n194_), .D(_abc_3576_new_n195_), .Y(_abc_3576_new_n204_));
OAI22X1 OAI22X1_3 ( .A(RMIN_REG_5_), .B(RMAX_REG_5_), .C(RMAX_REG_6_), .D(RMIN_REG_6_), .Y(_abc_3576_new_n205_));
OAI22X1 OAI22X1_4 ( .A(REG4_REG_1_), .B(DATA_IN_1_), .C(REG4_REG_2_), .D(DATA_IN_2_), .Y(_abc_3576_new_n217_));
OAI22X1 OAI22X1_5 ( .A(_abc_3576_new_n222_), .B(_abc_3576_new_n223_), .C(_abc_3576_new_n214_), .D(_abc_3576_new_n215_), .Y(_abc_3576_new_n224_));
OAI22X1 OAI22X1_6 ( .A(DATA_IN_6_), .B(REG4_REG_6_), .C(REG4_REG_5_), .D(DATA_IN_5_), .Y(_abc_3576_new_n226_));
OAI22X1 OAI22X1_7 ( .A(DATA_IN_7_), .B(REG4_REG_7_), .C(_abc_3576_new_n228_), .D(_abc_3576_new_n229_), .Y(_abc_3576_new_n230_));
OAI22X1 OAI22X1_8 ( .A(_abc_3576_new_n212_), .B(_abc_3576_new_n213_), .C(_abc_3576_new_n230_), .D(_abc_3576_new_n227_), .Y(_abc_3576_new_n231_));
OAI22X1 OAI22X1_9 ( .A(_abc_3576_new_n168_), .B(_abc_3576_new_n169_), .C(_abc_3576_new_n157_), .D(_abc_3576_new_n158_), .Y(_abc_3576_new_n267_));
OR2X2 OR2X2_1 ( .A(RESTART_bF_buf4), .B(REG4_REG_1_), .Y(_abc_3576_new_n179_));
OR2X2 OR2X2_2 ( .A(_abc_3576_new_n321_), .B(_abc_3576_new_n323_), .Y(_abc_3576_new_n328_));
OR2X2 OR2X2_3 ( .A(_abc_3576_new_n356_), .B(_abc_3576_new_n358_), .Y(_abc_3576_new_n359_));
OR2X2 OR2X2_4 ( .A(_abc_3576_new_n386_), .B(_abc_3576_new_n383_), .Y(_abc_3576_new_n387_));


endmodule