
module xtea(clock, reset, mode, \data_in1[0] , \data_in1[1] , \data_in1[2] , \data_in1[3] , \data_in1[4] , \data_in1[5] , \data_in1[6] , \data_in1[7] , \data_in1[8] , \data_in1[9] , \data_in1[10] , \data_in1[11] , \data_in1[12] , \data_in1[13] , \data_in1[14] , \data_in1[15] , \data_in1[16] , \data_in1[17] , \data_in1[18] , \data_in1[19] , \data_in1[20] , \data_in1[21] , \data_in1[22] , \data_in1[23] , \data_in1[24] , \data_in1[25] , \data_in1[26] , \data_in1[27] , \data_in1[28] , \data_in1[29] , \data_in1[30] , \data_in1[31] , \data_in2[0] , \data_in2[1] , \data_in2[2] , \data_in2[3] , \data_in2[4] , \data_in2[5] , \data_in2[6] , \data_in2[7] , \data_in2[8] , \data_in2[9] , \data_in2[10] , \data_in2[11] , \data_in2[12] , \data_in2[13] , \data_in2[14] , \data_in2[15] , \data_in2[16] , \data_in2[17] , \data_in2[18] , \data_in2[19] , \data_in2[20] , \data_in2[21] , \data_in2[22] , \data_in2[23] , \data_in2[24] , \data_in2[25] , \data_in2[26] , \data_in2[27] , \data_in2[28] , \data_in2[29] , \data_in2[30] , \data_in2[31] , \key_in[0] , \key_in[1] , \key_in[2] , \key_in[3] , \key_in[4] , \key_in[5] , \key_in[6] , \key_in[7] , \key_in[8] , \key_in[9] , \key_in[10] , \key_in[11] , \key_in[12] , \key_in[13] , \key_in[14] , \key_in[15] , \key_in[16] , \key_in[17] , \key_in[18] , \key_in[19] , \key_in[20] , \key_in[21] , \key_in[22] , \key_in[23] , \key_in[24] , \key_in[25] , \key_in[26] , \key_in[27] , \key_in[28] , \key_in[29] , \key_in[30] , \key_in[31] , \key_in[32] , \key_in[33] , \key_in[34] , \key_in[35] , \key_in[36] , \key_in[37] , \key_in[38] , \key_in[39] , \key_in[40] , \key_in[41] , \key_in[42] , \key_in[43] , \key_in[44] , \key_in[45] , \key_in[46] , \key_in[47] , \key_in[48] , \key_in[49] , \key_in[50] , \key_in[51] , \key_in[52] , \key_in[53] , \key_in[54] , \key_in[55] , \key_in[56] , \key_in[57] , \key_in[58] , \key_in[59] , \key_in[60] , \key_in[61] , \key_in[62] , \key_in[63] , \key_in[64] , \key_in[65] , \key_in[66] , \key_in[67] , \key_in[68] , \key_in[69] , \key_in[70] , \key_in[71] , \key_in[72] , \key_in[73] , \key_in[74] , \key_in[75] , \key_in[76] , \key_in[77] , \key_in[78] , \key_in[79] , \key_in[80] , \key_in[81] , \key_in[82] , \key_in[83] , \key_in[84] , \key_in[85] , \key_in[86] , \key_in[87] , \key_in[88] , \key_in[89] , \key_in[90] , \key_in[91] , \key_in[92] , \key_in[93] , \key_in[94] , \key_in[95] , \key_in[96] , \key_in[97] , \key_in[98] , \key_in[99] , \key_in[100] , \key_in[101] , \key_in[102] , \key_in[103] , \key_in[104] , \key_in[105] , \key_in[106] , \key_in[107] , \key_in[108] , \key_in[109] , \key_in[110] , \key_in[111] , \key_in[112] , \key_in[113] , \key_in[114] , \key_in[115] , \key_in[116] , \key_in[117] , \key_in[118] , \key_in[119] , \key_in[120] , \key_in[121] , \key_in[122] , \key_in[123] , \key_in[124] , \key_in[125] , \key_in[126] , \key_in[127] , \data_out1[0] , \data_out1[1] , \data_out1[2] , \data_out1[3] , \data_out1[4] , \data_out1[5] , \data_out1[6] , \data_out1[7] , \data_out1[8] , \data_out1[9] , \data_out1[10] , \data_out1[11] , \data_out1[12] , \data_out1[13] , \data_out1[14] , \data_out1[15] , \data_out1[16] , \data_out1[17] , \data_out1[18] , \data_out1[19] , \data_out1[20] , \data_out1[21] , \data_out1[22] , \data_out1[23] , \data_out1[24] , \data_out1[25] , \data_out1[26] , \data_out1[27] , \data_out1[28] , \data_out1[29] , \data_out1[30] , \data_out1[31] , \data_out2[0] , \data_out2[1] , \data_out2[2] , \data_out2[3] , \data_out2[4] , \data_out2[5] , \data_out2[6] , \data_out2[7] , \data_out2[8] , \data_out2[9] , \data_out2[10] , \data_out2[11] , \data_out2[12] , \data_out2[13] , \data_out2[14] , \data_out2[15] , \data_out2[16] , \data_out2[17] , \data_out2[18] , \data_out2[19] , \data_out2[20] , \data_out2[21] , \data_out2[22] , \data_out2[23] , \data_out2[24] , \data_out2[25] , \data_out2[26] , \data_out2[27] , \data_out2[28] , \data_out2[29] , \data_out2[30] , \data_out2[31] , all_done);
  wire _abc_10892_n1037;
  wire _abc_10892_n1125;
  wire _abc_10892_n6074;
  wire _abc_10892_n7323;
  wire _abc_10892_n7419;
  wire _abc_17692_n1000;
  wire _abc_17692_n10000;
  wire _abc_17692_n10001;
  wire _abc_17692_n10002;
  wire _abc_17692_n10003;
  wire _abc_17692_n10004;
  wire _abc_17692_n10005;
  wire _abc_17692_n10006;
  wire _abc_17692_n10007;
  wire _abc_17692_n10008;
  wire _abc_17692_n10009;
  wire _abc_17692_n1001;
  wire _abc_17692_n10010;
  wire _abc_17692_n10011;
  wire _abc_17692_n10012;
  wire _abc_17692_n10013;
  wire _abc_17692_n10014;
  wire _abc_17692_n10015;
  wire _abc_17692_n10016;
  wire _abc_17692_n10017;
  wire _abc_17692_n10018;
  wire _abc_17692_n10019;
  wire _abc_17692_n1002;
  wire _abc_17692_n10020;
  wire _abc_17692_n10021;
  wire _abc_17692_n10022;
  wire _abc_17692_n10023;
  wire _abc_17692_n10024;
  wire _abc_17692_n10025;
  wire _abc_17692_n10026;
  wire _abc_17692_n10027;
  wire _abc_17692_n10028;
  wire _abc_17692_n10029;
  wire _abc_17692_n1003;
  wire _abc_17692_n10030;
  wire _abc_17692_n10031;
  wire _abc_17692_n10032;
  wire _abc_17692_n10033;
  wire _abc_17692_n10034;
  wire _abc_17692_n10035;
  wire _abc_17692_n10036;
  wire _abc_17692_n10037;
  wire _abc_17692_n10038;
  wire _abc_17692_n10039;
  wire _abc_17692_n1004;
  wire _abc_17692_n10040;
  wire _abc_17692_n10041;
  wire _abc_17692_n10042;
  wire _abc_17692_n10043;
  wire _abc_17692_n10044;
  wire _abc_17692_n10045;
  wire _abc_17692_n10046;
  wire _abc_17692_n10047;
  wire _abc_17692_n10048;
  wire _abc_17692_n10049;
  wire _abc_17692_n1005;
  wire _abc_17692_n10050;
  wire _abc_17692_n10051;
  wire _abc_17692_n10052;
  wire _abc_17692_n10053;
  wire _abc_17692_n10054;
  wire _abc_17692_n10055;
  wire _abc_17692_n10056;
  wire _abc_17692_n10057;
  wire _abc_17692_n10058;
  wire _abc_17692_n10059;
  wire _abc_17692_n1006;
  wire _abc_17692_n10060;
  wire _abc_17692_n10061;
  wire _abc_17692_n10062;
  wire _abc_17692_n10063;
  wire _abc_17692_n10064;
  wire _abc_17692_n10065;
  wire _abc_17692_n10067;
  wire _abc_17692_n10068;
  wire _abc_17692_n10069;
  wire _abc_17692_n1007;
  wire _abc_17692_n10070;
  wire _abc_17692_n10071;
  wire _abc_17692_n10072;
  wire _abc_17692_n10073;
  wire _abc_17692_n10074;
  wire _abc_17692_n10075;
  wire _abc_17692_n10076;
  wire _abc_17692_n10077;
  wire _abc_17692_n10078;
  wire _abc_17692_n10079;
  wire _abc_17692_n1008;
  wire _abc_17692_n10080;
  wire _abc_17692_n10081;
  wire _abc_17692_n10082;
  wire _abc_17692_n10083;
  wire _abc_17692_n10084;
  wire _abc_17692_n10085;
  wire _abc_17692_n10086;
  wire _abc_17692_n10087;
  wire _abc_17692_n10088;
  wire _abc_17692_n10089;
  wire _abc_17692_n1009;
  wire _abc_17692_n10090;
  wire _abc_17692_n10091;
  wire _abc_17692_n10092;
  wire _abc_17692_n10093;
  wire _abc_17692_n10094;
  wire _abc_17692_n10095;
  wire _abc_17692_n10096;
  wire _abc_17692_n10097;
  wire _abc_17692_n10098;
  wire _abc_17692_n10099;
  wire _abc_17692_n1010;
  wire _abc_17692_n10100;
  wire _abc_17692_n10101;
  wire _abc_17692_n10102;
  wire _abc_17692_n10103;
  wire _abc_17692_n10104;
  wire _abc_17692_n10105;
  wire _abc_17692_n10106;
  wire _abc_17692_n10107;
  wire _abc_17692_n10108;
  wire _abc_17692_n10109;
  wire _abc_17692_n1011;
  wire _abc_17692_n10110;
  wire _abc_17692_n10111;
  wire _abc_17692_n10112;
  wire _abc_17692_n10113;
  wire _abc_17692_n10114;
  wire _abc_17692_n10115;
  wire _abc_17692_n10116;
  wire _abc_17692_n10117;
  wire _abc_17692_n10118;
  wire _abc_17692_n10119;
  wire _abc_17692_n1012;
  wire _abc_17692_n10120;
  wire _abc_17692_n10121;
  wire _abc_17692_n10122;
  wire _abc_17692_n10123;
  wire _abc_17692_n10124;
  wire _abc_17692_n10125;
  wire _abc_17692_n10126;
  wire _abc_17692_n10127;
  wire _abc_17692_n10128;
  wire _abc_17692_n10129;
  wire _abc_17692_n1013;
  wire _abc_17692_n10130;
  wire _abc_17692_n10131;
  wire _abc_17692_n10132;
  wire _abc_17692_n10133;
  wire _abc_17692_n10134;
  wire _abc_17692_n10135;
  wire _abc_17692_n10136;
  wire _abc_17692_n10137;
  wire _abc_17692_n10138;
  wire _abc_17692_n10139;
  wire _abc_17692_n1014;
  wire _abc_17692_n10140;
  wire _abc_17692_n10141;
  wire _abc_17692_n10142;
  wire _abc_17692_n10143;
  wire _abc_17692_n10144;
  wire _abc_17692_n10145;
  wire _abc_17692_n10146;
  wire _abc_17692_n10147;
  wire _abc_17692_n10148;
  wire _abc_17692_n10149;
  wire _abc_17692_n1015;
  wire _abc_17692_n10150;
  wire _abc_17692_n10151;
  wire _abc_17692_n10152;
  wire _abc_17692_n10153;
  wire _abc_17692_n10154;
  wire _abc_17692_n10155;
  wire _abc_17692_n10156;
  wire _abc_17692_n10157;
  wire _abc_17692_n10158;
  wire _abc_17692_n10159;
  wire _abc_17692_n1016;
  wire _abc_17692_n10160;
  wire _abc_17692_n10161;
  wire _abc_17692_n10162;
  wire _abc_17692_n10163;
  wire _abc_17692_n10164;
  wire _abc_17692_n10165;
  wire _abc_17692_n10166;
  wire _abc_17692_n10167;
  wire _abc_17692_n10168;
  wire _abc_17692_n10169;
  wire _abc_17692_n1017;
  wire _abc_17692_n10170;
  wire _abc_17692_n10171;
  wire _abc_17692_n10172;
  wire _abc_17692_n10173;
  wire _abc_17692_n10174;
  wire _abc_17692_n10175;
  wire _abc_17692_n10176;
  wire _abc_17692_n10177;
  wire _abc_17692_n10178;
  wire _abc_17692_n10179;
  wire _abc_17692_n1018;
  wire _abc_17692_n10180;
  wire _abc_17692_n10181;
  wire _abc_17692_n10182;
  wire _abc_17692_n10184;
  wire _abc_17692_n10185;
  wire _abc_17692_n10186;
  wire _abc_17692_n10187;
  wire _abc_17692_n10188;
  wire _abc_17692_n10189;
  wire _abc_17692_n1019;
  wire _abc_17692_n10190;
  wire _abc_17692_n10191;
  wire _abc_17692_n10192;
  wire _abc_17692_n10193;
  wire _abc_17692_n10194;
  wire _abc_17692_n10195;
  wire _abc_17692_n10196;
  wire _abc_17692_n10197;
  wire _abc_17692_n10198;
  wire _abc_17692_n10199;
  wire _abc_17692_n10200;
  wire _abc_17692_n10201;
  wire _abc_17692_n10202;
  wire _abc_17692_n10203;
  wire _abc_17692_n10204;
  wire _abc_17692_n10205;
  wire _abc_17692_n10206;
  wire _abc_17692_n10207;
  wire _abc_17692_n10208;
  wire _abc_17692_n10209;
  wire _abc_17692_n1021;
  wire _abc_17692_n10210;
  wire _abc_17692_n10211;
  wire _abc_17692_n10212;
  wire _abc_17692_n10213;
  wire _abc_17692_n10214;
  wire _abc_17692_n10215;
  wire _abc_17692_n10216;
  wire _abc_17692_n10217;
  wire _abc_17692_n10218;
  wire _abc_17692_n10219;
  wire _abc_17692_n1022;
  wire _abc_17692_n10220;
  wire _abc_17692_n10221;
  wire _abc_17692_n10222;
  wire _abc_17692_n10223;
  wire _abc_17692_n10224;
  wire _abc_17692_n10225;
  wire _abc_17692_n10226;
  wire _abc_17692_n10227;
  wire _abc_17692_n10228;
  wire _abc_17692_n10229;
  wire _abc_17692_n1023;
  wire _abc_17692_n10230;
  wire _abc_17692_n10231;
  wire _abc_17692_n10232;
  wire _abc_17692_n10233;
  wire _abc_17692_n10234;
  wire _abc_17692_n10235;
  wire _abc_17692_n10236;
  wire _abc_17692_n10237;
  wire _abc_17692_n10238;
  wire _abc_17692_n10239;
  wire _abc_17692_n1024;
  wire _abc_17692_n10240;
  wire _abc_17692_n10241;
  wire _abc_17692_n10242;
  wire _abc_17692_n10243;
  wire _abc_17692_n10244;
  wire _abc_17692_n10245;
  wire _abc_17692_n10246;
  wire _abc_17692_n10247;
  wire _abc_17692_n10248;
  wire _abc_17692_n10249;
  wire _abc_17692_n10250;
  wire _abc_17692_n10251;
  wire _abc_17692_n10252;
  wire _abc_17692_n10253;
  wire _abc_17692_n10254;
  wire _abc_17692_n10255;
  wire _abc_17692_n10256;
  wire _abc_17692_n10257;
  wire _abc_17692_n10258;
  wire _abc_17692_n10259;
  wire _abc_17692_n1025_1;
  wire _abc_17692_n1026;
  wire _abc_17692_n10260;
  wire _abc_17692_n10261;
  wire _abc_17692_n10262;
  wire _abc_17692_n10263;
  wire _abc_17692_n10264;
  wire _abc_17692_n10265;
  wire _abc_17692_n10266;
  wire _abc_17692_n10267;
  wire _abc_17692_n10268;
  wire _abc_17692_n10269;
  wire _abc_17692_n1027;
  wire _abc_17692_n10270;
  wire _abc_17692_n10271;
  wire _abc_17692_n10272;
  wire _abc_17692_n10273;
  wire _abc_17692_n10274;
  wire _abc_17692_n10275;
  wire _abc_17692_n10276;
  wire _abc_17692_n10277;
  wire _abc_17692_n10278;
  wire _abc_17692_n10279;
  wire _abc_17692_n10280;
  wire _abc_17692_n10281;
  wire _abc_17692_n10282;
  wire _abc_17692_n10283;
  wire _abc_17692_n10284;
  wire _abc_17692_n10285;
  wire _abc_17692_n10286;
  wire _abc_17692_n10287;
  wire _abc_17692_n10288;
  wire _abc_17692_n10289;
  wire _abc_17692_n1028_1;
  wire _abc_17692_n1029;
  wire _abc_17692_n10290;
  wire _abc_17692_n10291;
  wire _abc_17692_n10292;
  wire _abc_17692_n10293;
  wire _abc_17692_n10294;
  wire _abc_17692_n10295;
  wire _abc_17692_n10296;
  wire _abc_17692_n10297;
  wire _abc_17692_n10298;
  wire _abc_17692_n10299;
  wire _abc_17692_n1030;
  wire _abc_17692_n10300;
  wire _abc_17692_n10301;
  wire _abc_17692_n10302;
  wire _abc_17692_n10303;
  wire _abc_17692_n10304;
  wire _abc_17692_n10305;
  wire _abc_17692_n10306;
  wire _abc_17692_n10307;
  wire _abc_17692_n10308;
  wire _abc_17692_n10309;
  wire _abc_17692_n1031;
  wire _abc_17692_n10310;
  wire _abc_17692_n10311;
  wire _abc_17692_n10312;
  wire _abc_17692_n10313;
  wire _abc_17692_n10314;
  wire _abc_17692_n10315;
  wire _abc_17692_n10316;
  wire _abc_17692_n10317;
  wire _abc_17692_n10318;
  wire _abc_17692_n10319;
  wire _abc_17692_n1032;
  wire _abc_17692_n10320;
  wire _abc_17692_n10321;
  wire _abc_17692_n10322;
  wire _abc_17692_n10323;
  wire _abc_17692_n10324;
  wire _abc_17692_n10325;
  wire _abc_17692_n10326;
  wire _abc_17692_n10327;
  wire _abc_17692_n10328;
  wire _abc_17692_n10329;
  wire _abc_17692_n1033;
  wire _abc_17692_n10330;
  wire _abc_17692_n10331;
  wire _abc_17692_n10332;
  wire _abc_17692_n10333;
  wire _abc_17692_n10334;
  wire _abc_17692_n10335;
  wire _abc_17692_n10336;
  wire _abc_17692_n10337;
  wire _abc_17692_n10338;
  wire _abc_17692_n10339;
  wire _abc_17692_n1034;
  wire _abc_17692_n10340;
  wire _abc_17692_n10341;
  wire _abc_17692_n10342;
  wire _abc_17692_n10344;
  wire _abc_17692_n10345;
  wire _abc_17692_n10346;
  wire _abc_17692_n10347;
  wire _abc_17692_n10348;
  wire _abc_17692_n10349;
  wire _abc_17692_n10350;
  wire _abc_17692_n10351;
  wire _abc_17692_n10352;
  wire _abc_17692_n10353;
  wire _abc_17692_n10354;
  wire _abc_17692_n10355;
  wire _abc_17692_n10356;
  wire _abc_17692_n10357;
  wire _abc_17692_n10358;
  wire _abc_17692_n10359;
  wire _abc_17692_n1035_1;
  wire _abc_17692_n1036;
  wire _abc_17692_n10360;
  wire _abc_17692_n10361;
  wire _abc_17692_n10362;
  wire _abc_17692_n10363;
  wire _abc_17692_n10364;
  wire _abc_17692_n10365;
  wire _abc_17692_n10366;
  wire _abc_17692_n10367;
  wire _abc_17692_n10368;
  wire _abc_17692_n10369;
  wire _abc_17692_n1037;
  wire _abc_17692_n10370;
  wire _abc_17692_n10371;
  wire _abc_17692_n10372;
  wire _abc_17692_n10373;
  wire _abc_17692_n10374;
  wire _abc_17692_n10375;
  wire _abc_17692_n10376;
  wire _abc_17692_n10377;
  wire _abc_17692_n10378;
  wire _abc_17692_n10379;
  wire _abc_17692_n1038;
  wire _abc_17692_n10380;
  wire _abc_17692_n10381;
  wire _abc_17692_n10382;
  wire _abc_17692_n10383;
  wire _abc_17692_n10384;
  wire _abc_17692_n10385;
  wire _abc_17692_n10386;
  wire _abc_17692_n10387;
  wire _abc_17692_n10388;
  wire _abc_17692_n10389;
  wire _abc_17692_n1039;
  wire _abc_17692_n10390;
  wire _abc_17692_n10391;
  wire _abc_17692_n10392;
  wire _abc_17692_n10393;
  wire _abc_17692_n10394;
  wire _abc_17692_n10395;
  wire _abc_17692_n10396;
  wire _abc_17692_n10397;
  wire _abc_17692_n10398;
  wire _abc_17692_n10399;
  wire _abc_17692_n1040;
  wire _abc_17692_n10400;
  wire _abc_17692_n10401;
  wire _abc_17692_n10402;
  wire _abc_17692_n10403;
  wire _abc_17692_n10404;
  wire _abc_17692_n10405;
  wire _abc_17692_n10406;
  wire _abc_17692_n10407;
  wire _abc_17692_n10408;
  wire _abc_17692_n10409;
  wire _abc_17692_n1041;
  wire _abc_17692_n10410;
  wire _abc_17692_n10411;
  wire _abc_17692_n10412;
  wire _abc_17692_n10413;
  wire _abc_17692_n10414;
  wire _abc_17692_n10415;
  wire _abc_17692_n10416;
  wire _abc_17692_n10417;
  wire _abc_17692_n10418;
  wire _abc_17692_n10419;
  wire _abc_17692_n1042;
  wire _abc_17692_n10420;
  wire _abc_17692_n10421;
  wire _abc_17692_n10422;
  wire _abc_17692_n10423;
  wire _abc_17692_n10424;
  wire _abc_17692_n10425;
  wire _abc_17692_n10426;
  wire _abc_17692_n10427;
  wire _abc_17692_n10428;
  wire _abc_17692_n10429;
  wire _abc_17692_n1043;
  wire _abc_17692_n10430;
  wire _abc_17692_n10431;
  wire _abc_17692_n10432;
  wire _abc_17692_n10433;
  wire _abc_17692_n10434;
  wire _abc_17692_n10435;
  wire _abc_17692_n10436;
  wire _abc_17692_n10437;
  wire _abc_17692_n10438;
  wire _abc_17692_n10439;
  wire _abc_17692_n1044;
  wire _abc_17692_n10440;
  wire _abc_17692_n10441;
  wire _abc_17692_n10442;
  wire _abc_17692_n10443;
  wire _abc_17692_n10444;
  wire _abc_17692_n10445;
  wire _abc_17692_n10446;
  wire _abc_17692_n10447;
  wire _abc_17692_n10448;
  wire _abc_17692_n10449;
  wire _abc_17692_n1045;
  wire _abc_17692_n10450;
  wire _abc_17692_n10451;
  wire _abc_17692_n10452;
  wire _abc_17692_n10453;
  wire _abc_17692_n10454;
  wire _abc_17692_n10455;
  wire _abc_17692_n10456;
  wire _abc_17692_n10457;
  wire _abc_17692_n10458;
  wire _abc_17692_n10459;
  wire _abc_17692_n10460;
  wire _abc_17692_n10461;
  wire _abc_17692_n10462;
  wire _abc_17692_n10463;
  wire _abc_17692_n10464;
  wire _abc_17692_n10465;
  wire _abc_17692_n10466;
  wire _abc_17692_n10467;
  wire _abc_17692_n10468;
  wire _abc_17692_n10469;
  wire _abc_17692_n1047;
  wire _abc_17692_n10470;
  wire _abc_17692_n10472;
  wire _abc_17692_n10473;
  wire _abc_17692_n10474;
  wire _abc_17692_n10475;
  wire _abc_17692_n10476;
  wire _abc_17692_n10477;
  wire _abc_17692_n10478;
  wire _abc_17692_n10479;
  wire _abc_17692_n1048;
  wire _abc_17692_n10480;
  wire _abc_17692_n10481;
  wire _abc_17692_n10482;
  wire _abc_17692_n10483;
  wire _abc_17692_n10484;
  wire _abc_17692_n10485;
  wire _abc_17692_n10486;
  wire _abc_17692_n10487;
  wire _abc_17692_n10488;
  wire _abc_17692_n10489;
  wire _abc_17692_n1049;
  wire _abc_17692_n10490;
  wire _abc_17692_n10491;
  wire _abc_17692_n10492;
  wire _abc_17692_n10493;
  wire _abc_17692_n10494;
  wire _abc_17692_n10495;
  wire _abc_17692_n10496;
  wire _abc_17692_n10497;
  wire _abc_17692_n10498;
  wire _abc_17692_n10499;
  wire _abc_17692_n1050;
  wire _abc_17692_n10500;
  wire _abc_17692_n10501;
  wire _abc_17692_n10502;
  wire _abc_17692_n10503;
  wire _abc_17692_n10504;
  wire _abc_17692_n10505;
  wire _abc_17692_n10506;
  wire _abc_17692_n10507;
  wire _abc_17692_n10508;
  wire _abc_17692_n10509;
  wire _abc_17692_n1051;
  wire _abc_17692_n10510;
  wire _abc_17692_n10511;
  wire _abc_17692_n10512;
  wire _abc_17692_n10513;
  wire _abc_17692_n10514;
  wire _abc_17692_n10515;
  wire _abc_17692_n10516;
  wire _abc_17692_n10517;
  wire _abc_17692_n10518;
  wire _abc_17692_n10519;
  wire _abc_17692_n1052;
  wire _abc_17692_n10520;
  wire _abc_17692_n10521;
  wire _abc_17692_n10522;
  wire _abc_17692_n10523;
  wire _abc_17692_n10524;
  wire _abc_17692_n10525;
  wire _abc_17692_n10526;
  wire _abc_17692_n10527;
  wire _abc_17692_n10528;
  wire _abc_17692_n10529;
  wire _abc_17692_n1053;
  wire _abc_17692_n10530;
  wire _abc_17692_n10531;
  wire _abc_17692_n10532;
  wire _abc_17692_n10533;
  wire _abc_17692_n10534;
  wire _abc_17692_n10535;
  wire _abc_17692_n10536;
  wire _abc_17692_n10537;
  wire _abc_17692_n10538;
  wire _abc_17692_n10539;
  wire _abc_17692_n1054;
  wire _abc_17692_n10540;
  wire _abc_17692_n10541;
  wire _abc_17692_n10542;
  wire _abc_17692_n10543;
  wire _abc_17692_n10544;
  wire _abc_17692_n10545;
  wire _abc_17692_n10546;
  wire _abc_17692_n10547;
  wire _abc_17692_n10548;
  wire _abc_17692_n10549;
  wire _abc_17692_n1055;
  wire _abc_17692_n10550;
  wire _abc_17692_n10551;
  wire _abc_17692_n10552;
  wire _abc_17692_n10553;
  wire _abc_17692_n10554;
  wire _abc_17692_n10555;
  wire _abc_17692_n10556;
  wire _abc_17692_n10557;
  wire _abc_17692_n10558;
  wire _abc_17692_n10559;
  wire _abc_17692_n1056;
  wire _abc_17692_n10560;
  wire _abc_17692_n10561;
  wire _abc_17692_n10562;
  wire _abc_17692_n10563;
  wire _abc_17692_n10564;
  wire _abc_17692_n10565;
  wire _abc_17692_n10566;
  wire _abc_17692_n10567;
  wire _abc_17692_n10568;
  wire _abc_17692_n10569;
  wire _abc_17692_n10570;
  wire _abc_17692_n10571;
  wire _abc_17692_n10572;
  wire _abc_17692_n10573;
  wire _abc_17692_n10574;
  wire _abc_17692_n10575;
  wire _abc_17692_n10576;
  wire _abc_17692_n10577;
  wire _abc_17692_n10578;
  wire _abc_17692_n10579;
  wire _abc_17692_n1057_1;
  wire _abc_17692_n1058;
  wire _abc_17692_n10580;
  wire _abc_17692_n10581;
  wire _abc_17692_n10582;
  wire _abc_17692_n10583;
  wire _abc_17692_n10584;
  wire _abc_17692_n10585;
  wire _abc_17692_n10586;
  wire _abc_17692_n10587;
  wire _abc_17692_n10588;
  wire _abc_17692_n10589;
  wire _abc_17692_n1059;
  wire _abc_17692_n10590;
  wire _abc_17692_n10591;
  wire _abc_17692_n10592;
  wire _abc_17692_n10593;
  wire _abc_17692_n10594;
  wire _abc_17692_n10595;
  wire _abc_17692_n10596;
  wire _abc_17692_n10597;
  wire _abc_17692_n10598;
  wire _abc_17692_n10599;
  wire _abc_17692_n1060;
  wire _abc_17692_n10600;
  wire _abc_17692_n10601;
  wire _abc_17692_n10602;
  wire _abc_17692_n10603;
  wire _abc_17692_n10604;
  wire _abc_17692_n10605;
  wire _abc_17692_n10606;
  wire _abc_17692_n10607;
  wire _abc_17692_n10608;
  wire _abc_17692_n10609;
  wire _abc_17692_n1061;
  wire _abc_17692_n10610;
  wire _abc_17692_n10611;
  wire _abc_17692_n10612;
  wire _abc_17692_n10613;
  wire _abc_17692_n10614;
  wire _abc_17692_n10615;
  wire _abc_17692_n10616;
  wire _abc_17692_n10617;
  wire _abc_17692_n10618;
  wire _abc_17692_n10619;
  wire _abc_17692_n1062;
  wire _abc_17692_n10620;
  wire _abc_17692_n10621;
  wire _abc_17692_n10622;
  wire _abc_17692_n10623;
  wire _abc_17692_n10624;
  wire _abc_17692_n10625;
  wire _abc_17692_n10626;
  wire _abc_17692_n10627;
  wire _abc_17692_n10628;
  wire _abc_17692_n10629;
  wire _abc_17692_n1063;
  wire _abc_17692_n10630;
  wire _abc_17692_n10631;
  wire _abc_17692_n10632;
  wire _abc_17692_n10633;
  wire _abc_17692_n10634;
  wire _abc_17692_n10635;
  wire _abc_17692_n10636;
  wire _abc_17692_n10637;
  wire _abc_17692_n10638;
  wire _abc_17692_n10639;
  wire _abc_17692_n1064;
  wire _abc_17692_n10640;
  wire _abc_17692_n10641;
  wire _abc_17692_n10642;
  wire _abc_17692_n10643;
  wire _abc_17692_n10644;
  wire _abc_17692_n10645;
  wire _abc_17692_n10646;
  wire _abc_17692_n10647;
  wire _abc_17692_n10648;
  wire _abc_17692_n10649;
  wire _abc_17692_n1065;
  wire _abc_17692_n10650;
  wire _abc_17692_n10651;
  wire _abc_17692_n10652;
  wire _abc_17692_n10653;
  wire _abc_17692_n10654;
  wire _abc_17692_n10655;
  wire _abc_17692_n10656;
  wire _abc_17692_n10657;
  wire _abc_17692_n10658;
  wire _abc_17692_n10659;
  wire _abc_17692_n1066;
  wire _abc_17692_n10660;
  wire _abc_17692_n10661;
  wire _abc_17692_n10662;
  wire _abc_17692_n10663;
  wire _abc_17692_n10664;
  wire _abc_17692_n10665;
  wire _abc_17692_n10666;
  wire _abc_17692_n10667;
  wire _abc_17692_n10669;
  wire _abc_17692_n1067;
  wire _abc_17692_n10670;
  wire _abc_17692_n10671;
  wire _abc_17692_n10672;
  wire _abc_17692_n10673;
  wire _abc_17692_n10674;
  wire _abc_17692_n10675;
  wire _abc_17692_n10676;
  wire _abc_17692_n10677;
  wire _abc_17692_n10678;
  wire _abc_17692_n10679;
  wire _abc_17692_n1068;
  wire _abc_17692_n10680;
  wire _abc_17692_n10681;
  wire _abc_17692_n10682;
  wire _abc_17692_n10683;
  wire _abc_17692_n10684;
  wire _abc_17692_n10685;
  wire _abc_17692_n10686;
  wire _abc_17692_n10687;
  wire _abc_17692_n10688;
  wire _abc_17692_n10689;
  wire _abc_17692_n10690;
  wire _abc_17692_n10691;
  wire _abc_17692_n10692;
  wire _abc_17692_n10693;
  wire _abc_17692_n10694;
  wire _abc_17692_n10695;
  wire _abc_17692_n10696;
  wire _abc_17692_n10697;
  wire _abc_17692_n10698;
  wire _abc_17692_n10699;
  wire _abc_17692_n1070;
  wire _abc_17692_n10700;
  wire _abc_17692_n10701;
  wire _abc_17692_n10702;
  wire _abc_17692_n10703;
  wire _abc_17692_n10704;
  wire _abc_17692_n10705;
  wire _abc_17692_n10706;
  wire _abc_17692_n10707;
  wire _abc_17692_n10708;
  wire _abc_17692_n10709;
  wire _abc_17692_n1071;
  wire _abc_17692_n10710;
  wire _abc_17692_n10711;
  wire _abc_17692_n10712;
  wire _abc_17692_n10713;
  wire _abc_17692_n10714;
  wire _abc_17692_n10715;
  wire _abc_17692_n10716;
  wire _abc_17692_n10717;
  wire _abc_17692_n10718;
  wire _abc_17692_n10719;
  wire _abc_17692_n1072;
  wire _abc_17692_n10720;
  wire _abc_17692_n10721;
  wire _abc_17692_n10722;
  wire _abc_17692_n10723;
  wire _abc_17692_n10724;
  wire _abc_17692_n10725;
  wire _abc_17692_n10726;
  wire _abc_17692_n10727;
  wire _abc_17692_n10728;
  wire _abc_17692_n10729;
  wire _abc_17692_n1073;
  wire _abc_17692_n10730;
  wire _abc_17692_n10731;
  wire _abc_17692_n10732;
  wire _abc_17692_n10733;
  wire _abc_17692_n10734;
  wire _abc_17692_n10735;
  wire _abc_17692_n10736;
  wire _abc_17692_n10737;
  wire _abc_17692_n10738;
  wire _abc_17692_n10739;
  wire _abc_17692_n1074;
  wire _abc_17692_n10740;
  wire _abc_17692_n10741;
  wire _abc_17692_n10742;
  wire _abc_17692_n10743;
  wire _abc_17692_n10744;
  wire _abc_17692_n10745;
  wire _abc_17692_n10746;
  wire _abc_17692_n10747;
  wire _abc_17692_n10748;
  wire _abc_17692_n10749;
  wire _abc_17692_n1075;
  wire _abc_17692_n10750;
  wire _abc_17692_n10751;
  wire _abc_17692_n10752;
  wire _abc_17692_n10753;
  wire _abc_17692_n10754;
  wire _abc_17692_n10755;
  wire _abc_17692_n10756;
  wire _abc_17692_n10757;
  wire _abc_17692_n10758;
  wire _abc_17692_n10759;
  wire _abc_17692_n1076;
  wire _abc_17692_n10760;
  wire _abc_17692_n10761;
  wire _abc_17692_n10762;
  wire _abc_17692_n10763;
  wire _abc_17692_n10764;
  wire _abc_17692_n10765;
  wire _abc_17692_n10766;
  wire _abc_17692_n10767;
  wire _abc_17692_n10768;
  wire _abc_17692_n10769;
  wire _abc_17692_n1077;
  wire _abc_17692_n10770;
  wire _abc_17692_n10771;
  wire _abc_17692_n10772;
  wire _abc_17692_n10773;
  wire _abc_17692_n10774;
  wire _abc_17692_n10775;
  wire _abc_17692_n10776;
  wire _abc_17692_n10777;
  wire _abc_17692_n10778;
  wire _abc_17692_n10779;
  wire _abc_17692_n1078;
  wire _abc_17692_n10780;
  wire _abc_17692_n10781;
  wire _abc_17692_n10782;
  wire _abc_17692_n10783;
  wire _abc_17692_n10784;
  wire _abc_17692_n10785;
  wire _abc_17692_n10786;
  wire _abc_17692_n10787;
  wire _abc_17692_n10788;
  wire _abc_17692_n10789;
  wire _abc_17692_n1079;
  wire _abc_17692_n10790;
  wire _abc_17692_n10791;
  wire _abc_17692_n10792;
  wire _abc_17692_n10793;
  wire _abc_17692_n10795;
  wire _abc_17692_n10796;
  wire _abc_17692_n10797;
  wire _abc_17692_n10798;
  wire _abc_17692_n10799;
  wire _abc_17692_n1080;
  wire _abc_17692_n10800;
  wire _abc_17692_n10801;
  wire _abc_17692_n10802;
  wire _abc_17692_n10803;
  wire _abc_17692_n10804;
  wire _abc_17692_n10805;
  wire _abc_17692_n10806;
  wire _abc_17692_n10807;
  wire _abc_17692_n10808;
  wire _abc_17692_n10809;
  wire _abc_17692_n1081;
  wire _abc_17692_n10810;
  wire _abc_17692_n10811;
  wire _abc_17692_n10812;
  wire _abc_17692_n10813;
  wire _abc_17692_n10814;
  wire _abc_17692_n10815;
  wire _abc_17692_n10816;
  wire _abc_17692_n10817;
  wire _abc_17692_n10818;
  wire _abc_17692_n10819;
  wire _abc_17692_n1082;
  wire _abc_17692_n10820;
  wire _abc_17692_n10821;
  wire _abc_17692_n10822;
  wire _abc_17692_n10823;
  wire _abc_17692_n10824;
  wire _abc_17692_n10825;
  wire _abc_17692_n10826;
  wire _abc_17692_n10827;
  wire _abc_17692_n10828;
  wire _abc_17692_n10829;
  wire _abc_17692_n1083;
  wire _abc_17692_n10830;
  wire _abc_17692_n10831;
  wire _abc_17692_n10832;
  wire _abc_17692_n10833;
  wire _abc_17692_n10834;
  wire _abc_17692_n10835;
  wire _abc_17692_n10836;
  wire _abc_17692_n10837;
  wire _abc_17692_n10838;
  wire _abc_17692_n10839;
  wire _abc_17692_n1084;
  wire _abc_17692_n10840;
  wire _abc_17692_n10841;
  wire _abc_17692_n10842;
  wire _abc_17692_n10843;
  wire _abc_17692_n10844;
  wire _abc_17692_n10845;
  wire _abc_17692_n10846;
  wire _abc_17692_n10847;
  wire _abc_17692_n10848;
  wire _abc_17692_n10849;
  wire _abc_17692_n1085;
  wire _abc_17692_n10850;
  wire _abc_17692_n10851;
  wire _abc_17692_n10852;
  wire _abc_17692_n10853;
  wire _abc_17692_n10854;
  wire _abc_17692_n10855;
  wire _abc_17692_n10856;
  wire _abc_17692_n10857;
  wire _abc_17692_n10858;
  wire _abc_17692_n10859;
  wire _abc_17692_n1086;
  wire _abc_17692_n10860;
  wire _abc_17692_n10861;
  wire _abc_17692_n10862;
  wire _abc_17692_n10863;
  wire _abc_17692_n10864;
  wire _abc_17692_n10865;
  wire _abc_17692_n10866;
  wire _abc_17692_n10867;
  wire _abc_17692_n10868;
  wire _abc_17692_n10869;
  wire _abc_17692_n1087;
  wire _abc_17692_n10870;
  wire _abc_17692_n10871;
  wire _abc_17692_n10872;
  wire _abc_17692_n10873;
  wire _abc_17692_n10874;
  wire _abc_17692_n10875;
  wire _abc_17692_n10876;
  wire _abc_17692_n10877;
  wire _abc_17692_n10878;
  wire _abc_17692_n10879;
  wire _abc_17692_n1088;
  wire _abc_17692_n10880;
  wire _abc_17692_n10881;
  wire _abc_17692_n10882;
  wire _abc_17692_n10883;
  wire _abc_17692_n10884;
  wire _abc_17692_n10885;
  wire _abc_17692_n10886;
  wire _abc_17692_n10887;
  wire _abc_17692_n10888;
  wire _abc_17692_n10889;
  wire _abc_17692_n1089;
  wire _abc_17692_n10890;
  wire _abc_17692_n10891;
  wire _abc_17692_n10892;
  wire _abc_17692_n10893;
  wire _abc_17692_n10894;
  wire _abc_17692_n10895;
  wire _abc_17692_n10896;
  wire _abc_17692_n10897;
  wire _abc_17692_n10898;
  wire _abc_17692_n10899;
  wire _abc_17692_n1090;
  wire _abc_17692_n10900;
  wire _abc_17692_n10901;
  wire _abc_17692_n10902;
  wire _abc_17692_n10903;
  wire _abc_17692_n10904;
  wire _abc_17692_n10905;
  wire _abc_17692_n10906;
  wire _abc_17692_n10907;
  wire _abc_17692_n10908;
  wire _abc_17692_n10909;
  wire _abc_17692_n1091;
  wire _abc_17692_n10910;
  wire _abc_17692_n10911;
  wire _abc_17692_n10912;
  wire _abc_17692_n10913;
  wire _abc_17692_n10914;
  wire _abc_17692_n10915;
  wire _abc_17692_n10916;
  wire _abc_17692_n10917;
  wire _abc_17692_n10918;
  wire _abc_17692_n10919;
  wire _abc_17692_n1092;
  wire _abc_17692_n10920;
  wire _abc_17692_n10921;
  wire _abc_17692_n10922;
  wire _abc_17692_n10923;
  wire _abc_17692_n10924;
  wire _abc_17692_n10925;
  wire _abc_17692_n10926;
  wire _abc_17692_n10927;
  wire _abc_17692_n10928;
  wire _abc_17692_n10929;
  wire _abc_17692_n1093;
  wire _abc_17692_n10930;
  wire _abc_17692_n10931;
  wire _abc_17692_n10932;
  wire _abc_17692_n10933;
  wire _abc_17692_n10934;
  wire _abc_17692_n10935;
  wire _abc_17692_n10936;
  wire _abc_17692_n10937;
  wire _abc_17692_n10938;
  wire _abc_17692_n10939;
  wire _abc_17692_n1094;
  wire _abc_17692_n10940;
  wire _abc_17692_n10941;
  wire _abc_17692_n10942;
  wire _abc_17692_n10943;
  wire _abc_17692_n10944;
  wire _abc_17692_n10945;
  wire _abc_17692_n10946;
  wire _abc_17692_n10947;
  wire _abc_17692_n10948;
  wire _abc_17692_n10949;
  wire _abc_17692_n10950;
  wire _abc_17692_n10951;
  wire _abc_17692_n10952;
  wire _abc_17692_n10953;
  wire _abc_17692_n10955;
  wire _abc_17692_n10956;
  wire _abc_17692_n10957;
  wire _abc_17692_n10958;
  wire _abc_17692_n10959;
  wire _abc_17692_n1096;
  wire _abc_17692_n10960;
  wire _abc_17692_n10961;
  wire _abc_17692_n10962;
  wire _abc_17692_n10963;
  wire _abc_17692_n10964;
  wire _abc_17692_n10965;
  wire _abc_17692_n10966;
  wire _abc_17692_n10967;
  wire _abc_17692_n10968;
  wire _abc_17692_n10969;
  wire _abc_17692_n1097;
  wire _abc_17692_n10970;
  wire _abc_17692_n10971;
  wire _abc_17692_n10972;
  wire _abc_17692_n10973;
  wire _abc_17692_n10974;
  wire _abc_17692_n10975;
  wire _abc_17692_n10976;
  wire _abc_17692_n10977;
  wire _abc_17692_n10978;
  wire _abc_17692_n10979;
  wire _abc_17692_n1098;
  wire _abc_17692_n10980;
  wire _abc_17692_n10981;
  wire _abc_17692_n10982;
  wire _abc_17692_n10983;
  wire _abc_17692_n10984;
  wire _abc_17692_n10985;
  wire _abc_17692_n10986;
  wire _abc_17692_n10987;
  wire _abc_17692_n10988;
  wire _abc_17692_n10989;
  wire _abc_17692_n1099;
  wire _abc_17692_n10990;
  wire _abc_17692_n10991;
  wire _abc_17692_n10992;
  wire _abc_17692_n10993;
  wire _abc_17692_n10994;
  wire _abc_17692_n10995;
  wire _abc_17692_n10996;
  wire _abc_17692_n10997;
  wire _abc_17692_n10998;
  wire _abc_17692_n10999;
  wire _abc_17692_n1100;
  wire _abc_17692_n11000;
  wire _abc_17692_n11001;
  wire _abc_17692_n11002;
  wire _abc_17692_n11003;
  wire _abc_17692_n11004;
  wire _abc_17692_n11005;
  wire _abc_17692_n11006;
  wire _abc_17692_n11007;
  wire _abc_17692_n11008;
  wire _abc_17692_n11009;
  wire _abc_17692_n1101;
  wire _abc_17692_n11010;
  wire _abc_17692_n11011;
  wire _abc_17692_n11012;
  wire _abc_17692_n11013;
  wire _abc_17692_n11014;
  wire _abc_17692_n11015;
  wire _abc_17692_n11016;
  wire _abc_17692_n11017;
  wire _abc_17692_n11018;
  wire _abc_17692_n11019;
  wire _abc_17692_n1102;
  wire _abc_17692_n11020;
  wire _abc_17692_n11021;
  wire _abc_17692_n11022;
  wire _abc_17692_n11023;
  wire _abc_17692_n11024;
  wire _abc_17692_n11025;
  wire _abc_17692_n11026;
  wire _abc_17692_n11027;
  wire _abc_17692_n11028;
  wire _abc_17692_n11029;
  wire _abc_17692_n1103;
  wire _abc_17692_n11030;
  wire _abc_17692_n11031;
  wire _abc_17692_n11032;
  wire _abc_17692_n11033;
  wire _abc_17692_n11034;
  wire _abc_17692_n11035;
  wire _abc_17692_n11036;
  wire _abc_17692_n11037;
  wire _abc_17692_n11038;
  wire _abc_17692_n11039;
  wire _abc_17692_n11040;
  wire _abc_17692_n11041;
  wire _abc_17692_n11042;
  wire _abc_17692_n11043;
  wire _abc_17692_n11044;
  wire _abc_17692_n11045;
  wire _abc_17692_n11046;
  wire _abc_17692_n11047;
  wire _abc_17692_n11048;
  wire _abc_17692_n11049;
  wire _abc_17692_n1104_1;
  wire _abc_17692_n1105;
  wire _abc_17692_n11050;
  wire _abc_17692_n11051;
  wire _abc_17692_n11052;
  wire _abc_17692_n11053;
  wire _abc_17692_n11054;
  wire _abc_17692_n11055;
  wire _abc_17692_n11056;
  wire _abc_17692_n11057;
  wire _abc_17692_n11058;
  wire _abc_17692_n11059;
  wire _abc_17692_n1106;
  wire _abc_17692_n11060;
  wire _abc_17692_n11061;
  wire _abc_17692_n11062;
  wire _abc_17692_n11063;
  wire _abc_17692_n11064;
  wire _abc_17692_n11065;
  wire _abc_17692_n11066;
  wire _abc_17692_n11067;
  wire _abc_17692_n11068;
  wire _abc_17692_n11069;
  wire _abc_17692_n11070;
  wire _abc_17692_n11071;
  wire _abc_17692_n11072;
  wire _abc_17692_n11073;
  wire _abc_17692_n11074;
  wire _abc_17692_n11075;
  wire _abc_17692_n11076;
  wire _abc_17692_n11077;
  wire _abc_17692_n11078;
  wire _abc_17692_n11079;
  wire _abc_17692_n1107_1;
  wire _abc_17692_n1108;
  wire _abc_17692_n11080;
  wire _abc_17692_n11081;
  wire _abc_17692_n11082;
  wire _abc_17692_n11083;
  wire _abc_17692_n11085;
  wire _abc_17692_n11086;
  wire _abc_17692_n11087;
  wire _abc_17692_n11088;
  wire _abc_17692_n11089;
  wire _abc_17692_n1109;
  wire _abc_17692_n11090;
  wire _abc_17692_n11091;
  wire _abc_17692_n11092;
  wire _abc_17692_n11093;
  wire _abc_17692_n11094;
  wire _abc_17692_n11095;
  wire _abc_17692_n11096;
  wire _abc_17692_n11097;
  wire _abc_17692_n11098;
  wire _abc_17692_n11099;
  wire _abc_17692_n1110;
  wire _abc_17692_n11100;
  wire _abc_17692_n11101;
  wire _abc_17692_n11102;
  wire _abc_17692_n11103;
  wire _abc_17692_n11104;
  wire _abc_17692_n11105;
  wire _abc_17692_n11106;
  wire _abc_17692_n11107;
  wire _abc_17692_n11108;
  wire _abc_17692_n11109;
  wire _abc_17692_n1111;
  wire _abc_17692_n11110;
  wire _abc_17692_n11111;
  wire _abc_17692_n11112;
  wire _abc_17692_n11113;
  wire _abc_17692_n11114;
  wire _abc_17692_n11115;
  wire _abc_17692_n11116;
  wire _abc_17692_n11117;
  wire _abc_17692_n11118;
  wire _abc_17692_n11119;
  wire _abc_17692_n1112;
  wire _abc_17692_n11120;
  wire _abc_17692_n11121;
  wire _abc_17692_n11122;
  wire _abc_17692_n11123;
  wire _abc_17692_n11124;
  wire _abc_17692_n11125;
  wire _abc_17692_n11126;
  wire _abc_17692_n11127;
  wire _abc_17692_n11128;
  wire _abc_17692_n11129;
  wire _abc_17692_n1113;
  wire _abc_17692_n11130;
  wire _abc_17692_n11131;
  wire _abc_17692_n11132;
  wire _abc_17692_n11133;
  wire _abc_17692_n11134;
  wire _abc_17692_n11135;
  wire _abc_17692_n11136;
  wire _abc_17692_n11137;
  wire _abc_17692_n11138;
  wire _abc_17692_n11139;
  wire _abc_17692_n1114;
  wire _abc_17692_n11140;
  wire _abc_17692_n11141;
  wire _abc_17692_n11142;
  wire _abc_17692_n11143;
  wire _abc_17692_n11144;
  wire _abc_17692_n11145;
  wire _abc_17692_n11146;
  wire _abc_17692_n11147;
  wire _abc_17692_n11148;
  wire _abc_17692_n11149;
  wire _abc_17692_n11150;
  wire _abc_17692_n11151;
  wire _abc_17692_n11152;
  wire _abc_17692_n11153;
  wire _abc_17692_n11154;
  wire _abc_17692_n11155;
  wire _abc_17692_n11156;
  wire _abc_17692_n11157;
  wire _abc_17692_n11158;
  wire _abc_17692_n11159;
  wire _abc_17692_n1115_1;
  wire _abc_17692_n1116;
  wire _abc_17692_n11160;
  wire _abc_17692_n11161;
  wire _abc_17692_n11162;
  wire _abc_17692_n11163;
  wire _abc_17692_n11164;
  wire _abc_17692_n11165;
  wire _abc_17692_n11166;
  wire _abc_17692_n11167;
  wire _abc_17692_n11168;
  wire _abc_17692_n11169;
  wire _abc_17692_n1117;
  wire _abc_17692_n11170;
  wire _abc_17692_n11171;
  wire _abc_17692_n11172;
  wire _abc_17692_n11173;
  wire _abc_17692_n11174;
  wire _abc_17692_n11175;
  wire _abc_17692_n11176;
  wire _abc_17692_n11177;
  wire _abc_17692_n11178;
  wire _abc_17692_n11179;
  wire _abc_17692_n1118;
  wire _abc_17692_n11180;
  wire _abc_17692_n11181;
  wire _abc_17692_n11182;
  wire _abc_17692_n11183;
  wire _abc_17692_n11184;
  wire _abc_17692_n11185;
  wire _abc_17692_n11186;
  wire _abc_17692_n11187;
  wire _abc_17692_n11188;
  wire _abc_17692_n11189;
  wire _abc_17692_n1119;
  wire _abc_17692_n11190;
  wire _abc_17692_n11191;
  wire _abc_17692_n11192;
  wire _abc_17692_n11193;
  wire _abc_17692_n11194;
  wire _abc_17692_n11195;
  wire _abc_17692_n11196;
  wire _abc_17692_n11197;
  wire _abc_17692_n11198;
  wire _abc_17692_n11199;
  wire _abc_17692_n11200;
  wire _abc_17692_n11201;
  wire _abc_17692_n11202;
  wire _abc_17692_n11203;
  wire _abc_17692_n11204;
  wire _abc_17692_n11205;
  wire _abc_17692_n11206;
  wire _abc_17692_n11207;
  wire _abc_17692_n11208;
  wire _abc_17692_n11209;
  wire _abc_17692_n1121;
  wire _abc_17692_n11210;
  wire _abc_17692_n11211;
  wire _abc_17692_n11212;
  wire _abc_17692_n11213;
  wire _abc_17692_n11214;
  wire _abc_17692_n11215;
  wire _abc_17692_n11216;
  wire _abc_17692_n11217;
  wire _abc_17692_n11218;
  wire _abc_17692_n11219;
  wire _abc_17692_n1122;
  wire _abc_17692_n11220;
  wire _abc_17692_n11221;
  wire _abc_17692_n11222;
  wire _abc_17692_n11223;
  wire _abc_17692_n11224;
  wire _abc_17692_n11225;
  wire _abc_17692_n11226;
  wire _abc_17692_n11227;
  wire _abc_17692_n11228;
  wire _abc_17692_n11229;
  wire _abc_17692_n1123;
  wire _abc_17692_n11230;
  wire _abc_17692_n11231;
  wire _abc_17692_n11232;
  wire _abc_17692_n11233;
  wire _abc_17692_n11234;
  wire _abc_17692_n11235;
  wire _abc_17692_n11236;
  wire _abc_17692_n11237;
  wire _abc_17692_n11238;
  wire _abc_17692_n11239;
  wire _abc_17692_n1124;
  wire _abc_17692_n11240;
  wire _abc_17692_n11241;
  wire _abc_17692_n11242;
  wire _abc_17692_n11243;
  wire _abc_17692_n11244;
  wire _abc_17692_n11245;
  wire _abc_17692_n11246;
  wire _abc_17692_n11247;
  wire _abc_17692_n11248;
  wire _abc_17692_n11249;
  wire _abc_17692_n1125;
  wire _abc_17692_n11250;
  wire _abc_17692_n11251;
  wire _abc_17692_n11252;
  wire _abc_17692_n11253;
  wire _abc_17692_n11254;
  wire _abc_17692_n11255;
  wire _abc_17692_n11256;
  wire _abc_17692_n11257;
  wire _abc_17692_n11258;
  wire _abc_17692_n11259;
  wire _abc_17692_n1126;
  wire _abc_17692_n11260;
  wire _abc_17692_n11261;
  wire _abc_17692_n11262;
  wire _abc_17692_n11263;
  wire _abc_17692_n11264;
  wire _abc_17692_n11265;
  wire _abc_17692_n11266;
  wire _abc_17692_n11267;
  wire _abc_17692_n11268;
  wire _abc_17692_n11269;
  wire _abc_17692_n11270;
  wire _abc_17692_n11271;
  wire _abc_17692_n11272;
  wire _abc_17692_n11273;
  wire _abc_17692_n11274;
  wire _abc_17692_n11275;
  wire _abc_17692_n11276;
  wire _abc_17692_n11277;
  wire _abc_17692_n11278;
  wire _abc_17692_n11279;
  wire _abc_17692_n1127_1;
  wire _abc_17692_n1128;
  wire _abc_17692_n11280;
  wire _abc_17692_n11281;
  wire _abc_17692_n11282;
  wire _abc_17692_n11283;
  wire _abc_17692_n11284;
  wire _abc_17692_n11285;
  wire _abc_17692_n11286;
  wire _abc_17692_n11287;
  wire _abc_17692_n11288;
  wire _abc_17692_n11289;
  wire _abc_17692_n1129;
  wire _abc_17692_n11290;
  wire _abc_17692_n11291;
  wire _abc_17692_n11293;
  wire _abc_17692_n11294;
  wire _abc_17692_n11295;
  wire _abc_17692_n11296;
  wire _abc_17692_n11297;
  wire _abc_17692_n11298;
  wire _abc_17692_n11299;
  wire _abc_17692_n1130;
  wire _abc_17692_n11300;
  wire _abc_17692_n11301;
  wire _abc_17692_n11302;
  wire _abc_17692_n11303;
  wire _abc_17692_n11304;
  wire _abc_17692_n11305;
  wire _abc_17692_n11306;
  wire _abc_17692_n11307;
  wire _abc_17692_n11308;
  wire _abc_17692_n11309;
  wire _abc_17692_n1131;
  wire _abc_17692_n11310;
  wire _abc_17692_n11311;
  wire _abc_17692_n11312;
  wire _abc_17692_n11313;
  wire _abc_17692_n11314;
  wire _abc_17692_n11315;
  wire _abc_17692_n11316;
  wire _abc_17692_n11317;
  wire _abc_17692_n11318;
  wire _abc_17692_n11319;
  wire _abc_17692_n1132;
  wire _abc_17692_n11320;
  wire _abc_17692_n11321;
  wire _abc_17692_n11322;
  wire _abc_17692_n11323;
  wire _abc_17692_n11324;
  wire _abc_17692_n11325;
  wire _abc_17692_n11326;
  wire _abc_17692_n11327;
  wire _abc_17692_n11328;
  wire _abc_17692_n11329;
  wire _abc_17692_n1133;
  wire _abc_17692_n11330;
  wire _abc_17692_n11331;
  wire _abc_17692_n11332;
  wire _abc_17692_n11333;
  wire _abc_17692_n11334;
  wire _abc_17692_n11335;
  wire _abc_17692_n11336;
  wire _abc_17692_n11337;
  wire _abc_17692_n11338;
  wire _abc_17692_n11339;
  wire _abc_17692_n1134;
  wire _abc_17692_n11340;
  wire _abc_17692_n11341;
  wire _abc_17692_n11342;
  wire _abc_17692_n11343;
  wire _abc_17692_n11344;
  wire _abc_17692_n11345;
  wire _abc_17692_n11346;
  wire _abc_17692_n11347;
  wire _abc_17692_n11348;
  wire _abc_17692_n11349;
  wire _abc_17692_n1135;
  wire _abc_17692_n11350;
  wire _abc_17692_n11351;
  wire _abc_17692_n11352;
  wire _abc_17692_n11353;
  wire _abc_17692_n11354;
  wire _abc_17692_n11355;
  wire _abc_17692_n11356;
  wire _abc_17692_n11357;
  wire _abc_17692_n11358;
  wire _abc_17692_n11359;
  wire _abc_17692_n1136;
  wire _abc_17692_n11360;
  wire _abc_17692_n11361;
  wire _abc_17692_n11362;
  wire _abc_17692_n11363;
  wire _abc_17692_n11364;
  wire _abc_17692_n11365;
  wire _abc_17692_n11366;
  wire _abc_17692_n11367;
  wire _abc_17692_n11368;
  wire _abc_17692_n11369;
  wire _abc_17692_n1137;
  wire _abc_17692_n11370;
  wire _abc_17692_n11371;
  wire _abc_17692_n11372;
  wire _abc_17692_n11373;
  wire _abc_17692_n11374;
  wire _abc_17692_n11375;
  wire _abc_17692_n11376;
  wire _abc_17692_n11377;
  wire _abc_17692_n11378;
  wire _abc_17692_n11379;
  wire _abc_17692_n11380;
  wire _abc_17692_n11381;
  wire _abc_17692_n11382;
  wire _abc_17692_n11383;
  wire _abc_17692_n11384;
  wire _abc_17692_n11385;
  wire _abc_17692_n11386;
  wire _abc_17692_n11387;
  wire _abc_17692_n11388;
  wire _abc_17692_n11389;
  wire _abc_17692_n1138_1;
  wire _abc_17692_n1139;
  wire _abc_17692_n11390;
  wire _abc_17692_n11391;
  wire _abc_17692_n11392;
  wire _abc_17692_n11393;
  wire _abc_17692_n11394;
  wire _abc_17692_n11395;
  wire _abc_17692_n11396;
  wire _abc_17692_n11397;
  wire _abc_17692_n11398;
  wire _abc_17692_n11399;
  wire _abc_17692_n1140;
  wire _abc_17692_n11400;
  wire _abc_17692_n11401;
  wire _abc_17692_n11402;
  wire _abc_17692_n11403;
  wire _abc_17692_n11404;
  wire _abc_17692_n11405;
  wire _abc_17692_n11406;
  wire _abc_17692_n11407;
  wire _abc_17692_n11408;
  wire _abc_17692_n11409;
  wire _abc_17692_n1141;
  wire _abc_17692_n11410;
  wire _abc_17692_n11411;
  wire _abc_17692_n11412;
  wire _abc_17692_n11413;
  wire _abc_17692_n11414;
  wire _abc_17692_n11416;
  wire _abc_17692_n11417;
  wire _abc_17692_n11418;
  wire _abc_17692_n11419;
  wire _abc_17692_n1142;
  wire _abc_17692_n11420;
  wire _abc_17692_n11421;
  wire _abc_17692_n11422;
  wire _abc_17692_n11423;
  wire _abc_17692_n11424;
  wire _abc_17692_n11425;
  wire _abc_17692_n11426;
  wire _abc_17692_n11427;
  wire _abc_17692_n11428;
  wire _abc_17692_n11429;
  wire _abc_17692_n1143;
  wire _abc_17692_n11430;
  wire _abc_17692_n11431;
  wire _abc_17692_n11432;
  wire _abc_17692_n11433;
  wire _abc_17692_n11434;
  wire _abc_17692_n11435;
  wire _abc_17692_n11436;
  wire _abc_17692_n11437;
  wire _abc_17692_n11438;
  wire _abc_17692_n11439;
  wire _abc_17692_n1144;
  wire _abc_17692_n11440;
  wire _abc_17692_n11441;
  wire _abc_17692_n11442;
  wire _abc_17692_n11443;
  wire _abc_17692_n11444;
  wire _abc_17692_n11445;
  wire _abc_17692_n11446;
  wire _abc_17692_n11447;
  wire _abc_17692_n11448;
  wire _abc_17692_n11449;
  wire _abc_17692_n1145;
  wire _abc_17692_n11450;
  wire _abc_17692_n11451;
  wire _abc_17692_n11452;
  wire _abc_17692_n11453;
  wire _abc_17692_n11454;
  wire _abc_17692_n11455;
  wire _abc_17692_n11456;
  wire _abc_17692_n11457;
  wire _abc_17692_n11458;
  wire _abc_17692_n11459;
  wire _abc_17692_n1146;
  wire _abc_17692_n11460;
  wire _abc_17692_n11461;
  wire _abc_17692_n11462;
  wire _abc_17692_n11463;
  wire _abc_17692_n11464;
  wire _abc_17692_n11465;
  wire _abc_17692_n11466;
  wire _abc_17692_n11467;
  wire _abc_17692_n11468;
  wire _abc_17692_n11469;
  wire _abc_17692_n1147;
  wire _abc_17692_n11470;
  wire _abc_17692_n11471;
  wire _abc_17692_n11472;
  wire _abc_17692_n11473;
  wire _abc_17692_n11474;
  wire _abc_17692_n11475;
  wire _abc_17692_n11476;
  wire _abc_17692_n11477;
  wire _abc_17692_n11478;
  wire _abc_17692_n11479;
  wire _abc_17692_n1148;
  wire _abc_17692_n11480;
  wire _abc_17692_n11481;
  wire _abc_17692_n11482;
  wire _abc_17692_n11483;
  wire _abc_17692_n11484;
  wire _abc_17692_n11485;
  wire _abc_17692_n11486;
  wire _abc_17692_n11487;
  wire _abc_17692_n11488;
  wire _abc_17692_n11489;
  wire _abc_17692_n11490;
  wire _abc_17692_n11491;
  wire _abc_17692_n11492;
  wire _abc_17692_n11493;
  wire _abc_17692_n11494;
  wire _abc_17692_n11495;
  wire _abc_17692_n11496;
  wire _abc_17692_n11497;
  wire _abc_17692_n11498;
  wire _abc_17692_n11499;
  wire _abc_17692_n1150;
  wire _abc_17692_n11500;
  wire _abc_17692_n11501;
  wire _abc_17692_n11502;
  wire _abc_17692_n11503;
  wire _abc_17692_n11504;
  wire _abc_17692_n11505;
  wire _abc_17692_n11506;
  wire _abc_17692_n11507;
  wire _abc_17692_n11508;
  wire _abc_17692_n11509;
  wire _abc_17692_n1151;
  wire _abc_17692_n11510;
  wire _abc_17692_n11511;
  wire _abc_17692_n11512;
  wire _abc_17692_n11513;
  wire _abc_17692_n11514;
  wire _abc_17692_n11515;
  wire _abc_17692_n11516;
  wire _abc_17692_n11517;
  wire _abc_17692_n11518;
  wire _abc_17692_n11519;
  wire _abc_17692_n11520;
  wire _abc_17692_n11521;
  wire _abc_17692_n11522;
  wire _abc_17692_n11523;
  wire _abc_17692_n11524;
  wire _abc_17692_n11525;
  wire _abc_17692_n11526;
  wire _abc_17692_n11527;
  wire _abc_17692_n11528;
  wire _abc_17692_n11529;
  wire _abc_17692_n1152_1;
  wire _abc_17692_n1153;
  wire _abc_17692_n11530;
  wire _abc_17692_n11531;
  wire _abc_17692_n11532;
  wire _abc_17692_n11533;
  wire _abc_17692_n11534;
  wire _abc_17692_n11535;
  wire _abc_17692_n11536;
  wire _abc_17692_n11537;
  wire _abc_17692_n11538;
  wire _abc_17692_n11539;
  wire _abc_17692_n1154;
  wire _abc_17692_n11540;
  wire _abc_17692_n11541;
  wire _abc_17692_n11542;
  wire _abc_17692_n11543;
  wire _abc_17692_n11544;
  wire _abc_17692_n11545;
  wire _abc_17692_n11546;
  wire _abc_17692_n11547;
  wire _abc_17692_n11548;
  wire _abc_17692_n11549;
  wire _abc_17692_n1155;
  wire _abc_17692_n11550;
  wire _abc_17692_n11551;
  wire _abc_17692_n11552;
  wire _abc_17692_n11553;
  wire _abc_17692_n11554;
  wire _abc_17692_n11555;
  wire _abc_17692_n11556;
  wire _abc_17692_n11557;
  wire _abc_17692_n11558;
  wire _abc_17692_n11559;
  wire _abc_17692_n1156;
  wire _abc_17692_n11560;
  wire _abc_17692_n11561;
  wire _abc_17692_n11562;
  wire _abc_17692_n11563;
  wire _abc_17692_n11564;
  wire _abc_17692_n11565;
  wire _abc_17692_n11566;
  wire _abc_17692_n11567;
  wire _abc_17692_n11568;
  wire _abc_17692_n11569;
  wire _abc_17692_n1157;
  wire _abc_17692_n11570;
  wire _abc_17692_n11571;
  wire _abc_17692_n11572;
  wire _abc_17692_n11573;
  wire _abc_17692_n11574;
  wire _abc_17692_n11576;
  wire _abc_17692_n11577;
  wire _abc_17692_n11578;
  wire _abc_17692_n11579;
  wire _abc_17692_n1158;
  wire _abc_17692_n11580;
  wire _abc_17692_n11581;
  wire _abc_17692_n11582;
  wire _abc_17692_n11583;
  wire _abc_17692_n11584;
  wire _abc_17692_n11585;
  wire _abc_17692_n11586;
  wire _abc_17692_n11587;
  wire _abc_17692_n11588;
  wire _abc_17692_n11589;
  wire _abc_17692_n1159;
  wire _abc_17692_n11590;
  wire _abc_17692_n11591;
  wire _abc_17692_n11592;
  wire _abc_17692_n11593;
  wire _abc_17692_n11594;
  wire _abc_17692_n11595;
  wire _abc_17692_n11596;
  wire _abc_17692_n11597;
  wire _abc_17692_n11598;
  wire _abc_17692_n11599;
  wire _abc_17692_n1160;
  wire _abc_17692_n11600;
  wire _abc_17692_n11601;
  wire _abc_17692_n11602;
  wire _abc_17692_n11603;
  wire _abc_17692_n11604;
  wire _abc_17692_n11605;
  wire _abc_17692_n11606;
  wire _abc_17692_n11607;
  wire _abc_17692_n11608;
  wire _abc_17692_n11609;
  wire _abc_17692_n1161;
  wire _abc_17692_n11610;
  wire _abc_17692_n11611;
  wire _abc_17692_n11612;
  wire _abc_17692_n11613;
  wire _abc_17692_n11614;
  wire _abc_17692_n11615;
  wire _abc_17692_n11616;
  wire _abc_17692_n11617;
  wire _abc_17692_n11618;
  wire _abc_17692_n11619;
  wire _abc_17692_n1162;
  wire _abc_17692_n11620;
  wire _abc_17692_n11621;
  wire _abc_17692_n11622;
  wire _abc_17692_n11623;
  wire _abc_17692_n11624;
  wire _abc_17692_n11625;
  wire _abc_17692_n11626;
  wire _abc_17692_n11627;
  wire _abc_17692_n11628;
  wire _abc_17692_n11629;
  wire _abc_17692_n1163;
  wire _abc_17692_n11630;
  wire _abc_17692_n11631;
  wire _abc_17692_n11632;
  wire _abc_17692_n11633;
  wire _abc_17692_n11634;
  wire _abc_17692_n11635;
  wire _abc_17692_n11636;
  wire _abc_17692_n11637;
  wire _abc_17692_n11638;
  wire _abc_17692_n11639;
  wire _abc_17692_n1164;
  wire _abc_17692_n11640;
  wire _abc_17692_n11641;
  wire _abc_17692_n11642;
  wire _abc_17692_n11643;
  wire _abc_17692_n11644;
  wire _abc_17692_n11645;
  wire _abc_17692_n11646;
  wire _abc_17692_n11647;
  wire _abc_17692_n11648;
  wire _abc_17692_n11649;
  wire _abc_17692_n1165;
  wire _abc_17692_n11650;
  wire _abc_17692_n11651;
  wire _abc_17692_n11652;
  wire _abc_17692_n11653;
  wire _abc_17692_n11654;
  wire _abc_17692_n11655;
  wire _abc_17692_n11656;
  wire _abc_17692_n11657;
  wire _abc_17692_n11658;
  wire _abc_17692_n11659;
  wire _abc_17692_n1166;
  wire _abc_17692_n11660;
  wire _abc_17692_n11661;
  wire _abc_17692_n11662;
  wire _abc_17692_n11663;
  wire _abc_17692_n11664;
  wire _abc_17692_n11665;
  wire _abc_17692_n11666;
  wire _abc_17692_n11667;
  wire _abc_17692_n11668;
  wire _abc_17692_n11669;
  wire _abc_17692_n1167;
  wire _abc_17692_n11670;
  wire _abc_17692_n11671;
  wire _abc_17692_n11672;
  wire _abc_17692_n11673;
  wire _abc_17692_n11674;
  wire _abc_17692_n11675;
  wire _abc_17692_n11676;
  wire _abc_17692_n11677;
  wire _abc_17692_n11678;
  wire _abc_17692_n11679;
  wire _abc_17692_n1168;
  wire _abc_17692_n11680;
  wire _abc_17692_n11681;
  wire _abc_17692_n11682;
  wire _abc_17692_n11683;
  wire _abc_17692_n11684;
  wire _abc_17692_n11685;
  wire _abc_17692_n11686;
  wire _abc_17692_n11687;
  wire _abc_17692_n11688;
  wire _abc_17692_n11689;
  wire _abc_17692_n1169;
  wire _abc_17692_n11690;
  wire _abc_17692_n11691;
  wire _abc_17692_n11692;
  wire _abc_17692_n11693;
  wire _abc_17692_n11694;
  wire _abc_17692_n11695;
  wire _abc_17692_n11696;
  wire _abc_17692_n11697;
  wire _abc_17692_n11698;
  wire _abc_17692_n11699;
  wire _abc_17692_n1170;
  wire _abc_17692_n11700;
  wire _abc_17692_n11701;
  wire _abc_17692_n11702;
  wire _abc_17692_n11703;
  wire _abc_17692_n11704;
  wire _abc_17692_n11705;
  wire _abc_17692_n11706;
  wire _abc_17692_n11707;
  wire _abc_17692_n11708;
  wire _abc_17692_n1171;
  wire _abc_17692_n11710;
  wire _abc_17692_n11711;
  wire _abc_17692_n11712;
  wire _abc_17692_n11713;
  wire _abc_17692_n11714;
  wire _abc_17692_n11715;
  wire _abc_17692_n11716;
  wire _abc_17692_n11717;
  wire _abc_17692_n11718;
  wire _abc_17692_n11719;
  wire _abc_17692_n1172;
  wire _abc_17692_n11720;
  wire _abc_17692_n11721;
  wire _abc_17692_n11722;
  wire _abc_17692_n11723;
  wire _abc_17692_n11724;
  wire _abc_17692_n11725;
  wire _abc_17692_n11726;
  wire _abc_17692_n11727;
  wire _abc_17692_n11728;
  wire _abc_17692_n11729;
  wire _abc_17692_n1173;
  wire _abc_17692_n11730;
  wire _abc_17692_n11731;
  wire _abc_17692_n11732;
  wire _abc_17692_n11733;
  wire _abc_17692_n11734;
  wire _abc_17692_n11735;
  wire _abc_17692_n11736;
  wire _abc_17692_n11737;
  wire _abc_17692_n11738;
  wire _abc_17692_n11739;
  wire _abc_17692_n1174;
  wire _abc_17692_n11740;
  wire _abc_17692_n11741;
  wire _abc_17692_n11742;
  wire _abc_17692_n11743;
  wire _abc_17692_n11744;
  wire _abc_17692_n11745;
  wire _abc_17692_n11746;
  wire _abc_17692_n11747;
  wire _abc_17692_n11748;
  wire _abc_17692_n11749;
  wire _abc_17692_n1175;
  wire _abc_17692_n11750;
  wire _abc_17692_n11751;
  wire _abc_17692_n11752;
  wire _abc_17692_n11753;
  wire _abc_17692_n11754;
  wire _abc_17692_n11755;
  wire _abc_17692_n11756;
  wire _abc_17692_n11757;
  wire _abc_17692_n11758;
  wire _abc_17692_n11759;
  wire _abc_17692_n1176;
  wire _abc_17692_n11760;
  wire _abc_17692_n11761;
  wire _abc_17692_n11762;
  wire _abc_17692_n11763;
  wire _abc_17692_n11764;
  wire _abc_17692_n11765;
  wire _abc_17692_n11766;
  wire _abc_17692_n11767;
  wire _abc_17692_n11768;
  wire _abc_17692_n11769;
  wire _abc_17692_n1177;
  wire _abc_17692_n11770;
  wire _abc_17692_n11771;
  wire _abc_17692_n11772;
  wire _abc_17692_n11773;
  wire _abc_17692_n11774;
  wire _abc_17692_n11775;
  wire _abc_17692_n11776;
  wire _abc_17692_n11777;
  wire _abc_17692_n11778;
  wire _abc_17692_n11779;
  wire _abc_17692_n1178;
  wire _abc_17692_n11780;
  wire _abc_17692_n11781;
  wire _abc_17692_n11782;
  wire _abc_17692_n11783;
  wire _abc_17692_n11784;
  wire _abc_17692_n11785;
  wire _abc_17692_n11786;
  wire _abc_17692_n11787;
  wire _abc_17692_n11788;
  wire _abc_17692_n11789;
  wire _abc_17692_n11790;
  wire _abc_17692_n11791;
  wire _abc_17692_n11792;
  wire _abc_17692_n11793;
  wire _abc_17692_n11794;
  wire _abc_17692_n11795;
  wire _abc_17692_n11796;
  wire _abc_17692_n11797;
  wire _abc_17692_n11798;
  wire _abc_17692_n11799;
  wire _abc_17692_n1180;
  wire _abc_17692_n11800;
  wire _abc_17692_n11801;
  wire _abc_17692_n11802;
  wire _abc_17692_n11803;
  wire _abc_17692_n11804;
  wire _abc_17692_n11805;
  wire _abc_17692_n11806;
  wire _abc_17692_n11807;
  wire _abc_17692_n11808;
  wire _abc_17692_n11809;
  wire _abc_17692_n1181;
  wire _abc_17692_n11810;
  wire _abc_17692_n11811;
  wire _abc_17692_n11812;
  wire _abc_17692_n11813;
  wire _abc_17692_n11814;
  wire _abc_17692_n11815;
  wire _abc_17692_n11816;
  wire _abc_17692_n11817;
  wire _abc_17692_n11818;
  wire _abc_17692_n11819;
  wire _abc_17692_n1182;
  wire _abc_17692_n11820;
  wire _abc_17692_n11821;
  wire _abc_17692_n11822;
  wire _abc_17692_n11823;
  wire _abc_17692_n11824;
  wire _abc_17692_n11825;
  wire _abc_17692_n11826;
  wire _abc_17692_n11827;
  wire _abc_17692_n11828;
  wire _abc_17692_n11829;
  wire _abc_17692_n1183;
  wire _abc_17692_n11830;
  wire _abc_17692_n11831;
  wire _abc_17692_n11832;
  wire _abc_17692_n11833;
  wire _abc_17692_n11834;
  wire _abc_17692_n11835;
  wire _abc_17692_n11836;
  wire _abc_17692_n11837;
  wire _abc_17692_n11838;
  wire _abc_17692_n11839;
  wire _abc_17692_n1184;
  wire _abc_17692_n11840;
  wire _abc_17692_n11841;
  wire _abc_17692_n11842;
  wire _abc_17692_n11843;
  wire _abc_17692_n11844;
  wire _abc_17692_n11845;
  wire _abc_17692_n11846;
  wire _abc_17692_n11847;
  wire _abc_17692_n11848;
  wire _abc_17692_n11849;
  wire _abc_17692_n1185;
  wire _abc_17692_n11850;
  wire _abc_17692_n11851;
  wire _abc_17692_n11852;
  wire _abc_17692_n11853;
  wire _abc_17692_n11854;
  wire _abc_17692_n11855;
  wire _abc_17692_n11856;
  wire _abc_17692_n11857;
  wire _abc_17692_n11858;
  wire _abc_17692_n11859;
  wire _abc_17692_n1186;
  wire _abc_17692_n11860;
  wire _abc_17692_n11861;
  wire _abc_17692_n11862;
  wire _abc_17692_n11863;
  wire _abc_17692_n11864;
  wire _abc_17692_n11865;
  wire _abc_17692_n11866;
  wire _abc_17692_n11867;
  wire _abc_17692_n11868;
  wire _abc_17692_n11869;
  wire _abc_17692_n1187;
  wire _abc_17692_n11870;
  wire _abc_17692_n11871;
  wire _abc_17692_n11872;
  wire _abc_17692_n11873;
  wire _abc_17692_n11874;
  wire _abc_17692_n11875;
  wire _abc_17692_n11876;
  wire _abc_17692_n11877;
  wire _abc_17692_n11878;
  wire _abc_17692_n11879;
  wire _abc_17692_n1188;
  wire _abc_17692_n11880;
  wire _abc_17692_n11881;
  wire _abc_17692_n11882;
  wire _abc_17692_n11883;
  wire _abc_17692_n11884;
  wire _abc_17692_n11885;
  wire _abc_17692_n11886;
  wire _abc_17692_n11887;
  wire _abc_17692_n11888;
  wire _abc_17692_n11889;
  wire _abc_17692_n1189;
  wire _abc_17692_n11890;
  wire _abc_17692_n11891;
  wire _abc_17692_n11892;
  wire _abc_17692_n11893;
  wire _abc_17692_n11894;
  wire _abc_17692_n11895;
  wire _abc_17692_n11896;
  wire _abc_17692_n11897;
  wire _abc_17692_n11898;
  wire _abc_17692_n11899;
  wire _abc_17692_n1190;
  wire _abc_17692_n11900;
  wire _abc_17692_n11901;
  wire _abc_17692_n11902;
  wire _abc_17692_n11903;
  wire _abc_17692_n11904;
  wire _abc_17692_n11905;
  wire _abc_17692_n11906;
  wire _abc_17692_n11907;
  wire _abc_17692_n11908;
  wire _abc_17692_n11909;
  wire _abc_17692_n1191;
  wire _abc_17692_n11910;
  wire _abc_17692_n11911;
  wire _abc_17692_n11912;
  wire _abc_17692_n11913;
  wire _abc_17692_n11914;
  wire _abc_17692_n11915;
  wire _abc_17692_n11916;
  wire _abc_17692_n11917;
  wire _abc_17692_n11918;
  wire _abc_17692_n11919;
  wire _abc_17692_n11920;
  wire _abc_17692_n11921;
  wire _abc_17692_n11922;
  wire _abc_17692_n11924;
  wire _abc_17692_n11925;
  wire _abc_17692_n11926;
  wire _abc_17692_n11927;
  wire _abc_17692_n11928;
  wire _abc_17692_n11929;
  wire _abc_17692_n1192_1;
  wire _abc_17692_n1193;
  wire _abc_17692_n11930;
  wire _abc_17692_n11931;
  wire _abc_17692_n11932;
  wire _abc_17692_n11933;
  wire _abc_17692_n11934;
  wire _abc_17692_n11935;
  wire _abc_17692_n11936;
  wire _abc_17692_n11937;
  wire _abc_17692_n11938;
  wire _abc_17692_n11939;
  wire _abc_17692_n1194;
  wire _abc_17692_n11940;
  wire _abc_17692_n11941;
  wire _abc_17692_n11942;
  wire _abc_17692_n11943;
  wire _abc_17692_n11944;
  wire _abc_17692_n11945;
  wire _abc_17692_n11946;
  wire _abc_17692_n11947;
  wire _abc_17692_n11948;
  wire _abc_17692_n11949;
  wire _abc_17692_n11950;
  wire _abc_17692_n11951;
  wire _abc_17692_n11952;
  wire _abc_17692_n11953;
  wire _abc_17692_n11954;
  wire _abc_17692_n11955;
  wire _abc_17692_n11956;
  wire _abc_17692_n11957;
  wire _abc_17692_n11958;
  wire _abc_17692_n11959;
  wire _abc_17692_n1195_1;
  wire _abc_17692_n1196;
  wire _abc_17692_n11960;
  wire _abc_17692_n11961;
  wire _abc_17692_n11962;
  wire _abc_17692_n11963;
  wire _abc_17692_n11964;
  wire _abc_17692_n11965;
  wire _abc_17692_n11966;
  wire _abc_17692_n11967;
  wire _abc_17692_n11968;
  wire _abc_17692_n11969;
  wire _abc_17692_n1197;
  wire _abc_17692_n11970;
  wire _abc_17692_n11971;
  wire _abc_17692_n11972;
  wire _abc_17692_n11973;
  wire _abc_17692_n11974;
  wire _abc_17692_n11975;
  wire _abc_17692_n11976;
  wire _abc_17692_n11977;
  wire _abc_17692_n11978;
  wire _abc_17692_n11979;
  wire _abc_17692_n1198;
  wire _abc_17692_n11980;
  wire _abc_17692_n11981;
  wire _abc_17692_n11982;
  wire _abc_17692_n11983;
  wire _abc_17692_n11984;
  wire _abc_17692_n11985;
  wire _abc_17692_n11986;
  wire _abc_17692_n11987;
  wire _abc_17692_n11988;
  wire _abc_17692_n11989;
  wire _abc_17692_n1199;
  wire _abc_17692_n11990;
  wire _abc_17692_n11991;
  wire _abc_17692_n11992;
  wire _abc_17692_n11993;
  wire _abc_17692_n11994;
  wire _abc_17692_n11995;
  wire _abc_17692_n11996;
  wire _abc_17692_n11997;
  wire _abc_17692_n11998;
  wire _abc_17692_n11999;
  wire _abc_17692_n1200;
  wire _abc_17692_n12000;
  wire _abc_17692_n12001;
  wire _abc_17692_n12002;
  wire _abc_17692_n12003;
  wire _abc_17692_n12004;
  wire _abc_17692_n12005;
  wire _abc_17692_n12006;
  wire _abc_17692_n12007;
  wire _abc_17692_n12008;
  wire _abc_17692_n12009;
  wire _abc_17692_n1201;
  wire _abc_17692_n12010;
  wire _abc_17692_n12011;
  wire _abc_17692_n12012;
  wire _abc_17692_n12013;
  wire _abc_17692_n12014;
  wire _abc_17692_n12015;
  wire _abc_17692_n12016;
  wire _abc_17692_n12017;
  wire _abc_17692_n12018;
  wire _abc_17692_n12019;
  wire _abc_17692_n1202;
  wire _abc_17692_n12020;
  wire _abc_17692_n12021;
  wire _abc_17692_n12022;
  wire _abc_17692_n12023;
  wire _abc_17692_n12024;
  wire _abc_17692_n12025;
  wire _abc_17692_n12026;
  wire _abc_17692_n12027;
  wire _abc_17692_n12028;
  wire _abc_17692_n12029;
  wire _abc_17692_n12030;
  wire _abc_17692_n12031;
  wire _abc_17692_n12032;
  wire _abc_17692_n12033;
  wire _abc_17692_n12034;
  wire _abc_17692_n12035;
  wire _abc_17692_n12036;
  wire _abc_17692_n12037;
  wire _abc_17692_n12038;
  wire _abc_17692_n12039;
  wire _abc_17692_n1204;
  wire _abc_17692_n12040;
  wire _abc_17692_n12041;
  wire _abc_17692_n12042;
  wire _abc_17692_n12043;
  wire _abc_17692_n12044;
  wire _abc_17692_n12045;
  wire _abc_17692_n12046;
  wire _abc_17692_n12047;
  wire _abc_17692_n12048;
  wire _abc_17692_n12049;
  wire _abc_17692_n1205;
  wire _abc_17692_n12050;
  wire _abc_17692_n12051;
  wire _abc_17692_n12052;
  wire _abc_17692_n12053;
  wire _abc_17692_n12055;
  wire _abc_17692_n12056;
  wire _abc_17692_n12057;
  wire _abc_17692_n12058;
  wire _abc_17692_n12059;
  wire _abc_17692_n12060;
  wire _abc_17692_n12061;
  wire _abc_17692_n12062;
  wire _abc_17692_n12063;
  wire _abc_17692_n12064;
  wire _abc_17692_n12065;
  wire _abc_17692_n12066;
  wire _abc_17692_n12067;
  wire _abc_17692_n12068;
  wire _abc_17692_n12069;
  wire _abc_17692_n1206_1;
  wire _abc_17692_n1207;
  wire _abc_17692_n12070;
  wire _abc_17692_n12071;
  wire _abc_17692_n12072;
  wire _abc_17692_n12073;
  wire _abc_17692_n12074;
  wire _abc_17692_n12075;
  wire _abc_17692_n12076;
  wire _abc_17692_n12077;
  wire _abc_17692_n12078;
  wire _abc_17692_n12079;
  wire _abc_17692_n1208;
  wire _abc_17692_n12080;
  wire _abc_17692_n12081;
  wire _abc_17692_n12082;
  wire _abc_17692_n12083;
  wire _abc_17692_n12084;
  wire _abc_17692_n12085;
  wire _abc_17692_n12086;
  wire _abc_17692_n12087;
  wire _abc_17692_n12088;
  wire _abc_17692_n12089;
  wire _abc_17692_n1209;
  wire _abc_17692_n12090;
  wire _abc_17692_n12091;
  wire _abc_17692_n12092;
  wire _abc_17692_n12093;
  wire _abc_17692_n12094;
  wire _abc_17692_n12095;
  wire _abc_17692_n12096;
  wire _abc_17692_n12097;
  wire _abc_17692_n12098;
  wire _abc_17692_n12099;
  wire _abc_17692_n1210;
  wire _abc_17692_n12100;
  wire _abc_17692_n12101;
  wire _abc_17692_n12102;
  wire _abc_17692_n12103;
  wire _abc_17692_n12104;
  wire _abc_17692_n12105;
  wire _abc_17692_n12106;
  wire _abc_17692_n12107;
  wire _abc_17692_n12108;
  wire _abc_17692_n12109;
  wire _abc_17692_n1211;
  wire _abc_17692_n12110;
  wire _abc_17692_n12111;
  wire _abc_17692_n12112;
  wire _abc_17692_n12113;
  wire _abc_17692_n12114;
  wire _abc_17692_n12115;
  wire _abc_17692_n12116;
  wire _abc_17692_n12117;
  wire _abc_17692_n12118;
  wire _abc_17692_n12119;
  wire _abc_17692_n1212;
  wire _abc_17692_n12120;
  wire _abc_17692_n12121;
  wire _abc_17692_n12122;
  wire _abc_17692_n12123;
  wire _abc_17692_n12124;
  wire _abc_17692_n12125;
  wire _abc_17692_n12126;
  wire _abc_17692_n12127;
  wire _abc_17692_n12128;
  wire _abc_17692_n12129;
  wire _abc_17692_n1213;
  wire _abc_17692_n12130;
  wire _abc_17692_n12131;
  wire _abc_17692_n12132;
  wire _abc_17692_n12133;
  wire _abc_17692_n12134;
  wire _abc_17692_n12135;
  wire _abc_17692_n12136;
  wire _abc_17692_n12137;
  wire _abc_17692_n12138;
  wire _abc_17692_n12139;
  wire _abc_17692_n1214;
  wire _abc_17692_n12140;
  wire _abc_17692_n12141;
  wire _abc_17692_n12142;
  wire _abc_17692_n12143;
  wire _abc_17692_n12144;
  wire _abc_17692_n12145;
  wire _abc_17692_n12146;
  wire _abc_17692_n12147;
  wire _abc_17692_n12148;
  wire _abc_17692_n12149;
  wire _abc_17692_n1215;
  wire _abc_17692_n12150;
  wire _abc_17692_n12151;
  wire _abc_17692_n12152;
  wire _abc_17692_n12153;
  wire _abc_17692_n12154;
  wire _abc_17692_n12155;
  wire _abc_17692_n12156;
  wire _abc_17692_n12157;
  wire _abc_17692_n12158;
  wire _abc_17692_n12159;
  wire _abc_17692_n1216;
  wire _abc_17692_n12160;
  wire _abc_17692_n12161;
  wire _abc_17692_n12162;
  wire _abc_17692_n12163;
  wire _abc_17692_n12164;
  wire _abc_17692_n12165;
  wire _abc_17692_n12166;
  wire _abc_17692_n12167;
  wire _abc_17692_n12168;
  wire _abc_17692_n12169;
  wire _abc_17692_n1217;
  wire _abc_17692_n12170;
  wire _abc_17692_n12171;
  wire _abc_17692_n12172;
  wire _abc_17692_n12173;
  wire _abc_17692_n12174;
  wire _abc_17692_n12175;
  wire _abc_17692_n12176;
  wire _abc_17692_n12177;
  wire _abc_17692_n12178;
  wire _abc_17692_n12179;
  wire _abc_17692_n1218;
  wire _abc_17692_n12180;
  wire _abc_17692_n12181;
  wire _abc_17692_n12182;
  wire _abc_17692_n12183;
  wire _abc_17692_n12184;
  wire _abc_17692_n12185;
  wire _abc_17692_n12186;
  wire _abc_17692_n12187;
  wire _abc_17692_n12188;
  wire _abc_17692_n12189;
  wire _abc_17692_n1219;
  wire _abc_17692_n12190;
  wire _abc_17692_n12191;
  wire _abc_17692_n12192;
  wire _abc_17692_n12193;
  wire _abc_17692_n12194;
  wire _abc_17692_n12195;
  wire _abc_17692_n12196;
  wire _abc_17692_n12197;
  wire _abc_17692_n12198;
  wire _abc_17692_n12199;
  wire _abc_17692_n1220;
  wire _abc_17692_n12200;
  wire _abc_17692_n12201;
  wire _abc_17692_n12202;
  wire _abc_17692_n12203;
  wire _abc_17692_n12204;
  wire _abc_17692_n12205;
  wire _abc_17692_n12206;
  wire _abc_17692_n12207;
  wire _abc_17692_n12208;
  wire _abc_17692_n12209;
  wire _abc_17692_n1221;
  wire _abc_17692_n12210;
  wire _abc_17692_n12212;
  wire _abc_17692_n12213;
  wire _abc_17692_n12214;
  wire _abc_17692_n12215;
  wire _abc_17692_n12216;
  wire _abc_17692_n12217;
  wire _abc_17692_n12218;
  wire _abc_17692_n12219;
  wire _abc_17692_n1222;
  wire _abc_17692_n12220;
  wire _abc_17692_n12221;
  wire _abc_17692_n12222;
  wire _abc_17692_n12223;
  wire _abc_17692_n12224;
  wire _abc_17692_n12225;
  wire _abc_17692_n12226;
  wire _abc_17692_n12227;
  wire _abc_17692_n12228;
  wire _abc_17692_n12229;
  wire _abc_17692_n12230;
  wire _abc_17692_n12231;
  wire _abc_17692_n12232;
  wire _abc_17692_n12233;
  wire _abc_17692_n12234;
  wire _abc_17692_n12235;
  wire _abc_17692_n12236;
  wire _abc_17692_n12237;
  wire _abc_17692_n12238;
  wire _abc_17692_n12239;
  wire _abc_17692_n1223_1;
  wire _abc_17692_n1224;
  wire _abc_17692_n12240;
  wire _abc_17692_n12241;
  wire _abc_17692_n12242;
  wire _abc_17692_n12243;
  wire _abc_17692_n12244;
  wire _abc_17692_n12245;
  wire _abc_17692_n12246;
  wire _abc_17692_n12247;
  wire _abc_17692_n12248;
  wire _abc_17692_n12249;
  wire _abc_17692_n1225;
  wire _abc_17692_n12250;
  wire _abc_17692_n12251;
  wire _abc_17692_n12252;
  wire _abc_17692_n12253;
  wire _abc_17692_n12254;
  wire _abc_17692_n12255;
  wire _abc_17692_n12256;
  wire _abc_17692_n12257;
  wire _abc_17692_n12258;
  wire _abc_17692_n12259;
  wire _abc_17692_n1226;
  wire _abc_17692_n12260;
  wire _abc_17692_n12261;
  wire _abc_17692_n12262;
  wire _abc_17692_n12263;
  wire _abc_17692_n12264;
  wire _abc_17692_n12265;
  wire _abc_17692_n12266;
  wire _abc_17692_n12267;
  wire _abc_17692_n12268;
  wire _abc_17692_n12269;
  wire _abc_17692_n1227;
  wire _abc_17692_n12270;
  wire _abc_17692_n12271;
  wire _abc_17692_n12272;
  wire _abc_17692_n12273;
  wire _abc_17692_n12274;
  wire _abc_17692_n12275;
  wire _abc_17692_n12276;
  wire _abc_17692_n12277;
  wire _abc_17692_n12278;
  wire _abc_17692_n12279;
  wire _abc_17692_n1228;
  wire _abc_17692_n12280;
  wire _abc_17692_n12281;
  wire _abc_17692_n12282;
  wire _abc_17692_n12283;
  wire _abc_17692_n12284;
  wire _abc_17692_n12285;
  wire _abc_17692_n12286;
  wire _abc_17692_n12287;
  wire _abc_17692_n12288;
  wire _abc_17692_n12289;
  wire _abc_17692_n1229;
  wire _abc_17692_n12290;
  wire _abc_17692_n12291;
  wire _abc_17692_n12292;
  wire _abc_17692_n12293;
  wire _abc_17692_n12294;
  wire _abc_17692_n12295;
  wire _abc_17692_n12296;
  wire _abc_17692_n12297;
  wire _abc_17692_n12298;
  wire _abc_17692_n12299;
  wire _abc_17692_n1230;
  wire _abc_17692_n12300;
  wire _abc_17692_n12301;
  wire _abc_17692_n12302;
  wire _abc_17692_n12303;
  wire _abc_17692_n12304;
  wire _abc_17692_n12305;
  wire _abc_17692_n12306;
  wire _abc_17692_n12307;
  wire _abc_17692_n12308;
  wire _abc_17692_n12309;
  wire _abc_17692_n1231;
  wire _abc_17692_n12310;
  wire _abc_17692_n12311;
  wire _abc_17692_n12312;
  wire _abc_17692_n12313;
  wire _abc_17692_n12314;
  wire _abc_17692_n12315;
  wire _abc_17692_n12316;
  wire _abc_17692_n12317;
  wire _abc_17692_n12318;
  wire _abc_17692_n12319;
  wire _abc_17692_n1232;
  wire _abc_17692_n12320;
  wire _abc_17692_n12321;
  wire _abc_17692_n12322;
  wire _abc_17692_n12323;
  wire _abc_17692_n12324;
  wire _abc_17692_n12325;
  wire _abc_17692_n12326;
  wire _abc_17692_n12327;
  wire _abc_17692_n12328;
  wire _abc_17692_n12329;
  wire _abc_17692_n1233;
  wire _abc_17692_n12330;
  wire _abc_17692_n12331;
  wire _abc_17692_n12332;
  wire _abc_17692_n12333;
  wire _abc_17692_n12334;
  wire _abc_17692_n12335;
  wire _abc_17692_n12336;
  wire _abc_17692_n12337;
  wire _abc_17692_n12339;
  wire _abc_17692_n1234;
  wire _abc_17692_n12340;
  wire _abc_17692_n12341;
  wire _abc_17692_n12342;
  wire _abc_17692_n12343;
  wire _abc_17692_n12344;
  wire _abc_17692_n12345;
  wire _abc_17692_n12346;
  wire _abc_17692_n12347;
  wire _abc_17692_n12348;
  wire _abc_17692_n12349;
  wire _abc_17692_n1235;
  wire _abc_17692_n12350;
  wire _abc_17692_n12351;
  wire _abc_17692_n12352;
  wire _abc_17692_n12353;
  wire _abc_17692_n12354;
  wire _abc_17692_n12355;
  wire _abc_17692_n12356;
  wire _abc_17692_n12357;
  wire _abc_17692_n12358;
  wire _abc_17692_n12359;
  wire _abc_17692_n1236;
  wire _abc_17692_n12360;
  wire _abc_17692_n12361;
  wire _abc_17692_n12362;
  wire _abc_17692_n12363;
  wire _abc_17692_n12364;
  wire _abc_17692_n12365;
  wire _abc_17692_n12366;
  wire _abc_17692_n12367;
  wire _abc_17692_n12368;
  wire _abc_17692_n12369;
  wire _abc_17692_n1237;
  wire _abc_17692_n12370;
  wire _abc_17692_n12371;
  wire _abc_17692_n12372;
  wire _abc_17692_n12373;
  wire _abc_17692_n12374;
  wire _abc_17692_n12375;
  wire _abc_17692_n12376;
  wire _abc_17692_n12377;
  wire _abc_17692_n12378;
  wire _abc_17692_n12379;
  wire _abc_17692_n1238;
  wire _abc_17692_n12380;
  wire _abc_17692_n12381;
  wire _abc_17692_n12382;
  wire _abc_17692_n12383;
  wire _abc_17692_n12384;
  wire _abc_17692_n12385;
  wire _abc_17692_n12386;
  wire _abc_17692_n12387;
  wire _abc_17692_n12388;
  wire _abc_17692_n12389;
  wire _abc_17692_n1239;
  wire _abc_17692_n12390;
  wire _abc_17692_n12391;
  wire _abc_17692_n12392;
  wire _abc_17692_n12393;
  wire _abc_17692_n12394;
  wire _abc_17692_n12395;
  wire _abc_17692_n12396;
  wire _abc_17692_n12397;
  wire _abc_17692_n12398;
  wire _abc_17692_n12399;
  wire _abc_17692_n1240;
  wire _abc_17692_n12400;
  wire _abc_17692_n12401;
  wire _abc_17692_n12402;
  wire _abc_17692_n12403;
  wire _abc_17692_n12404;
  wire _abc_17692_n12405;
  wire _abc_17692_n12406;
  wire _abc_17692_n12407;
  wire _abc_17692_n12408;
  wire _abc_17692_n12409;
  wire _abc_17692_n12410;
  wire _abc_17692_n12411;
  wire _abc_17692_n12412;
  wire _abc_17692_n12413;
  wire _abc_17692_n12414;
  wire _abc_17692_n12415;
  wire _abc_17692_n12416;
  wire _abc_17692_n12417;
  wire _abc_17692_n12418;
  wire _abc_17692_n12419;
  wire _abc_17692_n1241_1;
  wire _abc_17692_n1242;
  wire _abc_17692_n12420;
  wire _abc_17692_n12421;
  wire _abc_17692_n12422;
  wire _abc_17692_n12423;
  wire _abc_17692_n12424;
  wire _abc_17692_n12425;
  wire _abc_17692_n12426;
  wire _abc_17692_n12427;
  wire _abc_17692_n12428;
  wire _abc_17692_n12429;
  wire _abc_17692_n12430;
  wire _abc_17692_n12431;
  wire _abc_17692_n12432;
  wire _abc_17692_n12433;
  wire _abc_17692_n12434;
  wire _abc_17692_n12435;
  wire _abc_17692_n12436;
  wire _abc_17692_n12437;
  wire _abc_17692_n12438;
  wire _abc_17692_n12439;
  wire _abc_17692_n1244;
  wire _abc_17692_n12440;
  wire _abc_17692_n12441;
  wire _abc_17692_n12442;
  wire _abc_17692_n12443;
  wire _abc_17692_n12444;
  wire _abc_17692_n12445;
  wire _abc_17692_n12446;
  wire _abc_17692_n12447;
  wire _abc_17692_n12448;
  wire _abc_17692_n12449;
  wire _abc_17692_n1245;
  wire _abc_17692_n12450;
  wire _abc_17692_n12451;
  wire _abc_17692_n12452;
  wire _abc_17692_n12453;
  wire _abc_17692_n12454;
  wire _abc_17692_n12455;
  wire _abc_17692_n12456;
  wire _abc_17692_n12457;
  wire _abc_17692_n12458;
  wire _abc_17692_n12459;
  wire _abc_17692_n1246;
  wire _abc_17692_n12460;
  wire _abc_17692_n12461;
  wire _abc_17692_n12462;
  wire _abc_17692_n12463;
  wire _abc_17692_n12464;
  wire _abc_17692_n12465;
  wire _abc_17692_n12466;
  wire _abc_17692_n12467;
  wire _abc_17692_n12468;
  wire _abc_17692_n12469;
  wire _abc_17692_n1247;
  wire _abc_17692_n12470;
  wire _abc_17692_n12471;
  wire _abc_17692_n12472;
  wire _abc_17692_n12473;
  wire _abc_17692_n12474;
  wire _abc_17692_n12475;
  wire _abc_17692_n12476;
  wire _abc_17692_n12477;
  wire _abc_17692_n12478;
  wire _abc_17692_n12479;
  wire _abc_17692_n1248;
  wire _abc_17692_n12480;
  wire _abc_17692_n12481;
  wire _abc_17692_n12482;
  wire _abc_17692_n12483;
  wire _abc_17692_n12484;
  wire _abc_17692_n12485;
  wire _abc_17692_n12486;
  wire _abc_17692_n12487;
  wire _abc_17692_n12488;
  wire _abc_17692_n12489;
  wire _abc_17692_n1249;
  wire _abc_17692_n12490;
  wire _abc_17692_n12491;
  wire _abc_17692_n12492;
  wire _abc_17692_n12493;
  wire _abc_17692_n12494;
  wire _abc_17692_n12495;
  wire _abc_17692_n12496;
  wire _abc_17692_n12497;
  wire _abc_17692_n12498;
  wire _abc_17692_n12499;
  wire _abc_17692_n1250;
  wire _abc_17692_n12500;
  wire _abc_17692_n12501;
  wire _abc_17692_n12502;
  wire _abc_17692_n12503;
  wire _abc_17692_n12504;
  wire _abc_17692_n12505;
  wire _abc_17692_n12506;
  wire _abc_17692_n12507;
  wire _abc_17692_n12508;
  wire _abc_17692_n12509;
  wire _abc_17692_n1251;
  wire _abc_17692_n12510;
  wire _abc_17692_n12511;
  wire _abc_17692_n12512;
  wire _abc_17692_n12513;
  wire _abc_17692_n12514;
  wire _abc_17692_n12515;
  wire _abc_17692_n12516;
  wire _abc_17692_n12517;
  wire _abc_17692_n12518;
  wire _abc_17692_n12519;
  wire _abc_17692_n1252;
  wire _abc_17692_n12520;
  wire _abc_17692_n12522;
  wire _abc_17692_n12523;
  wire _abc_17692_n12524;
  wire _abc_17692_n12525;
  wire _abc_17692_n12526;
  wire _abc_17692_n12527;
  wire _abc_17692_n12528;
  wire _abc_17692_n12529;
  wire _abc_17692_n1253;
  wire _abc_17692_n12530;
  wire _abc_17692_n12531;
  wire _abc_17692_n12532;
  wire _abc_17692_n12533;
  wire _abc_17692_n12534;
  wire _abc_17692_n12535;
  wire _abc_17692_n12536;
  wire _abc_17692_n12537;
  wire _abc_17692_n12538;
  wire _abc_17692_n12539;
  wire _abc_17692_n1254;
  wire _abc_17692_n12540;
  wire _abc_17692_n12541;
  wire _abc_17692_n12542;
  wire _abc_17692_n12543;
  wire _abc_17692_n12544;
  wire _abc_17692_n12545;
  wire _abc_17692_n12546;
  wire _abc_17692_n12547;
  wire _abc_17692_n12548;
  wire _abc_17692_n12549;
  wire _abc_17692_n1255;
  wire _abc_17692_n12550;
  wire _abc_17692_n12551;
  wire _abc_17692_n12552;
  wire _abc_17692_n12553;
  wire _abc_17692_n12554;
  wire _abc_17692_n12555;
  wire _abc_17692_n12556;
  wire _abc_17692_n12557;
  wire _abc_17692_n12558;
  wire _abc_17692_n12559;
  wire _abc_17692_n1256;
  wire _abc_17692_n12560;
  wire _abc_17692_n12561;
  wire _abc_17692_n12562;
  wire _abc_17692_n12563;
  wire _abc_17692_n12564;
  wire _abc_17692_n12565;
  wire _abc_17692_n12566;
  wire _abc_17692_n12567;
  wire _abc_17692_n12568;
  wire _abc_17692_n12569;
  wire _abc_17692_n1257;
  wire _abc_17692_n12570;
  wire _abc_17692_n12571;
  wire _abc_17692_n12572;
  wire _abc_17692_n12573;
  wire _abc_17692_n12574;
  wire _abc_17692_n12575;
  wire _abc_17692_n12576;
  wire _abc_17692_n12577;
  wire _abc_17692_n12578;
  wire _abc_17692_n12579;
  wire _abc_17692_n12580;
  wire _abc_17692_n12581;
  wire _abc_17692_n12582;
  wire _abc_17692_n12583;
  wire _abc_17692_n12584;
  wire _abc_17692_n12585;
  wire _abc_17692_n12586;
  wire _abc_17692_n12587;
  wire _abc_17692_n12588;
  wire _abc_17692_n12589;
  wire _abc_17692_n1258_1;
  wire _abc_17692_n1259;
  wire _abc_17692_n12590;
  wire _abc_17692_n12591;
  wire _abc_17692_n12592;
  wire _abc_17692_n12593;
  wire _abc_17692_n12594;
  wire _abc_17692_n12595;
  wire _abc_17692_n12596;
  wire _abc_17692_n12597;
  wire _abc_17692_n12598;
  wire _abc_17692_n12599;
  wire _abc_17692_n1260;
  wire _abc_17692_n12600;
  wire _abc_17692_n12601;
  wire _abc_17692_n12602;
  wire _abc_17692_n12603;
  wire _abc_17692_n12604;
  wire _abc_17692_n12605;
  wire _abc_17692_n12606;
  wire _abc_17692_n12607;
  wire _abc_17692_n12608;
  wire _abc_17692_n12609;
  wire _abc_17692_n1261;
  wire _abc_17692_n12610;
  wire _abc_17692_n12611;
  wire _abc_17692_n12612;
  wire _abc_17692_n12613;
  wire _abc_17692_n12614;
  wire _abc_17692_n12615;
  wire _abc_17692_n12616;
  wire _abc_17692_n12617;
  wire _abc_17692_n12618;
  wire _abc_17692_n12619;
  wire _abc_17692_n1262;
  wire _abc_17692_n12620;
  wire _abc_17692_n12621;
  wire _abc_17692_n12622;
  wire _abc_17692_n12623;
  wire _abc_17692_n12624;
  wire _abc_17692_n12625;
  wire _abc_17692_n12626;
  wire _abc_17692_n12627;
  wire _abc_17692_n12628;
  wire _abc_17692_n12629;
  wire _abc_17692_n1263;
  wire _abc_17692_n12630;
  wire _abc_17692_n12631;
  wire _abc_17692_n12632;
  wire _abc_17692_n12633;
  wire _abc_17692_n12634;
  wire _abc_17692_n12635;
  wire _abc_17692_n12636;
  wire _abc_17692_n12637;
  wire _abc_17692_n12638;
  wire _abc_17692_n12639;
  wire _abc_17692_n1264;
  wire _abc_17692_n12640;
  wire _abc_17692_n12641;
  wire _abc_17692_n12642;
  wire _abc_17692_n12643;
  wire _abc_17692_n12644;
  wire _abc_17692_n12645;
  wire _abc_17692_n12647;
  wire _abc_17692_n12648;
  wire _abc_17692_n12649;
  wire _abc_17692_n1265;
  wire _abc_17692_n12650;
  wire _abc_17692_n12651;
  wire _abc_17692_n12652;
  wire _abc_17692_n12653;
  wire _abc_17692_n12654;
  wire _abc_17692_n12655;
  wire _abc_17692_n12656;
  wire _abc_17692_n12657;
  wire _abc_17692_n12658;
  wire _abc_17692_n12659;
  wire _abc_17692_n1266;
  wire _abc_17692_n12660;
  wire _abc_17692_n12661;
  wire _abc_17692_n12662;
  wire _abc_17692_n12663;
  wire _abc_17692_n12664;
  wire _abc_17692_n12665;
  wire _abc_17692_n12666;
  wire _abc_17692_n12667;
  wire _abc_17692_n12668;
  wire _abc_17692_n12669;
  wire _abc_17692_n1267;
  wire _abc_17692_n12670;
  wire _abc_17692_n12671;
  wire _abc_17692_n12672;
  wire _abc_17692_n12673;
  wire _abc_17692_n12674;
  wire _abc_17692_n12675;
  wire _abc_17692_n12676;
  wire _abc_17692_n12677;
  wire _abc_17692_n12678;
  wire _abc_17692_n12679;
  wire _abc_17692_n1268;
  wire _abc_17692_n12680;
  wire _abc_17692_n12681;
  wire _abc_17692_n12682;
  wire _abc_17692_n12683;
  wire _abc_17692_n12684;
  wire _abc_17692_n12685;
  wire _abc_17692_n12686;
  wire _abc_17692_n12687;
  wire _abc_17692_n12688;
  wire _abc_17692_n12689;
  wire _abc_17692_n1269;
  wire _abc_17692_n12690;
  wire _abc_17692_n12691;
  wire _abc_17692_n12692;
  wire _abc_17692_n12693;
  wire _abc_17692_n12694;
  wire _abc_17692_n12695;
  wire _abc_17692_n12696;
  wire _abc_17692_n12697;
  wire _abc_17692_n12698;
  wire _abc_17692_n12699;
  wire _abc_17692_n1270;
  wire _abc_17692_n12700;
  wire _abc_17692_n12701;
  wire _abc_17692_n12702;
  wire _abc_17692_n12703;
  wire _abc_17692_n12704;
  wire _abc_17692_n12705;
  wire _abc_17692_n12706;
  wire _abc_17692_n12707;
  wire _abc_17692_n12708;
  wire _abc_17692_n12709;
  wire _abc_17692_n1271;
  wire _abc_17692_n12710;
  wire _abc_17692_n12711;
  wire _abc_17692_n12712;
  wire _abc_17692_n12713;
  wire _abc_17692_n12714;
  wire _abc_17692_n12715;
  wire _abc_17692_n12716;
  wire _abc_17692_n12717;
  wire _abc_17692_n12718;
  wire _abc_17692_n12719;
  wire _abc_17692_n1272;
  wire _abc_17692_n12720;
  wire _abc_17692_n12721;
  wire _abc_17692_n12722;
  wire _abc_17692_n12723;
  wire _abc_17692_n12724;
  wire _abc_17692_n12725;
  wire _abc_17692_n12726;
  wire _abc_17692_n12727;
  wire _abc_17692_n12728;
  wire _abc_17692_n12729;
  wire _abc_17692_n12730;
  wire _abc_17692_n12731;
  wire _abc_17692_n12732;
  wire _abc_17692_n12733;
  wire _abc_17692_n12734;
  wire _abc_17692_n12735;
  wire _abc_17692_n12736;
  wire _abc_17692_n12737;
  wire _abc_17692_n12738;
  wire _abc_17692_n12739;
  wire _abc_17692_n1274;
  wire _abc_17692_n12740;
  wire _abc_17692_n12741;
  wire _abc_17692_n12742;
  wire _abc_17692_n12743;
  wire _abc_17692_n12744;
  wire _abc_17692_n12745;
  wire _abc_17692_n12746;
  wire _abc_17692_n12747;
  wire _abc_17692_n12748;
  wire _abc_17692_n12749;
  wire _abc_17692_n1275;
  wire _abc_17692_n12750;
  wire _abc_17692_n12751;
  wire _abc_17692_n12752;
  wire _abc_17692_n12753;
  wire _abc_17692_n12754;
  wire _abc_17692_n12755;
  wire _abc_17692_n12756;
  wire _abc_17692_n12757;
  wire _abc_17692_n12758;
  wire _abc_17692_n12759;
  wire _abc_17692_n1276;
  wire _abc_17692_n12760;
  wire _abc_17692_n12761;
  wire _abc_17692_n12762;
  wire _abc_17692_n12763;
  wire _abc_17692_n12764;
  wire _abc_17692_n12765;
  wire _abc_17692_n12766;
  wire _abc_17692_n12767;
  wire _abc_17692_n12768;
  wire _abc_17692_n12769;
  wire _abc_17692_n1277;
  wire _abc_17692_n12770;
  wire _abc_17692_n12771;
  wire _abc_17692_n12772;
  wire _abc_17692_n12773;
  wire _abc_17692_n12774;
  wire _abc_17692_n12775;
  wire _abc_17692_n12776;
  wire _abc_17692_n12777;
  wire _abc_17692_n12778;
  wire _abc_17692_n12779;
  wire _abc_17692_n1278;
  wire _abc_17692_n12780;
  wire _abc_17692_n12781;
  wire _abc_17692_n12782;
  wire _abc_17692_n12783;
  wire _abc_17692_n12784;
  wire _abc_17692_n12785;
  wire _abc_17692_n12786;
  wire _abc_17692_n12787;
  wire _abc_17692_n12788;
  wire _abc_17692_n12789;
  wire _abc_17692_n1279;
  wire _abc_17692_n12790;
  wire _abc_17692_n12791;
  wire _abc_17692_n12792;
  wire _abc_17692_n12793;
  wire _abc_17692_n12794;
  wire _abc_17692_n12795;
  wire _abc_17692_n12796;
  wire _abc_17692_n12797;
  wire _abc_17692_n12798;
  wire _abc_17692_n12799;
  wire _abc_17692_n1280;
  wire _abc_17692_n12800;
  wire _abc_17692_n12801;
  wire _abc_17692_n12802;
  wire _abc_17692_n12803;
  wire _abc_17692_n12804;
  wire _abc_17692_n12805;
  wire _abc_17692_n12806;
  wire _abc_17692_n12807;
  wire _abc_17692_n12808;
  wire _abc_17692_n12809;
  wire _abc_17692_n1281;
  wire _abc_17692_n12810;
  wire _abc_17692_n12811;
  wire _abc_17692_n12812;
  wire _abc_17692_n12813;
  wire _abc_17692_n12814;
  wire _abc_17692_n12815;
  wire _abc_17692_n12816;
  wire _abc_17692_n12817;
  wire _abc_17692_n12818;
  wire _abc_17692_n12819;
  wire _abc_17692_n1282;
  wire _abc_17692_n12820;
  wire _abc_17692_n12821;
  wire _abc_17692_n12822;
  wire _abc_17692_n12823;
  wire _abc_17692_n12824;
  wire _abc_17692_n12825;
  wire _abc_17692_n12826;
  wire _abc_17692_n12827;
  wire _abc_17692_n12828;
  wire _abc_17692_n12829;
  wire _abc_17692_n1283;
  wire _abc_17692_n12830;
  wire _abc_17692_n12831;
  wire _abc_17692_n12832;
  wire _abc_17692_n12833;
  wire _abc_17692_n12834;
  wire _abc_17692_n12835;
  wire _abc_17692_n12836;
  wire _abc_17692_n12837;
  wire _abc_17692_n12838;
  wire _abc_17692_n12839;
  wire _abc_17692_n1284;
  wire _abc_17692_n12840;
  wire _abc_17692_n12842;
  wire _abc_17692_n12843;
  wire _abc_17692_n12844;
  wire _abc_17692_n12845;
  wire _abc_17692_n12846;
  wire _abc_17692_n12847;
  wire _abc_17692_n12848;
  wire _abc_17692_n12849;
  wire _abc_17692_n1285;
  wire _abc_17692_n12850;
  wire _abc_17692_n12851;
  wire _abc_17692_n12852;
  wire _abc_17692_n12853;
  wire _abc_17692_n12854;
  wire _abc_17692_n12855;
  wire _abc_17692_n12856;
  wire _abc_17692_n12857;
  wire _abc_17692_n12858;
  wire _abc_17692_n12859;
  wire _abc_17692_n1286;
  wire _abc_17692_n12860;
  wire _abc_17692_n12861;
  wire _abc_17692_n12862;
  wire _abc_17692_n12863;
  wire _abc_17692_n12864;
  wire _abc_17692_n12865;
  wire _abc_17692_n12866;
  wire _abc_17692_n12867;
  wire _abc_17692_n12868;
  wire _abc_17692_n12869;
  wire _abc_17692_n1287;
  wire _abc_17692_n12870;
  wire _abc_17692_n12871;
  wire _abc_17692_n12872;
  wire _abc_17692_n12873;
  wire _abc_17692_n12874;
  wire _abc_17692_n12875;
  wire _abc_17692_n12876;
  wire _abc_17692_n12877;
  wire _abc_17692_n12878;
  wire _abc_17692_n12879;
  wire _abc_17692_n1288;
  wire _abc_17692_n12880;
  wire _abc_17692_n12881;
  wire _abc_17692_n12882;
  wire _abc_17692_n12883;
  wire _abc_17692_n12884;
  wire _abc_17692_n12885;
  wire _abc_17692_n12886;
  wire _abc_17692_n12887;
  wire _abc_17692_n12888;
  wire _abc_17692_n12889;
  wire _abc_17692_n1289;
  wire _abc_17692_n12890;
  wire _abc_17692_n12891;
  wire _abc_17692_n12892;
  wire _abc_17692_n12893;
  wire _abc_17692_n12894;
  wire _abc_17692_n12895;
  wire _abc_17692_n12896;
  wire _abc_17692_n12897;
  wire _abc_17692_n12898;
  wire _abc_17692_n12899;
  wire _abc_17692_n1290;
  wire _abc_17692_n12900;
  wire _abc_17692_n12901;
  wire _abc_17692_n12902;
  wire _abc_17692_n12903;
  wire _abc_17692_n12904;
  wire _abc_17692_n12905;
  wire _abc_17692_n12906;
  wire _abc_17692_n12907;
  wire _abc_17692_n12908;
  wire _abc_17692_n12909;
  wire _abc_17692_n1291;
  wire _abc_17692_n12910;
  wire _abc_17692_n12911;
  wire _abc_17692_n12912;
  wire _abc_17692_n12913;
  wire _abc_17692_n12914;
  wire _abc_17692_n12915;
  wire _abc_17692_n12916;
  wire _abc_17692_n12917;
  wire _abc_17692_n12918;
  wire _abc_17692_n12919;
  wire _abc_17692_n1292;
  wire _abc_17692_n12920;
  wire _abc_17692_n12921;
  wire _abc_17692_n12922;
  wire _abc_17692_n12923;
  wire _abc_17692_n12924;
  wire _abc_17692_n12925;
  wire _abc_17692_n12926;
  wire _abc_17692_n12927;
  wire _abc_17692_n12928;
  wire _abc_17692_n12929;
  wire _abc_17692_n1293;
  wire _abc_17692_n12930;
  wire _abc_17692_n12931;
  wire _abc_17692_n12932;
  wire _abc_17692_n12933;
  wire _abc_17692_n12934;
  wire _abc_17692_n12935;
  wire _abc_17692_n12936;
  wire _abc_17692_n12937;
  wire _abc_17692_n12938;
  wire _abc_17692_n12939;
  wire _abc_17692_n1294;
  wire _abc_17692_n12941;
  wire _abc_17692_n12942;
  wire _abc_17692_n12943;
  wire _abc_17692_n12944;
  wire _abc_17692_n12945;
  wire _abc_17692_n12946;
  wire _abc_17692_n12947;
  wire _abc_17692_n12948;
  wire _abc_17692_n1295;
  wire _abc_17692_n12950;
  wire _abc_17692_n12951;
  wire _abc_17692_n12952;
  wire _abc_17692_n12953;
  wire _abc_17692_n12955;
  wire _abc_17692_n1296;
  wire _abc_17692_n1297;
  wire _abc_17692_n1298;
  wire _abc_17692_n1299;
  wire _abc_17692_n1300;
  wire _abc_17692_n1301;
  wire _abc_17692_n1303;
  wire _abc_17692_n1304;
  wire _abc_17692_n1305;
  wire _abc_17692_n1306;
  wire _abc_17692_n1307;
  wire _abc_17692_n1308_1;
  wire _abc_17692_n1309;
  wire _abc_17692_n1310;
  wire _abc_17692_n1311_1;
  wire _abc_17692_n1312;
  wire _abc_17692_n1313;
  wire _abc_17692_n1314;
  wire _abc_17692_n1315;
  wire _abc_17692_n1316;
  wire _abc_17692_n1317;
  wire _abc_17692_n1318;
  wire _abc_17692_n1319;
  wire _abc_17692_n1320_1;
  wire _abc_17692_n1321;
  wire _abc_17692_n1322;
  wire _abc_17692_n1323;
  wire _abc_17692_n1324;
  wire _abc_17692_n1326;
  wire _abc_17692_n1327;
  wire _abc_17692_n1328;
  wire _abc_17692_n1329;
  wire _abc_17692_n1330;
  wire _abc_17692_n1331_1;
  wire _abc_17692_n1332;
  wire _abc_17692_n1333;
  wire _abc_17692_n1334;
  wire _abc_17692_n1335;
  wire _abc_17692_n1336;
  wire _abc_17692_n1337;
  wire _abc_17692_n1338;
  wire _abc_17692_n1339;
  wire _abc_17692_n1340;
  wire _abc_17692_n1341;
  wire _abc_17692_n1342;
  wire _abc_17692_n1343_1;
  wire _abc_17692_n1344;
  wire _abc_17692_n1345;
  wire _abc_17692_n1346;
  wire _abc_17692_n1347;
  wire _abc_17692_n1348;
  wire _abc_17692_n1349;
  wire _abc_17692_n1350;
  wire _abc_17692_n1351;
  wire _abc_17692_n1352;
  wire _abc_17692_n1353;
  wire _abc_17692_n1354;
  wire _abc_17692_n1355_1;
  wire _abc_17692_n1356;
  wire _abc_17692_n1357;
  wire _abc_17692_n1358;
  wire _abc_17692_n1359;
  wire _abc_17692_n1360;
  wire _abc_17692_n1361;
  wire _abc_17692_n1362;
  wire _abc_17692_n1363;
  wire _abc_17692_n1364;
  wire _abc_17692_n1365;
  wire _abc_17692_n1366;
  wire _abc_17692_n1367;
  wire _abc_17692_n1369;
  wire _abc_17692_n1370;
  wire _abc_17692_n1371;
  wire _abc_17692_n1372;
  wire _abc_17692_n1373;
  wire _abc_17692_n1374;
  wire _abc_17692_n1375;
  wire _abc_17692_n1376;
  wire _abc_17692_n1377;
  wire _abc_17692_n1378;
  wire _abc_17692_n1379;
  wire _abc_17692_n1380;
  wire _abc_17692_n1381;
  wire _abc_17692_n1382;
  wire _abc_17692_n1383;
  wire _abc_17692_n1384;
  wire _abc_17692_n1385;
  wire _abc_17692_n1386;
  wire _abc_17692_n1387;
  wire _abc_17692_n1388;
  wire _abc_17692_n1389_1;
  wire _abc_17692_n1390;
  wire _abc_17692_n1391;
  wire _abc_17692_n1392_1;
  wire _abc_17692_n1393;
  wire _abc_17692_n1394;
  wire _abc_17692_n1395;
  wire _abc_17692_n1396;
  wire _abc_17692_n1398;
  wire _abc_17692_n1399;
  wire _abc_17692_n1400;
  wire _abc_17692_n1401;
  wire _abc_17692_n1402;
  wire _abc_17692_n1403_1;
  wire _abc_17692_n1404;
  wire _abc_17692_n1405;
  wire _abc_17692_n1406;
  wire _abc_17692_n1407;
  wire _abc_17692_n1408;
  wire _abc_17692_n1409;
  wire _abc_17692_n1410;
  wire _abc_17692_n1411;
  wire _abc_17692_n1412;
  wire _abc_17692_n1413;
  wire _abc_17692_n1414;
  wire _abc_17692_n1415;
  wire _abc_17692_n1416;
  wire _abc_17692_n1417;
  wire _abc_17692_n1418;
  wire _abc_17692_n1419;
  wire _abc_17692_n1420;
  wire _abc_17692_n1421_1;
  wire _abc_17692_n1422;
  wire _abc_17692_n1423;
  wire _abc_17692_n1424;
  wire _abc_17692_n1425;
  wire _abc_17692_n1426;
  wire _abc_17692_n1427;
  wire _abc_17692_n1428;
  wire _abc_17692_n1430;
  wire _abc_17692_n1431;
  wire _abc_17692_n1432;
  wire _abc_17692_n1433;
  wire _abc_17692_n1434;
  wire _abc_17692_n1435;
  wire _abc_17692_n1436;
  wire _abc_17692_n1437;
  wire _abc_17692_n1438;
  wire _abc_17692_n1439;
  wire _abc_17692_n1440;
  wire _abc_17692_n1441_1;
  wire _abc_17692_n1442;
  wire _abc_17692_n1443;
  wire _abc_17692_n1444;
  wire _abc_17692_n1445;
  wire _abc_17692_n1446;
  wire _abc_17692_n1447;
  wire _abc_17692_n1448;
  wire _abc_17692_n1449;
  wire _abc_17692_n1450;
  wire _abc_17692_n1451;
  wire _abc_17692_n1452;
  wire _abc_17692_n1453;
  wire _abc_17692_n1454;
  wire _abc_17692_n1456;
  wire _abc_17692_n1457;
  wire _abc_17692_n1458;
  wire _abc_17692_n1459_1;
  wire _abc_17692_n1460;
  wire _abc_17692_n1461;
  wire _abc_17692_n1462;
  wire _abc_17692_n1463;
  wire _abc_17692_n1464;
  wire _abc_17692_n1465;
  wire _abc_17692_n1466;
  wire _abc_17692_n1467;
  wire _abc_17692_n1468;
  wire _abc_17692_n1469;
  wire _abc_17692_n1470;
  wire _abc_17692_n1471;
  wire _abc_17692_n1472;
  wire _abc_17692_n1473;
  wire _abc_17692_n1474;
  wire _abc_17692_n1475;
  wire _abc_17692_n1476;
  wire _abc_17692_n1477;
  wire _abc_17692_n1478;
  wire _abc_17692_n1479;
  wire _abc_17692_n1480;
  wire _abc_17692_n1481;
  wire _abc_17692_n1482;
  wire _abc_17692_n1483;
  wire _abc_17692_n1484;
  wire _abc_17692_n1485;
  wire _abc_17692_n1486;
  wire _abc_17692_n1487;
  wire _abc_17692_n1488;
  wire _abc_17692_n1489;
  wire _abc_17692_n1490;
  wire _abc_17692_n1491;
  wire _abc_17692_n1492;
  wire _abc_17692_n1494;
  wire _abc_17692_n1495;
  wire _abc_17692_n1496;
  wire _abc_17692_n1497;
  wire _abc_17692_n1498;
  wire _abc_17692_n1499;
  wire _abc_17692_n1500;
  wire _abc_17692_n1501;
  wire _abc_17692_n1502;
  wire _abc_17692_n1503;
  wire _abc_17692_n1504;
  wire _abc_17692_n1505;
  wire _abc_17692_n1506;
  wire _abc_17692_n1507;
  wire _abc_17692_n1508;
  wire _abc_17692_n1509;
  wire _abc_17692_n1510;
  wire _abc_17692_n1511;
  wire _abc_17692_n1512;
  wire _abc_17692_n1513;
  wire _abc_17692_n1514;
  wire _abc_17692_n1515;
  wire _abc_17692_n1516;
  wire _abc_17692_n1517_1;
  wire _abc_17692_n1518;
  wire _abc_17692_n1519;
  wire _abc_17692_n1520_1;
  wire _abc_17692_n1521;
  wire _abc_17692_n1522;
  wire _abc_17692_n1524;
  wire _abc_17692_n1525;
  wire _abc_17692_n1526_1;
  wire _abc_17692_n1527;
  wire _abc_17692_n1528;
  wire _abc_17692_n1529;
  wire _abc_17692_n1530;
  wire _abc_17692_n1531;
  wire _abc_17692_n1532;
  wire _abc_17692_n1533;
  wire _abc_17692_n1534;
  wire _abc_17692_n1535;
  wire _abc_17692_n1536;
  wire _abc_17692_n1537;
  wire _abc_17692_n1538_1;
  wire _abc_17692_n1539;
  wire _abc_17692_n1540;
  wire _abc_17692_n1541;
  wire _abc_17692_n1542;
  wire _abc_17692_n1543;
  wire _abc_17692_n1544;
  wire _abc_17692_n1545;
  wire _abc_17692_n1546;
  wire _abc_17692_n1547;
  wire _abc_17692_n1548;
  wire _abc_17692_n1549;
  wire _abc_17692_n1550_1;
  wire _abc_17692_n1551;
  wire _abc_17692_n1552;
  wire _abc_17692_n1553;
  wire _abc_17692_n1555;
  wire _abc_17692_n1556;
  wire _abc_17692_n1557;
  wire _abc_17692_n1558;
  wire _abc_17692_n1559;
  wire _abc_17692_n1560;
  wire _abc_17692_n1561;
  wire _abc_17692_n1562_1;
  wire _abc_17692_n1563;
  wire _abc_17692_n1564;
  wire _abc_17692_n1565;
  wire _abc_17692_n1566;
  wire _abc_17692_n1567;
  wire _abc_17692_n1568;
  wire _abc_17692_n1569;
  wire _abc_17692_n1570;
  wire _abc_17692_n1571;
  wire _abc_17692_n1572;
  wire _abc_17692_n1573;
  wire _abc_17692_n1574;
  wire _abc_17692_n1575;
  wire _abc_17692_n1576;
  wire _abc_17692_n1577;
  wire _abc_17692_n1578;
  wire _abc_17692_n1579;
  wire _abc_17692_n1581;
  wire _abc_17692_n1582;
  wire _abc_17692_n1583;
  wire _abc_17692_n1584;
  wire _abc_17692_n1585;
  wire _abc_17692_n1586;
  wire _abc_17692_n1587;
  wire _abc_17692_n1588;
  wire _abc_17692_n1589;
  wire _abc_17692_n1590;
  wire _abc_17692_n1591;
  wire _abc_17692_n1592;
  wire _abc_17692_n1593;
  wire _abc_17692_n1594;
  wire _abc_17692_n1595_1;
  wire _abc_17692_n1596;
  wire _abc_17692_n1597;
  wire _abc_17692_n1598_1;
  wire _abc_17692_n1599;
  wire _abc_17692_n1600;
  wire _abc_17692_n1601;
  wire _abc_17692_n1602;
  wire _abc_17692_n1603;
  wire _abc_17692_n1604;
  wire _abc_17692_n1605;
  wire _abc_17692_n1606;
  wire _abc_17692_n1607;
  wire _abc_17692_n1608;
  wire _abc_17692_n1609;
  wire _abc_17692_n1610;
  wire _abc_17692_n1611;
  wire _abc_17692_n1612;
  wire _abc_17692_n1613_1;
  wire _abc_17692_n1614;
  wire _abc_17692_n1615;
  wire _abc_17692_n1616;
  wire _abc_17692_n1617;
  wire _abc_17692_n1618;
  wire _abc_17692_n1619;
  wire _abc_17692_n1620;
  wire _abc_17692_n1622;
  wire _abc_17692_n1623;
  wire _abc_17692_n1624;
  wire _abc_17692_n1625;
  wire _abc_17692_n1626;
  wire _abc_17692_n1627;
  wire _abc_17692_n1628;
  wire _abc_17692_n1629;
  wire _abc_17692_n1630;
  wire _abc_17692_n1631;
  wire _abc_17692_n1632;
  wire _abc_17692_n1633;
  wire _abc_17692_n1634;
  wire _abc_17692_n1635;
  wire _abc_17692_n1636_1;
  wire _abc_17692_n1637;
  wire _abc_17692_n1638;
  wire _abc_17692_n1639;
  wire _abc_17692_n1640;
  wire _abc_17692_n1641;
  wire _abc_17692_n1642;
  wire _abc_17692_n1643;
  wire _abc_17692_n1644;
  wire _abc_17692_n1645;
  wire _abc_17692_n1646;
  wire _abc_17692_n1647;
  wire _abc_17692_n1648;
  wire _abc_17692_n1649;
  wire _abc_17692_n1651;
  wire _abc_17692_n1652;
  wire _abc_17692_n1653;
  wire _abc_17692_n1654;
  wire _abc_17692_n1655;
  wire _abc_17692_n1656;
  wire _abc_17692_n1657;
  wire _abc_17692_n1658;
  wire _abc_17692_n1659;
  wire _abc_17692_n1660_1;
  wire _abc_17692_n1661;
  wire _abc_17692_n1662;
  wire _abc_17692_n1663;
  wire _abc_17692_n1664;
  wire _abc_17692_n1665;
  wire _abc_17692_n1666;
  wire _abc_17692_n1667;
  wire _abc_17692_n1668;
  wire _abc_17692_n1669;
  wire _abc_17692_n1670;
  wire _abc_17692_n1671;
  wire _abc_17692_n1672;
  wire _abc_17692_n1673;
  wire _abc_17692_n1674;
  wire _abc_17692_n1675;
  wire _abc_17692_n1676;
  wire _abc_17692_n1677;
  wire _abc_17692_n1678;
  wire _abc_17692_n1679;
  wire _abc_17692_n1680;
  wire _abc_17692_n1682;
  wire _abc_17692_n1683;
  wire _abc_17692_n1684;
  wire _abc_17692_n1685_1;
  wire _abc_17692_n1686;
  wire _abc_17692_n1687;
  wire _abc_17692_n1688;
  wire _abc_17692_n1689;
  wire _abc_17692_n1690;
  wire _abc_17692_n1691;
  wire _abc_17692_n1692;
  wire _abc_17692_n1693;
  wire _abc_17692_n1694;
  wire _abc_17692_n1695;
  wire _abc_17692_n1696;
  wire _abc_17692_n1697;
  wire _abc_17692_n1698;
  wire _abc_17692_n1699;
  wire _abc_17692_n1700;
  wire _abc_17692_n1701;
  wire _abc_17692_n1702;
  wire _abc_17692_n1703;
  wire _abc_17692_n1704;
  wire _abc_17692_n1705;
  wire _abc_17692_n1706;
  wire _abc_17692_n1707;
  wire _abc_17692_n1708;
  wire _abc_17692_n1709;
  wire _abc_17692_n1710;
  wire _abc_17692_n1712;
  wire _abc_17692_n1713;
  wire _abc_17692_n1714;
  wire _abc_17692_n1715;
  wire _abc_17692_n1716;
  wire _abc_17692_n1717;
  wire _abc_17692_n1718;
  wire _abc_17692_n1719;
  wire _abc_17692_n1720;
  wire _abc_17692_n1721;
  wire _abc_17692_n1722;
  wire _abc_17692_n1723;
  wire _abc_17692_n1724;
  wire _abc_17692_n1725;
  wire _abc_17692_n1726;
  wire _abc_17692_n1727;
  wire _abc_17692_n1728;
  wire _abc_17692_n1729;
  wire _abc_17692_n1730;
  wire _abc_17692_n1731;
  wire _abc_17692_n1732;
  wire _abc_17692_n1733;
  wire _abc_17692_n1734;
  wire _abc_17692_n1735;
  wire _abc_17692_n1736;
  wire _abc_17692_n1738;
  wire _abc_17692_n1739;
  wire _abc_17692_n1740;
  wire _abc_17692_n1741;
  wire _abc_17692_n1742;
  wire _abc_17692_n1743;
  wire _abc_17692_n1744;
  wire _abc_17692_n1745;
  wire _abc_17692_n1746;
  wire _abc_17692_n1747;
  wire _abc_17692_n1748;
  wire _abc_17692_n1749;
  wire _abc_17692_n1750;
  wire _abc_17692_n1751;
  wire _abc_17692_n1752;
  wire _abc_17692_n1753;
  wire _abc_17692_n1754;
  wire _abc_17692_n1755_1;
  wire _abc_17692_n1756;
  wire _abc_17692_n1757;
  wire _abc_17692_n1758_1;
  wire _abc_17692_n1759;
  wire _abc_17692_n1760;
  wire _abc_17692_n1761;
  wire _abc_17692_n1763;
  wire _abc_17692_n1764;
  wire _abc_17692_n1765;
  wire _abc_17692_n1766;
  wire _abc_17692_n1767;
  wire _abc_17692_n1768;
  wire _abc_17692_n1769;
  wire _abc_17692_n1770;
  wire _abc_17692_n1771;
  wire _abc_17692_n1772;
  wire _abc_17692_n1773;
  wire _abc_17692_n1774;
  wire _abc_17692_n1775_1;
  wire _abc_17692_n1776;
  wire _abc_17692_n1777;
  wire _abc_17692_n1778;
  wire _abc_17692_n1779;
  wire _abc_17692_n1780;
  wire _abc_17692_n1781;
  wire _abc_17692_n1782;
  wire _abc_17692_n1783;
  wire _abc_17692_n1784;
  wire _abc_17692_n1785;
  wire _abc_17692_n1786;
  wire _abc_17692_n1787;
  wire _abc_17692_n1788_1;
  wire _abc_17692_n1790;
  wire _abc_17692_n1791;
  wire _abc_17692_n1792;
  wire _abc_17692_n1793;
  wire _abc_17692_n1794;
  wire _abc_17692_n1795;
  wire _abc_17692_n1796;
  wire _abc_17692_n1797;
  wire _abc_17692_n1798;
  wire _abc_17692_n1799;
  wire _abc_17692_n1800;
  wire _abc_17692_n1801;
  wire _abc_17692_n1802;
  wire _abc_17692_n1803;
  wire _abc_17692_n1804_1;
  wire _abc_17692_n1805;
  wire _abc_17692_n1806;
  wire _abc_17692_n1807;
  wire _abc_17692_n1808;
  wire _abc_17692_n1809;
  wire _abc_17692_n1810;
  wire _abc_17692_n1811;
  wire _abc_17692_n1812;
  wire _abc_17692_n1814;
  wire _abc_17692_n1815_1;
  wire _abc_17692_n1816;
  wire _abc_17692_n1817;
  wire _abc_17692_n1818;
  wire _abc_17692_n1819;
  wire _abc_17692_n1820;
  wire _abc_17692_n1821;
  wire _abc_17692_n1822;
  wire _abc_17692_n1823;
  wire _abc_17692_n1824;
  wire _abc_17692_n1825;
  wire _abc_17692_n1826;
  wire _abc_17692_n1827;
  wire _abc_17692_n1828;
  wire _abc_17692_n1829;
  wire _abc_17692_n1830;
  wire _abc_17692_n1830_bF_buf0;
  wire _abc_17692_n1830_bF_buf1;
  wire _abc_17692_n1830_bF_buf10;
  wire _abc_17692_n1830_bF_buf2;
  wire _abc_17692_n1830_bF_buf3;
  wire _abc_17692_n1830_bF_buf4;
  wire _abc_17692_n1830_bF_buf5;
  wire _abc_17692_n1830_bF_buf6;
  wire _abc_17692_n1830_bF_buf7;
  wire _abc_17692_n1830_bF_buf8;
  wire _abc_17692_n1830_bF_buf9;
  wire _abc_17692_n1831;
  wire _abc_17692_n1832;
  wire _abc_17692_n1833;
  wire _abc_17692_n1834;
  wire _abc_17692_n1835;
  wire _abc_17692_n1836;
  wire _abc_17692_n1837;
  wire _abc_17692_n1838;
  wire _abc_17692_n1839;
  wire _abc_17692_n1840;
  wire _abc_17692_n1841;
  wire _abc_17692_n1842;
  wire _abc_17692_n1843;
  wire _abc_17692_n1844;
  wire _abc_17692_n1845;
  wire _abc_17692_n1846;
  wire _abc_17692_n1846_bF_buf0;
  wire _abc_17692_n1846_bF_buf1;
  wire _abc_17692_n1846_bF_buf10;
  wire _abc_17692_n1846_bF_buf2;
  wire _abc_17692_n1846_bF_buf3;
  wire _abc_17692_n1846_bF_buf4;
  wire _abc_17692_n1846_bF_buf5;
  wire _abc_17692_n1846_bF_buf6;
  wire _abc_17692_n1846_bF_buf7;
  wire _abc_17692_n1846_bF_buf8;
  wire _abc_17692_n1846_bF_buf9;
  wire _abc_17692_n1847;
  wire _abc_17692_n1848;
  wire _abc_17692_n1849;
  wire _abc_17692_n1850;
  wire _abc_17692_n1851;
  wire _abc_17692_n1852_1;
  wire _abc_17692_n1853;
  wire _abc_17692_n1854;
  wire _abc_17692_n1855_1;
  wire _abc_17692_n1856;
  wire _abc_17692_n1857;
  wire _abc_17692_n1858;
  wire _abc_17692_n1859;
  wire _abc_17692_n1860;
  wire _abc_17692_n1861;
  wire _abc_17692_n1862;
  wire _abc_17692_n1863;
  wire _abc_17692_n1863_bF_buf0;
  wire _abc_17692_n1863_bF_buf1;
  wire _abc_17692_n1863_bF_buf10;
  wire _abc_17692_n1863_bF_buf2;
  wire _abc_17692_n1863_bF_buf3;
  wire _abc_17692_n1863_bF_buf4;
  wire _abc_17692_n1863_bF_buf5;
  wire _abc_17692_n1863_bF_buf6;
  wire _abc_17692_n1863_bF_buf7;
  wire _abc_17692_n1863_bF_buf8;
  wire _abc_17692_n1863_bF_buf9;
  wire _abc_17692_n1864;
  wire _abc_17692_n1865;
  wire _abc_17692_n1866;
  wire _abc_17692_n1867_1;
  wire _abc_17692_n1868;
  wire _abc_17692_n1869;
  wire _abc_17692_n1870;
  wire _abc_17692_n1871;
  wire _abc_17692_n1872;
  wire _abc_17692_n1873;
  wire _abc_17692_n1874;
  wire _abc_17692_n1875;
  wire _abc_17692_n1876;
  wire _abc_17692_n1877;
  wire _abc_17692_n1877_bF_buf0;
  wire _abc_17692_n1877_bF_buf1;
  wire _abc_17692_n1877_bF_buf10;
  wire _abc_17692_n1877_bF_buf2;
  wire _abc_17692_n1877_bF_buf3;
  wire _abc_17692_n1877_bF_buf4;
  wire _abc_17692_n1877_bF_buf5;
  wire _abc_17692_n1877_bF_buf6;
  wire _abc_17692_n1877_bF_buf7;
  wire _abc_17692_n1877_bF_buf8;
  wire _abc_17692_n1877_bF_buf9;
  wire _abc_17692_n1878;
  wire _abc_17692_n1879;
  wire _abc_17692_n1880;
  wire _abc_17692_n1881;
  wire _abc_17692_n1882;
  wire _abc_17692_n1883;
  wire _abc_17692_n1884_1;
  wire _abc_17692_n1885;
  wire _abc_17692_n1885_bF_buf0;
  wire _abc_17692_n1885_bF_buf1;
  wire _abc_17692_n1885_bF_buf2;
  wire _abc_17692_n1885_bF_buf3;
  wire _abc_17692_n1885_bF_buf4;
  wire _abc_17692_n1886;
  wire _abc_17692_n1887;
  wire _abc_17692_n1888;
  wire _abc_17692_n1890;
  wire _abc_17692_n1891;
  wire _abc_17692_n1892;
  wire _abc_17692_n1893;
  wire _abc_17692_n1894;
  wire _abc_17692_n1895;
  wire _abc_17692_n1896;
  wire _abc_17692_n1897;
  wire _abc_17692_n1898;
  wire _abc_17692_n1899;
  wire _abc_17692_n1900;
  wire _abc_17692_n1901_1;
  wire _abc_17692_n1902;
  wire _abc_17692_n1903;
  wire _abc_17692_n1904;
  wire _abc_17692_n1905;
  wire _abc_17692_n1906;
  wire _abc_17692_n1907;
  wire _abc_17692_n1908;
  wire _abc_17692_n1909;
  wire _abc_17692_n1910;
  wire _abc_17692_n1911;
  wire _abc_17692_n1912;
  wire _abc_17692_n1913;
  wire _abc_17692_n1914;
  wire _abc_17692_n1915;
  wire _abc_17692_n1916;
  wire _abc_17692_n1917;
  wire _abc_17692_n1918;
  wire _abc_17692_n1919_1;
  wire _abc_17692_n1920;
  wire _abc_17692_n1921;
  wire _abc_17692_n1922;
  wire _abc_17692_n1923;
  wire _abc_17692_n1924;
  wire _abc_17692_n1925;
  wire _abc_17692_n1926;
  wire _abc_17692_n1927;
  wire _abc_17692_n1928;
  wire _abc_17692_n1929;
  wire _abc_17692_n1930;
  wire _abc_17692_n1931;
  wire _abc_17692_n1932;
  wire _abc_17692_n1933;
  wire _abc_17692_n1934;
  wire _abc_17692_n1935;
  wire _abc_17692_n1936;
  wire _abc_17692_n1937;
  wire _abc_17692_n1938;
  wire _abc_17692_n1939;
  wire _abc_17692_n1940;
  wire _abc_17692_n1941;
  wire _abc_17692_n1942;
  wire _abc_17692_n1943;
  wire _abc_17692_n1944;
  wire _abc_17692_n1945;
  wire _abc_17692_n1946;
  wire _abc_17692_n1947;
  wire _abc_17692_n1948;
  wire _abc_17692_n1949;
  wire _abc_17692_n1950;
  wire _abc_17692_n1951;
  wire _abc_17692_n1952;
  wire _abc_17692_n1953;
  wire _abc_17692_n1954;
  wire _abc_17692_n1955;
  wire _abc_17692_n1956;
  wire _abc_17692_n1957;
  wire _abc_17692_n1958;
  wire _abc_17692_n1959;
  wire _abc_17692_n1960;
  wire _abc_17692_n1961;
  wire _abc_17692_n1962;
  wire _abc_17692_n1963;
  wire _abc_17692_n1964;
  wire _abc_17692_n1965;
  wire _abc_17692_n1966;
  wire _abc_17692_n1967;
  wire _abc_17692_n1968;
  wire _abc_17692_n1969;
  wire _abc_17692_n1970;
  wire _abc_17692_n1971_1;
  wire _abc_17692_n1972;
  wire _abc_17692_n1973;
  wire _abc_17692_n1974_1;
  wire _abc_17692_n1975;
  wire _abc_17692_n1976;
  wire _abc_17692_n1977;
  wire _abc_17692_n1978;
  wire _abc_17692_n1979;
  wire _abc_17692_n1980;
  wire _abc_17692_n1981_1;
  wire _abc_17692_n1982;
  wire _abc_17692_n1983;
  wire _abc_17692_n1984;
  wire _abc_17692_n1985;
  wire _abc_17692_n1986;
  wire _abc_17692_n1987;
  wire _abc_17692_n1988;
  wire _abc_17692_n1989;
  wire _abc_17692_n1990;
  wire _abc_17692_n1991;
  wire _abc_17692_n1992;
  wire _abc_17692_n1993_1;
  wire _abc_17692_n1994;
  wire _abc_17692_n1995;
  wire _abc_17692_n1996;
  wire _abc_17692_n1997;
  wire _abc_17692_n1998;
  wire _abc_17692_n1999;
  wire _abc_17692_n2000;
  wire _abc_17692_n2001;
  wire _abc_17692_n2002;
  wire _abc_17692_n2003;
  wire _abc_17692_n2004_1;
  wire _abc_17692_n2005;
  wire _abc_17692_n2006;
  wire _abc_17692_n2007;
  wire _abc_17692_n2008;
  wire _abc_17692_n2009;
  wire _abc_17692_n2010;
  wire _abc_17692_n2011;
  wire _abc_17692_n2012;
  wire _abc_17692_n2013;
  wire _abc_17692_n2014;
  wire _abc_17692_n2015;
  wire _abc_17692_n2016_1;
  wire _abc_17692_n2017;
  wire _abc_17692_n2018;
  wire _abc_17692_n2019;
  wire _abc_17692_n2020;
  wire _abc_17692_n2021;
  wire _abc_17692_n2022;
  wire _abc_17692_n2023;
  wire _abc_17692_n2024;
  wire _abc_17692_n2025;
  wire _abc_17692_n2026;
  wire _abc_17692_n2027;
  wire _abc_17692_n2028;
  wire _abc_17692_n2029;
  wire _abc_17692_n2030;
  wire _abc_17692_n2031;
  wire _abc_17692_n2032;
  wire _abc_17692_n2033;
  wire _abc_17692_n2034;
  wire _abc_17692_n2035;
  wire _abc_17692_n2036;
  wire _abc_17692_n2037;
  wire _abc_17692_n2038;
  wire _abc_17692_n2039;
  wire _abc_17692_n2040;
  wire _abc_17692_n2041;
  wire _abc_17692_n2042;
  wire _abc_17692_n2043;
  wire _abc_17692_n2044;
  wire _abc_17692_n2045;
  wire _abc_17692_n2046;
  wire _abc_17692_n2047;
  wire _abc_17692_n2048;
  wire _abc_17692_n2049_1;
  wire _abc_17692_n2050;
  wire _abc_17692_n2051;
  wire _abc_17692_n2052_1;
  wire _abc_17692_n2053;
  wire _abc_17692_n2054;
  wire _abc_17692_n2055;
  wire _abc_17692_n2056;
  wire _abc_17692_n2057;
  wire _abc_17692_n2058;
  wire _abc_17692_n2060;
  wire _abc_17692_n2061;
  wire _abc_17692_n2062_1;
  wire _abc_17692_n2063;
  wire _abc_17692_n2064;
  wire _abc_17692_n2065;
  wire _abc_17692_n2066;
  wire _abc_17692_n2067;
  wire _abc_17692_n2068;
  wire _abc_17692_n2069;
  wire _abc_17692_n2070;
  wire _abc_17692_n2071;
  wire _abc_17692_n2072;
  wire _abc_17692_n2073;
  wire _abc_17692_n2074;
  wire _abc_17692_n2075;
  wire _abc_17692_n2076;
  wire _abc_17692_n2077;
  wire _abc_17692_n2078;
  wire _abc_17692_n2079;
  wire _abc_17692_n2080;
  wire _abc_17692_n2081;
  wire _abc_17692_n2082;
  wire _abc_17692_n2083;
  wire _abc_17692_n2084;
  wire _abc_17692_n2085;
  wire _abc_17692_n2086;
  wire _abc_17692_n2087_1;
  wire _abc_17692_n2088;
  wire _abc_17692_n2089;
  wire _abc_17692_n2090;
  wire _abc_17692_n2091;
  wire _abc_17692_n2092;
  wire _abc_17692_n2093;
  wire _abc_17692_n2094;
  wire _abc_17692_n2095;
  wire _abc_17692_n2096;
  wire _abc_17692_n2097;
  wire _abc_17692_n2098;
  wire _abc_17692_n2099;
  wire _abc_17692_n2100;
  wire _abc_17692_n2101;
  wire _abc_17692_n2102;
  wire _abc_17692_n2103;
  wire _abc_17692_n2104;
  wire _abc_17692_n2105;
  wire _abc_17692_n2106;
  wire _abc_17692_n2107;
  wire _abc_17692_n2108;
  wire _abc_17692_n2109;
  wire _abc_17692_n2110;
  wire _abc_17692_n2111;
  wire _abc_17692_n2112_1;
  wire _abc_17692_n2113;
  wire _abc_17692_n2114;
  wire _abc_17692_n2115;
  wire _abc_17692_n2116;
  wire _abc_17692_n2117;
  wire _abc_17692_n2118;
  wire _abc_17692_n2119;
  wire _abc_17692_n2120;
  wire _abc_17692_n2121;
  wire _abc_17692_n2122;
  wire _abc_17692_n2123;
  wire _abc_17692_n2124;
  wire _abc_17692_n2125;
  wire _abc_17692_n2126;
  wire _abc_17692_n2127;
  wire _abc_17692_n2128;
  wire _abc_17692_n2129;
  wire _abc_17692_n2130;
  wire _abc_17692_n2131;
  wire _abc_17692_n2132;
  wire _abc_17692_n2133;
  wire _abc_17692_n2134;
  wire _abc_17692_n2135;
  wire _abc_17692_n2136;
  wire _abc_17692_n2137_1;
  wire _abc_17692_n2138;
  wire _abc_17692_n2139;
  wire _abc_17692_n2140;
  wire _abc_17692_n2141;
  wire _abc_17692_n2142;
  wire _abc_17692_n2143;
  wire _abc_17692_n2144;
  wire _abc_17692_n2145;
  wire _abc_17692_n2146;
  wire _abc_17692_n2147;
  wire _abc_17692_n2148;
  wire _abc_17692_n2149;
  wire _abc_17692_n2150;
  wire _abc_17692_n2151;
  wire _abc_17692_n2152;
  wire _abc_17692_n2153;
  wire _abc_17692_n2154;
  wire _abc_17692_n2155;
  wire _abc_17692_n2156;
  wire _abc_17692_n2157;
  wire _abc_17692_n2158;
  wire _abc_17692_n2159;
  wire _abc_17692_n2160;
  wire _abc_17692_n2161;
  wire _abc_17692_n2162;
  wire _abc_17692_n2163;
  wire _abc_17692_n2164;
  wire _abc_17692_n2165;
  wire _abc_17692_n2166;
  wire _abc_17692_n2167;
  wire _abc_17692_n2168;
  wire _abc_17692_n2169;
  wire _abc_17692_n2170;
  wire _abc_17692_n2171;
  wire _abc_17692_n2172;
  wire _abc_17692_n2173;
  wire _abc_17692_n2174;
  wire _abc_17692_n2175;
  wire _abc_17692_n2176;
  wire _abc_17692_n2177;
  wire _abc_17692_n2178;
  wire _abc_17692_n2179;
  wire _abc_17692_n2180;
  wire _abc_17692_n2181;
  wire _abc_17692_n2182;
  wire _abc_17692_n2183;
  wire _abc_17692_n2184;
  wire _abc_17692_n2185;
  wire _abc_17692_n2186;
  wire _abc_17692_n2187;
  wire _abc_17692_n2188;
  wire _abc_17692_n2189;
  wire _abc_17692_n2190;
  wire _abc_17692_n2191;
  wire _abc_17692_n2192;
  wire _abc_17692_n2193;
  wire _abc_17692_n2194;
  wire _abc_17692_n2195;
  wire _abc_17692_n2196;
  wire _abc_17692_n2197;
  wire _abc_17692_n2198;
  wire _abc_17692_n2199;
  wire _abc_17692_n2200;
  wire _abc_17692_n2201;
  wire _abc_17692_n2202;
  wire _abc_17692_n2203;
  wire _abc_17692_n2204;
  wire _abc_17692_n2205;
  wire _abc_17692_n2206;
  wire _abc_17692_n2207;
  wire _abc_17692_n2208;
  wire _abc_17692_n2209;
  wire _abc_17692_n2210;
  wire _abc_17692_n2211_1;
  wire _abc_17692_n2212;
  wire _abc_17692_n2213;
  wire _abc_17692_n2214_1;
  wire _abc_17692_n2215;
  wire _abc_17692_n2216;
  wire _abc_17692_n2217;
  wire _abc_17692_n2218;
  wire _abc_17692_n2219;
  wire _abc_17692_n2220;
  wire _abc_17692_n2221;
  wire _abc_17692_n2222;
  wire _abc_17692_n2223;
  wire _abc_17692_n2224;
  wire _abc_17692_n2225;
  wire _abc_17692_n2226_1;
  wire _abc_17692_n2227;
  wire _abc_17692_n2228;
  wire _abc_17692_n2229;
  wire _abc_17692_n2230;
  wire _abc_17692_n2231;
  wire _abc_17692_n2232;
  wire _abc_17692_n2233;
  wire _abc_17692_n2234;
  wire _abc_17692_n2235;
  wire _abc_17692_n2236;
  wire _abc_17692_n2237;
  wire _abc_17692_n2238;
  wire _abc_17692_n2239;
  wire _abc_17692_n2240;
  wire _abc_17692_n2241;
  wire _abc_17692_n2242_1;
  wire _abc_17692_n2243;
  wire _abc_17692_n2244;
  wire _abc_17692_n2246;
  wire _abc_17692_n2247;
  wire _abc_17692_n2248;
  wire _abc_17692_n2249;
  wire _abc_17692_n2250;
  wire _abc_17692_n2251;
  wire _abc_17692_n2252;
  wire _abc_17692_n2253;
  wire _abc_17692_n2254;
  wire _abc_17692_n2255;
  wire _abc_17692_n2256;
  wire _abc_17692_n2257_1;
  wire _abc_17692_n2258;
  wire _abc_17692_n2259;
  wire _abc_17692_n2260;
  wire _abc_17692_n2261;
  wire _abc_17692_n2262;
  wire _abc_17692_n2263;
  wire _abc_17692_n2264;
  wire _abc_17692_n2265;
  wire _abc_17692_n2266;
  wire _abc_17692_n2267;
  wire _abc_17692_n2268;
  wire _abc_17692_n2269;
  wire _abc_17692_n2270;
  wire _abc_17692_n2271;
  wire _abc_17692_n2272;
  wire _abc_17692_n2273;
  wire _abc_17692_n2274;
  wire _abc_17692_n2275;
  wire _abc_17692_n2276;
  wire _abc_17692_n2277;
  wire _abc_17692_n2278_1;
  wire _abc_17692_n2279;
  wire _abc_17692_n2280;
  wire _abc_17692_n2281;
  wire _abc_17692_n2282;
  wire _abc_17692_n2283;
  wire _abc_17692_n2284;
  wire _abc_17692_n2285;
  wire _abc_17692_n2286;
  wire _abc_17692_n2287;
  wire _abc_17692_n2288;
  wire _abc_17692_n2289;
  wire _abc_17692_n2290;
  wire _abc_17692_n2291;
  wire _abc_17692_n2292;
  wire _abc_17692_n2293;
  wire _abc_17692_n2294;
  wire _abc_17692_n2295;
  wire _abc_17692_n2296;
  wire _abc_17692_n2297;
  wire _abc_17692_n2298;
  wire _abc_17692_n2299;
  wire _abc_17692_n2300;
  wire _abc_17692_n2301;
  wire _abc_17692_n2302;
  wire _abc_17692_n2303;
  wire _abc_17692_n2304;
  wire _abc_17692_n2305;
  wire _abc_17692_n2306;
  wire _abc_17692_n2307;
  wire _abc_17692_n2308;
  wire _abc_17692_n2309;
  wire _abc_17692_n2310;
  wire _abc_17692_n2311;
  wire _abc_17692_n2312;
  wire _abc_17692_n2313;
  wire _abc_17692_n2314;
  wire _abc_17692_n2315;
  wire _abc_17692_n2316;
  wire _abc_17692_n2317;
  wire _abc_17692_n2318;
  wire _abc_17692_n2319;
  wire _abc_17692_n2320;
  wire _abc_17692_n2321;
  wire _abc_17692_n2322;
  wire _abc_17692_n2323;
  wire _abc_17692_n2324;
  wire _abc_17692_n2325;
  wire _abc_17692_n2326_1;
  wire _abc_17692_n2327;
  wire _abc_17692_n2328;
  wire _abc_17692_n2329_1;
  wire _abc_17692_n2330;
  wire _abc_17692_n2331;
  wire _abc_17692_n2332;
  wire _abc_17692_n2333;
  wire _abc_17692_n2334;
  wire _abc_17692_n2335;
  wire _abc_17692_n2336;
  wire _abc_17692_n2337;
  wire _abc_17692_n2338;
  wire _abc_17692_n2339;
  wire _abc_17692_n2340_1;
  wire _abc_17692_n2341;
  wire _abc_17692_n2342;
  wire _abc_17692_n2343;
  wire _abc_17692_n2344;
  wire _abc_17692_n2345;
  wire _abc_17692_n2346;
  wire _abc_17692_n2347;
  wire _abc_17692_n2348;
  wire _abc_17692_n2349;
  wire _abc_17692_n2350;
  wire _abc_17692_n2351;
  wire _abc_17692_n2352;
  wire _abc_17692_n2353;
  wire _abc_17692_n2354;
  wire _abc_17692_n2355;
  wire _abc_17692_n2356;
  wire _abc_17692_n2357;
  wire _abc_17692_n2358;
  wire _abc_17692_n2359;
  wire _abc_17692_n2360;
  wire _abc_17692_n2361_1;
  wire _abc_17692_n2362;
  wire _abc_17692_n2363;
  wire _abc_17692_n2364;
  wire _abc_17692_n2365;
  wire _abc_17692_n2366;
  wire _abc_17692_n2367;
  wire _abc_17692_n2368;
  wire _abc_17692_n2369;
  wire _abc_17692_n2370;
  wire _abc_17692_n2371;
  wire _abc_17692_n2372;
  wire _abc_17692_n2373;
  wire _abc_17692_n2374;
  wire _abc_17692_n2375;
  wire _abc_17692_n2376;
  wire _abc_17692_n2377;
  wire _abc_17692_n2378;
  wire _abc_17692_n2379;
  wire _abc_17692_n2380_1;
  wire _abc_17692_n2381;
  wire _abc_17692_n2382;
  wire _abc_17692_n2383;
  wire _abc_17692_n2384;
  wire _abc_17692_n2385;
  wire _abc_17692_n2386;
  wire _abc_17692_n2387;
  wire _abc_17692_n2388;
  wire _abc_17692_n2389;
  wire _abc_17692_n2390;
  wire _abc_17692_n2391;
  wire _abc_17692_n2392;
  wire _abc_17692_n2393;
  wire _abc_17692_n2394;
  wire _abc_17692_n2395;
  wire _abc_17692_n2396;
  wire _abc_17692_n2397;
  wire _abc_17692_n2398;
  wire _abc_17692_n2399_1;
  wire _abc_17692_n2400;
  wire _abc_17692_n2401;
  wire _abc_17692_n2402;
  wire _abc_17692_n2403;
  wire _abc_17692_n2404;
  wire _abc_17692_n2405;
  wire _abc_17692_n2406;
  wire _abc_17692_n2407;
  wire _abc_17692_n2408;
  wire _abc_17692_n2409;
  wire _abc_17692_n2410;
  wire _abc_17692_n2411;
  wire _abc_17692_n2412;
  wire _abc_17692_n2413;
  wire _abc_17692_n2414;
  wire _abc_17692_n2415;
  wire _abc_17692_n2416;
  wire _abc_17692_n2417;
  wire _abc_17692_n2418;
  wire _abc_17692_n2419;
  wire _abc_17692_n2420;
  wire _abc_17692_n2421;
  wire _abc_17692_n2422;
  wire _abc_17692_n2423;
  wire _abc_17692_n2424;
  wire _abc_17692_n2425;
  wire _abc_17692_n2426;
  wire _abc_17692_n2427;
  wire _abc_17692_n2428;
  wire _abc_17692_n2429;
  wire _abc_17692_n2430;
  wire _abc_17692_n2431;
  wire _abc_17692_n2433;
  wire _abc_17692_n2434;
  wire _abc_17692_n2435;
  wire _abc_17692_n2436;
  wire _abc_17692_n2437;
  wire _abc_17692_n2438;
  wire _abc_17692_n2439;
  wire _abc_17692_n2440;
  wire _abc_17692_n2441;
  wire _abc_17692_n2442;
  wire _abc_17692_n2443;
  wire _abc_17692_n2444;
  wire _abc_17692_n2445;
  wire _abc_17692_n2446;
  wire _abc_17692_n2447;
  wire _abc_17692_n2448;
  wire _abc_17692_n2449;
  wire _abc_17692_n2450;
  wire _abc_17692_n2451;
  wire _abc_17692_n2452;
  wire _abc_17692_n2453;
  wire _abc_17692_n2454;
  wire _abc_17692_n2455;
  wire _abc_17692_n2456;
  wire _abc_17692_n2457;
  wire _abc_17692_n2458;
  wire _abc_17692_n2459_1;
  wire _abc_17692_n2460;
  wire _abc_17692_n2461;
  wire _abc_17692_n2462_1;
  wire _abc_17692_n2463;
  wire _abc_17692_n2464;
  wire _abc_17692_n2465;
  wire _abc_17692_n2466;
  wire _abc_17692_n2467;
  wire _abc_17692_n2468;
  wire _abc_17692_n2469_1;
  wire _abc_17692_n2470;
  wire _abc_17692_n2471;
  wire _abc_17692_n2472;
  wire _abc_17692_n2473;
  wire _abc_17692_n2474;
  wire _abc_17692_n2475;
  wire _abc_17692_n2476;
  wire _abc_17692_n2477;
  wire _abc_17692_n2478;
  wire _abc_17692_n2479_1;
  wire _abc_17692_n2480;
  wire _abc_17692_n2481;
  wire _abc_17692_n2482;
  wire _abc_17692_n2483;
  wire _abc_17692_n2484;
  wire _abc_17692_n2485;
  wire _abc_17692_n2486;
  wire _abc_17692_n2487;
  wire _abc_17692_n2488;
  wire _abc_17692_n2489;
  wire _abc_17692_n2490_1;
  wire _abc_17692_n2491;
  wire _abc_17692_n2492;
  wire _abc_17692_n2493;
  wire _abc_17692_n2494;
  wire _abc_17692_n2495;
  wire _abc_17692_n2496;
  wire _abc_17692_n2497;
  wire _abc_17692_n2498;
  wire _abc_17692_n2499;
  wire _abc_17692_n2500_1;
  wire _abc_17692_n2501;
  wire _abc_17692_n2502;
  wire _abc_17692_n2503;
  wire _abc_17692_n2504;
  wire _abc_17692_n2505;
  wire _abc_17692_n2506;
  wire _abc_17692_n2507;
  wire _abc_17692_n2508;
  wire _abc_17692_n2509;
  wire _abc_17692_n2510;
  wire _abc_17692_n2511;
  wire _abc_17692_n2512;
  wire _abc_17692_n2513;
  wire _abc_17692_n2514;
  wire _abc_17692_n2515;
  wire _abc_17692_n2516;
  wire _abc_17692_n2517;
  wire _abc_17692_n2518;
  wire _abc_17692_n2519;
  wire _abc_17692_n2520;
  wire _abc_17692_n2521;
  wire _abc_17692_n2522;
  wire _abc_17692_n2523;
  wire _abc_17692_n2524;
  wire _abc_17692_n2525;
  wire _abc_17692_n2526;
  wire _abc_17692_n2527;
  wire _abc_17692_n2528;
  wire _abc_17692_n2529;
  wire _abc_17692_n2530;
  wire _abc_17692_n2531;
  wire _abc_17692_n2532;
  wire _abc_17692_n2533;
  wire _abc_17692_n2534;
  wire _abc_17692_n2535_1;
  wire _abc_17692_n2536;
  wire _abc_17692_n2537;
  wire _abc_17692_n2538_1;
  wire _abc_17692_n2539;
  wire _abc_17692_n2540;
  wire _abc_17692_n2541;
  wire _abc_17692_n2542;
  wire _abc_17692_n2543;
  wire _abc_17692_n2544;
  wire _abc_17692_n2545;
  wire _abc_17692_n2546;
  wire _abc_17692_n2547;
  wire _abc_17692_n2548;
  wire _abc_17692_n2549;
  wire _abc_17692_n2550;
  wire _abc_17692_n2551;
  wire _abc_17692_n2552_1;
  wire _abc_17692_n2553;
  wire _abc_17692_n2554;
  wire _abc_17692_n2555;
  wire _abc_17692_n2556;
  wire _abc_17692_n2557;
  wire _abc_17692_n2558;
  wire _abc_17692_n2559;
  wire _abc_17692_n2560;
  wire _abc_17692_n2561;
  wire _abc_17692_n2562;
  wire _abc_17692_n2563;
  wire _abc_17692_n2564;
  wire _abc_17692_n2565;
  wire _abc_17692_n2566;
  wire _abc_17692_n2567;
  wire _abc_17692_n2568;
  wire _abc_17692_n2569;
  wire _abc_17692_n2570;
  wire _abc_17692_n2571;
  wire _abc_17692_n2572;
  wire _abc_17692_n2573;
  wire _abc_17692_n2574;
  wire _abc_17692_n2575;
  wire _abc_17692_n2576;
  wire _abc_17692_n2577;
  wire _abc_17692_n2578;
  wire _abc_17692_n2579;
  wire _abc_17692_n2580;
  wire _abc_17692_n2581_1;
  wire _abc_17692_n2582;
  wire _abc_17692_n2583;
  wire _abc_17692_n2584;
  wire _abc_17692_n2585;
  wire _abc_17692_n2586;
  wire _abc_17692_n2587;
  wire _abc_17692_n2588;
  wire _abc_17692_n2589;
  wire _abc_17692_n2590;
  wire _abc_17692_n2591;
  wire _abc_17692_n2592;
  wire _abc_17692_n2593;
  wire _abc_17692_n2594;
  wire _abc_17692_n2595;
  wire _abc_17692_n2596;
  wire _abc_17692_n2597;
  wire _abc_17692_n2598;
  wire _abc_17692_n2599;
  wire _abc_17692_n2600;
  wire _abc_17692_n2601;
  wire _abc_17692_n2602;
  wire _abc_17692_n2603;
  wire _abc_17692_n2604;
  wire _abc_17692_n2605;
  wire _abc_17692_n2606;
  wire _abc_17692_n2607;
  wire _abc_17692_n2608_1;
  wire _abc_17692_n2609;
  wire _abc_17692_n2610;
  wire _abc_17692_n2611;
  wire _abc_17692_n2612;
  wire _abc_17692_n2613;
  wire _abc_17692_n2614;
  wire _abc_17692_n2615;
  wire _abc_17692_n2616;
  wire _abc_17692_n2617;
  wire _abc_17692_n2618;
  wire _abc_17692_n2619;
  wire _abc_17692_n2620;
  wire _abc_17692_n2621;
  wire _abc_17692_n2622;
  wire _abc_17692_n2623;
  wire _abc_17692_n2624;
  wire _abc_17692_n2625;
  wire _abc_17692_n2626;
  wire _abc_17692_n2627;
  wire _abc_17692_n2628;
  wire _abc_17692_n2629;
  wire _abc_17692_n2630;
  wire _abc_17692_n2631;
  wire _abc_17692_n2633;
  wire _abc_17692_n2634_1;
  wire _abc_17692_n2635;
  wire _abc_17692_n2636;
  wire _abc_17692_n2637;
  wire _abc_17692_n2638;
  wire _abc_17692_n2639;
  wire _abc_17692_n2640;
  wire _abc_17692_n2641;
  wire _abc_17692_n2642;
  wire _abc_17692_n2643;
  wire _abc_17692_n2644;
  wire _abc_17692_n2645;
  wire _abc_17692_n2646;
  wire _abc_17692_n2647;
  wire _abc_17692_n2648;
  wire _abc_17692_n2649;
  wire _abc_17692_n2650;
  wire _abc_17692_n2651;
  wire _abc_17692_n2652;
  wire _abc_17692_n2653;
  wire _abc_17692_n2654;
  wire _abc_17692_n2655;
  wire _abc_17692_n2656;
  wire _abc_17692_n2657;
  wire _abc_17692_n2658;
  wire _abc_17692_n2659;
  wire _abc_17692_n2660;
  wire _abc_17692_n2661;
  wire _abc_17692_n2662;
  wire _abc_17692_n2663;
  wire _abc_17692_n2664;
  wire _abc_17692_n2665;
  wire _abc_17692_n2666;
  wire _abc_17692_n2667;
  wire _abc_17692_n2668;
  wire _abc_17692_n2669;
  wire _abc_17692_n2670;
  wire _abc_17692_n2671;
  wire _abc_17692_n2672;
  wire _abc_17692_n2673;
  wire _abc_17692_n2674;
  wire _abc_17692_n2675;
  wire _abc_17692_n2676;
  wire _abc_17692_n2677;
  wire _abc_17692_n2678;
  wire _abc_17692_n2679;
  wire _abc_17692_n2680;
  wire _abc_17692_n2681;
  wire _abc_17692_n2682;
  wire _abc_17692_n2683;
  wire _abc_17692_n2684;
  wire _abc_17692_n2685;
  wire _abc_17692_n2686;
  wire _abc_17692_n2687;
  wire _abc_17692_n2688;
  wire _abc_17692_n2689;
  wire _abc_17692_n2690;
  wire _abc_17692_n2691;
  wire _abc_17692_n2692;
  wire _abc_17692_n2693;
  wire _abc_17692_n2694;
  wire _abc_17692_n2695;
  wire _abc_17692_n2696;
  wire _abc_17692_n2697;
  wire _abc_17692_n2698;
  wire _abc_17692_n2699;
  wire _abc_17692_n2700;
  wire _abc_17692_n2701;
  wire _abc_17692_n2702;
  wire _abc_17692_n2703;
  wire _abc_17692_n2704;
  wire _abc_17692_n2705;
  wire _abc_17692_n2706;
  wire _abc_17692_n2707;
  wire _abc_17692_n2708;
  wire _abc_17692_n2709;
  wire _abc_17692_n2710;
  wire _abc_17692_n2711;
  wire _abc_17692_n2712;
  wire _abc_17692_n2713_1;
  wire _abc_17692_n2714;
  wire _abc_17692_n2715;
  wire _abc_17692_n2716_1;
  wire _abc_17692_n2717;
  wire _abc_17692_n2718;
  wire _abc_17692_n2719;
  wire _abc_17692_n2720;
  wire _abc_17692_n2721;
  wire _abc_17692_n2722;
  wire _abc_17692_n2723_1;
  wire _abc_17692_n2724;
  wire _abc_17692_n2725;
  wire _abc_17692_n2726;
  wire _abc_17692_n2727;
  wire _abc_17692_n2728;
  wire _abc_17692_n2729;
  wire _abc_17692_n2730;
  wire _abc_17692_n2731;
  wire _abc_17692_n2732;
  wire _abc_17692_n2733;
  wire _abc_17692_n2734_1;
  wire _abc_17692_n2735;
  wire _abc_17692_n2736;
  wire _abc_17692_n2737;
  wire _abc_17692_n2738;
  wire _abc_17692_n2739;
  wire _abc_17692_n2740;
  wire _abc_17692_n2741;
  wire _abc_17692_n2742;
  wire _abc_17692_n2743;
  wire _abc_17692_n2744;
  wire _abc_17692_n2745_1;
  wire _abc_17692_n2746;
  wire _abc_17692_n2747;
  wire _abc_17692_n2748;
  wire _abc_17692_n2749;
  wire _abc_17692_n2750;
  wire _abc_17692_n2751;
  wire _abc_17692_n2752;
  wire _abc_17692_n2753;
  wire _abc_17692_n2754;
  wire _abc_17692_n2755;
  wire _abc_17692_n2756;
  wire _abc_17692_n2757_1;
  wire _abc_17692_n2758;
  wire _abc_17692_n2759;
  wire _abc_17692_n2760;
  wire _abc_17692_n2761;
  wire _abc_17692_n2762;
  wire _abc_17692_n2763;
  wire _abc_17692_n2764;
  wire _abc_17692_n2765;
  wire _abc_17692_n2766;
  wire _abc_17692_n2767;
  wire _abc_17692_n2768;
  wire _abc_17692_n2769;
  wire _abc_17692_n2770;
  wire _abc_17692_n2771;
  wire _abc_17692_n2772;
  wire _abc_17692_n2773;
  wire _abc_17692_n2774;
  wire _abc_17692_n2775;
  wire _abc_17692_n2776;
  wire _abc_17692_n2777;
  wire _abc_17692_n2778;
  wire _abc_17692_n2779;
  wire _abc_17692_n2780;
  wire _abc_17692_n2781;
  wire _abc_17692_n2782;
  wire _abc_17692_n2783;
  wire _abc_17692_n2784;
  wire _abc_17692_n2785;
  wire _abc_17692_n2786;
  wire _abc_17692_n2787;
  wire _abc_17692_n2788;
  wire _abc_17692_n2789;
  wire _abc_17692_n2790;
  wire _abc_17692_n2791;
  wire _abc_17692_n2792;
  wire _abc_17692_n2793;
  wire _abc_17692_n2794;
  wire _abc_17692_n2795;
  wire _abc_17692_n2796;
  wire _abc_17692_n2797_1;
  wire _abc_17692_n2798;
  wire _abc_17692_n2799;
  wire _abc_17692_n2800_1;
  wire _abc_17692_n2801;
  wire _abc_17692_n2802;
  wire _abc_17692_n2803;
  wire _abc_17692_n2804;
  wire _abc_17692_n2805;
  wire _abc_17692_n2806;
  wire _abc_17692_n2807;
  wire _abc_17692_n2808;
  wire _abc_17692_n2809;
  wire _abc_17692_n2810;
  wire _abc_17692_n2811;
  wire _abc_17692_n2812_1;
  wire _abc_17692_n2813;
  wire _abc_17692_n2814;
  wire _abc_17692_n2816;
  wire _abc_17692_n2817;
  wire _abc_17692_n2818;
  wire _abc_17692_n2819;
  wire _abc_17692_n2820;
  wire _abc_17692_n2821;
  wire _abc_17692_n2822;
  wire _abc_17692_n2823;
  wire _abc_17692_n2824;
  wire _abc_17692_n2825;
  wire _abc_17692_n2826;
  wire _abc_17692_n2827;
  wire _abc_17692_n2828;
  wire _abc_17692_n2829;
  wire _abc_17692_n2830_1;
  wire _abc_17692_n2831;
  wire _abc_17692_n2832;
  wire _abc_17692_n2833;
  wire _abc_17692_n2834;
  wire _abc_17692_n2835;
  wire _abc_17692_n2836;
  wire _abc_17692_n2837;
  wire _abc_17692_n2838;
  wire _abc_17692_n2839;
  wire _abc_17692_n2840;
  wire _abc_17692_n2841;
  wire _abc_17692_n2842;
  wire _abc_17692_n2843;
  wire _abc_17692_n2844;
  wire _abc_17692_n2845;
  wire _abc_17692_n2846;
  wire _abc_17692_n2847;
  wire _abc_17692_n2848;
  wire _abc_17692_n2849_1;
  wire _abc_17692_n2850;
  wire _abc_17692_n2851;
  wire _abc_17692_n2852;
  wire _abc_17692_n2853;
  wire _abc_17692_n2854;
  wire _abc_17692_n2855;
  wire _abc_17692_n2856;
  wire _abc_17692_n2857;
  wire _abc_17692_n2858;
  wire _abc_17692_n2859;
  wire _abc_17692_n2860;
  wire _abc_17692_n2861;
  wire _abc_17692_n2862;
  wire _abc_17692_n2863;
  wire _abc_17692_n2864;
  wire _abc_17692_n2865;
  wire _abc_17692_n2866;
  wire _abc_17692_n2867_1;
  wire _abc_17692_n2868;
  wire _abc_17692_n2869;
  wire _abc_17692_n2870;
  wire _abc_17692_n2871;
  wire _abc_17692_n2872;
  wire _abc_17692_n2873;
  wire _abc_17692_n2874;
  wire _abc_17692_n2875;
  wire _abc_17692_n2876;
  wire _abc_17692_n2877;
  wire _abc_17692_n2878;
  wire _abc_17692_n2879;
  wire _abc_17692_n2880;
  wire _abc_17692_n2881;
  wire _abc_17692_n2882;
  wire _abc_17692_n2883;
  wire _abc_17692_n2884;
  wire _abc_17692_n2885;
  wire _abc_17692_n2886;
  wire _abc_17692_n2887;
  wire _abc_17692_n2888;
  wire _abc_17692_n2889;
  wire _abc_17692_n2890;
  wire _abc_17692_n2891;
  wire _abc_17692_n2892;
  wire _abc_17692_n2893;
  wire _abc_17692_n2894;
  wire _abc_17692_n2895;
  wire _abc_17692_n2896;
  wire _abc_17692_n2897;
  wire _abc_17692_n2898;
  wire _abc_17692_n2899;
  wire _abc_17692_n2900;
  wire _abc_17692_n2901;
  wire _abc_17692_n2902;
  wire _abc_17692_n2903;
  wire _abc_17692_n2904;
  wire _abc_17692_n2905;
  wire _abc_17692_n2906;
  wire _abc_17692_n2907;
  wire _abc_17692_n2908;
  wire _abc_17692_n2909;
  wire _abc_17692_n2910;
  wire _abc_17692_n2911;
  wire _abc_17692_n2912;
  wire _abc_17692_n2913;
  wire _abc_17692_n2914;
  wire _abc_17692_n2915;
  wire _abc_17692_n2916_1;
  wire _abc_17692_n2917;
  wire _abc_17692_n2918;
  wire _abc_17692_n2919_1;
  wire _abc_17692_n2920;
  wire _abc_17692_n2921;
  wire _abc_17692_n2922;
  wire _abc_17692_n2923;
  wire _abc_17692_n2924;
  wire _abc_17692_n2925;
  wire _abc_17692_n2926_1;
  wire _abc_17692_n2927;
  wire _abc_17692_n2928;
  wire _abc_17692_n2929;
  wire _abc_17692_n2930;
  wire _abc_17692_n2931;
  wire _abc_17692_n2932;
  wire _abc_17692_n2933;
  wire _abc_17692_n2934;
  wire _abc_17692_n2935;
  wire _abc_17692_n2936;
  wire _abc_17692_n2937;
  wire _abc_17692_n2938_1;
  wire _abc_17692_n2939;
  wire _abc_17692_n2940;
  wire _abc_17692_n2941;
  wire _abc_17692_n2942;
  wire _abc_17692_n2943;
  wire _abc_17692_n2944;
  wire _abc_17692_n2945;
  wire _abc_17692_n2946;
  wire _abc_17692_n2947;
  wire _abc_17692_n2948;
  wire _abc_17692_n2949_1;
  wire _abc_17692_n2950;
  wire _abc_17692_n2951;
  wire _abc_17692_n2952;
  wire _abc_17692_n2953;
  wire _abc_17692_n2954;
  wire _abc_17692_n2955;
  wire _abc_17692_n2956;
  wire _abc_17692_n2957;
  wire _abc_17692_n2958;
  wire _abc_17692_n2959;
  wire _abc_17692_n2960_1;
  wire _abc_17692_n2961;
  wire _abc_17692_n2962;
  wire _abc_17692_n2963;
  wire _abc_17692_n2964;
  wire _abc_17692_n2965;
  wire _abc_17692_n2966;
  wire _abc_17692_n2967;
  wire _abc_17692_n2968;
  wire _abc_17692_n2969;
  wire _abc_17692_n2970;
  wire _abc_17692_n2971;
  wire _abc_17692_n2972;
  wire _abc_17692_n2973;
  wire _abc_17692_n2974;
  wire _abc_17692_n2975;
  wire _abc_17692_n2976;
  wire _abc_17692_n2977;
  wire _abc_17692_n2978;
  wire _abc_17692_n2979;
  wire _abc_17692_n2980;
  wire _abc_17692_n2981;
  wire _abc_17692_n2982;
  wire _abc_17692_n2983;
  wire _abc_17692_n2984;
  wire _abc_17692_n2985;
  wire _abc_17692_n2986;
  wire _abc_17692_n2987;
  wire _abc_17692_n2988;
  wire _abc_17692_n2989;
  wire _abc_17692_n2990;
  wire _abc_17692_n2991;
  wire _abc_17692_n2992;
  wire _abc_17692_n2993;
  wire _abc_17692_n2994;
  wire _abc_17692_n2995_1;
  wire _abc_17692_n2996;
  wire _abc_17692_n2997;
  wire _abc_17692_n2998_1;
  wire _abc_17692_n2999;
  wire _abc_17692_n3000;
  wire _abc_17692_n3001;
  wire _abc_17692_n3002;
  wire _abc_17692_n3003;
  wire _abc_17692_n3004;
  wire _abc_17692_n3005;
  wire _abc_17692_n3006;
  wire _abc_17692_n3007;
  wire _abc_17692_n3008;
  wire _abc_17692_n3009_1;
  wire _abc_17692_n3010;
  wire _abc_17692_n3011;
  wire _abc_17692_n3012;
  wire _abc_17692_n3013;
  wire _abc_17692_n3014;
  wire _abc_17692_n3015;
  wire _abc_17692_n3016;
  wire _abc_17692_n3017;
  wire _abc_17692_n3018;
  wire _abc_17692_n3019;
  wire _abc_17692_n3020;
  wire _abc_17692_n3021;
  wire _abc_17692_n3023;
  wire _abc_17692_n3024;
  wire _abc_17692_n3025;
  wire _abc_17692_n3026;
  wire _abc_17692_n3027;
  wire _abc_17692_n3028;
  wire _abc_17692_n3029;
  wire _abc_17692_n3030;
  wire _abc_17692_n3031;
  wire _abc_17692_n3032;
  wire _abc_17692_n3033;
  wire _abc_17692_n3034_1;
  wire _abc_17692_n3035;
  wire _abc_17692_n3036;
  wire _abc_17692_n3037;
  wire _abc_17692_n3038;
  wire _abc_17692_n3039;
  wire _abc_17692_n3040;
  wire _abc_17692_n3041;
  wire _abc_17692_n3042;
  wire _abc_17692_n3043;
  wire _abc_17692_n3044;
  wire _abc_17692_n3045;
  wire _abc_17692_n3046;
  wire _abc_17692_n3047;
  wire _abc_17692_n3048;
  wire _abc_17692_n3049;
  wire _abc_17692_n3050;
  wire _abc_17692_n3051;
  wire _abc_17692_n3052;
  wire _abc_17692_n3053;
  wire _abc_17692_n3054;
  wire _abc_17692_n3055;
  wire _abc_17692_n3056;
  wire _abc_17692_n3057;
  wire _abc_17692_n3058_1;
  wire _abc_17692_n3059;
  wire _abc_17692_n3060;
  wire _abc_17692_n3061;
  wire _abc_17692_n3062;
  wire _abc_17692_n3063;
  wire _abc_17692_n3064;
  wire _abc_17692_n3065;
  wire _abc_17692_n3066;
  wire _abc_17692_n3067;
  wire _abc_17692_n3068;
  wire _abc_17692_n3069;
  wire _abc_17692_n3070;
  wire _abc_17692_n3071;
  wire _abc_17692_n3072;
  wire _abc_17692_n3073;
  wire _abc_17692_n3074;
  wire _abc_17692_n3075;
  wire _abc_17692_n3076;
  wire _abc_17692_n3077;
  wire _abc_17692_n3078;
  wire _abc_17692_n3079;
  wire _abc_17692_n3080_1;
  wire _abc_17692_n3081;
  wire _abc_17692_n3082;
  wire _abc_17692_n3083;
  wire _abc_17692_n3084;
  wire _abc_17692_n3085;
  wire _abc_17692_n3086;
  wire _abc_17692_n3087;
  wire _abc_17692_n3088;
  wire _abc_17692_n3089;
  wire _abc_17692_n3090;
  wire _abc_17692_n3091;
  wire _abc_17692_n3092;
  wire _abc_17692_n3093;
  wire _abc_17692_n3094;
  wire _abc_17692_n3095;
  wire _abc_17692_n3096;
  wire _abc_17692_n3097;
  wire _abc_17692_n3098;
  wire _abc_17692_n3099;
  wire _abc_17692_n3100;
  wire _abc_17692_n3101;
  wire _abc_17692_n3102;
  wire _abc_17692_n3103;
  wire _abc_17692_n3104;
  wire _abc_17692_n3105;
  wire _abc_17692_n3106;
  wire _abc_17692_n3107;
  wire _abc_17692_n3108;
  wire _abc_17692_n3109;
  wire _abc_17692_n3110;
  wire _abc_17692_n3111;
  wire _abc_17692_n3112;
  wire _abc_17692_n3113;
  wire _abc_17692_n3114;
  wire _abc_17692_n3115;
  wire _abc_17692_n3116;
  wire _abc_17692_n3117;
  wire _abc_17692_n3118;
  wire _abc_17692_n3119;
  wire _abc_17692_n3120;
  wire _abc_17692_n3121;
  wire _abc_17692_n3122;
  wire _abc_17692_n3123;
  wire _abc_17692_n3124;
  wire _abc_17692_n3125;
  wire _abc_17692_n3126;
  wire _abc_17692_n3127;
  wire _abc_17692_n3128;
  wire _abc_17692_n3129;
  wire _abc_17692_n3130;
  wire _abc_17692_n3131;
  wire _abc_17692_n3132;
  wire _abc_17692_n3133;
  wire _abc_17692_n3134;
  wire _abc_17692_n3135;
  wire _abc_17692_n3136;
  wire _abc_17692_n3137;
  wire _abc_17692_n3138;
  wire _abc_17692_n3139;
  wire _abc_17692_n3140;
  wire _abc_17692_n3141_1;
  wire _abc_17692_n3142;
  wire _abc_17692_n3143;
  wire _abc_17692_n3144_1;
  wire _abc_17692_n3145;
  wire _abc_17692_n3146;
  wire _abc_17692_n3147;
  wire _abc_17692_n3148;
  wire _abc_17692_n3149;
  wire _abc_17692_n3150;
  wire _abc_17692_n3151;
  wire _abc_17692_n3152;
  wire _abc_17692_n3153_1;
  wire _abc_17692_n3154;
  wire _abc_17692_n3155;
  wire _abc_17692_n3156;
  wire _abc_17692_n3157;
  wire _abc_17692_n3158;
  wire _abc_17692_n3159;
  wire _abc_17692_n3160;
  wire _abc_17692_n3161;
  wire _abc_17692_n3162;
  wire _abc_17692_n3163;
  wire _abc_17692_n3164;
  wire _abc_17692_n3165;
  wire _abc_17692_n3166_1;
  wire _abc_17692_n3167;
  wire _abc_17692_n3168;
  wire _abc_17692_n3169;
  wire _abc_17692_n3170;
  wire _abc_17692_n3171;
  wire _abc_17692_n3172;
  wire _abc_17692_n3173;
  wire _abc_17692_n3174;
  wire _abc_17692_n3175;
  wire _abc_17692_n3176;
  wire _abc_17692_n3177;
  wire _abc_17692_n3178_1;
  wire _abc_17692_n3179;
  wire _abc_17692_n3180;
  wire _abc_17692_n3181;
  wire _abc_17692_n3182;
  wire _abc_17692_n3183;
  wire _abc_17692_n3184;
  wire _abc_17692_n3185;
  wire _abc_17692_n3186;
  wire _abc_17692_n3187;
  wire _abc_17692_n3188;
  wire _abc_17692_n3189_1;
  wire _abc_17692_n3190;
  wire _abc_17692_n3191;
  wire _abc_17692_n3192;
  wire _abc_17692_n3193;
  wire _abc_17692_n3194;
  wire _abc_17692_n3195;
  wire _abc_17692_n3196;
  wire _abc_17692_n3198;
  wire _abc_17692_n3199;
  wire _abc_17692_n3200;
  wire _abc_17692_n3201;
  wire _abc_17692_n3202;
  wire _abc_17692_n3203;
  wire _abc_17692_n3204;
  wire _abc_17692_n3205;
  wire _abc_17692_n3206;
  wire _abc_17692_n3207;
  wire _abc_17692_n3208;
  wire _abc_17692_n3209;
  wire _abc_17692_n3210;
  wire _abc_17692_n3211;
  wire _abc_17692_n3212;
  wire _abc_17692_n3213;
  wire _abc_17692_n3214;
  wire _abc_17692_n3215;
  wire _abc_17692_n3216;
  wire _abc_17692_n3217;
  wire _abc_17692_n3218;
  wire _abc_17692_n3219;
  wire _abc_17692_n3220;
  wire _abc_17692_n3221;
  wire _abc_17692_n3222;
  wire _abc_17692_n3223;
  wire _abc_17692_n3224_1;
  wire _abc_17692_n3225;
  wire _abc_17692_n3226;
  wire _abc_17692_n3227_1;
  wire _abc_17692_n3228;
  wire _abc_17692_n3229;
  wire _abc_17692_n3230;
  wire _abc_17692_n3231;
  wire _abc_17692_n3232;
  wire _abc_17692_n3233;
  wire _abc_17692_n3234;
  wire _abc_17692_n3235;
  wire _abc_17692_n3236;
  wire _abc_17692_n3237;
  wire _abc_17692_n3238;
  wire _abc_17692_n3239;
  wire _abc_17692_n3240_1;
  wire _abc_17692_n3241;
  wire _abc_17692_n3242;
  wire _abc_17692_n3243;
  wire _abc_17692_n3244;
  wire _abc_17692_n3245;
  wire _abc_17692_n3246;
  wire _abc_17692_n3247;
  wire _abc_17692_n3248;
  wire _abc_17692_n3249;
  wire _abc_17692_n3250;
  wire _abc_17692_n3251;
  wire _abc_17692_n3252;
  wire _abc_17692_n3253;
  wire _abc_17692_n3254;
  wire _abc_17692_n3255;
  wire _abc_17692_n3256;
  wire _abc_17692_n3257;
  wire _abc_17692_n3258_1;
  wire _abc_17692_n3259;
  wire _abc_17692_n3260;
  wire _abc_17692_n3261;
  wire _abc_17692_n3262;
  wire _abc_17692_n3263;
  wire _abc_17692_n3264;
  wire _abc_17692_n3265;
  wire _abc_17692_n3266;
  wire _abc_17692_n3267;
  wire _abc_17692_n3268;
  wire _abc_17692_n3269;
  wire _abc_17692_n3270;
  wire _abc_17692_n3271;
  wire _abc_17692_n3272;
  wire _abc_17692_n3273;
  wire _abc_17692_n3274;
  wire _abc_17692_n3275;
  wire _abc_17692_n3276;
  wire _abc_17692_n3277;
  wire _abc_17692_n3278_1;
  wire _abc_17692_n3279;
  wire _abc_17692_n3280;
  wire _abc_17692_n3281;
  wire _abc_17692_n3282;
  wire _abc_17692_n3283;
  wire _abc_17692_n3284;
  wire _abc_17692_n3285;
  wire _abc_17692_n3286;
  wire _abc_17692_n3287;
  wire _abc_17692_n3288;
  wire _abc_17692_n3289;
  wire _abc_17692_n3290;
  wire _abc_17692_n3291;
  wire _abc_17692_n3292;
  wire _abc_17692_n3293;
  wire _abc_17692_n3294;
  wire _abc_17692_n3295_1;
  wire _abc_17692_n3296;
  wire _abc_17692_n3297;
  wire _abc_17692_n3298;
  wire _abc_17692_n3299;
  wire _abc_17692_n3300;
  wire _abc_17692_n3301;
  wire _abc_17692_n3302;
  wire _abc_17692_n3303;
  wire _abc_17692_n3304;
  wire _abc_17692_n3305;
  wire _abc_17692_n3306;
  wire _abc_17692_n3307;
  wire _abc_17692_n3308;
  wire _abc_17692_n3309;
  wire _abc_17692_n3310;
  wire _abc_17692_n3311;
  wire _abc_17692_n3312;
  wire _abc_17692_n3313;
  wire _abc_17692_n3314;
  wire _abc_17692_n3315;
  wire _abc_17692_n3316;
  wire _abc_17692_n3317;
  wire _abc_17692_n3318;
  wire _abc_17692_n3319;
  wire _abc_17692_n3320;
  wire _abc_17692_n3321;
  wire _abc_17692_n3322;
  wire _abc_17692_n3323;
  wire _abc_17692_n3324;
  wire _abc_17692_n3325;
  wire _abc_17692_n3326;
  wire _abc_17692_n3327;
  wire _abc_17692_n3328;
  wire _abc_17692_n3329;
  wire _abc_17692_n3330;
  wire _abc_17692_n3331;
  wire _abc_17692_n3332;
  wire _abc_17692_n3333;
  wire _abc_17692_n3334;
  wire _abc_17692_n3335;
  wire _abc_17692_n3336;
  wire _abc_17692_n3337;
  wire _abc_17692_n3338;
  wire _abc_17692_n3339;
  wire _abc_17692_n3340;
  wire _abc_17692_n3341;
  wire _abc_17692_n3342;
  wire _abc_17692_n3343;
  wire _abc_17692_n3344;
  wire _abc_17692_n3345;
  wire _abc_17692_n3346_1;
  wire _abc_17692_n3347;
  wire _abc_17692_n3348;
  wire _abc_17692_n3349_1;
  wire _abc_17692_n3350;
  wire _abc_17692_n3351;
  wire _abc_17692_n3352;
  wire _abc_17692_n3353;
  wire _abc_17692_n3354;
  wire _abc_17692_n3355_1;
  wire _abc_17692_n3356;
  wire _abc_17692_n3357;
  wire _abc_17692_n3358;
  wire _abc_17692_n3359;
  wire _abc_17692_n3360;
  wire _abc_17692_n3361;
  wire _abc_17692_n3362;
  wire _abc_17692_n3363;
  wire _abc_17692_n3364;
  wire _abc_17692_n3365;
  wire _abc_17692_n3366_1;
  wire _abc_17692_n3367;
  wire _abc_17692_n3368;
  wire _abc_17692_n3369;
  wire _abc_17692_n3370;
  wire _abc_17692_n3371;
  wire _abc_17692_n3372;
  wire _abc_17692_n3373;
  wire _abc_17692_n3374;
  wire _abc_17692_n3375;
  wire _abc_17692_n3376_1;
  wire _abc_17692_n3377;
  wire _abc_17692_n3378;
  wire _abc_17692_n3379;
  wire _abc_17692_n3380;
  wire _abc_17692_n3381;
  wire _abc_17692_n3382;
  wire _abc_17692_n3383;
  wire _abc_17692_n3384;
  wire _abc_17692_n3385;
  wire _abc_17692_n3386;
  wire _abc_17692_n3387;
  wire _abc_17692_n3388_1;
  wire _abc_17692_n3389;
  wire _abc_17692_n3390;
  wire _abc_17692_n3391;
  wire _abc_17692_n3392;
  wire _abc_17692_n3393;
  wire _abc_17692_n3394;
  wire _abc_17692_n3395;
  wire _abc_17692_n3396;
  wire _abc_17692_n3397;
  wire _abc_17692_n3398;
  wire _abc_17692_n3399;
  wire _abc_17692_n3400;
  wire _abc_17692_n3401;
  wire _abc_17692_n3402;
  wire _abc_17692_n3403;
  wire _abc_17692_n3404;
  wire _abc_17692_n3405;
  wire _abc_17692_n3406;
  wire _abc_17692_n3407;
  wire _abc_17692_n3408;
  wire _abc_17692_n3409;
  wire _abc_17692_n3410;
  wire _abc_17692_n3411;
  wire _abc_17692_n3412;
  wire _abc_17692_n3413;
  wire _abc_17692_n3414;
  wire _abc_17692_n3415;
  wire _abc_17692_n3416;
  wire _abc_17692_n3417;
  wire _abc_17692_n3418;
  wire _abc_17692_n3419;
  wire _abc_17692_n3420;
  wire _abc_17692_n3421;
  wire _abc_17692_n3422;
  wire _abc_17692_n3423;
  wire _abc_17692_n3424_1;
  wire _abc_17692_n3425;
  wire _abc_17692_n3426;
  wire _abc_17692_n3427_1;
  wire _abc_17692_n3428;
  wire _abc_17692_n3429;
  wire _abc_17692_n3430;
  wire _abc_17692_n3431;
  wire _abc_17692_n3432;
  wire _abc_17692_n3433;
  wire _abc_17692_n3434;
  wire _abc_17692_n3435;
  wire _abc_17692_n3437;
  wire _abc_17692_n3438;
  wire _abc_17692_n3439;
  wire _abc_17692_n3440;
  wire _abc_17692_n3441;
  wire _abc_17692_n3442;
  wire _abc_17692_n3443;
  wire _abc_17692_n3444_1;
  wire _abc_17692_n3445;
  wire _abc_17692_n3446;
  wire _abc_17692_n3447;
  wire _abc_17692_n3448;
  wire _abc_17692_n3449;
  wire _abc_17692_n3450;
  wire _abc_17692_n3451;
  wire _abc_17692_n3452;
  wire _abc_17692_n3453;
  wire _abc_17692_n3454;
  wire _abc_17692_n3455;
  wire _abc_17692_n3456;
  wire _abc_17692_n3457;
  wire _abc_17692_n3458;
  wire _abc_17692_n3459;
  wire _abc_17692_n3460;
  wire _abc_17692_n3461;
  wire _abc_17692_n3462;
  wire _abc_17692_n3463;
  wire _abc_17692_n3464;
  wire _abc_17692_n3465;
  wire _abc_17692_n3466;
  wire _abc_17692_n3467;
  wire _abc_17692_n3468;
  wire _abc_17692_n3469;
  wire _abc_17692_n3470;
  wire _abc_17692_n3471;
  wire _abc_17692_n3472_1;
  wire _abc_17692_n3473;
  wire _abc_17692_n3474;
  wire _abc_17692_n3475;
  wire _abc_17692_n3476;
  wire _abc_17692_n3477;
  wire _abc_17692_n3478;
  wire _abc_17692_n3479;
  wire _abc_17692_n3480;
  wire _abc_17692_n3481;
  wire _abc_17692_n3482;
  wire _abc_17692_n3483;
  wire _abc_17692_n3484;
  wire _abc_17692_n3485;
  wire _abc_17692_n3486;
  wire _abc_17692_n3487;
  wire _abc_17692_n3488;
  wire _abc_17692_n3489;
  wire _abc_17692_n3490;
  wire _abc_17692_n3491;
  wire _abc_17692_n3492;
  wire _abc_17692_n3493;
  wire _abc_17692_n3494;
  wire _abc_17692_n3495;
  wire _abc_17692_n3496;
  wire _abc_17692_n3497;
  wire _abc_17692_n3498;
  wire _abc_17692_n3499;
  wire _abc_17692_n3500;
  wire _abc_17692_n3501;
  wire _abc_17692_n3502;
  wire _abc_17692_n3503_1;
  wire _abc_17692_n3504;
  wire _abc_17692_n3505;
  wire _abc_17692_n3506;
  wire _abc_17692_n3507;
  wire _abc_17692_n3508;
  wire _abc_17692_n3509;
  wire _abc_17692_n3510;
  wire _abc_17692_n3511;
  wire _abc_17692_n3512;
  wire _abc_17692_n3513;
  wire _abc_17692_n3514;
  wire _abc_17692_n3515;
  wire _abc_17692_n3516;
  wire _abc_17692_n3517;
  wire _abc_17692_n3518;
  wire _abc_17692_n3519;
  wire _abc_17692_n3520;
  wire _abc_17692_n3521;
  wire _abc_17692_n3522;
  wire _abc_17692_n3523;
  wire _abc_17692_n3524;
  wire _abc_17692_n3525;
  wire _abc_17692_n3526;
  wire _abc_17692_n3527;
  wire _abc_17692_n3528;
  wire _abc_17692_n3529;
  wire _abc_17692_n3530;
  wire _abc_17692_n3531;
  wire _abc_17692_n3532;
  wire _abc_17692_n3533_1;
  wire _abc_17692_n3534;
  wire _abc_17692_n3535;
  wire _abc_17692_n3536;
  wire _abc_17692_n3537;
  wire _abc_17692_n3538;
  wire _abc_17692_n3539;
  wire _abc_17692_n3540;
  wire _abc_17692_n3541;
  wire _abc_17692_n3542;
  wire _abc_17692_n3543;
  wire _abc_17692_n3544;
  wire _abc_17692_n3545;
  wire _abc_17692_n3546;
  wire _abc_17692_n3547;
  wire _abc_17692_n3548;
  wire _abc_17692_n3549;
  wire _abc_17692_n3550;
  wire _abc_17692_n3551;
  wire _abc_17692_n3552;
  wire _abc_17692_n3553;
  wire _abc_17692_n3554;
  wire _abc_17692_n3555;
  wire _abc_17692_n3556;
  wire _abc_17692_n3557;
  wire _abc_17692_n3558;
  wire _abc_17692_n3559;
  wire _abc_17692_n3560;
  wire _abc_17692_n3561;
  wire _abc_17692_n3562;
  wire _abc_17692_n3563;
  wire _abc_17692_n3564;
  wire _abc_17692_n3565;
  wire _abc_17692_n3566;
  wire _abc_17692_n3567;
  wire _abc_17692_n3568;
  wire _abc_17692_n3569;
  wire _abc_17692_n3570;
  wire _abc_17692_n3571;
  wire _abc_17692_n3572;
  wire _abc_17692_n3573;
  wire _abc_17692_n3574;
  wire _abc_17692_n3575;
  wire _abc_17692_n3576;
  wire _abc_17692_n3577;
  wire _abc_17692_n3578;
  wire _abc_17692_n3579;
  wire _abc_17692_n3580;
  wire _abc_17692_n3581;
  wire _abc_17692_n3582;
  wire _abc_17692_n3583;
  wire _abc_17692_n3584;
  wire _abc_17692_n3585;
  wire _abc_17692_n3586;
  wire _abc_17692_n3587;
  wire _abc_17692_n3588;
  wire _abc_17692_n3589;
  wire _abc_17692_n3590;
  wire _abc_17692_n3591;
  wire _abc_17692_n3592;
  wire _abc_17692_n3593;
  wire _abc_17692_n3594;
  wire _abc_17692_n3595;
  wire _abc_17692_n3596;
  wire _abc_17692_n3597;
  wire _abc_17692_n3598;
  wire _abc_17692_n3599;
  wire _abc_17692_n3600;
  wire _abc_17692_n3601;
  wire _abc_17692_n3602;
  wire _abc_17692_n3603;
  wire _abc_17692_n3604;
  wire _abc_17692_n3606;
  wire _abc_17692_n3607;
  wire _abc_17692_n3608;
  wire _abc_17692_n3609;
  wire _abc_17692_n3610;
  wire _abc_17692_n3611;
  wire _abc_17692_n3612;
  wire _abc_17692_n3613;
  wire _abc_17692_n3614;
  wire _abc_17692_n3615;
  wire _abc_17692_n3616;
  wire _abc_17692_n3617;
  wire _abc_17692_n3618_1;
  wire _abc_17692_n3619;
  wire _abc_17692_n3620;
  wire _abc_17692_n3621_1;
  wire _abc_17692_n3622;
  wire _abc_17692_n3623;
  wire _abc_17692_n3624;
  wire _abc_17692_n3625;
  wire _abc_17692_n3626;
  wire _abc_17692_n3627;
  wire _abc_17692_n3628;
  wire _abc_17692_n3629;
  wire _abc_17692_n3630_1;
  wire _abc_17692_n3631;
  wire _abc_17692_n3632;
  wire _abc_17692_n3633;
  wire _abc_17692_n3634;
  wire _abc_17692_n3635;
  wire _abc_17692_n3636;
  wire _abc_17692_n3637;
  wire _abc_17692_n3638;
  wire _abc_17692_n3639;
  wire _abc_17692_n3640_1;
  wire _abc_17692_n3641;
  wire _abc_17692_n3642;
  wire _abc_17692_n3643;
  wire _abc_17692_n3644;
  wire _abc_17692_n3645;
  wire _abc_17692_n3646;
  wire _abc_17692_n3647;
  wire _abc_17692_n3648;
  wire _abc_17692_n3649;
  wire _abc_17692_n3650_1;
  wire _abc_17692_n3651;
  wire _abc_17692_n3652;
  wire _abc_17692_n3653;
  wire _abc_17692_n3654;
  wire _abc_17692_n3655;
  wire _abc_17692_n3656;
  wire _abc_17692_n3657;
  wire _abc_17692_n3658;
  wire _abc_17692_n3659;
  wire _abc_17692_n3660;
  wire _abc_17692_n3661_1;
  wire _abc_17692_n3662;
  wire _abc_17692_n3663;
  wire _abc_17692_n3664;
  wire _abc_17692_n3665;
  wire _abc_17692_n3666;
  wire _abc_17692_n3667;
  wire _abc_17692_n3668;
  wire _abc_17692_n3669;
  wire _abc_17692_n3670;
  wire _abc_17692_n3671;
  wire _abc_17692_n3672;
  wire _abc_17692_n3673;
  wire _abc_17692_n3674;
  wire _abc_17692_n3675;
  wire _abc_17692_n3676;
  wire _abc_17692_n3677;
  wire _abc_17692_n3678;
  wire _abc_17692_n3679;
  wire _abc_17692_n3680;
  wire _abc_17692_n3681;
  wire _abc_17692_n3682;
  wire _abc_17692_n3683;
  wire _abc_17692_n3684;
  wire _abc_17692_n3685;
  wire _abc_17692_n3686;
  wire _abc_17692_n3687;
  wire _abc_17692_n3688;
  wire _abc_17692_n3689;
  wire _abc_17692_n3690;
  wire _abc_17692_n3691;
  wire _abc_17692_n3692;
  wire _abc_17692_n3693;
  wire _abc_17692_n3694;
  wire _abc_17692_n3695;
  wire _abc_17692_n3696_1;
  wire _abc_17692_n3697;
  wire _abc_17692_n3698;
  wire _abc_17692_n3699_1;
  wire _abc_17692_n3700;
  wire _abc_17692_n3701;
  wire _abc_17692_n3702;
  wire _abc_17692_n3703;
  wire _abc_17692_n3704;
  wire _abc_17692_n3705;
  wire _abc_17692_n3706;
  wire _abc_17692_n3707;
  wire _abc_17692_n3708;
  wire _abc_17692_n3709;
  wire _abc_17692_n3710;
  wire _abc_17692_n3711;
  wire _abc_17692_n3712_1;
  wire _abc_17692_n3713;
  wire _abc_17692_n3714;
  wire _abc_17692_n3715;
  wire _abc_17692_n3716;
  wire _abc_17692_n3717;
  wire _abc_17692_n3718;
  wire _abc_17692_n3719;
  wire _abc_17692_n3720;
  wire _abc_17692_n3721;
  wire _abc_17692_n3722;
  wire _abc_17692_n3723;
  wire _abc_17692_n3724;
  wire _abc_17692_n3725;
  wire _abc_17692_n3726;
  wire _abc_17692_n3727;
  wire _abc_17692_n3728;
  wire _abc_17692_n3729;
  wire _abc_17692_n3730;
  wire _abc_17692_n3731;
  wire _abc_17692_n3732;
  wire _abc_17692_n3733_1;
  wire _abc_17692_n3734;
  wire _abc_17692_n3735;
  wire _abc_17692_n3736;
  wire _abc_17692_n3737;
  wire _abc_17692_n3738;
  wire _abc_17692_n3739;
  wire _abc_17692_n3740;
  wire _abc_17692_n3741;
  wire _abc_17692_n3742;
  wire _abc_17692_n3743;
  wire _abc_17692_n3744;
  wire _abc_17692_n3745;
  wire _abc_17692_n3746;
  wire _abc_17692_n3747;
  wire _abc_17692_n3748;
  wire _abc_17692_n3749;
  wire _abc_17692_n3750;
  wire _abc_17692_n3751;
  wire _abc_17692_n3752;
  wire _abc_17692_n3753;
  wire _abc_17692_n3754_1;
  wire _abc_17692_n3755;
  wire _abc_17692_n3756;
  wire _abc_17692_n3757;
  wire _abc_17692_n3758;
  wire _abc_17692_n3759;
  wire _abc_17692_n3760;
  wire _abc_17692_n3761;
  wire _abc_17692_n3762;
  wire _abc_17692_n3763;
  wire _abc_17692_n3764;
  wire _abc_17692_n3765;
  wire _abc_17692_n3766;
  wire _abc_17692_n3767;
  wire _abc_17692_n3768;
  wire _abc_17692_n3769;
  wire _abc_17692_n3770;
  wire _abc_17692_n3771;
  wire _abc_17692_n3772;
  wire _abc_17692_n3773;
  wire _abc_17692_n3774;
  wire _abc_17692_n3775;
  wire _abc_17692_n3776_1;
  wire _abc_17692_n3777;
  wire _abc_17692_n3778;
  wire _abc_17692_n3779;
  wire _abc_17692_n3780;
  wire _abc_17692_n3781;
  wire _abc_17692_n3782;
  wire _abc_17692_n3783;
  wire _abc_17692_n3784;
  wire _abc_17692_n3785;
  wire _abc_17692_n3786;
  wire _abc_17692_n3787;
  wire _abc_17692_n3788;
  wire _abc_17692_n3789;
  wire _abc_17692_n3790;
  wire _abc_17692_n3791;
  wire _abc_17692_n3792;
  wire _abc_17692_n3793;
  wire _abc_17692_n3794;
  wire _abc_17692_n3795;
  wire _abc_17692_n3796;
  wire _abc_17692_n3797;
  wire _abc_17692_n3798;
  wire _abc_17692_n3799;
  wire _abc_17692_n3800;
  wire _abc_17692_n3801;
  wire _abc_17692_n3802;
  wire _abc_17692_n3803;
  wire _abc_17692_n3804;
  wire _abc_17692_n3805;
  wire _abc_17692_n3806;
  wire _abc_17692_n3807;
  wire _abc_17692_n3808;
  wire _abc_17692_n3809;
  wire _abc_17692_n3810;
  wire _abc_17692_n3811;
  wire _abc_17692_n3812;
  wire _abc_17692_n3813;
  wire _abc_17692_n3814;
  wire _abc_17692_n3815;
  wire _abc_17692_n3816;
  wire _abc_17692_n3817;
  wire _abc_17692_n3818;
  wire _abc_17692_n3819;
  wire _abc_17692_n3820;
  wire _abc_17692_n3821;
  wire _abc_17692_n3822;
  wire _abc_17692_n3823;
  wire _abc_17692_n3824;
  wire _abc_17692_n3825;
  wire _abc_17692_n3826;
  wire _abc_17692_n3827;
  wire _abc_17692_n3828;
  wire _abc_17692_n3829;
  wire _abc_17692_n3830;
  wire _abc_17692_n3831;
  wire _abc_17692_n3832;
  wire _abc_17692_n3833;
  wire _abc_17692_n3834_1;
  wire _abc_17692_n3835;
  wire _abc_17692_n3836;
  wire _abc_17692_n3837_1;
  wire _abc_17692_n3838;
  wire _abc_17692_n3839;
  wire _abc_17692_n3840;
  wire _abc_17692_n3841;
  wire _abc_17692_n3842;
  wire _abc_17692_n3843_1;
  wire _abc_17692_n3844;
  wire _abc_17692_n3845;
  wire _abc_17692_n3846;
  wire _abc_17692_n3847;
  wire _abc_17692_n3848;
  wire _abc_17692_n3849;
  wire _abc_17692_n3850;
  wire _abc_17692_n3851;
  wire _abc_17692_n3852;
  wire _abc_17692_n3853;
  wire _abc_17692_n3854;
  wire _abc_17692_n3855_1;
  wire _abc_17692_n3856;
  wire _abc_17692_n3857;
  wire _abc_17692_n3858;
  wire _abc_17692_n3859;
  wire _abc_17692_n3860;
  wire _abc_17692_n3861;
  wire _abc_17692_n3862;
  wire _abc_17692_n3863;
  wire _abc_17692_n3865;
  wire _abc_17692_n3866_1;
  wire _abc_17692_n3867;
  wire _abc_17692_n3868;
  wire _abc_17692_n3869;
  wire _abc_17692_n3870;
  wire _abc_17692_n3871;
  wire _abc_17692_n3872;
  wire _abc_17692_n3873;
  wire _abc_17692_n3874;
  wire _abc_17692_n3875;
  wire _abc_17692_n3876;
  wire _abc_17692_n3877_1;
  wire _abc_17692_n3878;
  wire _abc_17692_n3879;
  wire _abc_17692_n3880;
  wire _abc_17692_n3881;
  wire _abc_17692_n3882;
  wire _abc_17692_n3883;
  wire _abc_17692_n3884;
  wire _abc_17692_n3885;
  wire _abc_17692_n3886;
  wire _abc_17692_n3887;
  wire _abc_17692_n3888;
  wire _abc_17692_n3889;
  wire _abc_17692_n3890;
  wire _abc_17692_n3891;
  wire _abc_17692_n3892;
  wire _abc_17692_n3893;
  wire _abc_17692_n3894;
  wire _abc_17692_n3895;
  wire _abc_17692_n3896;
  wire _abc_17692_n3897;
  wire _abc_17692_n3898;
  wire _abc_17692_n3899;
  wire _abc_17692_n3900;
  wire _abc_17692_n3901;
  wire _abc_17692_n3902;
  wire _abc_17692_n3903;
  wire _abc_17692_n3904;
  wire _abc_17692_n3905;
  wire _abc_17692_n3906;
  wire _abc_17692_n3907;
  wire _abc_17692_n3908;
  wire _abc_17692_n3909;
  wire _abc_17692_n3910;
  wire _abc_17692_n3911;
  wire _abc_17692_n3912_1;
  wire _abc_17692_n3913;
  wire _abc_17692_n3914;
  wire _abc_17692_n3915_1;
  wire _abc_17692_n3916;
  wire _abc_17692_n3917;
  wire _abc_17692_n3918;
  wire _abc_17692_n3919;
  wire _abc_17692_n3920;
  wire _abc_17692_n3921;
  wire _abc_17692_n3922;
  wire _abc_17692_n3923;
  wire _abc_17692_n3924;
  wire _abc_17692_n3925;
  wire _abc_17692_n3926;
  wire _abc_17692_n3927;
  wire _abc_17692_n3928;
  wire _abc_17692_n3929;
  wire _abc_17692_n3930_1;
  wire _abc_17692_n3931;
  wire _abc_17692_n3932;
  wire _abc_17692_n3933;
  wire _abc_17692_n3934;
  wire _abc_17692_n3935;
  wire _abc_17692_n3936;
  wire _abc_17692_n3937;
  wire _abc_17692_n3938;
  wire _abc_17692_n3939;
  wire _abc_17692_n3940;
  wire _abc_17692_n3941;
  wire _abc_17692_n3942;
  wire _abc_17692_n3943;
  wire _abc_17692_n3944;
  wire _abc_17692_n3945;
  wire _abc_17692_n3946;
  wire _abc_17692_n3947;
  wire _abc_17692_n3948;
  wire _abc_17692_n3949;
  wire _abc_17692_n3950;
  wire _abc_17692_n3951;
  wire _abc_17692_n3952;
  wire _abc_17692_n3953;
  wire _abc_17692_n3954_1;
  wire _abc_17692_n3955;
  wire _abc_17692_n3956;
  wire _abc_17692_n3957;
  wire _abc_17692_n3958;
  wire _abc_17692_n3959;
  wire _abc_17692_n3960;
  wire _abc_17692_n3961;
  wire _abc_17692_n3962;
  wire _abc_17692_n3963;
  wire _abc_17692_n3964;
  wire _abc_17692_n3965;
  wire _abc_17692_n3966;
  wire _abc_17692_n3967;
  wire _abc_17692_n3968;
  wire _abc_17692_n3969;
  wire _abc_17692_n3970;
  wire _abc_17692_n3971;
  wire _abc_17692_n3972;
  wire _abc_17692_n3973;
  wire _abc_17692_n3974;
  wire _abc_17692_n3975;
  wire _abc_17692_n3976;
  wire _abc_17692_n3977;
  wire _abc_17692_n3978_1;
  wire _abc_17692_n3979;
  wire _abc_17692_n3980;
  wire _abc_17692_n3981;
  wire _abc_17692_n3982;
  wire _abc_17692_n3983;
  wire _abc_17692_n3984;
  wire _abc_17692_n3985;
  wire _abc_17692_n3986;
  wire _abc_17692_n3987;
  wire _abc_17692_n3988;
  wire _abc_17692_n3989;
  wire _abc_17692_n3990;
  wire _abc_17692_n3991;
  wire _abc_17692_n3992;
  wire _abc_17692_n3993;
  wire _abc_17692_n3994;
  wire _abc_17692_n3995;
  wire _abc_17692_n3996;
  wire _abc_17692_n3997;
  wire _abc_17692_n3998;
  wire _abc_17692_n3999;
  wire _abc_17692_n4000;
  wire _abc_17692_n4001;
  wire _abc_17692_n4002_1;
  wire _abc_17692_n4003;
  wire _abc_17692_n4004;
  wire _abc_17692_n4005;
  wire _abc_17692_n4006;
  wire _abc_17692_n4007;
  wire _abc_17692_n4008;
  wire _abc_17692_n4009;
  wire _abc_17692_n4010;
  wire _abc_17692_n4011;
  wire _abc_17692_n4012;
  wire _abc_17692_n4013;
  wire _abc_17692_n4014;
  wire _abc_17692_n4015;
  wire _abc_17692_n4016;
  wire _abc_17692_n4017;
  wire _abc_17692_n4018;
  wire _abc_17692_n4019;
  wire _abc_17692_n4020;
  wire _abc_17692_n4021;
  wire _abc_17692_n4022;
  wire _abc_17692_n4023;
  wire _abc_17692_n4024;
  wire _abc_17692_n4025;
  wire _abc_17692_n4026;
  wire _abc_17692_n4027;
  wire _abc_17692_n4028;
  wire _abc_17692_n4029;
  wire _abc_17692_n4030;
  wire _abc_17692_n4031;
  wire _abc_17692_n4032;
  wire _abc_17692_n4033;
  wire _abc_17692_n4034;
  wire _abc_17692_n4035;
  wire _abc_17692_n4036;
  wire _abc_17692_n4037;
  wire _abc_17692_n4038;
  wire _abc_17692_n4039;
  wire _abc_17692_n4040;
  wire _abc_17692_n4041;
  wire _abc_17692_n4042;
  wire _abc_17692_n4043;
  wire _abc_17692_n4044;
  wire _abc_17692_n4045;
  wire _abc_17692_n4047;
  wire _abc_17692_n4047_bF_buf0;
  wire _abc_17692_n4047_bF_buf1;
  wire _abc_17692_n4047_bF_buf2;
  wire _abc_17692_n4047_bF_buf3;
  wire _abc_17692_n4047_bF_buf4;
  wire _abc_17692_n4048;
  wire _abc_17692_n4049;
  wire _abc_17692_n4050;
  wire _abc_17692_n4051;
  wire _abc_17692_n4052;
  wire _abc_17692_n4053;
  wire _abc_17692_n4054;
  wire _abc_17692_n4055;
  wire _abc_17692_n4056;
  wire _abc_17692_n4057;
  wire _abc_17692_n4058;
  wire _abc_17692_n4059;
  wire _abc_17692_n4060;
  wire _abc_17692_n4061;
  wire _abc_17692_n4062;
  wire _abc_17692_n4063;
  wire _abc_17692_n4064_1;
  wire _abc_17692_n4065;
  wire _abc_17692_n4066;
  wire _abc_17692_n4067_1;
  wire _abc_17692_n4068;
  wire _abc_17692_n4069;
  wire _abc_17692_n4070;
  wire _abc_17692_n4071;
  wire _abc_17692_n4072;
  wire _abc_17692_n4073_1;
  wire _abc_17692_n4074;
  wire _abc_17692_n4075;
  wire _abc_17692_n4076;
  wire _abc_17692_n4077;
  wire _abc_17692_n4078;
  wire _abc_17692_n4079;
  wire _abc_17692_n4080;
  wire _abc_17692_n4081;
  wire _abc_17692_n4082;
  wire _abc_17692_n4083;
  wire _abc_17692_n4084_1;
  wire _abc_17692_n4085;
  wire _abc_17692_n4086;
  wire _abc_17692_n4087;
  wire _abc_17692_n4088;
  wire _abc_17692_n4089;
  wire _abc_17692_n4090;
  wire _abc_17692_n4091;
  wire _abc_17692_n4092;
  wire _abc_17692_n4093;
  wire _abc_17692_n4094;
  wire _abc_17692_n4095;
  wire _abc_17692_n4096_1;
  wire _abc_17692_n4097;
  wire _abc_17692_n4098;
  wire _abc_17692_n4099;
  wire _abc_17692_n4100;
  wire _abc_17692_n4101;
  wire _abc_17692_n4102;
  wire _abc_17692_n4103;
  wire _abc_17692_n4104;
  wire _abc_17692_n4105;
  wire _abc_17692_n4106;
  wire _abc_17692_n4107_1;
  wire _abc_17692_n4108;
  wire _abc_17692_n4109;
  wire _abc_17692_n4110;
  wire _abc_17692_n4111;
  wire _abc_17692_n4112;
  wire _abc_17692_n4113;
  wire _abc_17692_n4114;
  wire _abc_17692_n4115;
  wire _abc_17692_n4116;
  wire _abc_17692_n4117;
  wire _abc_17692_n4118;
  wire _abc_17692_n4119;
  wire _abc_17692_n4120;
  wire _abc_17692_n4121;
  wire _abc_17692_n4122;
  wire _abc_17692_n4123;
  wire _abc_17692_n4124;
  wire _abc_17692_n4125;
  wire _abc_17692_n4126;
  wire _abc_17692_n4127;
  wire _abc_17692_n4128;
  wire _abc_17692_n4129;
  wire _abc_17692_n4130;
  wire _abc_17692_n4131;
  wire _abc_17692_n4132;
  wire _abc_17692_n4133;
  wire _abc_17692_n4134;
  wire _abc_17692_n4135;
  wire _abc_17692_n4136;
  wire _abc_17692_n4137;
  wire _abc_17692_n4138;
  wire _abc_17692_n4139;
  wire _abc_17692_n4140_1;
  wire _abc_17692_n4141;
  wire _abc_17692_n4142;
  wire _abc_17692_n4143_1;
  wire _abc_17692_n4144;
  wire _abc_17692_n4145;
  wire _abc_17692_n4146;
  wire _abc_17692_n4147;
  wire _abc_17692_n4148;
  wire _abc_17692_n4149;
  wire _abc_17692_n4150;
  wire _abc_17692_n4151;
  wire _abc_17692_n4152_1;
  wire _abc_17692_n4153;
  wire _abc_17692_n4154;
  wire _abc_17692_n4155;
  wire _abc_17692_n4156;
  wire _abc_17692_n4157;
  wire _abc_17692_n4158;
  wire _abc_17692_n4159;
  wire _abc_17692_n4160;
  wire _abc_17692_n4161;
  wire _abc_17692_n4162;
  wire _abc_17692_n4163;
  wire _abc_17692_n4164;
  wire _abc_17692_n4165;
  wire _abc_17692_n4166;
  wire _abc_17692_n4167;
  wire _abc_17692_n4168;
  wire _abc_17692_n4169_1;
  wire _abc_17692_n4170;
  wire _abc_17692_n4171;
  wire _abc_17692_n4172;
  wire _abc_17692_n4173;
  wire _abc_17692_n4174;
  wire _abc_17692_n4175;
  wire _abc_17692_n4176;
  wire _abc_17692_n4177;
  wire _abc_17692_n4178;
  wire _abc_17692_n4179;
  wire _abc_17692_n4180;
  wire _abc_17692_n4181;
  wire _abc_17692_n4182;
  wire _abc_17692_n4183;
  wire _abc_17692_n4184;
  wire _abc_17692_n4185;
  wire _abc_17692_n4186_1;
  wire _abc_17692_n4187;
  wire _abc_17692_n4188;
  wire _abc_17692_n4189;
  wire _abc_17692_n4190;
  wire _abc_17692_n4191;
  wire _abc_17692_n4192;
  wire _abc_17692_n4193;
  wire _abc_17692_n4194;
  wire _abc_17692_n4195;
  wire _abc_17692_n4196;
  wire _abc_17692_n4197;
  wire _abc_17692_n4198;
  wire _abc_17692_n4199;
  wire _abc_17692_n4200;
  wire _abc_17692_n4201;
  wire _abc_17692_n4202_1;
  wire _abc_17692_n4203;
  wire _abc_17692_n4204;
  wire _abc_17692_n4205;
  wire _abc_17692_n4206;
  wire _abc_17692_n4207;
  wire _abc_17692_n4208;
  wire _abc_17692_n4209;
  wire _abc_17692_n4210;
  wire _abc_17692_n4211;
  wire _abc_17692_n4212;
  wire _abc_17692_n4213;
  wire _abc_17692_n4214;
  wire _abc_17692_n4215;
  wire _abc_17692_n4216;
  wire _abc_17692_n4217;
  wire _abc_17692_n4218;
  wire _abc_17692_n4219;
  wire _abc_17692_n4220;
  wire _abc_17692_n4221;
  wire _abc_17692_n4222;
  wire _abc_17692_n4223;
  wire _abc_17692_n4224;
  wire _abc_17692_n4225;
  wire _abc_17692_n4226;
  wire _abc_17692_n4227;
  wire _abc_17692_n4228;
  wire _abc_17692_n4229;
  wire _abc_17692_n4230;
  wire _abc_17692_n4231;
  wire _abc_17692_n4232;
  wire _abc_17692_n4233;
  wire _abc_17692_n4234;
  wire _abc_17692_n4235;
  wire _abc_17692_n4236;
  wire _abc_17692_n4237;
  wire _abc_17692_n4238;
  wire _abc_17692_n4239;
  wire _abc_17692_n4240;
  wire _abc_17692_n4241;
  wire _abc_17692_n4242;
  wire _abc_17692_n4243;
  wire _abc_17692_n4244;
  wire _abc_17692_n4245;
  wire _abc_17692_n4246;
  wire _abc_17692_n4247;
  wire _abc_17692_n4248;
  wire _abc_17692_n4249;
  wire _abc_17692_n4250_1;
  wire _abc_17692_n4251;
  wire _abc_17692_n4252;
  wire _abc_17692_n4253_1;
  wire _abc_17692_n4254;
  wire _abc_17692_n4255;
  wire _abc_17692_n4256;
  wire _abc_17692_n4257;
  wire _abc_17692_n4258_1;
  wire _abc_17692_n4259;
  wire _abc_17692_n4260;
  wire _abc_17692_n4261;
  wire _abc_17692_n4262;
  wire _abc_17692_n4263;
  wire _abc_17692_n4264;
  wire _abc_17692_n4265;
  wire _abc_17692_n4266;
  wire _abc_17692_n4267;
  wire _abc_17692_n4268;
  wire _abc_17692_n4269_1;
  wire _abc_17692_n4270;
  wire _abc_17692_n4271;
  wire _abc_17692_n4272;
  wire _abc_17692_n4273;
  wire _abc_17692_n4274;
  wire _abc_17692_n4275;
  wire _abc_17692_n4276;
  wire _abc_17692_n4277;
  wire _abc_17692_n4278;
  wire _abc_17692_n4279_1;
  wire _abc_17692_n4280;
  wire _abc_17692_n4281;
  wire _abc_17692_n4282;
  wire _abc_17692_n4283;
  wire _abc_17692_n4284;
  wire _abc_17692_n4285;
  wire _abc_17692_n4286;
  wire _abc_17692_n4287;
  wire _abc_17692_n4288;
  wire _abc_17692_n4289_1;
  wire _abc_17692_n4290;
  wire _abc_17692_n4291;
  wire _abc_17692_n4292;
  wire _abc_17692_n4293;
  wire _abc_17692_n4294;
  wire _abc_17692_n4295;
  wire _abc_17692_n4296;
  wire _abc_17692_n4297;
  wire _abc_17692_n4298;
  wire _abc_17692_n4299;
  wire _abc_17692_n4300;
  wire _abc_17692_n4301;
  wire _abc_17692_n4302;
  wire _abc_17692_n4303;
  wire _abc_17692_n4304;
  wire _abc_17692_n4305;
  wire _abc_17692_n4306;
  wire _abc_17692_n4307;
  wire _abc_17692_n4308;
  wire _abc_17692_n4309;
  wire _abc_17692_n4310;
  wire _abc_17692_n4311;
  wire _abc_17692_n4312;
  wire _abc_17692_n4313;
  wire _abc_17692_n4314;
  wire _abc_17692_n4315;
  wire _abc_17692_n4316;
  wire _abc_17692_n4317_1;
  wire _abc_17692_n4318;
  wire _abc_17692_n4319;
  wire _abc_17692_n4321;
  wire _abc_17692_n4322;
  wire _abc_17692_n4323;
  wire _abc_17692_n4324;
  wire _abc_17692_n4325;
  wire _abc_17692_n4326;
  wire _abc_17692_n4327;
  wire _abc_17692_n4328;
  wire _abc_17692_n4329;
  wire _abc_17692_n4330;
  wire _abc_17692_n4331;
  wire _abc_17692_n4332;
  wire _abc_17692_n4333;
  wire _abc_17692_n4334;
  wire _abc_17692_n4335;
  wire _abc_17692_n4336;
  wire _abc_17692_n4337;
  wire _abc_17692_n4338;
  wire _abc_17692_n4339;
  wire _abc_17692_n4340;
  wire _abc_17692_n4341;
  wire _abc_17692_n4342;
  wire _abc_17692_n4343;
  wire _abc_17692_n4344_1;
  wire _abc_17692_n4345;
  wire _abc_17692_n4346;
  wire _abc_17692_n4347_1;
  wire _abc_17692_n4348;
  wire _abc_17692_n4349;
  wire _abc_17692_n4350;
  wire _abc_17692_n4351;
  wire _abc_17692_n4352;
  wire _abc_17692_n4353;
  wire _abc_17692_n4354;
  wire _abc_17692_n4355;
  wire _abc_17692_n4356;
  wire _abc_17692_n4357;
  wire _abc_17692_n4358;
  wire _abc_17692_n4359;
  wire _abc_17692_n4360;
  wire _abc_17692_n4361;
  wire _abc_17692_n4362;
  wire _abc_17692_n4363;
  wire _abc_17692_n4364;
  wire _abc_17692_n4365;
  wire _abc_17692_n4366;
  wire _abc_17692_n4367;
  wire _abc_17692_n4368;
  wire _abc_17692_n4369;
  wire _abc_17692_n4370;
  wire _abc_17692_n4371;
  wire _abc_17692_n4372;
  wire _abc_17692_n4373;
  wire _abc_17692_n4374;
  wire _abc_17692_n4375;
  wire _abc_17692_n4376;
  wire _abc_17692_n4377;
  wire _abc_17692_n4378;
  wire _abc_17692_n4379;
  wire _abc_17692_n4380;
  wire _abc_17692_n4381;
  wire _abc_17692_n4382;
  wire _abc_17692_n4383;
  wire _abc_17692_n4384;
  wire _abc_17692_n4385;
  wire _abc_17692_n4386;
  wire _abc_17692_n4387;
  wire _abc_17692_n4388;
  wire _abc_17692_n4389_1;
  wire _abc_17692_n4390;
  wire _abc_17692_n4391;
  wire _abc_17692_n4392_1;
  wire _abc_17692_n4393;
  wire _abc_17692_n4394;
  wire _abc_17692_n4395;
  wire _abc_17692_n4396;
  wire _abc_17692_n4397;
  wire _abc_17692_n4398;
  wire _abc_17692_n4399;
  wire _abc_17692_n4400;
  wire _abc_17692_n4401;
  wire _abc_17692_n4402;
  wire _abc_17692_n4403;
  wire _abc_17692_n4404;
  wire _abc_17692_n4405;
  wire _abc_17692_n4406;
  wire _abc_17692_n4407;
  wire _abc_17692_n4408;
  wire _abc_17692_n4409;
  wire _abc_17692_n4410;
  wire _abc_17692_n4411;
  wire _abc_17692_n4412;
  wire _abc_17692_n4413;
  wire _abc_17692_n4414;
  wire _abc_17692_n4415;
  wire _abc_17692_n4416;
  wire _abc_17692_n4417;
  wire _abc_17692_n4418;
  wire _abc_17692_n4419;
  wire _abc_17692_n4420;
  wire _abc_17692_n4421;
  wire _abc_17692_n4422;
  wire _abc_17692_n4423;
  wire _abc_17692_n4424;
  wire _abc_17692_n4425;
  wire _abc_17692_n4426;
  wire _abc_17692_n4427;
  wire _abc_17692_n4428;
  wire _abc_17692_n4429;
  wire _abc_17692_n4430;
  wire _abc_17692_n4431;
  wire _abc_17692_n4432;
  wire _abc_17692_n4433;
  wire _abc_17692_n4434;
  wire _abc_17692_n4435;
  wire _abc_17692_n4436;
  wire _abc_17692_n4437;
  wire _abc_17692_n4438;
  wire _abc_17692_n4439;
  wire _abc_17692_n4440;
  wire _abc_17692_n4441;
  wire _abc_17692_n4442;
  wire _abc_17692_n4443;
  wire _abc_17692_n4444_1;
  wire _abc_17692_n4445;
  wire _abc_17692_n4446;
  wire _abc_17692_n4447_1;
  wire _abc_17692_n4448;
  wire _abc_17692_n4449;
  wire _abc_17692_n4450;
  wire _abc_17692_n4451;
  wire _abc_17692_n4452;
  wire _abc_17692_n4453;
  wire _abc_17692_n4454;
  wire _abc_17692_n4455;
  wire _abc_17692_n4456;
  wire _abc_17692_n4457;
  wire _abc_17692_n4458;
  wire _abc_17692_n4459;
  wire _abc_17692_n4460;
  wire _abc_17692_n4461;
  wire _abc_17692_n4462;
  wire _abc_17692_n4463;
  wire _abc_17692_n4464;
  wire _abc_17692_n4465;
  wire _abc_17692_n4466;
  wire _abc_17692_n4467;
  wire _abc_17692_n4468;
  wire _abc_17692_n4469;
  wire _abc_17692_n4470;
  wire _abc_17692_n4471;
  wire _abc_17692_n4472;
  wire _abc_17692_n4473;
  wire _abc_17692_n4474;
  wire _abc_17692_n4475;
  wire _abc_17692_n4476;
  wire _abc_17692_n4477;
  wire _abc_17692_n4478;
  wire _abc_17692_n4479;
  wire _abc_17692_n4480;
  wire _abc_17692_n4481;
  wire _abc_17692_n4482;
  wire _abc_17692_n4483;
  wire _abc_17692_n4484;
  wire _abc_17692_n4485;
  wire _abc_17692_n4486;
  wire _abc_17692_n4488;
  wire _abc_17692_n4489;
  wire _abc_17692_n4490;
  wire _abc_17692_n4491;
  wire _abc_17692_n4492;
  wire _abc_17692_n4493;
  wire _abc_17692_n4494;
  wire _abc_17692_n4495;
  wire _abc_17692_n4496;
  wire _abc_17692_n4497;
  wire _abc_17692_n4498;
  wire _abc_17692_n4499;
  wire _abc_17692_n4500;
  wire _abc_17692_n4501;
  wire _abc_17692_n4502;
  wire _abc_17692_n4503;
  wire _abc_17692_n4504;
  wire _abc_17692_n4505;
  wire _abc_17692_n4506;
  wire _abc_17692_n4507_1;
  wire _abc_17692_n4508;
  wire _abc_17692_n4509;
  wire _abc_17692_n4510_1;
  wire _abc_17692_n4511;
  wire _abc_17692_n4512;
  wire _abc_17692_n4513;
  wire _abc_17692_n4514;
  wire _abc_17692_n4515;
  wire _abc_17692_n4516;
  wire _abc_17692_n4517;
  wire _abc_17692_n4518;
  wire _abc_17692_n4519;
  wire _abc_17692_n4520;
  wire _abc_17692_n4521;
  wire _abc_17692_n4522;
  wire _abc_17692_n4523;
  wire _abc_17692_n4524;
  wire _abc_17692_n4525;
  wire _abc_17692_n4526;
  wire _abc_17692_n4527;
  wire _abc_17692_n4528;
  wire _abc_17692_n4529;
  wire _abc_17692_n4530;
  wire _abc_17692_n4531;
  wire _abc_17692_n4532;
  wire _abc_17692_n4533;
  wire _abc_17692_n4534;
  wire _abc_17692_n4535;
  wire _abc_17692_n4536;
  wire _abc_17692_n4537;
  wire _abc_17692_n4538;
  wire _abc_17692_n4539;
  wire _abc_17692_n4540;
  wire _abc_17692_n4541;
  wire _abc_17692_n4542;
  wire _abc_17692_n4543;
  wire _abc_17692_n4544;
  wire _abc_17692_n4545;
  wire _abc_17692_n4546;
  wire _abc_17692_n4547;
  wire _abc_17692_n4548;
  wire _abc_17692_n4549;
  wire _abc_17692_n4550;
  wire _abc_17692_n4551;
  wire _abc_17692_n4552;
  wire _abc_17692_n4553;
  wire _abc_17692_n4554;
  wire _abc_17692_n4555;
  wire _abc_17692_n4556;
  wire _abc_17692_n4557;
  wire _abc_17692_n4558;
  wire _abc_17692_n4559;
  wire _abc_17692_n4560;
  wire _abc_17692_n4561;
  wire _abc_17692_n4562;
  wire _abc_17692_n4563;
  wire _abc_17692_n4564;
  wire _abc_17692_n4565;
  wire _abc_17692_n4566;
  wire _abc_17692_n4567;
  wire _abc_17692_n4568;
  wire _abc_17692_n4569;
  wire _abc_17692_n4570;
  wire _abc_17692_n4571;
  wire _abc_17692_n4572;
  wire _abc_17692_n4573;
  wire _abc_17692_n4574;
  wire _abc_17692_n4575;
  wire _abc_17692_n4576;
  wire _abc_17692_n4577;
  wire _abc_17692_n4578;
  wire _abc_17692_n4579;
  wire _abc_17692_n4580;
  wire _abc_17692_n4581;
  wire _abc_17692_n4582;
  wire _abc_17692_n4583;
  wire _abc_17692_n4584_1;
  wire _abc_17692_n4585;
  wire _abc_17692_n4586;
  wire _abc_17692_n4587_1;
  wire _abc_17692_n4588;
  wire _abc_17692_n4589;
  wire _abc_17692_n4590;
  wire _abc_17692_n4591;
  wire _abc_17692_n4592;
  wire _abc_17692_n4593;
  wire _abc_17692_n4594;
  wire _abc_17692_n4595;
  wire _abc_17692_n4596;
  wire _abc_17692_n4597;
  wire _abc_17692_n4598;
  wire _abc_17692_n4599;
  wire _abc_17692_n4600;
  wire _abc_17692_n4601;
  wire _abc_17692_n4602;
  wire _abc_17692_n4603;
  wire _abc_17692_n4604;
  wire _abc_17692_n4605;
  wire _abc_17692_n4606;
  wire _abc_17692_n4607;
  wire _abc_17692_n4608;
  wire _abc_17692_n4609;
  wire _abc_17692_n4610;
  wire _abc_17692_n4611;
  wire _abc_17692_n4612;
  wire _abc_17692_n4613;
  wire _abc_17692_n4614;
  wire _abc_17692_n4615;
  wire _abc_17692_n4616;
  wire _abc_17692_n4617;
  wire _abc_17692_n4618;
  wire _abc_17692_n4619;
  wire _abc_17692_n4620;
  wire _abc_17692_n4621;
  wire _abc_17692_n4622;
  wire _abc_17692_n4623;
  wire _abc_17692_n4624;
  wire _abc_17692_n4625;
  wire _abc_17692_n4626;
  wire _abc_17692_n4627;
  wire _abc_17692_n4628;
  wire _abc_17692_n4629;
  wire _abc_17692_n4630;
  wire _abc_17692_n4631;
  wire _abc_17692_n4632;
  wire _abc_17692_n4633;
  wire _abc_17692_n4634;
  wire _abc_17692_n4635;
  wire _abc_17692_n4636;
  wire _abc_17692_n4637;
  wire _abc_17692_n4638;
  wire _abc_17692_n4639;
  wire _abc_17692_n4640;
  wire _abc_17692_n4641;
  wire _abc_17692_n4642;
  wire _abc_17692_n4643_1;
  wire _abc_17692_n4644;
  wire _abc_17692_n4645;
  wire _abc_17692_n4646_1;
  wire _abc_17692_n4647;
  wire _abc_17692_n4648;
  wire _abc_17692_n4649;
  wire _abc_17692_n4650;
  wire _abc_17692_n4651;
  wire _abc_17692_n4652;
  wire _abc_17692_n4653;
  wire _abc_17692_n4654;
  wire _abc_17692_n4655;
  wire _abc_17692_n4656;
  wire _abc_17692_n4657;
  wire _abc_17692_n4658;
  wire _abc_17692_n4659;
  wire _abc_17692_n4660;
  wire _abc_17692_n4661;
  wire _abc_17692_n4662;
  wire _abc_17692_n4663;
  wire _abc_17692_n4664;
  wire _abc_17692_n4665;
  wire _abc_17692_n4666;
  wire _abc_17692_n4667;
  wire _abc_17692_n4668;
  wire _abc_17692_n4669;
  wire _abc_17692_n4670;
  wire _abc_17692_n4671;
  wire _abc_17692_n4672;
  wire _abc_17692_n4673;
  wire _abc_17692_n4674;
  wire _abc_17692_n4675;
  wire _abc_17692_n4676;
  wire _abc_17692_n4677;
  wire _abc_17692_n4678;
  wire _abc_17692_n4679;
  wire _abc_17692_n4680;
  wire _abc_17692_n4681;
  wire _abc_17692_n4682;
  wire _abc_17692_n4683;
  wire _abc_17692_n4684;
  wire _abc_17692_n4685;
  wire _abc_17692_n4686;
  wire _abc_17692_n4687;
  wire _abc_17692_n4688;
  wire _abc_17692_n4689;
  wire _abc_17692_n4690;
  wire _abc_17692_n4691;
  wire _abc_17692_n4692;
  wire _abc_17692_n4693;
  wire _abc_17692_n4694;
  wire _abc_17692_n4695;
  wire _abc_17692_n4696;
  wire _abc_17692_n4697;
  wire _abc_17692_n4698;
  wire _abc_17692_n4699;
  wire _abc_17692_n4700;
  wire _abc_17692_n4701;
  wire _abc_17692_n4702;
  wire _abc_17692_n4703;
  wire _abc_17692_n4704;
  wire _abc_17692_n4705;
  wire _abc_17692_n4706;
  wire _abc_17692_n4707;
  wire _abc_17692_n4708;
  wire _abc_17692_n4709;
  wire _abc_17692_n4710;
  wire _abc_17692_n4711;
  wire _abc_17692_n4712;
  wire _abc_17692_n4713;
  wire _abc_17692_n4714;
  wire _abc_17692_n4715;
  wire _abc_17692_n4716;
  wire _abc_17692_n4717;
  wire _abc_17692_n4718;
  wire _abc_17692_n4719;
  wire _abc_17692_n4720;
  wire _abc_17692_n4721;
  wire _abc_17692_n4722;
  wire _abc_17692_n4723;
  wire _abc_17692_n4724;
  wire _abc_17692_n4725;
  wire _abc_17692_n4726;
  wire _abc_17692_n4727;
  wire _abc_17692_n4729;
  wire _abc_17692_n4730;
  wire _abc_17692_n4731;
  wire _abc_17692_n4732;
  wire _abc_17692_n4733;
  wire _abc_17692_n4734;
  wire _abc_17692_n4735_1;
  wire _abc_17692_n4736;
  wire _abc_17692_n4737;
  wire _abc_17692_n4738_1;
  wire _abc_17692_n4739;
  wire _abc_17692_n4740;
  wire _abc_17692_n4741;
  wire _abc_17692_n4742;
  wire _abc_17692_n4743;
  wire _abc_17692_n4744;
  wire _abc_17692_n4745;
  wire _abc_17692_n4746;
  wire _abc_17692_n4747;
  wire _abc_17692_n4748;
  wire _abc_17692_n4749;
  wire _abc_17692_n4750;
  wire _abc_17692_n4751;
  wire _abc_17692_n4752;
  wire _abc_17692_n4753;
  wire _abc_17692_n4754;
  wire _abc_17692_n4755;
  wire _abc_17692_n4756;
  wire _abc_17692_n4757;
  wire _abc_17692_n4758;
  wire _abc_17692_n4759;
  wire _abc_17692_n4760;
  wire _abc_17692_n4761;
  wire _abc_17692_n4762;
  wire _abc_17692_n4763;
  wire _abc_17692_n4764;
  wire _abc_17692_n4765;
  wire _abc_17692_n4766;
  wire _abc_17692_n4767;
  wire _abc_17692_n4768;
  wire _abc_17692_n4769;
  wire _abc_17692_n4770;
  wire _abc_17692_n4771;
  wire _abc_17692_n4772;
  wire _abc_17692_n4773;
  wire _abc_17692_n4774;
  wire _abc_17692_n4775;
  wire _abc_17692_n4776;
  wire _abc_17692_n4777;
  wire _abc_17692_n4778;
  wire _abc_17692_n4779;
  wire _abc_17692_n4780;
  wire _abc_17692_n4781;
  wire _abc_17692_n4782;
  wire _abc_17692_n4783;
  wire _abc_17692_n4784;
  wire _abc_17692_n4785;
  wire _abc_17692_n4786;
  wire _abc_17692_n4787;
  wire _abc_17692_n4788;
  wire _abc_17692_n4789_1;
  wire _abc_17692_n4790;
  wire _abc_17692_n4791;
  wire _abc_17692_n4792_1;
  wire _abc_17692_n4793;
  wire _abc_17692_n4794;
  wire _abc_17692_n4795;
  wire _abc_17692_n4796;
  wire _abc_17692_n4797;
  wire _abc_17692_n4798;
  wire _abc_17692_n4799;
  wire _abc_17692_n4800;
  wire _abc_17692_n4801;
  wire _abc_17692_n4802;
  wire _abc_17692_n4803;
  wire _abc_17692_n4804;
  wire _abc_17692_n4805;
  wire _abc_17692_n4806;
  wire _abc_17692_n4807;
  wire _abc_17692_n4808;
  wire _abc_17692_n4809;
  wire _abc_17692_n4810;
  wire _abc_17692_n4811;
  wire _abc_17692_n4812;
  wire _abc_17692_n4813;
  wire _abc_17692_n4814;
  wire _abc_17692_n4815;
  wire _abc_17692_n4816;
  wire _abc_17692_n4817;
  wire _abc_17692_n4818;
  wire _abc_17692_n4819;
  wire _abc_17692_n4820;
  wire _abc_17692_n4821;
  wire _abc_17692_n4822;
  wire _abc_17692_n4823;
  wire _abc_17692_n4824;
  wire _abc_17692_n4825;
  wire _abc_17692_n4826;
  wire _abc_17692_n4827;
  wire _abc_17692_n4828;
  wire _abc_17692_n4829;
  wire _abc_17692_n4830;
  wire _abc_17692_n4831;
  wire _abc_17692_n4832;
  wire _abc_17692_n4833;
  wire _abc_17692_n4834;
  wire _abc_17692_n4835;
  wire _abc_17692_n4836;
  wire _abc_17692_n4837;
  wire _abc_17692_n4838;
  wire _abc_17692_n4839;
  wire _abc_17692_n4840;
  wire _abc_17692_n4841;
  wire _abc_17692_n4842;
  wire _abc_17692_n4843;
  wire _abc_17692_n4844;
  wire _abc_17692_n4845;
  wire _abc_17692_n4846;
  wire _abc_17692_n4847;
  wire _abc_17692_n4848;
  wire _abc_17692_n4849;
  wire _abc_17692_n4850;
  wire _abc_17692_n4851;
  wire _abc_17692_n4852;
  wire _abc_17692_n4853;
  wire _abc_17692_n4854;
  wire _abc_17692_n4855;
  wire _abc_17692_n4856;
  wire _abc_17692_n4857;
  wire _abc_17692_n4858;
  wire _abc_17692_n4859;
  wire _abc_17692_n4860;
  wire _abc_17692_n4861;
  wire _abc_17692_n4862;
  wire _abc_17692_n4863;
  wire _abc_17692_n4864;
  wire _abc_17692_n4865;
  wire _abc_17692_n4866;
  wire _abc_17692_n4867;
  wire _abc_17692_n4868;
  wire _abc_17692_n4869;
  wire _abc_17692_n4870;
  wire _abc_17692_n4871;
  wire _abc_17692_n4872;
  wire _abc_17692_n4873;
  wire _abc_17692_n4874;
  wire _abc_17692_n4875;
  wire _abc_17692_n4876;
  wire _abc_17692_n4877;
  wire _abc_17692_n4878;
  wire _abc_17692_n4879;
  wire _abc_17692_n4880;
  wire _abc_17692_n4881;
  wire _abc_17692_n4882;
  wire _abc_17692_n4883;
  wire _abc_17692_n4884;
  wire _abc_17692_n4885;
  wire _abc_17692_n4886;
  wire _abc_17692_n4887;
  wire _abc_17692_n4888;
  wire _abc_17692_n4889;
  wire _abc_17692_n4890;
  wire _abc_17692_n4891;
  wire _abc_17692_n4892;
  wire _abc_17692_n4893_1;
  wire _abc_17692_n4894;
  wire _abc_17692_n4895;
  wire _abc_17692_n4896_1;
  wire _abc_17692_n4897;
  wire _abc_17692_n4898;
  wire _abc_17692_n4899;
  wire _abc_17692_n4900;
  wire _abc_17692_n4901;
  wire _abc_17692_n4902;
  wire _abc_17692_n4903;
  wire _abc_17692_n4904;
  wire _abc_17692_n4905;
  wire _abc_17692_n4906;
  wire _abc_17692_n4907;
  wire _abc_17692_n4908;
  wire _abc_17692_n4909;
  wire _abc_17692_n4910;
  wire _abc_17692_n4911;
  wire _abc_17692_n4912;
  wire _abc_17692_n4914;
  wire _abc_17692_n4915;
  wire _abc_17692_n4916;
  wire _abc_17692_n4917;
  wire _abc_17692_n4918;
  wire _abc_17692_n4919;
  wire _abc_17692_n4920;
  wire _abc_17692_n4921;
  wire _abc_17692_n4922;
  wire _abc_17692_n4923;
  wire _abc_17692_n4924;
  wire _abc_17692_n4925;
  wire _abc_17692_n4926;
  wire _abc_17692_n4927;
  wire _abc_17692_n4928;
  wire _abc_17692_n4929;
  wire _abc_17692_n4930;
  wire _abc_17692_n4931;
  wire _abc_17692_n4932;
  wire _abc_17692_n4933;
  wire _abc_17692_n4934;
  wire _abc_17692_n4935;
  wire _abc_17692_n4936;
  wire _abc_17692_n4937;
  wire _abc_17692_n4938;
  wire _abc_17692_n4939;
  wire _abc_17692_n4940;
  wire _abc_17692_n4941;
  wire _abc_17692_n4942;
  wire _abc_17692_n4943;
  wire _abc_17692_n4944;
  wire _abc_17692_n4945;
  wire _abc_17692_n4946;
  wire _abc_17692_n4947;
  wire _abc_17692_n4948;
  wire _abc_17692_n4949;
  wire _abc_17692_n4950;
  wire _abc_17692_n4951;
  wire _abc_17692_n4952;
  wire _abc_17692_n4953;
  wire _abc_17692_n4954;
  wire _abc_17692_n4955;
  wire _abc_17692_n4956;
  wire _abc_17692_n4957;
  wire _abc_17692_n4958;
  wire _abc_17692_n4959;
  wire _abc_17692_n4960;
  wire _abc_17692_n4961;
  wire _abc_17692_n4962;
  wire _abc_17692_n4963_1;
  wire _abc_17692_n4964;
  wire _abc_17692_n4965;
  wire _abc_17692_n4966_1;
  wire _abc_17692_n4967;
  wire _abc_17692_n4968;
  wire _abc_17692_n4969;
  wire _abc_17692_n4970;
  wire _abc_17692_n4971;
  wire _abc_17692_n4972;
  wire _abc_17692_n4973;
  wire _abc_17692_n4974;
  wire _abc_17692_n4975;
  wire _abc_17692_n4976;
  wire _abc_17692_n4977;
  wire _abc_17692_n4978;
  wire _abc_17692_n4979;
  wire _abc_17692_n4980;
  wire _abc_17692_n4981;
  wire _abc_17692_n4982;
  wire _abc_17692_n4983;
  wire _abc_17692_n4984;
  wire _abc_17692_n4985;
  wire _abc_17692_n4986;
  wire _abc_17692_n4987;
  wire _abc_17692_n4988;
  wire _abc_17692_n4989;
  wire _abc_17692_n4990;
  wire _abc_17692_n4991;
  wire _abc_17692_n4992;
  wire _abc_17692_n4993;
  wire _abc_17692_n4994;
  wire _abc_17692_n4995;
  wire _abc_17692_n4996;
  wire _abc_17692_n4997;
  wire _abc_17692_n4998;
  wire _abc_17692_n4999;
  wire _abc_17692_n5000;
  wire _abc_17692_n5001;
  wire _abc_17692_n5002;
  wire _abc_17692_n5003;
  wire _abc_17692_n5004;
  wire _abc_17692_n5005;
  wire _abc_17692_n5006;
  wire _abc_17692_n5007;
  wire _abc_17692_n5008;
  wire _abc_17692_n5009;
  wire _abc_17692_n5010;
  wire _abc_17692_n5011;
  wire _abc_17692_n5012;
  wire _abc_17692_n5013;
  wire _abc_17692_n5014;
  wire _abc_17692_n5015;
  wire _abc_17692_n5016;
  wire _abc_17692_n5017;
  wire _abc_17692_n5018;
  wire _abc_17692_n5019;
  wire _abc_17692_n5020;
  wire _abc_17692_n5021;
  wire _abc_17692_n5022;
  wire _abc_17692_n5023;
  wire _abc_17692_n5024;
  wire _abc_17692_n5025;
  wire _abc_17692_n5026;
  wire _abc_17692_n5027;
  wire _abc_17692_n5028;
  wire _abc_17692_n5029;
  wire _abc_17692_n5030;
  wire _abc_17692_n5031;
  wire _abc_17692_n5032;
  wire _abc_17692_n5033;
  wire _abc_17692_n5034;
  wire _abc_17692_n5035;
  wire _abc_17692_n5036;
  wire _abc_17692_n5037;
  wire _abc_17692_n5038;
  wire _abc_17692_n5039;
  wire _abc_17692_n5040;
  wire _abc_17692_n5041;
  wire _abc_17692_n5042;
  wire _abc_17692_n5043;
  wire _abc_17692_n5044_1;
  wire _abc_17692_n5045;
  wire _abc_17692_n5046;
  wire _abc_17692_n5047_1;
  wire _abc_17692_n5048;
  wire _abc_17692_n5049;
  wire _abc_17692_n5050;
  wire _abc_17692_n5051;
  wire _abc_17692_n5052;
  wire _abc_17692_n5053;
  wire _abc_17692_n5054;
  wire _abc_17692_n5055;
  wire _abc_17692_n5056;
  wire _abc_17692_n5057;
  wire _abc_17692_n5058;
  wire _abc_17692_n5059;
  wire _abc_17692_n5060;
  wire _abc_17692_n5061;
  wire _abc_17692_n5062;
  wire _abc_17692_n5063;
  wire _abc_17692_n5064;
  wire _abc_17692_n5065;
  wire _abc_17692_n5066;
  wire _abc_17692_n5067;
  wire _abc_17692_n5068;
  wire _abc_17692_n5069;
  wire _abc_17692_n5070;
  wire _abc_17692_n5071;
  wire _abc_17692_n5072;
  wire _abc_17692_n5073;
  wire _abc_17692_n5074;
  wire _abc_17692_n5075;
  wire _abc_17692_n5076;
  wire _abc_17692_n5077;
  wire _abc_17692_n5078;
  wire _abc_17692_n5079;
  wire _abc_17692_n5080;
  wire _abc_17692_n5081;
  wire _abc_17692_n5082;
  wire _abc_17692_n5083;
  wire _abc_17692_n5084;
  wire _abc_17692_n5085;
  wire _abc_17692_n5086;
  wire _abc_17692_n5087;
  wire _abc_17692_n5088;
  wire _abc_17692_n5089;
  wire _abc_17692_n5090;
  wire _abc_17692_n5091;
  wire _abc_17692_n5092;
  wire _abc_17692_n5093;
  wire _abc_17692_n5094;
  wire _abc_17692_n5095;
  wire _abc_17692_n5096;
  wire _abc_17692_n5097_1;
  wire _abc_17692_n5098;
  wire _abc_17692_n5099;
  wire _abc_17692_n5100_1;
  wire _abc_17692_n5101;
  wire _abc_17692_n5102;
  wire _abc_17692_n5103;
  wire _abc_17692_n5104;
  wire _abc_17692_n5105;
  wire _abc_17692_n5106;
  wire _abc_17692_n5107;
  wire _abc_17692_n5108;
  wire _abc_17692_n5109;
  wire _abc_17692_n5110;
  wire _abc_17692_n5111;
  wire _abc_17692_n5112;
  wire _abc_17692_n5113;
  wire _abc_17692_n5114;
  wire _abc_17692_n5115;
  wire _abc_17692_n5116;
  wire _abc_17692_n5117;
  wire _abc_17692_n5118;
  wire _abc_17692_n5119;
  wire _abc_17692_n5120;
  wire _abc_17692_n5121;
  wire _abc_17692_n5122;
  wire _abc_17692_n5123;
  wire _abc_17692_n5124;
  wire _abc_17692_n5125;
  wire _abc_17692_n5126;
  wire _abc_17692_n5127;
  wire _abc_17692_n5128;
  wire _abc_17692_n5129;
  wire _abc_17692_n5130;
  wire _abc_17692_n5131;
  wire _abc_17692_n5132;
  wire _abc_17692_n5133;
  wire _abc_17692_n5134;
  wire _abc_17692_n5135;
  wire _abc_17692_n5136;
  wire _abc_17692_n5137;
  wire _abc_17692_n5138;
  wire _abc_17692_n5139;
  wire _abc_17692_n5140;
  wire _abc_17692_n5141;
  wire _abc_17692_n5142;
  wire _abc_17692_n5143;
  wire _abc_17692_n5144;
  wire _abc_17692_n5145;
  wire _abc_17692_n5146;
  wire _abc_17692_n5147;
  wire _abc_17692_n5148;
  wire _abc_17692_n5149;
  wire _abc_17692_n5150;
  wire _abc_17692_n5151;
  wire _abc_17692_n5152;
  wire _abc_17692_n5153;
  wire _abc_17692_n5154;
  wire _abc_17692_n5155;
  wire _abc_17692_n5156;
  wire _abc_17692_n5157;
  wire _abc_17692_n5158;
  wire _abc_17692_n5159;
  wire _abc_17692_n5160;
  wire _abc_17692_n5161;
  wire _abc_17692_n5162;
  wire _abc_17692_n5163;
  wire _abc_17692_n5164;
  wire _abc_17692_n5165;
  wire _abc_17692_n5166;
  wire _abc_17692_n5167;
  wire _abc_17692_n5168;
  wire _abc_17692_n5169;
  wire _abc_17692_n5170;
  wire _abc_17692_n5171;
  wire _abc_17692_n5172;
  wire _abc_17692_n5173;
  wire _abc_17692_n5174;
  wire _abc_17692_n5175;
  wire _abc_17692_n5176;
  wire _abc_17692_n5177;
  wire _abc_17692_n5178;
  wire _abc_17692_n5179;
  wire _abc_17692_n5180;
  wire _abc_17692_n5181;
  wire _abc_17692_n5182;
  wire _abc_17692_n5183;
  wire _abc_17692_n5184;
  wire _abc_17692_n5185;
  wire _abc_17692_n5186;
  wire _abc_17692_n5187;
  wire _abc_17692_n5188;
  wire _abc_17692_n5189;
  wire _abc_17692_n5190;
  wire _abc_17692_n5191;
  wire _abc_17692_n5192;
  wire _abc_17692_n5193;
  wire _abc_17692_n5194;
  wire _abc_17692_n5195;
  wire _abc_17692_n5196;
  wire _abc_17692_n5197;
  wire _abc_17692_n5198;
  wire _abc_17692_n5199;
  wire _abc_17692_n5200;
  wire _abc_17692_n5202;
  wire _abc_17692_n5203;
  wire _abc_17692_n5204;
  wire _abc_17692_n5205;
  wire _abc_17692_n5206;
  wire _abc_17692_n5207;
  wire _abc_17692_n5208;
  wire _abc_17692_n5209;
  wire _abc_17692_n5210;
  wire _abc_17692_n5211;
  wire _abc_17692_n5212_1;
  wire _abc_17692_n5213;
  wire _abc_17692_n5214;
  wire _abc_17692_n5215_1;
  wire _abc_17692_n5216;
  wire _abc_17692_n5217;
  wire _abc_17692_n5218;
  wire _abc_17692_n5219;
  wire _abc_17692_n5220;
  wire _abc_17692_n5221;
  wire _abc_17692_n5222;
  wire _abc_17692_n5223;
  wire _abc_17692_n5224;
  wire _abc_17692_n5225;
  wire _abc_17692_n5226;
  wire _abc_17692_n5227;
  wire _abc_17692_n5228;
  wire _abc_17692_n5229;
  wire _abc_17692_n5230;
  wire _abc_17692_n5231;
  wire _abc_17692_n5232;
  wire _abc_17692_n5233;
  wire _abc_17692_n5234;
  wire _abc_17692_n5235;
  wire _abc_17692_n5236;
  wire _abc_17692_n5237;
  wire _abc_17692_n5238;
  wire _abc_17692_n5239;
  wire _abc_17692_n5240;
  wire _abc_17692_n5241;
  wire _abc_17692_n5242;
  wire _abc_17692_n5243;
  wire _abc_17692_n5244;
  wire _abc_17692_n5245;
  wire _abc_17692_n5246;
  wire _abc_17692_n5247;
  wire _abc_17692_n5248;
  wire _abc_17692_n5249;
  wire _abc_17692_n5250;
  wire _abc_17692_n5251;
  wire _abc_17692_n5252;
  wire _abc_17692_n5253;
  wire _abc_17692_n5254;
  wire _abc_17692_n5255;
  wire _abc_17692_n5256;
  wire _abc_17692_n5257;
  wire _abc_17692_n5258;
  wire _abc_17692_n5259;
  wire _abc_17692_n5260;
  wire _abc_17692_n5261;
  wire _abc_17692_n5262;
  wire _abc_17692_n5263;
  wire _abc_17692_n5264;
  wire _abc_17692_n5265;
  wire _abc_17692_n5266;
  wire _abc_17692_n5267;
  wire _abc_17692_n5268;
  wire _abc_17692_n5269;
  wire _abc_17692_n5270;
  wire _abc_17692_n5271;
  wire _abc_17692_n5272;
  wire _abc_17692_n5273;
  wire _abc_17692_n5274;
  wire _abc_17692_n5275_1;
  wire _abc_17692_n5276;
  wire _abc_17692_n5277;
  wire _abc_17692_n5278_1;
  wire _abc_17692_n5279;
  wire _abc_17692_n5280;
  wire _abc_17692_n5281;
  wire _abc_17692_n5282;
  wire _abc_17692_n5283;
  wire _abc_17692_n5284;
  wire _abc_17692_n5285;
  wire _abc_17692_n5286;
  wire _abc_17692_n5287;
  wire _abc_17692_n5288;
  wire _abc_17692_n5289;
  wire _abc_17692_n5290;
  wire _abc_17692_n5291;
  wire _abc_17692_n5292;
  wire _abc_17692_n5293;
  wire _abc_17692_n5294;
  wire _abc_17692_n5295;
  wire _abc_17692_n5296;
  wire _abc_17692_n5297;
  wire _abc_17692_n5298;
  wire _abc_17692_n5299;
  wire _abc_17692_n5300;
  wire _abc_17692_n5301;
  wire _abc_17692_n5302;
  wire _abc_17692_n5303;
  wire _abc_17692_n5304;
  wire _abc_17692_n5305;
  wire _abc_17692_n5306;
  wire _abc_17692_n5307;
  wire _abc_17692_n5308;
  wire _abc_17692_n5309;
  wire _abc_17692_n5310;
  wire _abc_17692_n5311;
  wire _abc_17692_n5312;
  wire _abc_17692_n5313;
  wire _abc_17692_n5314;
  wire _abc_17692_n5315;
  wire _abc_17692_n5316;
  wire _abc_17692_n5317;
  wire _abc_17692_n5318;
  wire _abc_17692_n5319;
  wire _abc_17692_n5320;
  wire _abc_17692_n5321;
  wire _abc_17692_n5322;
  wire _abc_17692_n5323;
  wire _abc_17692_n5324;
  wire _abc_17692_n5325;
  wire _abc_17692_n5326;
  wire _abc_17692_n5327;
  wire _abc_17692_n5328;
  wire _abc_17692_n5329;
  wire _abc_17692_n5330;
  wire _abc_17692_n5331;
  wire _abc_17692_n5332;
  wire _abc_17692_n5333;
  wire _abc_17692_n5334;
  wire _abc_17692_n5335;
  wire _abc_17692_n5336;
  wire _abc_17692_n5337;
  wire _abc_17692_n5338;
  wire _abc_17692_n5339;
  wire _abc_17692_n5340;
  wire _abc_17692_n5341;
  wire _abc_17692_n5342;
  wire _abc_17692_n5343;
  wire _abc_17692_n5344;
  wire _abc_17692_n5345;
  wire _abc_17692_n5346;
  wire _abc_17692_n5347;
  wire _abc_17692_n5348;
  wire _abc_17692_n5349;
  wire _abc_17692_n5350;
  wire _abc_17692_n5351;
  wire _abc_17692_n5352;
  wire _abc_17692_n5353;
  wire _abc_17692_n5354;
  wire _abc_17692_n5355;
  wire _abc_17692_n5356;
  wire _abc_17692_n5357;
  wire _abc_17692_n5358;
  wire _abc_17692_n5359;
  wire _abc_17692_n5360;
  wire _abc_17692_n5361;
  wire _abc_17692_n5362;
  wire _abc_17692_n5363;
  wire _abc_17692_n5364;
  wire _abc_17692_n5365;
  wire _abc_17692_n5366_1;
  wire _abc_17692_n5367;
  wire _abc_17692_n5368;
  wire _abc_17692_n5369_1;
  wire _abc_17692_n5370;
  wire _abc_17692_n5371;
  wire _abc_17692_n5372;
  wire _abc_17692_n5373;
  wire _abc_17692_n5374;
  wire _abc_17692_n5376;
  wire _abc_17692_n5377;
  wire _abc_17692_n5378;
  wire _abc_17692_n5379;
  wire _abc_17692_n5380;
  wire _abc_17692_n5381;
  wire _abc_17692_n5382;
  wire _abc_17692_n5383;
  wire _abc_17692_n5384;
  wire _abc_17692_n5385;
  wire _abc_17692_n5386;
  wire _abc_17692_n5387;
  wire _abc_17692_n5388;
  wire _abc_17692_n5389;
  wire _abc_17692_n5390;
  wire _abc_17692_n5391;
  wire _abc_17692_n5392;
  wire _abc_17692_n5393;
  wire _abc_17692_n5394;
  wire _abc_17692_n5395;
  wire _abc_17692_n5396;
  wire _abc_17692_n5397;
  wire _abc_17692_n5398;
  wire _abc_17692_n5399;
  wire _abc_17692_n5400;
  wire _abc_17692_n5401;
  wire _abc_17692_n5402;
  wire _abc_17692_n5403;
  wire _abc_17692_n5404;
  wire _abc_17692_n5405;
  wire _abc_17692_n5406;
  wire _abc_17692_n5407;
  wire _abc_17692_n5408;
  wire _abc_17692_n5409;
  wire _abc_17692_n5410;
  wire _abc_17692_n5411;
  wire _abc_17692_n5412;
  wire _abc_17692_n5413;
  wire _abc_17692_n5414;
  wire _abc_17692_n5415;
  wire _abc_17692_n5416;
  wire _abc_17692_n5417;
  wire _abc_17692_n5418;
  wire _abc_17692_n5419;
  wire _abc_17692_n5420_1;
  wire _abc_17692_n5421;
  wire _abc_17692_n5422;
  wire _abc_17692_n5423_1;
  wire _abc_17692_n5424;
  wire _abc_17692_n5425;
  wire _abc_17692_n5426;
  wire _abc_17692_n5427;
  wire _abc_17692_n5428;
  wire _abc_17692_n5429;
  wire _abc_17692_n5430;
  wire _abc_17692_n5431;
  wire _abc_17692_n5432;
  wire _abc_17692_n5433;
  wire _abc_17692_n5434;
  wire _abc_17692_n5435;
  wire _abc_17692_n5436;
  wire _abc_17692_n5437;
  wire _abc_17692_n5438;
  wire _abc_17692_n5439;
  wire _abc_17692_n5440;
  wire _abc_17692_n5441;
  wire _abc_17692_n5442;
  wire _abc_17692_n5443;
  wire _abc_17692_n5444;
  wire _abc_17692_n5445;
  wire _abc_17692_n5446;
  wire _abc_17692_n5447;
  wire _abc_17692_n5448;
  wire _abc_17692_n5449;
  wire _abc_17692_n5450;
  wire _abc_17692_n5451;
  wire _abc_17692_n5452;
  wire _abc_17692_n5453;
  wire _abc_17692_n5454;
  wire _abc_17692_n5455;
  wire _abc_17692_n5456;
  wire _abc_17692_n5457;
  wire _abc_17692_n5458;
  wire _abc_17692_n5459;
  wire _abc_17692_n5460;
  wire _abc_17692_n5461;
  wire _abc_17692_n5462;
  wire _abc_17692_n5463;
  wire _abc_17692_n5464;
  wire _abc_17692_n5465;
  wire _abc_17692_n5466;
  wire _abc_17692_n5467;
  wire _abc_17692_n5468;
  wire _abc_17692_n5469;
  wire _abc_17692_n5470;
  wire _abc_17692_n5471;
  wire _abc_17692_n5472;
  wire _abc_17692_n5473;
  wire _abc_17692_n5474;
  wire _abc_17692_n5475;
  wire _abc_17692_n5476;
  wire _abc_17692_n5477;
  wire _abc_17692_n5478;
  wire _abc_17692_n5479;
  wire _abc_17692_n5480;
  wire _abc_17692_n5481;
  wire _abc_17692_n5482;
  wire _abc_17692_n5483;
  wire _abc_17692_n5484;
  wire _abc_17692_n5485;
  wire _abc_17692_n5486;
  wire _abc_17692_n5487;
  wire _abc_17692_n5488;
  wire _abc_17692_n5489;
  wire _abc_17692_n5490;
  wire _abc_17692_n5491;
  wire _abc_17692_n5492;
  wire _abc_17692_n5493;
  wire _abc_17692_n5494;
  wire _abc_17692_n5495;
  wire _abc_17692_n5496;
  wire _abc_17692_n5497;
  wire _abc_17692_n5498;
  wire _abc_17692_n5499;
  wire _abc_17692_n5500;
  wire _abc_17692_n5501;
  wire _abc_17692_n5502;
  wire _abc_17692_n5503;
  wire _abc_17692_n5504;
  wire _abc_17692_n5505;
  wire _abc_17692_n5506;
  wire _abc_17692_n5507;
  wire _abc_17692_n5508;
  wire _abc_17692_n5509;
  wire _abc_17692_n5510;
  wire _abc_17692_n5511;
  wire _abc_17692_n5512;
  wire _abc_17692_n5513;
  wire _abc_17692_n5514;
  wire _abc_17692_n5515;
  wire _abc_17692_n5516;
  wire _abc_17692_n5517;
  wire _abc_17692_n5518;
  wire _abc_17692_n5519;
  wire _abc_17692_n5520;
  wire _abc_17692_n5521;
  wire _abc_17692_n5522;
  wire _abc_17692_n5523;
  wire _abc_17692_n5524;
  wire _abc_17692_n5525;
  wire _abc_17692_n5526;
  wire _abc_17692_n5527;
  wire _abc_17692_n5528;
  wire _abc_17692_n5529;
  wire _abc_17692_n5530;
  wire _abc_17692_n5531;
  wire _abc_17692_n5532;
  wire _abc_17692_n5533;
  wire _abc_17692_n5534;
  wire _abc_17692_n5535;
  wire _abc_17692_n5536;
  wire _abc_17692_n5537;
  wire _abc_17692_n5538;
  wire _abc_17692_n5539;
  wire _abc_17692_n5540;
  wire _abc_17692_n5541;
  wire _abc_17692_n5542;
  wire _abc_17692_n5543;
  wire _abc_17692_n5544;
  wire _abc_17692_n5545_1;
  wire _abc_17692_n5546;
  wire _abc_17692_n5547;
  wire _abc_17692_n5548_1;
  wire _abc_17692_n5549;
  wire _abc_17692_n5550;
  wire _abc_17692_n5551;
  wire _abc_17692_n5552;
  wire _abc_17692_n5553;
  wire _abc_17692_n5554;
  wire _abc_17692_n5555;
  wire _abc_17692_n5556;
  wire _abc_17692_n5557;
  wire _abc_17692_n5558;
  wire _abc_17692_n5559;
  wire _abc_17692_n5560;
  wire _abc_17692_n5561;
  wire _abc_17692_n5562;
  wire _abc_17692_n5563;
  wire _abc_17692_n5564;
  wire _abc_17692_n5565;
  wire _abc_17692_n5566;
  wire _abc_17692_n5567;
  wire _abc_17692_n5568;
  wire _abc_17692_n5569;
  wire _abc_17692_n5570;
  wire _abc_17692_n5571;
  wire _abc_17692_n5572;
  wire _abc_17692_n5573;
  wire _abc_17692_n5574;
  wire _abc_17692_n5575;
  wire _abc_17692_n5576;
  wire _abc_17692_n5577;
  wire _abc_17692_n5578;
  wire _abc_17692_n5579;
  wire _abc_17692_n5580;
  wire _abc_17692_n5581;
  wire _abc_17692_n5582;
  wire _abc_17692_n5583;
  wire _abc_17692_n5584;
  wire _abc_17692_n5585;
  wire _abc_17692_n5586;
  wire _abc_17692_n5587;
  wire _abc_17692_n5588;
  wire _abc_17692_n5589;
  wire _abc_17692_n5590;
  wire _abc_17692_n5591;
  wire _abc_17692_n5592;
  wire _abc_17692_n5593;
  wire _abc_17692_n5595;
  wire _abc_17692_n5596;
  wire _abc_17692_n5597;
  wire _abc_17692_n5598;
  wire _abc_17692_n5599;
  wire _abc_17692_n5600;
  wire _abc_17692_n5601;
  wire _abc_17692_n5602;
  wire _abc_17692_n5603;
  wire _abc_17692_n5604;
  wire _abc_17692_n5605;
  wire _abc_17692_n5606;
  wire _abc_17692_n5607;
  wire _abc_17692_n5608_1;
  wire _abc_17692_n5609;
  wire _abc_17692_n5610;
  wire _abc_17692_n5611_1;
  wire _abc_17692_n5612;
  wire _abc_17692_n5613;
  wire _abc_17692_n5614;
  wire _abc_17692_n5615;
  wire _abc_17692_n5616;
  wire _abc_17692_n5617;
  wire _abc_17692_n5618;
  wire _abc_17692_n5619;
  wire _abc_17692_n5620;
  wire _abc_17692_n5621;
  wire _abc_17692_n5622;
  wire _abc_17692_n5623;
  wire _abc_17692_n5624;
  wire _abc_17692_n5625;
  wire _abc_17692_n5626;
  wire _abc_17692_n5627;
  wire _abc_17692_n5628;
  wire _abc_17692_n5629;
  wire _abc_17692_n5630;
  wire _abc_17692_n5631;
  wire _abc_17692_n5632;
  wire _abc_17692_n5633;
  wire _abc_17692_n5634;
  wire _abc_17692_n5635;
  wire _abc_17692_n5636;
  wire _abc_17692_n5637;
  wire _abc_17692_n5638;
  wire _abc_17692_n5639;
  wire _abc_17692_n5640;
  wire _abc_17692_n5641;
  wire _abc_17692_n5642;
  wire _abc_17692_n5643;
  wire _abc_17692_n5644;
  wire _abc_17692_n5645;
  wire _abc_17692_n5646;
  wire _abc_17692_n5647;
  wire _abc_17692_n5648;
  wire _abc_17692_n5649;
  wire _abc_17692_n5650;
  wire _abc_17692_n5651;
  wire _abc_17692_n5652;
  wire _abc_17692_n5653;
  wire _abc_17692_n5654;
  wire _abc_17692_n5655;
  wire _abc_17692_n5656;
  wire _abc_17692_n5657;
  wire _abc_17692_n5658;
  wire _abc_17692_n5659;
  wire _abc_17692_n5660;
  wire _abc_17692_n5661;
  wire _abc_17692_n5662;
  wire _abc_17692_n5663;
  wire _abc_17692_n5664;
  wire _abc_17692_n5665;
  wire _abc_17692_n5666;
  wire _abc_17692_n5667;
  wire _abc_17692_n5668;
  wire _abc_17692_n5669;
  wire _abc_17692_n5670;
  wire _abc_17692_n5671;
  wire _abc_17692_n5672;
  wire _abc_17692_n5673;
  wire _abc_17692_n5674;
  wire _abc_17692_n5675;
  wire _abc_17692_n5676;
  wire _abc_17692_n5677;
  wire _abc_17692_n5678;
  wire _abc_17692_n5679;
  wire _abc_17692_n5680;
  wire _abc_17692_n5681;
  wire _abc_17692_n5682;
  wire _abc_17692_n5683;
  wire _abc_17692_n5684;
  wire _abc_17692_n5685;
  wire _abc_17692_n5686;
  wire _abc_17692_n5687;
  wire _abc_17692_n5688;
  wire _abc_17692_n5689;
  wire _abc_17692_n5690;
  wire _abc_17692_n5691;
  wire _abc_17692_n5692_1;
  wire _abc_17692_n5693;
  wire _abc_17692_n5694;
  wire _abc_17692_n5695_1;
  wire _abc_17692_n5696;
  wire _abc_17692_n5697;
  wire _abc_17692_n5698;
  wire _abc_17692_n5699;
  wire _abc_17692_n5700;
  wire _abc_17692_n5701;
  wire _abc_17692_n5702;
  wire _abc_17692_n5703;
  wire _abc_17692_n5704;
  wire _abc_17692_n5705;
  wire _abc_17692_n5706;
  wire _abc_17692_n5707;
  wire _abc_17692_n5708;
  wire _abc_17692_n5709;
  wire _abc_17692_n5710;
  wire _abc_17692_n5711;
  wire _abc_17692_n5712;
  wire _abc_17692_n5713;
  wire _abc_17692_n5714;
  wire _abc_17692_n5715;
  wire _abc_17692_n5716;
  wire _abc_17692_n5717;
  wire _abc_17692_n5718;
  wire _abc_17692_n5719;
  wire _abc_17692_n5720;
  wire _abc_17692_n5721;
  wire _abc_17692_n5722;
  wire _abc_17692_n5723;
  wire _abc_17692_n5724;
  wire _abc_17692_n5725;
  wire _abc_17692_n5726;
  wire _abc_17692_n5727;
  wire _abc_17692_n5728;
  wire _abc_17692_n5729;
  wire _abc_17692_n5730;
  wire _abc_17692_n5731;
  wire _abc_17692_n5732;
  wire _abc_17692_n5733;
  wire _abc_17692_n5734;
  wire _abc_17692_n5735;
  wire _abc_17692_n5736;
  wire _abc_17692_n5737;
  wire _abc_17692_n5738;
  wire _abc_17692_n5739;
  wire _abc_17692_n5740;
  wire _abc_17692_n5741;
  wire _abc_17692_n5742;
  wire _abc_17692_n5743;
  wire _abc_17692_n5744;
  wire _abc_17692_n5745_1;
  wire _abc_17692_n5746;
  wire _abc_17692_n5747;
  wire _abc_17692_n5748_1;
  wire _abc_17692_n5749;
  wire _abc_17692_n5750;
  wire _abc_17692_n5751;
  wire _abc_17692_n5752;
  wire _abc_17692_n5753;
  wire _abc_17692_n5754;
  wire _abc_17692_n5755;
  wire _abc_17692_n5756;
  wire _abc_17692_n5757;
  wire _abc_17692_n5758;
  wire _abc_17692_n5759;
  wire _abc_17692_n5760;
  wire _abc_17692_n5761;
  wire _abc_17692_n5762;
  wire _abc_17692_n5763;
  wire _abc_17692_n5764;
  wire _abc_17692_n5765;
  wire _abc_17692_n5766;
  wire _abc_17692_n5767;
  wire _abc_17692_n5769;
  wire _abc_17692_n5770;
  wire _abc_17692_n5771;
  wire _abc_17692_n5772;
  wire _abc_17692_n5773;
  wire _abc_17692_n5774;
  wire _abc_17692_n5775;
  wire _abc_17692_n5776;
  wire _abc_17692_n5777;
  wire _abc_17692_n5778;
  wire _abc_17692_n5779;
  wire _abc_17692_n5780;
  wire _abc_17692_n5781;
  wire _abc_17692_n5782;
  wire _abc_17692_n5783;
  wire _abc_17692_n5784;
  wire _abc_17692_n5785;
  wire _abc_17692_n5786;
  wire _abc_17692_n5787;
  wire _abc_17692_n5788;
  wire _abc_17692_n5789;
  wire _abc_17692_n5790;
  wire _abc_17692_n5791;
  wire _abc_17692_n5792;
  wire _abc_17692_n5793;
  wire _abc_17692_n5794;
  wire _abc_17692_n5795;
  wire _abc_17692_n5796;
  wire _abc_17692_n5797;
  wire _abc_17692_n5798;
  wire _abc_17692_n5799;
  wire _abc_17692_n5800;
  wire _abc_17692_n5801;
  wire _abc_17692_n5802;
  wire _abc_17692_n5803;
  wire _abc_17692_n5804;
  wire _abc_17692_n5805;
  wire _abc_17692_n5806;
  wire _abc_17692_n5807;
  wire _abc_17692_n5808;
  wire _abc_17692_n5809;
  wire _abc_17692_n5810;
  wire _abc_17692_n5811;
  wire _abc_17692_n5812;
  wire _abc_17692_n5813;
  wire _abc_17692_n5814;
  wire _abc_17692_n5815;
  wire _abc_17692_n5816;
  wire _abc_17692_n5817;
  wire _abc_17692_n5818;
  wire _abc_17692_n5819;
  wire _abc_17692_n5820;
  wire _abc_17692_n5821;
  wire _abc_17692_n5822;
  wire _abc_17692_n5823;
  wire _abc_17692_n5824;
  wire _abc_17692_n5825;
  wire _abc_17692_n5826;
  wire _abc_17692_n5827;
  wire _abc_17692_n5828;
  wire _abc_17692_n5829;
  wire _abc_17692_n5830;
  wire _abc_17692_n5831;
  wire _abc_17692_n5832;
  wire _abc_17692_n5833;
  wire _abc_17692_n5834;
  wire _abc_17692_n5835;
  wire _abc_17692_n5836;
  wire _abc_17692_n5837;
  wire _abc_17692_n5838;
  wire _abc_17692_n5839;
  wire _abc_17692_n5840;
  wire _abc_17692_n5841;
  wire _abc_17692_n5842;
  wire _abc_17692_n5843_1;
  wire _abc_17692_n5844;
  wire _abc_17692_n5845;
  wire _abc_17692_n5846_1;
  wire _abc_17692_n5847;
  wire _abc_17692_n5848;
  wire _abc_17692_n5849;
  wire _abc_17692_n5850;
  wire _abc_17692_n5851;
  wire _abc_17692_n5852;
  wire _abc_17692_n5853;
  wire _abc_17692_n5854;
  wire _abc_17692_n5855;
  wire _abc_17692_n5856;
  wire _abc_17692_n5857;
  wire _abc_17692_n5858;
  wire _abc_17692_n5859;
  wire _abc_17692_n5860;
  wire _abc_17692_n5861;
  wire _abc_17692_n5862;
  wire _abc_17692_n5863;
  wire _abc_17692_n5864;
  wire _abc_17692_n5865;
  wire _abc_17692_n5866;
  wire _abc_17692_n5867;
  wire _abc_17692_n5868;
  wire _abc_17692_n5869;
  wire _abc_17692_n5870;
  wire _abc_17692_n5871;
  wire _abc_17692_n5872;
  wire _abc_17692_n5873;
  wire _abc_17692_n5874;
  wire _abc_17692_n5875;
  wire _abc_17692_n5876;
  wire _abc_17692_n5877;
  wire _abc_17692_n5878;
  wire _abc_17692_n5879;
  wire _abc_17692_n5880;
  wire _abc_17692_n5881;
  wire _abc_17692_n5882;
  wire _abc_17692_n5883;
  wire _abc_17692_n5884;
  wire _abc_17692_n5885;
  wire _abc_17692_n5886;
  wire _abc_17692_n5887;
  wire _abc_17692_n5888;
  wire _abc_17692_n5889;
  wire _abc_17692_n5890;
  wire _abc_17692_n5891;
  wire _abc_17692_n5892;
  wire _abc_17692_n5893;
  wire _abc_17692_n5894;
  wire _abc_17692_n5895;
  wire _abc_17692_n5896;
  wire _abc_17692_n5897;
  wire _abc_17692_n5898;
  wire _abc_17692_n5899;
  wire _abc_17692_n5900_1;
  wire _abc_17692_n5901;
  wire _abc_17692_n5902;
  wire _abc_17692_n5903_1;
  wire _abc_17692_n5904;
  wire _abc_17692_n5905;
  wire _abc_17692_n5906;
  wire _abc_17692_n5907;
  wire _abc_17692_n5908;
  wire _abc_17692_n5909;
  wire _abc_17692_n5910;
  wire _abc_17692_n5911;
  wire _abc_17692_n5912;
  wire _abc_17692_n5913;
  wire _abc_17692_n5914;
  wire _abc_17692_n5915;
  wire _abc_17692_n5916;
  wire _abc_17692_n5917;
  wire _abc_17692_n5918;
  wire _abc_17692_n5919;
  wire _abc_17692_n5920;
  wire _abc_17692_n5921;
  wire _abc_17692_n5922;
  wire _abc_17692_n5923;
  wire _abc_17692_n5924;
  wire _abc_17692_n5925;
  wire _abc_17692_n5926;
  wire _abc_17692_n5927;
  wire _abc_17692_n5928;
  wire _abc_17692_n5929;
  wire _abc_17692_n5930;
  wire _abc_17692_n5931;
  wire _abc_17692_n5932;
  wire _abc_17692_n5933;
  wire _abc_17692_n5934;
  wire _abc_17692_n5935;
  wire _abc_17692_n5936;
  wire _abc_17692_n5937;
  wire _abc_17692_n5938;
  wire _abc_17692_n5939;
  wire _abc_17692_n5940;
  wire _abc_17692_n5941;
  wire _abc_17692_n5942;
  wire _abc_17692_n5943;
  wire _abc_17692_n5944;
  wire _abc_17692_n5945;
  wire _abc_17692_n5946;
  wire _abc_17692_n5947;
  wire _abc_17692_n5948;
  wire _abc_17692_n5949;
  wire _abc_17692_n5950;
  wire _abc_17692_n5951;
  wire _abc_17692_n5952;
  wire _abc_17692_n5953;
  wire _abc_17692_n5954;
  wire _abc_17692_n5955;
  wire _abc_17692_n5956;
  wire _abc_17692_n5957;
  wire _abc_17692_n5958;
  wire _abc_17692_n5959;
  wire _abc_17692_n5960;
  wire _abc_17692_n5961;
  wire _abc_17692_n5962;
  wire _abc_17692_n5963;
  wire _abc_17692_n5964;
  wire _abc_17692_n5965;
  wire _abc_17692_n5966;
  wire _abc_17692_n5967;
  wire _abc_17692_n5968;
  wire _abc_17692_n5969;
  wire _abc_17692_n5970;
  wire _abc_17692_n5971;
  wire _abc_17692_n5972;
  wire _abc_17692_n5973;
  wire _abc_17692_n5974;
  wire _abc_17692_n5975;
  wire _abc_17692_n5976;
  wire _abc_17692_n5977;
  wire _abc_17692_n5978;
  wire _abc_17692_n5979;
  wire _abc_17692_n5980;
  wire _abc_17692_n5981_1;
  wire _abc_17692_n5982;
  wire _abc_17692_n5983;
  wire _abc_17692_n5984_1;
  wire _abc_17692_n5985;
  wire _abc_17692_n5986;
  wire _abc_17692_n5987;
  wire _abc_17692_n5988;
  wire _abc_17692_n5989;
  wire _abc_17692_n5990;
  wire _abc_17692_n5991;
  wire _abc_17692_n5992;
  wire _abc_17692_n5993;
  wire _abc_17692_n5994;
  wire _abc_17692_n5995;
  wire _abc_17692_n5996;
  wire _abc_17692_n5997;
  wire _abc_17692_n5998;
  wire _abc_17692_n5999;
  wire _abc_17692_n6000;
  wire _abc_17692_n6001;
  wire _abc_17692_n6002;
  wire _abc_17692_n6003;
  wire _abc_17692_n6004;
  wire _abc_17692_n6005;
  wire _abc_17692_n6006;
  wire _abc_17692_n6007;
  wire _abc_17692_n6008;
  wire _abc_17692_n6009;
  wire _abc_17692_n6010;
  wire _abc_17692_n6011;
  wire _abc_17692_n6012;
  wire _abc_17692_n6013;
  wire _abc_17692_n6014;
  wire _abc_17692_n6015;
  wire _abc_17692_n6016;
  wire _abc_17692_n6017;
  wire _abc_17692_n6018;
  wire _abc_17692_n6019;
  wire _abc_17692_n6020;
  wire _abc_17692_n6021;
  wire _abc_17692_n6022;
  wire _abc_17692_n6023;
  wire _abc_17692_n6024;
  wire _abc_17692_n6025;
  wire _abc_17692_n6026;
  wire _abc_17692_n6027;
  wire _abc_17692_n6028;
  wire _abc_17692_n6029;
  wire _abc_17692_n6030;
  wire _abc_17692_n6031;
  wire _abc_17692_n6032;
  wire _abc_17692_n6033;
  wire _abc_17692_n6034;
  wire _abc_17692_n6035;
  wire _abc_17692_n6036;
  wire _abc_17692_n6037;
  wire _abc_17692_n6038_1;
  wire _abc_17692_n6039;
  wire _abc_17692_n6040;
  wire _abc_17692_n6041_1;
  wire _abc_17692_n6042;
  wire _abc_17692_n6043;
  wire _abc_17692_n6044;
  wire _abc_17692_n6045;
  wire _abc_17692_n6046;
  wire _abc_17692_n6047;
  wire _abc_17692_n6048;
  wire _abc_17692_n6049;
  wire _abc_17692_n6050;
  wire _abc_17692_n6051;
  wire _abc_17692_n6052;
  wire _abc_17692_n6053;
  wire _abc_17692_n6054;
  wire _abc_17692_n6055;
  wire _abc_17692_n6056;
  wire _abc_17692_n6057;
  wire _abc_17692_n6058;
  wire _abc_17692_n6059;
  wire _abc_17692_n6060;
  wire _abc_17692_n6062;
  wire _abc_17692_n6063;
  wire _abc_17692_n6064;
  wire _abc_17692_n6065;
  wire _abc_17692_n6066;
  wire _abc_17692_n6067;
  wire _abc_17692_n6068;
  wire _abc_17692_n6069;
  wire _abc_17692_n6070;
  wire _abc_17692_n6071;
  wire _abc_17692_n6072;
  wire _abc_17692_n6073;
  wire _abc_17692_n6074;
  wire _abc_17692_n6075;
  wire _abc_17692_n6076;
  wire _abc_17692_n6077;
  wire _abc_17692_n6078;
  wire _abc_17692_n6079;
  wire _abc_17692_n6080;
  wire _abc_17692_n6081;
  wire _abc_17692_n6082;
  wire _abc_17692_n6083;
  wire _abc_17692_n6084;
  wire _abc_17692_n6085;
  wire _abc_17692_n6086;
  wire _abc_17692_n6087;
  wire _abc_17692_n6088;
  wire _abc_17692_n6089;
  wire _abc_17692_n6090;
  wire _abc_17692_n6091;
  wire _abc_17692_n6092;
  wire _abc_17692_n6093;
  wire _abc_17692_n6094;
  wire _abc_17692_n6095;
  wire _abc_17692_n6096;
  wire _abc_17692_n6097;
  wire _abc_17692_n6098;
  wire _abc_17692_n6099;
  wire _abc_17692_n6100;
  wire _abc_17692_n6101;
  wire _abc_17692_n6102;
  wire _abc_17692_n6103;
  wire _abc_17692_n6104;
  wire _abc_17692_n6105;
  wire _abc_17692_n6106;
  wire _abc_17692_n6107;
  wire _abc_17692_n6108;
  wire _abc_17692_n6109;
  wire _abc_17692_n6110;
  wire _abc_17692_n6111;
  wire _abc_17692_n6112;
  wire _abc_17692_n6113;
  wire _abc_17692_n6114;
  wire _abc_17692_n6115;
  wire _abc_17692_n6116;
  wire _abc_17692_n6117;
  wire _abc_17692_n6118;
  wire _abc_17692_n6119;
  wire _abc_17692_n6120;
  wire _abc_17692_n6121;
  wire _abc_17692_n6122;
  wire _abc_17692_n6123;
  wire _abc_17692_n6124;
  wire _abc_17692_n6125;
  wire _abc_17692_n6126;
  wire _abc_17692_n6127;
  wire _abc_17692_n6128;
  wire _abc_17692_n6129;
  wire _abc_17692_n6130;
  wire _abc_17692_n6131;
  wire _abc_17692_n6132;
  wire _abc_17692_n6133;
  wire _abc_17692_n6134;
  wire _abc_17692_n6135;
  wire _abc_17692_n6136;
  wire _abc_17692_n6137;
  wire _abc_17692_n6138;
  wire _abc_17692_n6139;
  wire _abc_17692_n6140;
  wire _abc_17692_n6141;
  wire _abc_17692_n6142;
  wire _abc_17692_n6143;
  wire _abc_17692_n6144;
  wire _abc_17692_n6145;
  wire _abc_17692_n6146;
  wire _abc_17692_n6147;
  wire _abc_17692_n6148;
  wire _abc_17692_n6149;
  wire _abc_17692_n6150;
  wire _abc_17692_n6151;
  wire _abc_17692_n6152;
  wire _abc_17692_n6153;
  wire _abc_17692_n6154;
  wire _abc_17692_n6155;
  wire _abc_17692_n6156;
  wire _abc_17692_n6157;
  wire _abc_17692_n6158;
  wire _abc_17692_n6159;
  wire _abc_17692_n6160;
  wire _abc_17692_n6161;
  wire _abc_17692_n6162;
  wire _abc_17692_n6163;
  wire _abc_17692_n6164;
  wire _abc_17692_n6165;
  wire _abc_17692_n6166_1;
  wire _abc_17692_n6167;
  wire _abc_17692_n6168;
  wire _abc_17692_n6169_1;
  wire _abc_17692_n6170;
  wire _abc_17692_n6171;
  wire _abc_17692_n6172;
  wire _abc_17692_n6173;
  wire _abc_17692_n6174;
  wire _abc_17692_n6175;
  wire _abc_17692_n6176;
  wire _abc_17692_n6177;
  wire _abc_17692_n6178;
  wire _abc_17692_n6179;
  wire _abc_17692_n6180;
  wire _abc_17692_n6181;
  wire _abc_17692_n6182;
  wire _abc_17692_n6183;
  wire _abc_17692_n6184;
  wire _abc_17692_n6185;
  wire _abc_17692_n6186;
  wire _abc_17692_n6187;
  wire _abc_17692_n6188;
  wire _abc_17692_n6189;
  wire _abc_17692_n6190;
  wire _abc_17692_n6191;
  wire _abc_17692_n6192;
  wire _abc_17692_n6193;
  wire _abc_17692_n6194;
  wire _abc_17692_n6195;
  wire _abc_17692_n6196;
  wire _abc_17692_n6197;
  wire _abc_17692_n6198;
  wire _abc_17692_n6199;
  wire _abc_17692_n6200;
  wire _abc_17692_n6201;
  wire _abc_17692_n6202;
  wire _abc_17692_n6203;
  wire _abc_17692_n6204;
  wire _abc_17692_n6205;
  wire _abc_17692_n6206;
  wire _abc_17692_n6207;
  wire _abc_17692_n6208;
  wire _abc_17692_n6209;
  wire _abc_17692_n6210;
  wire _abc_17692_n6211;
  wire _abc_17692_n6212;
  wire _abc_17692_n6213;
  wire _abc_17692_n6214;
  wire _abc_17692_n6215;
  wire _abc_17692_n6216;
  wire _abc_17692_n6217;
  wire _abc_17692_n6218;
  wire _abc_17692_n6219;
  wire _abc_17692_n6220;
  wire _abc_17692_n6221;
  wire _abc_17692_n6222_1;
  wire _abc_17692_n6223;
  wire _abc_17692_n6224;
  wire _abc_17692_n6225_1;
  wire _abc_17692_n6226;
  wire _abc_17692_n6227;
  wire _abc_17692_n6228;
  wire _abc_17692_n6229;
  wire _abc_17692_n623;
  wire _abc_17692_n6230;
  wire _abc_17692_n6231;
  wire _abc_17692_n6232;
  wire _abc_17692_n6233;
  wire _abc_17692_n6234;
  wire _abc_17692_n6236;
  wire _abc_17692_n6237;
  wire _abc_17692_n6238;
  wire _abc_17692_n6239;
  wire _abc_17692_n624;
  wire _abc_17692_n6240;
  wire _abc_17692_n6241;
  wire _abc_17692_n6242;
  wire _abc_17692_n6243;
  wire _abc_17692_n6244;
  wire _abc_17692_n6245;
  wire _abc_17692_n6246;
  wire _abc_17692_n6247;
  wire _abc_17692_n6248;
  wire _abc_17692_n6249;
  wire _abc_17692_n6250;
  wire _abc_17692_n6251;
  wire _abc_17692_n6252;
  wire _abc_17692_n6253;
  wire _abc_17692_n6254;
  wire _abc_17692_n6255;
  wire _abc_17692_n6256;
  wire _abc_17692_n6257;
  wire _abc_17692_n6258;
  wire _abc_17692_n6259;
  wire _abc_17692_n626;
  wire _abc_17692_n6260;
  wire _abc_17692_n6261;
  wire _abc_17692_n6262;
  wire _abc_17692_n6263;
  wire _abc_17692_n6264;
  wire _abc_17692_n6265;
  wire _abc_17692_n6266;
  wire _abc_17692_n6267;
  wire _abc_17692_n6268;
  wire _abc_17692_n6269;
  wire _abc_17692_n627;
  wire _abc_17692_n6270;
  wire _abc_17692_n6271;
  wire _abc_17692_n6272;
  wire _abc_17692_n6273;
  wire _abc_17692_n6274;
  wire _abc_17692_n6275;
  wire _abc_17692_n6276;
  wire _abc_17692_n6277;
  wire _abc_17692_n6278;
  wire _abc_17692_n6279;
  wire _abc_17692_n628;
  wire _abc_17692_n6280;
  wire _abc_17692_n6281;
  wire _abc_17692_n6282;
  wire _abc_17692_n6283;
  wire _abc_17692_n6284;
  wire _abc_17692_n6285;
  wire _abc_17692_n6286;
  wire _abc_17692_n6287;
  wire _abc_17692_n6288;
  wire _abc_17692_n6289;
  wire _abc_17692_n629;
  wire _abc_17692_n6290;
  wire _abc_17692_n6291;
  wire _abc_17692_n6292;
  wire _abc_17692_n6293;
  wire _abc_17692_n6294;
  wire _abc_17692_n6295;
  wire _abc_17692_n6296;
  wire _abc_17692_n6297;
  wire _abc_17692_n6298;
  wire _abc_17692_n6299;
  wire _abc_17692_n6300;
  wire _abc_17692_n6301;
  wire _abc_17692_n6302;
  wire _abc_17692_n6303;
  wire _abc_17692_n6304;
  wire _abc_17692_n6305;
  wire _abc_17692_n6306;
  wire _abc_17692_n6307;
  wire _abc_17692_n6308;
  wire _abc_17692_n6309;
  wire _abc_17692_n631;
  wire _abc_17692_n6310;
  wire _abc_17692_n6311;
  wire _abc_17692_n6312;
  wire _abc_17692_n6313;
  wire _abc_17692_n6314;
  wire _abc_17692_n6315;
  wire _abc_17692_n6316_1;
  wire _abc_17692_n6317;
  wire _abc_17692_n6318;
  wire _abc_17692_n6319_1;
  wire _abc_17692_n632;
  wire _abc_17692_n6320;
  wire _abc_17692_n6321;
  wire _abc_17692_n6322;
  wire _abc_17692_n6323;
  wire _abc_17692_n6324;
  wire _abc_17692_n6325;
  wire _abc_17692_n6326;
  wire _abc_17692_n6327;
  wire _abc_17692_n6328;
  wire _abc_17692_n6329;
  wire _abc_17692_n633;
  wire _abc_17692_n6330;
  wire _abc_17692_n6331;
  wire _abc_17692_n6332;
  wire _abc_17692_n6333;
  wire _abc_17692_n6334;
  wire _abc_17692_n6335;
  wire _abc_17692_n6336;
  wire _abc_17692_n6337;
  wire _abc_17692_n6338;
  wire _abc_17692_n6339;
  wire _abc_17692_n6340;
  wire _abc_17692_n6341;
  wire _abc_17692_n6342;
  wire _abc_17692_n6343;
  wire _abc_17692_n6344;
  wire _abc_17692_n6345;
  wire _abc_17692_n6346;
  wire _abc_17692_n6347;
  wire _abc_17692_n6348;
  wire _abc_17692_n6349;
  wire _abc_17692_n6350;
  wire _abc_17692_n6351;
  wire _abc_17692_n6352;
  wire _abc_17692_n6353;
  wire _abc_17692_n6354;
  wire _abc_17692_n6355;
  wire _abc_17692_n6356;
  wire _abc_17692_n6357;
  wire _abc_17692_n6358;
  wire _abc_17692_n6359;
  wire _abc_17692_n6360;
  wire _abc_17692_n6361;
  wire _abc_17692_n6362;
  wire _abc_17692_n6363;
  wire _abc_17692_n6364;
  wire _abc_17692_n6365;
  wire _abc_17692_n6366;
  wire _abc_17692_n6367;
  wire _abc_17692_n6368;
  wire _abc_17692_n6369;
  wire _abc_17692_n6370;
  wire _abc_17692_n6371_1;
  wire _abc_17692_n6372;
  wire _abc_17692_n6373;
  wire _abc_17692_n6374_1;
  wire _abc_17692_n6375;
  wire _abc_17692_n6376;
  wire _abc_17692_n6377;
  wire _abc_17692_n6378;
  wire _abc_17692_n6379;
  wire _abc_17692_n6380;
  wire _abc_17692_n6381;
  wire _abc_17692_n6382;
  wire _abc_17692_n6383;
  wire _abc_17692_n6384;
  wire _abc_17692_n6385;
  wire _abc_17692_n6386;
  wire _abc_17692_n6387;
  wire _abc_17692_n6388;
  wire _abc_17692_n6389;
  wire _abc_17692_n6390;
  wire _abc_17692_n6391;
  wire _abc_17692_n6392;
  wire _abc_17692_n6393;
  wire _abc_17692_n6394;
  wire _abc_17692_n6395;
  wire _abc_17692_n6396;
  wire _abc_17692_n6397;
  wire _abc_17692_n6398;
  wire _abc_17692_n6399;
  wire _abc_17692_n6400;
  wire _abc_17692_n6401;
  wire _abc_17692_n6402;
  wire _abc_17692_n6403;
  wire _abc_17692_n6404;
  wire _abc_17692_n6405;
  wire _abc_17692_n6406;
  wire _abc_17692_n6407;
  wire _abc_17692_n6408;
  wire _abc_17692_n6409;
  wire _abc_17692_n6410;
  wire _abc_17692_n6411;
  wire _abc_17692_n6412;
  wire _abc_17692_n6413;
  wire _abc_17692_n6414;
  wire _abc_17692_n6415;
  wire _abc_17692_n6416;
  wire _abc_17692_n6417;
  wire _abc_17692_n6418;
  wire _abc_17692_n6419;
  wire _abc_17692_n6420;
  wire _abc_17692_n6421;
  wire _abc_17692_n6422;
  wire _abc_17692_n6423;
  wire _abc_17692_n6424;
  wire _abc_17692_n6425;
  wire _abc_17692_n6426;
  wire _abc_17692_n6427;
  wire _abc_17692_n6428;
  wire _abc_17692_n6429;
  wire _abc_17692_n6430;
  wire _abc_17692_n6431;
  wire _abc_17692_n6432;
  wire _abc_17692_n6433;
  wire _abc_17692_n6434;
  wire _abc_17692_n6435;
  wire _abc_17692_n6436;
  wire _abc_17692_n6437;
  wire _abc_17692_n6438;
  wire _abc_17692_n6439;
  wire _abc_17692_n6440;
  wire _abc_17692_n6441;
  wire _abc_17692_n6442;
  wire _abc_17692_n6443;
  wire _abc_17692_n6444;
  wire _abc_17692_n6445;
  wire _abc_17692_n6446;
  wire _abc_17692_n6447;
  wire _abc_17692_n6448;
  wire _abc_17692_n6449;
  wire _abc_17692_n6450;
  wire _abc_17692_n6451;
  wire _abc_17692_n6452;
  wire _abc_17692_n6453;
  wire _abc_17692_n6454;
  wire _abc_17692_n6455;
  wire _abc_17692_n6456;
  wire _abc_17692_n6457;
  wire _abc_17692_n6458;
  wire _abc_17692_n6459;
  wire _abc_17692_n6460;
  wire _abc_17692_n6461;
  wire _abc_17692_n6462;
  wire _abc_17692_n6463;
  wire _abc_17692_n6464;
  wire _abc_17692_n6466;
  wire _abc_17692_n6467;
  wire _abc_17692_n6468_1;
  wire _abc_17692_n6469;
  wire _abc_17692_n6470;
  wire _abc_17692_n6471;
  wire _abc_17692_n6472;
  wire _abc_17692_n6473;
  wire _abc_17692_n6474;
  wire _abc_17692_n6475;
  wire _abc_17692_n6476;
  wire _abc_17692_n6477;
  wire _abc_17692_n6478;
  wire _abc_17692_n6479;
  wire _abc_17692_n6480;
  wire _abc_17692_n6481;
  wire _abc_17692_n6482;
  wire _abc_17692_n6483;
  wire _abc_17692_n6484;
  wire _abc_17692_n6485;
  wire _abc_17692_n6486;
  wire _abc_17692_n6487;
  wire _abc_17692_n6488;
  wire _abc_17692_n6489;
  wire _abc_17692_n6490;
  wire _abc_17692_n6491;
  wire _abc_17692_n6492;
  wire _abc_17692_n6493;
  wire _abc_17692_n6494;
  wire _abc_17692_n6495;
  wire _abc_17692_n6496;
  wire _abc_17692_n6497;
  wire _abc_17692_n6498;
  wire _abc_17692_n6499;
  wire _abc_17692_n6500;
  wire _abc_17692_n6501;
  wire _abc_17692_n6502;
  wire _abc_17692_n6503;
  wire _abc_17692_n6504;
  wire _abc_17692_n6505;
  wire _abc_17692_n6506;
  wire _abc_17692_n6507;
  wire _abc_17692_n6508;
  wire _abc_17692_n6509;
  wire _abc_17692_n6510;
  wire _abc_17692_n6511;
  wire _abc_17692_n6512;
  wire _abc_17692_n6513;
  wire _abc_17692_n6514;
  wire _abc_17692_n6515;
  wire _abc_17692_n6516;
  wire _abc_17692_n6517;
  wire _abc_17692_n6518;
  wire _abc_17692_n6519;
  wire _abc_17692_n6520;
  wire _abc_17692_n6521;
  wire _abc_17692_n6522;
  wire _abc_17692_n6523_1;
  wire _abc_17692_n6524;
  wire _abc_17692_n6525;
  wire _abc_17692_n6526_1;
  wire _abc_17692_n6527;
  wire _abc_17692_n6528;
  wire _abc_17692_n6529;
  wire _abc_17692_n6530;
  wire _abc_17692_n6531;
  wire _abc_17692_n6532;
  wire _abc_17692_n6533;
  wire _abc_17692_n6534;
  wire _abc_17692_n6535;
  wire _abc_17692_n6536;
  wire _abc_17692_n6537;
  wire _abc_17692_n6538;
  wire _abc_17692_n6539;
  wire _abc_17692_n6540;
  wire _abc_17692_n6541;
  wire _abc_17692_n6542;
  wire _abc_17692_n6543;
  wire _abc_17692_n6544;
  wire _abc_17692_n6545;
  wire _abc_17692_n6546;
  wire _abc_17692_n6547;
  wire _abc_17692_n6548;
  wire _abc_17692_n6549;
  wire _abc_17692_n6550;
  wire _abc_17692_n6551;
  wire _abc_17692_n6552;
  wire _abc_17692_n6553;
  wire _abc_17692_n6554;
  wire _abc_17692_n6555;
  wire _abc_17692_n6556;
  wire _abc_17692_n6557;
  wire _abc_17692_n6558;
  wire _abc_17692_n6559;
  wire _abc_17692_n6560;
  wire _abc_17692_n6561;
  wire _abc_17692_n6562;
  wire _abc_17692_n6563;
  wire _abc_17692_n6564;
  wire _abc_17692_n6565;
  wire _abc_17692_n6566;
  wire _abc_17692_n6567;
  wire _abc_17692_n6568;
  wire _abc_17692_n6569;
  wire _abc_17692_n6570;
  wire _abc_17692_n6571;
  wire _abc_17692_n6572;
  wire _abc_17692_n6573;
  wire _abc_17692_n6574;
  wire _abc_17692_n6575;
  wire _abc_17692_n6576;
  wire _abc_17692_n6577;
  wire _abc_17692_n6578;
  wire _abc_17692_n6579;
  wire _abc_17692_n6580;
  wire _abc_17692_n6581;
  wire _abc_17692_n6582;
  wire _abc_17692_n6583;
  wire _abc_17692_n6584;
  wire _abc_17692_n6585;
  wire _abc_17692_n6586;
  wire _abc_17692_n6587;
  wire _abc_17692_n6588;
  wire _abc_17692_n6589;
  wire _abc_17692_n6590;
  wire _abc_17692_n6591;
  wire _abc_17692_n6592;
  wire _abc_17692_n6593;
  wire _abc_17692_n6594;
  wire _abc_17692_n6595;
  wire _abc_17692_n6596;
  wire _abc_17692_n6597_1;
  wire _abc_17692_n6598;
  wire _abc_17692_n6599;
  wire _abc_17692_n6600_1;
  wire _abc_17692_n6601;
  wire _abc_17692_n6602;
  wire _abc_17692_n6603;
  wire _abc_17692_n6604;
  wire _abc_17692_n6605;
  wire _abc_17692_n6606;
  wire _abc_17692_n6607;
  wire _abc_17692_n6608;
  wire _abc_17692_n6609;
  wire _abc_17692_n6610;
  wire _abc_17692_n6611;
  wire _abc_17692_n6612;
  wire _abc_17692_n6613;
  wire _abc_17692_n6614;
  wire _abc_17692_n6615;
  wire _abc_17692_n6616;
  wire _abc_17692_n6617;
  wire _abc_17692_n6618;
  wire _abc_17692_n6619;
  wire _abc_17692_n6620;
  wire _abc_17692_n6621;
  wire _abc_17692_n6622;
  wire _abc_17692_n6623;
  wire _abc_17692_n6624;
  wire _abc_17692_n6625;
  wire _abc_17692_n6626;
  wire _abc_17692_n6627;
  wire _abc_17692_n6628;
  wire _abc_17692_n6629;
  wire _abc_17692_n6630;
  wire _abc_17692_n6631;
  wire _abc_17692_n6632;
  wire _abc_17692_n6633;
  wire _abc_17692_n6634;
  wire _abc_17692_n6635;
  wire _abc_17692_n6636;
  wire _abc_17692_n6637;
  wire _abc_17692_n6638;
  wire _abc_17692_n6639;
  wire _abc_17692_n6640;
  wire _abc_17692_n6641;
  wire _abc_17692_n6642;
  wire _abc_17692_n6643;
  wire _abc_17692_n6644_1;
  wire _abc_17692_n6645;
  wire _abc_17692_n6646;
  wire _abc_17692_n6647_1;
  wire _abc_17692_n6648;
  wire _abc_17692_n6649;
  wire _abc_17692_n6650;
  wire _abc_17692_n6651;
  wire _abc_17692_n6652_1;
  wire _abc_17692_n6653;
  wire _abc_17692_n6654_1;
  wire _abc_17692_n6655;
  wire _abc_17692_n6657_1;
  wire _abc_17692_n6658_1;
  wire _abc_17692_n6659_1;
  wire _abc_17692_n6660;
  wire _abc_17692_n6660_1;
  wire _abc_17692_n6660_bF_buf0;
  wire _abc_17692_n6660_bF_buf1;
  wire _abc_17692_n6660_bF_buf10;
  wire _abc_17692_n6660_bF_buf11;
  wire _abc_17692_n6660_bF_buf12;
  wire _abc_17692_n6660_bF_buf13;
  wire _abc_17692_n6660_bF_buf2;
  wire _abc_17692_n6660_bF_buf3;
  wire _abc_17692_n6660_bF_buf4;
  wire _abc_17692_n6660_bF_buf5;
  wire _abc_17692_n6660_bF_buf6;
  wire _abc_17692_n6660_bF_buf7;
  wire _abc_17692_n6660_bF_buf8;
  wire _abc_17692_n6660_bF_buf9;
  wire _abc_17692_n6661;
  wire _abc_17692_n6662;
  wire _abc_17692_n6663;
  wire _abc_17692_n6664;
  wire _abc_17692_n6665;
  wire _abc_17692_n6666;
  wire _abc_17692_n6667;
  wire _abc_17692_n6668;
  wire _abc_17692_n6669;
  wire _abc_17692_n667;
  wire _abc_17692_n6670;
  wire _abc_17692_n6671;
  wire _abc_17692_n6672;
  wire _abc_17692_n6673;
  wire _abc_17692_n6674;
  wire _abc_17692_n6675;
  wire _abc_17692_n6676;
  wire _abc_17692_n6677;
  wire _abc_17692_n6678;
  wire _abc_17692_n6679;
  wire _abc_17692_n668;
  wire _abc_17692_n6680;
  wire _abc_17692_n6681;
  wire _abc_17692_n6682;
  wire _abc_17692_n6683;
  wire _abc_17692_n6684;
  wire _abc_17692_n6685;
  wire _abc_17692_n6686;
  wire _abc_17692_n6687;
  wire _abc_17692_n6688;
  wire _abc_17692_n6689;
  wire _abc_17692_n669;
  wire _abc_17692_n6690;
  wire _abc_17692_n6691;
  wire _abc_17692_n6692;
  wire _abc_17692_n6693;
  wire _abc_17692_n6694;
  wire _abc_17692_n6695;
  wire _abc_17692_n6696;
  wire _abc_17692_n6697;
  wire _abc_17692_n6698;
  wire _abc_17692_n6699;
  wire _abc_17692_n6700;
  wire _abc_17692_n6701;
  wire _abc_17692_n6702;
  wire _abc_17692_n6703;
  wire _abc_17692_n6704;
  wire _abc_17692_n6705;
  wire _abc_17692_n6706;
  wire _abc_17692_n6707;
  wire _abc_17692_n6708;
  wire _abc_17692_n6709;
  wire _abc_17692_n671;
  wire _abc_17692_n6710;
  wire _abc_17692_n6711;
  wire _abc_17692_n6712;
  wire _abc_17692_n6713;
  wire _abc_17692_n6714;
  wire _abc_17692_n6715;
  wire _abc_17692_n6716;
  wire _abc_17692_n6717;
  wire _abc_17692_n6718;
  wire _abc_17692_n6719;
  wire _abc_17692_n672;
  wire _abc_17692_n6720;
  wire _abc_17692_n6721;
  wire _abc_17692_n6722;
  wire _abc_17692_n6723;
  wire _abc_17692_n6724;
  wire _abc_17692_n6725;
  wire _abc_17692_n6726;
  wire _abc_17692_n6727;
  wire _abc_17692_n6728;
  wire _abc_17692_n6729;
  wire _abc_17692_n673;
  wire _abc_17692_n6730;
  wire _abc_17692_n6731;
  wire _abc_17692_n6732;
  wire _abc_17692_n6733;
  wire _abc_17692_n6734;
  wire _abc_17692_n6735;
  wire _abc_17692_n6736;
  wire _abc_17692_n6737;
  wire _abc_17692_n6738;
  wire _abc_17692_n6739;
  wire _abc_17692_n6740;
  wire _abc_17692_n6741;
  wire _abc_17692_n6742;
  wire _abc_17692_n6743;
  wire _abc_17692_n6744;
  wire _abc_17692_n6745;
  wire _abc_17692_n6746;
  wire _abc_17692_n6747;
  wire _abc_17692_n6748;
  wire _abc_17692_n6749;
  wire _abc_17692_n675;
  wire _abc_17692_n6750;
  wire _abc_17692_n6751;
  wire _abc_17692_n6752;
  wire _abc_17692_n6753;
  wire _abc_17692_n6754;
  wire _abc_17692_n6755;
  wire _abc_17692_n6756;
  wire _abc_17692_n6757;
  wire _abc_17692_n6758;
  wire _abc_17692_n6759;
  wire _abc_17692_n6760;
  wire _abc_17692_n6761;
  wire _abc_17692_n6762;
  wire _abc_17692_n6763;
  wire _abc_17692_n6764;
  wire _abc_17692_n6765;
  wire _abc_17692_n6766;
  wire _abc_17692_n6767;
  wire _abc_17692_n6768;
  wire _abc_17692_n6769;
  wire _abc_17692_n676_1;
  wire _abc_17692_n6770;
  wire _abc_17692_n6771;
  wire _abc_17692_n6772;
  wire _abc_17692_n6773;
  wire _abc_17692_n6774;
  wire _abc_17692_n6775;
  wire _abc_17692_n6776;
  wire _abc_17692_n6777;
  wire _abc_17692_n6778;
  wire _abc_17692_n6779;
  wire _abc_17692_n677_1;
  wire _abc_17692_n6780;
  wire _abc_17692_n6781;
  wire _abc_17692_n6782;
  wire _abc_17692_n6783;
  wire _abc_17692_n6784;
  wire _abc_17692_n6785;
  wire _abc_17692_n6786;
  wire _abc_17692_n6787;
  wire _abc_17692_n6788;
  wire _abc_17692_n6789;
  wire _abc_17692_n679;
  wire _abc_17692_n6790;
  wire _abc_17692_n6791;
  wire _abc_17692_n6792;
  wire _abc_17692_n6793;
  wire _abc_17692_n6794;
  wire _abc_17692_n6795;
  wire _abc_17692_n6796;
  wire _abc_17692_n6797;
  wire _abc_17692_n6798;
  wire _abc_17692_n6799;
  wire _abc_17692_n680;
  wire _abc_17692_n6800;
  wire _abc_17692_n6801;
  wire _abc_17692_n6802;
  wire _abc_17692_n6803;
  wire _abc_17692_n6804;
  wire _abc_17692_n6805;
  wire _abc_17692_n6806;
  wire _abc_17692_n6807;
  wire _abc_17692_n6808;
  wire _abc_17692_n6809;
  wire _abc_17692_n681;
  wire _abc_17692_n6810;
  wire _abc_17692_n6811;
  wire _abc_17692_n6812;
  wire _abc_17692_n6813;
  wire _abc_17692_n6814;
  wire _abc_17692_n6815;
  wire _abc_17692_n6816;
  wire _abc_17692_n6817;
  wire _abc_17692_n6818;
  wire _abc_17692_n6819;
  wire _abc_17692_n6820;
  wire _abc_17692_n6821;
  wire _abc_17692_n6822;
  wire _abc_17692_n6823;
  wire _abc_17692_n6824;
  wire _abc_17692_n6825;
  wire _abc_17692_n6826;
  wire _abc_17692_n6827;
  wire _abc_17692_n6828;
  wire _abc_17692_n6829;
  wire _abc_17692_n683;
  wire _abc_17692_n6830;
  wire _abc_17692_n6831;
  wire _abc_17692_n6832;
  wire _abc_17692_n6833;
  wire _abc_17692_n6834;
  wire _abc_17692_n6835;
  wire _abc_17692_n6836;
  wire _abc_17692_n6837;
  wire _abc_17692_n6838;
  wire _abc_17692_n6839;
  wire _abc_17692_n684;
  wire _abc_17692_n6840;
  wire _abc_17692_n6841;
  wire _abc_17692_n6842;
  wire _abc_17692_n6843;
  wire _abc_17692_n6844;
  wire _abc_17692_n6845;
  wire _abc_17692_n6846;
  wire _abc_17692_n6847;
  wire _abc_17692_n6848;
  wire _abc_17692_n6849;
  wire _abc_17692_n685;
  wire _abc_17692_n6850;
  wire _abc_17692_n6851;
  wire _abc_17692_n6852;
  wire _abc_17692_n6853;
  wire _abc_17692_n6854;
  wire _abc_17692_n6855;
  wire _abc_17692_n6856;
  wire _abc_17692_n6857;
  wire _abc_17692_n6858;
  wire _abc_17692_n6859;
  wire _abc_17692_n6860;
  wire _abc_17692_n6861;
  wire _abc_17692_n6862;
  wire _abc_17692_n6863;
  wire _abc_17692_n6864;
  wire _abc_17692_n6865;
  wire _abc_17692_n6866;
  wire _abc_17692_n6867;
  wire _abc_17692_n6868;
  wire _abc_17692_n6869;
  wire _abc_17692_n687;
  wire _abc_17692_n6870;
  wire _abc_17692_n6871;
  wire _abc_17692_n6872;
  wire _abc_17692_n6873;
  wire _abc_17692_n6874;
  wire _abc_17692_n6875;
  wire _abc_17692_n6876;
  wire _abc_17692_n6877;
  wire _abc_17692_n6878;
  wire _abc_17692_n6879;
  wire _abc_17692_n688;
  wire _abc_17692_n6880;
  wire _abc_17692_n6881;
  wire _abc_17692_n6882;
  wire _abc_17692_n6883;
  wire _abc_17692_n6884;
  wire _abc_17692_n6885;
  wire _abc_17692_n6886;
  wire _abc_17692_n6887;
  wire _abc_17692_n6888;
  wire _abc_17692_n6889;
  wire _abc_17692_n689;
  wire _abc_17692_n6890;
  wire _abc_17692_n6891;
  wire _abc_17692_n6892;
  wire _abc_17692_n6893;
  wire _abc_17692_n6894;
  wire _abc_17692_n6895;
  wire _abc_17692_n6896;
  wire _abc_17692_n6897;
  wire _abc_17692_n6898;
  wire _abc_17692_n6899;
  wire _abc_17692_n6900;
  wire _abc_17692_n6901;
  wire _abc_17692_n6902;
  wire _abc_17692_n6903;
  wire _abc_17692_n6904;
  wire _abc_17692_n6905;
  wire _abc_17692_n6906;
  wire _abc_17692_n6907;
  wire _abc_17692_n6908;
  wire _abc_17692_n6909;
  wire _abc_17692_n691;
  wire _abc_17692_n6910;
  wire _abc_17692_n6911;
  wire _abc_17692_n6912;
  wire _abc_17692_n6913;
  wire _abc_17692_n6914;
  wire _abc_17692_n6915;
  wire _abc_17692_n6916;
  wire _abc_17692_n6917;
  wire _abc_17692_n6918;
  wire _abc_17692_n6919;
  wire _abc_17692_n6920;
  wire _abc_17692_n6921;
  wire _abc_17692_n6922;
  wire _abc_17692_n6923;
  wire _abc_17692_n6924;
  wire _abc_17692_n6925;
  wire _abc_17692_n6926;
  wire _abc_17692_n6927;
  wire _abc_17692_n6928;
  wire _abc_17692_n6929;
  wire _abc_17692_n692_1;
  wire _abc_17692_n6930;
  wire _abc_17692_n6931;
  wire _abc_17692_n6932;
  wire _abc_17692_n6933;
  wire _abc_17692_n6934;
  wire _abc_17692_n6935;
  wire _abc_17692_n6936;
  wire _abc_17692_n6937;
  wire _abc_17692_n6938;
  wire _abc_17692_n6939;
  wire _abc_17692_n693_1;
  wire _abc_17692_n6940;
  wire _abc_17692_n6941;
  wire _abc_17692_n6942;
  wire _abc_17692_n6943;
  wire _abc_17692_n6944;
  wire _abc_17692_n6945;
  wire _abc_17692_n6946;
  wire _abc_17692_n6947;
  wire _abc_17692_n6948;
  wire _abc_17692_n6949;
  wire _abc_17692_n695;
  wire _abc_17692_n6950;
  wire _abc_17692_n6952;
  wire _abc_17692_n6953;
  wire _abc_17692_n6954;
  wire _abc_17692_n6955;
  wire _abc_17692_n6956;
  wire _abc_17692_n6957;
  wire _abc_17692_n6958;
  wire _abc_17692_n6959;
  wire _abc_17692_n696;
  wire _abc_17692_n6960;
  wire _abc_17692_n6961;
  wire _abc_17692_n6962;
  wire _abc_17692_n6963;
  wire _abc_17692_n6964;
  wire _abc_17692_n6965;
  wire _abc_17692_n6966;
  wire _abc_17692_n6967;
  wire _abc_17692_n6968;
  wire _abc_17692_n6969;
  wire _abc_17692_n697;
  wire _abc_17692_n6970;
  wire _abc_17692_n6971;
  wire _abc_17692_n6972;
  wire _abc_17692_n6973;
  wire _abc_17692_n6974;
  wire _abc_17692_n6975;
  wire _abc_17692_n6976;
  wire _abc_17692_n6977;
  wire _abc_17692_n6978;
  wire _abc_17692_n6979;
  wire _abc_17692_n6980;
  wire _abc_17692_n6981;
  wire _abc_17692_n6982;
  wire _abc_17692_n6983;
  wire _abc_17692_n6984;
  wire _abc_17692_n6985;
  wire _abc_17692_n6986;
  wire _abc_17692_n6987;
  wire _abc_17692_n6988;
  wire _abc_17692_n6989;
  wire _abc_17692_n699;
  wire _abc_17692_n6990;
  wire _abc_17692_n6991;
  wire _abc_17692_n6992;
  wire _abc_17692_n6993;
  wire _abc_17692_n6994;
  wire _abc_17692_n6995;
  wire _abc_17692_n6996;
  wire _abc_17692_n6997;
  wire _abc_17692_n6998;
  wire _abc_17692_n6999;
  wire _abc_17692_n700;
  wire _abc_17692_n7000;
  wire _abc_17692_n7001;
  wire _abc_17692_n7002;
  wire _abc_17692_n7003;
  wire _abc_17692_n7004;
  wire _abc_17692_n7005;
  wire _abc_17692_n7006;
  wire _abc_17692_n7007;
  wire _abc_17692_n7008;
  wire _abc_17692_n7009;
  wire _abc_17692_n701;
  wire _abc_17692_n7010;
  wire _abc_17692_n7011;
  wire _abc_17692_n7012;
  wire _abc_17692_n7013;
  wire _abc_17692_n7014;
  wire _abc_17692_n7015;
  wire _abc_17692_n7016;
  wire _abc_17692_n7017;
  wire _abc_17692_n7018;
  wire _abc_17692_n7019;
  wire _abc_17692_n702;
  wire _abc_17692_n7020;
  wire _abc_17692_n7021;
  wire _abc_17692_n7022;
  wire _abc_17692_n7023;
  wire _abc_17692_n7024;
  wire _abc_17692_n7025;
  wire _abc_17692_n7026;
  wire _abc_17692_n7027;
  wire _abc_17692_n7028;
  wire _abc_17692_n7029;
  wire _abc_17692_n703;
  wire _abc_17692_n7030;
  wire _abc_17692_n7031;
  wire _abc_17692_n7032;
  wire _abc_17692_n7033;
  wire _abc_17692_n7034;
  wire _abc_17692_n7035;
  wire _abc_17692_n7036;
  wire _abc_17692_n7037;
  wire _abc_17692_n7038;
  wire _abc_17692_n7039;
  wire _abc_17692_n704;
  wire _abc_17692_n7040;
  wire _abc_17692_n7041;
  wire _abc_17692_n7042;
  wire _abc_17692_n7043;
  wire _abc_17692_n7044;
  wire _abc_17692_n7045;
  wire _abc_17692_n7046;
  wire _abc_17692_n7047;
  wire _abc_17692_n7048;
  wire _abc_17692_n7049;
  wire _abc_17692_n705;
  wire _abc_17692_n7050;
  wire _abc_17692_n7051;
  wire _abc_17692_n7052;
  wire _abc_17692_n7053;
  wire _abc_17692_n7054;
  wire _abc_17692_n7055;
  wire _abc_17692_n7056;
  wire _abc_17692_n7057;
  wire _abc_17692_n7058;
  wire _abc_17692_n7059;
  wire _abc_17692_n706;
  wire _abc_17692_n7060;
  wire _abc_17692_n7061;
  wire _abc_17692_n7062;
  wire _abc_17692_n7063;
  wire _abc_17692_n7064;
  wire _abc_17692_n7065;
  wire _abc_17692_n7066;
  wire _abc_17692_n7067;
  wire _abc_17692_n7068;
  wire _abc_17692_n7069;
  wire _abc_17692_n7070;
  wire _abc_17692_n7071;
  wire _abc_17692_n7072;
  wire _abc_17692_n7073;
  wire _abc_17692_n7074;
  wire _abc_17692_n7075;
  wire _abc_17692_n7076;
  wire _abc_17692_n7077;
  wire _abc_17692_n7078;
  wire _abc_17692_n7079;
  wire _abc_17692_n708;
  wire _abc_17692_n7080;
  wire _abc_17692_n7081;
  wire _abc_17692_n7082;
  wire _abc_17692_n7083;
  wire _abc_17692_n7084;
  wire _abc_17692_n7085;
  wire _abc_17692_n7086;
  wire _abc_17692_n7087;
  wire _abc_17692_n7088;
  wire _abc_17692_n7089;
  wire _abc_17692_n709;
  wire _abc_17692_n7090;
  wire _abc_17692_n7091;
  wire _abc_17692_n7092;
  wire _abc_17692_n7093;
  wire _abc_17692_n7094;
  wire _abc_17692_n7095;
  wire _abc_17692_n7096;
  wire _abc_17692_n7097;
  wire _abc_17692_n7098;
  wire _abc_17692_n7099;
  wire _abc_17692_n710;
  wire _abc_17692_n7100;
  wire _abc_17692_n7101;
  wire _abc_17692_n7102;
  wire _abc_17692_n7103;
  wire _abc_17692_n7104;
  wire _abc_17692_n7105;
  wire _abc_17692_n7106;
  wire _abc_17692_n7107;
  wire _abc_17692_n7108;
  wire _abc_17692_n7109;
  wire _abc_17692_n711;
  wire _abc_17692_n7110;
  wire _abc_17692_n7111;
  wire _abc_17692_n7112;
  wire _abc_17692_n7113;
  wire _abc_17692_n7114;
  wire _abc_17692_n7115;
  wire _abc_17692_n7116;
  wire _abc_17692_n7117;
  wire _abc_17692_n7118;
  wire _abc_17692_n7119;
  wire _abc_17692_n712;
  wire _abc_17692_n7120;
  wire _abc_17692_n7121;
  wire _abc_17692_n7122;
  wire _abc_17692_n7123;
  wire _abc_17692_n7124;
  wire _abc_17692_n7125;
  wire _abc_17692_n7126;
  wire _abc_17692_n7128;
  wire _abc_17692_n7129;
  wire _abc_17692_n713;
  wire _abc_17692_n7130;
  wire _abc_17692_n7131;
  wire _abc_17692_n7132;
  wire _abc_17692_n7133;
  wire _abc_17692_n7134;
  wire _abc_17692_n7135;
  wire _abc_17692_n7136;
  wire _abc_17692_n7137;
  wire _abc_17692_n7138;
  wire _abc_17692_n7139;
  wire _abc_17692_n7140;
  wire _abc_17692_n7141;
  wire _abc_17692_n7142;
  wire _abc_17692_n7143;
  wire _abc_17692_n7144;
  wire _abc_17692_n7145;
  wire _abc_17692_n7146;
  wire _abc_17692_n7147;
  wire _abc_17692_n7148;
  wire _abc_17692_n7149;
  wire _abc_17692_n714_1;
  wire _abc_17692_n7150;
  wire _abc_17692_n7151;
  wire _abc_17692_n7152;
  wire _abc_17692_n7153;
  wire _abc_17692_n7154;
  wire _abc_17692_n7155;
  wire _abc_17692_n7156;
  wire _abc_17692_n7157;
  wire _abc_17692_n7158;
  wire _abc_17692_n7159;
  wire _abc_17692_n715_1;
  wire _abc_17692_n716;
  wire _abc_17692_n7160;
  wire _abc_17692_n7161;
  wire _abc_17692_n7162;
  wire _abc_17692_n7163;
  wire _abc_17692_n7164;
  wire _abc_17692_n7165;
  wire _abc_17692_n7166;
  wire _abc_17692_n7167;
  wire _abc_17692_n7168;
  wire _abc_17692_n7169;
  wire _abc_17692_n717;
  wire _abc_17692_n7170;
  wire _abc_17692_n7171;
  wire _abc_17692_n7172;
  wire _abc_17692_n7173;
  wire _abc_17692_n7174;
  wire _abc_17692_n7175;
  wire _abc_17692_n7176;
  wire _abc_17692_n7177;
  wire _abc_17692_n7178;
  wire _abc_17692_n7179;
  wire _abc_17692_n718;
  wire _abc_17692_n7180;
  wire _abc_17692_n7181;
  wire _abc_17692_n7182;
  wire _abc_17692_n7183;
  wire _abc_17692_n7184;
  wire _abc_17692_n7185;
  wire _abc_17692_n7186;
  wire _abc_17692_n7187;
  wire _abc_17692_n7188;
  wire _abc_17692_n7189;
  wire _abc_17692_n719;
  wire _abc_17692_n7190;
  wire _abc_17692_n7191;
  wire _abc_17692_n7192;
  wire _abc_17692_n7193;
  wire _abc_17692_n7194;
  wire _abc_17692_n7195;
  wire _abc_17692_n7196;
  wire _abc_17692_n7197;
  wire _abc_17692_n7198;
  wire _abc_17692_n7199;
  wire _abc_17692_n720;
  wire _abc_17692_n7200;
  wire _abc_17692_n7201;
  wire _abc_17692_n7202;
  wire _abc_17692_n7203;
  wire _abc_17692_n7204;
  wire _abc_17692_n7205;
  wire _abc_17692_n7206;
  wire _abc_17692_n7207;
  wire _abc_17692_n7208;
  wire _abc_17692_n7209;
  wire _abc_17692_n721;
  wire _abc_17692_n7210;
  wire _abc_17692_n7211;
  wire _abc_17692_n7212;
  wire _abc_17692_n7213;
  wire _abc_17692_n7214;
  wire _abc_17692_n7215;
  wire _abc_17692_n7216;
  wire _abc_17692_n7217;
  wire _abc_17692_n7218;
  wire _abc_17692_n7219;
  wire _abc_17692_n722;
  wire _abc_17692_n7220;
  wire _abc_17692_n7221;
  wire _abc_17692_n7222;
  wire _abc_17692_n7223;
  wire _abc_17692_n7224;
  wire _abc_17692_n7225;
  wire _abc_17692_n7226;
  wire _abc_17692_n7227;
  wire _abc_17692_n7228;
  wire _abc_17692_n7229;
  wire _abc_17692_n722_bF_buf0;
  wire _abc_17692_n722_bF_buf1;
  wire _abc_17692_n722_bF_buf2;
  wire _abc_17692_n722_bF_buf3;
  wire _abc_17692_n723;
  wire _abc_17692_n7230;
  wire _abc_17692_n7231;
  wire _abc_17692_n7232;
  wire _abc_17692_n7233;
  wire _abc_17692_n7234;
  wire _abc_17692_n7235;
  wire _abc_17692_n7236;
  wire _abc_17692_n7237;
  wire _abc_17692_n7238;
  wire _abc_17692_n7239;
  wire _abc_17692_n724;
  wire _abc_17692_n7240;
  wire _abc_17692_n7241;
  wire _abc_17692_n7242;
  wire _abc_17692_n7243;
  wire _abc_17692_n7244;
  wire _abc_17692_n7245;
  wire _abc_17692_n7246;
  wire _abc_17692_n7247;
  wire _abc_17692_n7248;
  wire _abc_17692_n7249;
  wire _abc_17692_n725;
  wire _abc_17692_n7250;
  wire _abc_17692_n7251;
  wire _abc_17692_n7252;
  wire _abc_17692_n7253;
  wire _abc_17692_n7254;
  wire _abc_17692_n7255;
  wire _abc_17692_n7256;
  wire _abc_17692_n7257;
  wire _abc_17692_n7258;
  wire _abc_17692_n7259;
  wire _abc_17692_n725_bF_buf0;
  wire _abc_17692_n725_bF_buf1;
  wire _abc_17692_n725_bF_buf2;
  wire _abc_17692_n725_bF_buf3;
  wire _abc_17692_n725_bF_buf4;
  wire _abc_17692_n725_bF_buf5;
  wire _abc_17692_n725_bF_buf6;
  wire _abc_17692_n725_bF_buf7;
  wire _abc_17692_n726;
  wire _abc_17692_n7260;
  wire _abc_17692_n7261;
  wire _abc_17692_n7262;
  wire _abc_17692_n7263;
  wire _abc_17692_n7264;
  wire _abc_17692_n7265;
  wire _abc_17692_n7266;
  wire _abc_17692_n7267;
  wire _abc_17692_n7268;
  wire _abc_17692_n7269;
  wire _abc_17692_n727;
  wire _abc_17692_n7270;
  wire _abc_17692_n7271;
  wire _abc_17692_n7272;
  wire _abc_17692_n7273;
  wire _abc_17692_n7274;
  wire _abc_17692_n7275;
  wire _abc_17692_n7276;
  wire _abc_17692_n7277;
  wire _abc_17692_n7278;
  wire _abc_17692_n7279;
  wire _abc_17692_n727_bF_buf0;
  wire _abc_17692_n727_bF_buf1;
  wire _abc_17692_n727_bF_buf2;
  wire _abc_17692_n727_bF_buf3;
  wire _abc_17692_n727_bF_buf4;
  wire _abc_17692_n727_bF_buf5;
  wire _abc_17692_n727_bF_buf6;
  wire _abc_17692_n727_bF_buf7;
  wire _abc_17692_n728;
  wire _abc_17692_n7280;
  wire _abc_17692_n7281;
  wire _abc_17692_n7282;
  wire _abc_17692_n7283;
  wire _abc_17692_n7284;
  wire _abc_17692_n7285;
  wire _abc_17692_n7286;
  wire _abc_17692_n7287;
  wire _abc_17692_n7288;
  wire _abc_17692_n7289;
  wire _abc_17692_n7290;
  wire _abc_17692_n7291;
  wire _abc_17692_n7292;
  wire _abc_17692_n7293;
  wire _abc_17692_n7294;
  wire _abc_17692_n7295;
  wire _abc_17692_n7296;
  wire _abc_17692_n7297;
  wire _abc_17692_n7298;
  wire _abc_17692_n7299;
  wire _abc_17692_n7300;
  wire _abc_17692_n7301;
  wire _abc_17692_n7302;
  wire _abc_17692_n7303;
  wire _abc_17692_n7304;
  wire _abc_17692_n7305;
  wire _abc_17692_n7306;
  wire _abc_17692_n7307;
  wire _abc_17692_n7308;
  wire _abc_17692_n7309;
  wire _abc_17692_n730_1;
  wire _abc_17692_n7310;
  wire _abc_17692_n7311;
  wire _abc_17692_n7312;
  wire _abc_17692_n7313;
  wire _abc_17692_n7314;
  wire _abc_17692_n7315;
  wire _abc_17692_n7316;
  wire _abc_17692_n7317;
  wire _abc_17692_n7318;
  wire _abc_17692_n7319;
  wire _abc_17692_n731_1;
  wire _abc_17692_n7320;
  wire _abc_17692_n7321;
  wire _abc_17692_n7322;
  wire _abc_17692_n7323;
  wire _abc_17692_n7324;
  wire _abc_17692_n7325;
  wire _abc_17692_n7326;
  wire _abc_17692_n7327;
  wire _abc_17692_n7328;
  wire _abc_17692_n7329;
  wire _abc_17692_n733;
  wire _abc_17692_n7330;
  wire _abc_17692_n7331;
  wire _abc_17692_n7332;
  wire _abc_17692_n7333;
  wire _abc_17692_n7334;
  wire _abc_17692_n7335;
  wire _abc_17692_n7336;
  wire _abc_17692_n7337;
  wire _abc_17692_n7338;
  wire _abc_17692_n7339;
  wire _abc_17692_n734;
  wire _abc_17692_n7340;
  wire _abc_17692_n7341;
  wire _abc_17692_n7342;
  wire _abc_17692_n7343;
  wire _abc_17692_n7344;
  wire _abc_17692_n7345;
  wire _abc_17692_n7346;
  wire _abc_17692_n7347;
  wire _abc_17692_n7348;
  wire _abc_17692_n7349;
  wire _abc_17692_n7350;
  wire _abc_17692_n7351;
  wire _abc_17692_n7352;
  wire _abc_17692_n7354;
  wire _abc_17692_n7355;
  wire _abc_17692_n7356;
  wire _abc_17692_n7357;
  wire _abc_17692_n7358;
  wire _abc_17692_n7359;
  wire _abc_17692_n736;
  wire _abc_17692_n7360;
  wire _abc_17692_n7361;
  wire _abc_17692_n7362;
  wire _abc_17692_n7363;
  wire _abc_17692_n7364;
  wire _abc_17692_n7365;
  wire _abc_17692_n7366;
  wire _abc_17692_n7367;
  wire _abc_17692_n7368;
  wire _abc_17692_n7369;
  wire _abc_17692_n737;
  wire _abc_17692_n7370;
  wire _abc_17692_n7371;
  wire _abc_17692_n7372;
  wire _abc_17692_n7373;
  wire _abc_17692_n7374;
  wire _abc_17692_n7375;
  wire _abc_17692_n7376;
  wire _abc_17692_n7377;
  wire _abc_17692_n7378;
  wire _abc_17692_n7379;
  wire _abc_17692_n7380;
  wire _abc_17692_n7381;
  wire _abc_17692_n7382;
  wire _abc_17692_n7383;
  wire _abc_17692_n7384;
  wire _abc_17692_n7385;
  wire _abc_17692_n7386;
  wire _abc_17692_n7387;
  wire _abc_17692_n7388;
  wire _abc_17692_n7389;
  wire _abc_17692_n739;
  wire _abc_17692_n7390;
  wire _abc_17692_n7391;
  wire _abc_17692_n7392;
  wire _abc_17692_n7393;
  wire _abc_17692_n7394;
  wire _abc_17692_n7395;
  wire _abc_17692_n7396;
  wire _abc_17692_n7397;
  wire _abc_17692_n7398;
  wire _abc_17692_n7399;
  wire _abc_17692_n740;
  wire _abc_17692_n7400;
  wire _abc_17692_n7401;
  wire _abc_17692_n7402;
  wire _abc_17692_n7403;
  wire _abc_17692_n7404;
  wire _abc_17692_n7405;
  wire _abc_17692_n7406;
  wire _abc_17692_n7407;
  wire _abc_17692_n7408;
  wire _abc_17692_n7409;
  wire _abc_17692_n7410;
  wire _abc_17692_n7411;
  wire _abc_17692_n7412;
  wire _abc_17692_n7413;
  wire _abc_17692_n7414;
  wire _abc_17692_n7415;
  wire _abc_17692_n7416;
  wire _abc_17692_n7417;
  wire _abc_17692_n7418;
  wire _abc_17692_n7419;
  wire _abc_17692_n742;
  wire _abc_17692_n7420;
  wire _abc_17692_n7421;
  wire _abc_17692_n7422;
  wire _abc_17692_n7423;
  wire _abc_17692_n7424;
  wire _abc_17692_n7425;
  wire _abc_17692_n7426;
  wire _abc_17692_n7427;
  wire _abc_17692_n7428;
  wire _abc_17692_n7429;
  wire _abc_17692_n743;
  wire _abc_17692_n7430;
  wire _abc_17692_n7431;
  wire _abc_17692_n7432;
  wire _abc_17692_n7433;
  wire _abc_17692_n7434;
  wire _abc_17692_n7435;
  wire _abc_17692_n7436;
  wire _abc_17692_n7437;
  wire _abc_17692_n7438;
  wire _abc_17692_n7439;
  wire _abc_17692_n7440;
  wire _abc_17692_n7441;
  wire _abc_17692_n7442;
  wire _abc_17692_n7443;
  wire _abc_17692_n7444;
  wire _abc_17692_n7445;
  wire _abc_17692_n7446;
  wire _abc_17692_n7447;
  wire _abc_17692_n7448;
  wire _abc_17692_n7449;
  wire _abc_17692_n745;
  wire _abc_17692_n7450;
  wire _abc_17692_n7451;
  wire _abc_17692_n7452;
  wire _abc_17692_n7453;
  wire _abc_17692_n7454;
  wire _abc_17692_n7455;
  wire _abc_17692_n7456;
  wire _abc_17692_n7457;
  wire _abc_17692_n7458;
  wire _abc_17692_n7459;
  wire _abc_17692_n746;
  wire _abc_17692_n7460;
  wire _abc_17692_n7461;
  wire _abc_17692_n7462;
  wire _abc_17692_n7463;
  wire _abc_17692_n7464;
  wire _abc_17692_n7465;
  wire _abc_17692_n7466;
  wire _abc_17692_n7467;
  wire _abc_17692_n7468;
  wire _abc_17692_n7469;
  wire _abc_17692_n7470;
  wire _abc_17692_n7471;
  wire _abc_17692_n7472;
  wire _abc_17692_n7473;
  wire _abc_17692_n7474;
  wire _abc_17692_n7475;
  wire _abc_17692_n7476;
  wire _abc_17692_n7477;
  wire _abc_17692_n7478;
  wire _abc_17692_n7479;
  wire _abc_17692_n748;
  wire _abc_17692_n7480;
  wire _abc_17692_n7481;
  wire _abc_17692_n7482;
  wire _abc_17692_n7483;
  wire _abc_17692_n7484;
  wire _abc_17692_n7485;
  wire _abc_17692_n7486;
  wire _abc_17692_n7487;
  wire _abc_17692_n7488;
  wire _abc_17692_n7489;
  wire _abc_17692_n749;
  wire _abc_17692_n7490;
  wire _abc_17692_n7491;
  wire _abc_17692_n7492;
  wire _abc_17692_n7493;
  wire _abc_17692_n7494;
  wire _abc_17692_n7495;
  wire _abc_17692_n7496;
  wire _abc_17692_n7497;
  wire _abc_17692_n7498;
  wire _abc_17692_n7499;
  wire _abc_17692_n7500;
  wire _abc_17692_n7501;
  wire _abc_17692_n7502;
  wire _abc_17692_n7503;
  wire _abc_17692_n7504;
  wire _abc_17692_n7505;
  wire _abc_17692_n7506;
  wire _abc_17692_n7507;
  wire _abc_17692_n7508;
  wire _abc_17692_n7509;
  wire _abc_17692_n7510;
  wire _abc_17692_n7511;
  wire _abc_17692_n7512;
  wire _abc_17692_n7513;
  wire _abc_17692_n7514;
  wire _abc_17692_n7515;
  wire _abc_17692_n7516;
  wire _abc_17692_n7517;
  wire _abc_17692_n7518;
  wire _abc_17692_n7519;
  wire _abc_17692_n751_1;
  wire _abc_17692_n752;
  wire _abc_17692_n7520;
  wire _abc_17692_n7521;
  wire _abc_17692_n7522;
  wire _abc_17692_n7523;
  wire _abc_17692_n7524;
  wire _abc_17692_n7525;
  wire _abc_17692_n7526;
  wire _abc_17692_n7527;
  wire _abc_17692_n7528;
  wire _abc_17692_n7529;
  wire _abc_17692_n7530;
  wire _abc_17692_n7531;
  wire _abc_17692_n7532;
  wire _abc_17692_n7533;
  wire _abc_17692_n7535;
  wire _abc_17692_n7536;
  wire _abc_17692_n7537;
  wire _abc_17692_n7538;
  wire _abc_17692_n7539;
  wire _abc_17692_n754;
  wire _abc_17692_n7540;
  wire _abc_17692_n7541;
  wire _abc_17692_n7542;
  wire _abc_17692_n7543;
  wire _abc_17692_n7544;
  wire _abc_17692_n7545;
  wire _abc_17692_n7546;
  wire _abc_17692_n7547;
  wire _abc_17692_n7548;
  wire _abc_17692_n7549;
  wire _abc_17692_n755;
  wire _abc_17692_n7550;
  wire _abc_17692_n7551;
  wire _abc_17692_n7552;
  wire _abc_17692_n7553;
  wire _abc_17692_n7554;
  wire _abc_17692_n7555;
  wire _abc_17692_n7556;
  wire _abc_17692_n7557;
  wire _abc_17692_n7558;
  wire _abc_17692_n7559;
  wire _abc_17692_n7560;
  wire _abc_17692_n7561;
  wire _abc_17692_n7562;
  wire _abc_17692_n7563;
  wire _abc_17692_n7564;
  wire _abc_17692_n7565;
  wire _abc_17692_n7566;
  wire _abc_17692_n7567;
  wire _abc_17692_n7568;
  wire _abc_17692_n7569;
  wire _abc_17692_n757;
  wire _abc_17692_n7570;
  wire _abc_17692_n7571;
  wire _abc_17692_n7572;
  wire _abc_17692_n7573;
  wire _abc_17692_n7574;
  wire _abc_17692_n7575;
  wire _abc_17692_n7576;
  wire _abc_17692_n7577;
  wire _abc_17692_n7578;
  wire _abc_17692_n7579;
  wire _abc_17692_n758;
  wire _abc_17692_n7580;
  wire _abc_17692_n7581;
  wire _abc_17692_n7582;
  wire _abc_17692_n7583;
  wire _abc_17692_n7584;
  wire _abc_17692_n7585;
  wire _abc_17692_n7586;
  wire _abc_17692_n7587;
  wire _abc_17692_n7588;
  wire _abc_17692_n7589;
  wire _abc_17692_n7590;
  wire _abc_17692_n7591;
  wire _abc_17692_n7592;
  wire _abc_17692_n7593;
  wire _abc_17692_n7594;
  wire _abc_17692_n7595;
  wire _abc_17692_n7596;
  wire _abc_17692_n7597;
  wire _abc_17692_n7598;
  wire _abc_17692_n7599;
  wire _abc_17692_n760;
  wire _abc_17692_n7600;
  wire _abc_17692_n7601;
  wire _abc_17692_n7602;
  wire _abc_17692_n7603;
  wire _abc_17692_n7604;
  wire _abc_17692_n7605;
  wire _abc_17692_n7606;
  wire _abc_17692_n7607;
  wire _abc_17692_n7608;
  wire _abc_17692_n7609;
  wire _abc_17692_n761;
  wire _abc_17692_n7610;
  wire _abc_17692_n7611;
  wire _abc_17692_n7612;
  wire _abc_17692_n7613;
  wire _abc_17692_n7614;
  wire _abc_17692_n7615;
  wire _abc_17692_n7616;
  wire _abc_17692_n7617;
  wire _abc_17692_n7618;
  wire _abc_17692_n7619;
  wire _abc_17692_n7620;
  wire _abc_17692_n7621;
  wire _abc_17692_n7622;
  wire _abc_17692_n7623;
  wire _abc_17692_n7624;
  wire _abc_17692_n7625;
  wire _abc_17692_n7626;
  wire _abc_17692_n7627;
  wire _abc_17692_n7628;
  wire _abc_17692_n7629;
  wire _abc_17692_n763;
  wire _abc_17692_n7630;
  wire _abc_17692_n7631;
  wire _abc_17692_n7632;
  wire _abc_17692_n7633;
  wire _abc_17692_n7634;
  wire _abc_17692_n7635;
  wire _abc_17692_n7636;
  wire _abc_17692_n7637;
  wire _abc_17692_n7638;
  wire _abc_17692_n7639;
  wire _abc_17692_n764;
  wire _abc_17692_n7640;
  wire _abc_17692_n7641;
  wire _abc_17692_n7642;
  wire _abc_17692_n7643;
  wire _abc_17692_n7644;
  wire _abc_17692_n7645;
  wire _abc_17692_n7646;
  wire _abc_17692_n7647;
  wire _abc_17692_n7648;
  wire _abc_17692_n7649;
  wire _abc_17692_n7650;
  wire _abc_17692_n7651;
  wire _abc_17692_n7652;
  wire _abc_17692_n7653;
  wire _abc_17692_n7654;
  wire _abc_17692_n7655;
  wire _abc_17692_n7656;
  wire _abc_17692_n7657;
  wire _abc_17692_n7658;
  wire _abc_17692_n7659;
  wire _abc_17692_n7660;
  wire _abc_17692_n7661;
  wire _abc_17692_n7662;
  wire _abc_17692_n7663;
  wire _abc_17692_n7664;
  wire _abc_17692_n7665;
  wire _abc_17692_n7666;
  wire _abc_17692_n7667;
  wire _abc_17692_n7668;
  wire _abc_17692_n7669;
  wire _abc_17692_n766_1;
  wire _abc_17692_n767;
  wire _abc_17692_n7670;
  wire _abc_17692_n7671;
  wire _abc_17692_n7672;
  wire _abc_17692_n7673;
  wire _abc_17692_n7674;
  wire _abc_17692_n7675;
  wire _abc_17692_n7676;
  wire _abc_17692_n7677;
  wire _abc_17692_n7678;
  wire _abc_17692_n7679;
  wire _abc_17692_n7680;
  wire _abc_17692_n7681;
  wire _abc_17692_n7682;
  wire _abc_17692_n7683;
  wire _abc_17692_n7684;
  wire _abc_17692_n7685;
  wire _abc_17692_n7686;
  wire _abc_17692_n7687;
  wire _abc_17692_n7688;
  wire _abc_17692_n7689;
  wire _abc_17692_n769;
  wire _abc_17692_n7690;
  wire _abc_17692_n7691;
  wire _abc_17692_n7692;
  wire _abc_17692_n7693;
  wire _abc_17692_n7694;
  wire _abc_17692_n7695;
  wire _abc_17692_n7696;
  wire _abc_17692_n7697;
  wire _abc_17692_n7698;
  wire _abc_17692_n7699;
  wire _abc_17692_n770;
  wire _abc_17692_n7700;
  wire _abc_17692_n7701;
  wire _abc_17692_n7702;
  wire _abc_17692_n7703;
  wire _abc_17692_n7704;
  wire _abc_17692_n7705;
  wire _abc_17692_n7706;
  wire _abc_17692_n7707;
  wire _abc_17692_n7708;
  wire _abc_17692_n7709;
  wire _abc_17692_n7710;
  wire _abc_17692_n7711;
  wire _abc_17692_n7712;
  wire _abc_17692_n7713;
  wire _abc_17692_n7714;
  wire _abc_17692_n7715;
  wire _abc_17692_n7716;
  wire _abc_17692_n7717;
  wire _abc_17692_n7718;
  wire _abc_17692_n7719;
  wire _abc_17692_n772;
  wire _abc_17692_n7720;
  wire _abc_17692_n7721;
  wire _abc_17692_n7722;
  wire _abc_17692_n7723;
  wire _abc_17692_n7724;
  wire _abc_17692_n7725;
  wire _abc_17692_n7726;
  wire _abc_17692_n7727;
  wire _abc_17692_n7728;
  wire _abc_17692_n7729;
  wire _abc_17692_n773;
  wire _abc_17692_n7730;
  wire _abc_17692_n7731;
  wire _abc_17692_n7732;
  wire _abc_17692_n7733;
  wire _abc_17692_n7734;
  wire _abc_17692_n7735;
  wire _abc_17692_n7736;
  wire _abc_17692_n7737;
  wire _abc_17692_n7738;
  wire _abc_17692_n7739;
  wire _abc_17692_n7740;
  wire _abc_17692_n7741;
  wire _abc_17692_n7742;
  wire _abc_17692_n7743;
  wire _abc_17692_n7744;
  wire _abc_17692_n7745;
  wire _abc_17692_n7746;
  wire _abc_17692_n7747;
  wire _abc_17692_n7748;
  wire _abc_17692_n7749;
  wire _abc_17692_n775;
  wire _abc_17692_n7750;
  wire _abc_17692_n7751;
  wire _abc_17692_n7752;
  wire _abc_17692_n7753;
  wire _abc_17692_n7754;
  wire _abc_17692_n7755;
  wire _abc_17692_n7756;
  wire _abc_17692_n7757;
  wire _abc_17692_n7758;
  wire _abc_17692_n7759;
  wire _abc_17692_n776;
  wire _abc_17692_n7760;
  wire _abc_17692_n7761;
  wire _abc_17692_n7762;
  wire _abc_17692_n7763;
  wire _abc_17692_n7764;
  wire _abc_17692_n7765;
  wire _abc_17692_n7766;
  wire _abc_17692_n7767;
  wire _abc_17692_n7768;
  wire _abc_17692_n7769;
  wire _abc_17692_n7770;
  wire _abc_17692_n7771;
  wire _abc_17692_n7772;
  wire _abc_17692_n7773;
  wire _abc_17692_n7774;
  wire _abc_17692_n7775;
  wire _abc_17692_n7776;
  wire _abc_17692_n7777;
  wire _abc_17692_n7778;
  wire _abc_17692_n7779;
  wire _abc_17692_n778;
  wire _abc_17692_n7780;
  wire _abc_17692_n7781;
  wire _abc_17692_n7783;
  wire _abc_17692_n7784;
  wire _abc_17692_n7785;
  wire _abc_17692_n7786;
  wire _abc_17692_n7787;
  wire _abc_17692_n7788;
  wire _abc_17692_n7789;
  wire _abc_17692_n779;
  wire _abc_17692_n7790;
  wire _abc_17692_n7791;
  wire _abc_17692_n7792;
  wire _abc_17692_n7793;
  wire _abc_17692_n7794;
  wire _abc_17692_n7795;
  wire _abc_17692_n7796;
  wire _abc_17692_n7797;
  wire _abc_17692_n7798;
  wire _abc_17692_n7799;
  wire _abc_17692_n7800;
  wire _abc_17692_n7801;
  wire _abc_17692_n7802;
  wire _abc_17692_n7803;
  wire _abc_17692_n7804;
  wire _abc_17692_n7805;
  wire _abc_17692_n7806;
  wire _abc_17692_n7807;
  wire _abc_17692_n7808;
  wire _abc_17692_n7809;
  wire _abc_17692_n781;
  wire _abc_17692_n7810;
  wire _abc_17692_n7811;
  wire _abc_17692_n7812;
  wire _abc_17692_n7813;
  wire _abc_17692_n7814;
  wire _abc_17692_n7815;
  wire _abc_17692_n7816;
  wire _abc_17692_n7817;
  wire _abc_17692_n7818;
  wire _abc_17692_n7819;
  wire _abc_17692_n782;
  wire _abc_17692_n7820;
  wire _abc_17692_n7821;
  wire _abc_17692_n7822;
  wire _abc_17692_n7823;
  wire _abc_17692_n7824;
  wire _abc_17692_n7825;
  wire _abc_17692_n7826;
  wire _abc_17692_n7827;
  wire _abc_17692_n7828;
  wire _abc_17692_n7829;
  wire _abc_17692_n7830;
  wire _abc_17692_n7831;
  wire _abc_17692_n7832;
  wire _abc_17692_n7833;
  wire _abc_17692_n7834;
  wire _abc_17692_n7835;
  wire _abc_17692_n7836;
  wire _abc_17692_n7837;
  wire _abc_17692_n7838;
  wire _abc_17692_n7839;
  wire _abc_17692_n784;
  wire _abc_17692_n7840;
  wire _abc_17692_n7841;
  wire _abc_17692_n7842;
  wire _abc_17692_n7843;
  wire _abc_17692_n7844;
  wire _abc_17692_n7845;
  wire _abc_17692_n7846;
  wire _abc_17692_n7847;
  wire _abc_17692_n7848;
  wire _abc_17692_n7849;
  wire _abc_17692_n785;
  wire _abc_17692_n7850;
  wire _abc_17692_n7851;
  wire _abc_17692_n7852;
  wire _abc_17692_n7853;
  wire _abc_17692_n7854;
  wire _abc_17692_n7855;
  wire _abc_17692_n7856;
  wire _abc_17692_n7857;
  wire _abc_17692_n7858;
  wire _abc_17692_n7859;
  wire _abc_17692_n7860;
  wire _abc_17692_n7861;
  wire _abc_17692_n7862;
  wire _abc_17692_n7863;
  wire _abc_17692_n7864;
  wire _abc_17692_n7865;
  wire _abc_17692_n7866;
  wire _abc_17692_n7867;
  wire _abc_17692_n7868;
  wire _abc_17692_n7869;
  wire _abc_17692_n787;
  wire _abc_17692_n7870;
  wire _abc_17692_n7871;
  wire _abc_17692_n7872;
  wire _abc_17692_n7873;
  wire _abc_17692_n7874;
  wire _abc_17692_n7875;
  wire _abc_17692_n7876;
  wire _abc_17692_n7877;
  wire _abc_17692_n7878;
  wire _abc_17692_n7879;
  wire _abc_17692_n788;
  wire _abc_17692_n7880;
  wire _abc_17692_n7881;
  wire _abc_17692_n7882;
  wire _abc_17692_n7883;
  wire _abc_17692_n7884;
  wire _abc_17692_n7885;
  wire _abc_17692_n7886;
  wire _abc_17692_n7887;
  wire _abc_17692_n7888;
  wire _abc_17692_n7889;
  wire _abc_17692_n7890;
  wire _abc_17692_n7891;
  wire _abc_17692_n7892;
  wire _abc_17692_n7893;
  wire _abc_17692_n7894;
  wire _abc_17692_n7895;
  wire _abc_17692_n7896;
  wire _abc_17692_n7897;
  wire _abc_17692_n7898;
  wire _abc_17692_n7899;
  wire _abc_17692_n790;
  wire _abc_17692_n7900;
  wire _abc_17692_n7901;
  wire _abc_17692_n7902;
  wire _abc_17692_n7903;
  wire _abc_17692_n7904;
  wire _abc_17692_n7905;
  wire _abc_17692_n7906;
  wire _abc_17692_n7907;
  wire _abc_17692_n7908;
  wire _abc_17692_n7909;
  wire _abc_17692_n791;
  wire _abc_17692_n7910;
  wire _abc_17692_n7911;
  wire _abc_17692_n7912;
  wire _abc_17692_n7913;
  wire _abc_17692_n7914;
  wire _abc_17692_n7915;
  wire _abc_17692_n7916;
  wire _abc_17692_n7917;
  wire _abc_17692_n7918;
  wire _abc_17692_n7919;
  wire _abc_17692_n7920;
  wire _abc_17692_n7921;
  wire _abc_17692_n7922;
  wire _abc_17692_n7923;
  wire _abc_17692_n7924;
  wire _abc_17692_n7925;
  wire _abc_17692_n7926;
  wire _abc_17692_n7927;
  wire _abc_17692_n7928;
  wire _abc_17692_n7929;
  wire _abc_17692_n793;
  wire _abc_17692_n7930;
  wire _abc_17692_n7931;
  wire _abc_17692_n7932;
  wire _abc_17692_n7933;
  wire _abc_17692_n7934;
  wire _abc_17692_n7935;
  wire _abc_17692_n7936;
  wire _abc_17692_n7937;
  wire _abc_17692_n7938;
  wire _abc_17692_n7939;
  wire _abc_17692_n794;
  wire _abc_17692_n7940;
  wire _abc_17692_n7941;
  wire _abc_17692_n7942;
  wire _abc_17692_n7943;
  wire _abc_17692_n7944;
  wire _abc_17692_n7945;
  wire _abc_17692_n7946;
  wire _abc_17692_n7947;
  wire _abc_17692_n7948;
  wire _abc_17692_n7949;
  wire _abc_17692_n7950;
  wire _abc_17692_n7951;
  wire _abc_17692_n7952;
  wire _abc_17692_n7953;
  wire _abc_17692_n7954;
  wire _abc_17692_n7955;
  wire _abc_17692_n7956;
  wire _abc_17692_n7957;
  wire _abc_17692_n7958;
  wire _abc_17692_n796;
  wire _abc_17692_n7960;
  wire _abc_17692_n7961;
  wire _abc_17692_n7962;
  wire _abc_17692_n7963;
  wire _abc_17692_n7964;
  wire _abc_17692_n7965;
  wire _abc_17692_n7966;
  wire _abc_17692_n7967;
  wire _abc_17692_n7968;
  wire _abc_17692_n7969;
  wire _abc_17692_n797;
  wire _abc_17692_n7970;
  wire _abc_17692_n7971;
  wire _abc_17692_n7972;
  wire _abc_17692_n7973;
  wire _abc_17692_n7974;
  wire _abc_17692_n7975;
  wire _abc_17692_n7976;
  wire _abc_17692_n7977;
  wire _abc_17692_n7978;
  wire _abc_17692_n7979;
  wire _abc_17692_n7980;
  wire _abc_17692_n7981;
  wire _abc_17692_n7982;
  wire _abc_17692_n7983;
  wire _abc_17692_n7984;
  wire _abc_17692_n7985;
  wire _abc_17692_n7986;
  wire _abc_17692_n7987;
  wire _abc_17692_n7988;
  wire _abc_17692_n7989;
  wire _abc_17692_n7990;
  wire _abc_17692_n7991;
  wire _abc_17692_n7992;
  wire _abc_17692_n7993;
  wire _abc_17692_n7994;
  wire _abc_17692_n7995;
  wire _abc_17692_n7996;
  wire _abc_17692_n7997;
  wire _abc_17692_n7998;
  wire _abc_17692_n7999;
  wire _abc_17692_n799_1;
  wire _abc_17692_n800;
  wire _abc_17692_n8000;
  wire _abc_17692_n8001;
  wire _abc_17692_n8002;
  wire _abc_17692_n8003;
  wire _abc_17692_n8004;
  wire _abc_17692_n8005;
  wire _abc_17692_n8006;
  wire _abc_17692_n8007;
  wire _abc_17692_n8008;
  wire _abc_17692_n8009;
  wire _abc_17692_n8010;
  wire _abc_17692_n8011;
  wire _abc_17692_n8012;
  wire _abc_17692_n8013;
  wire _abc_17692_n8014;
  wire _abc_17692_n8015;
  wire _abc_17692_n8016;
  wire _abc_17692_n8017;
  wire _abc_17692_n8018;
  wire _abc_17692_n8019;
  wire _abc_17692_n802;
  wire _abc_17692_n8020;
  wire _abc_17692_n8021;
  wire _abc_17692_n8022;
  wire _abc_17692_n8023;
  wire _abc_17692_n8024;
  wire _abc_17692_n8025;
  wire _abc_17692_n8026;
  wire _abc_17692_n8027;
  wire _abc_17692_n8028;
  wire _abc_17692_n8029;
  wire _abc_17692_n803;
  wire _abc_17692_n8030;
  wire _abc_17692_n8031;
  wire _abc_17692_n8032;
  wire _abc_17692_n8033;
  wire _abc_17692_n8034;
  wire _abc_17692_n8035;
  wire _abc_17692_n8036;
  wire _abc_17692_n8037;
  wire _abc_17692_n8038;
  wire _abc_17692_n8039;
  wire _abc_17692_n8040;
  wire _abc_17692_n8041;
  wire _abc_17692_n8042;
  wire _abc_17692_n8043;
  wire _abc_17692_n8044;
  wire _abc_17692_n8045;
  wire _abc_17692_n8046;
  wire _abc_17692_n8047;
  wire _abc_17692_n8048;
  wire _abc_17692_n8049;
  wire _abc_17692_n805;
  wire _abc_17692_n8050;
  wire _abc_17692_n8051;
  wire _abc_17692_n8052;
  wire _abc_17692_n8053;
  wire _abc_17692_n8054;
  wire _abc_17692_n8055;
  wire _abc_17692_n8056;
  wire _abc_17692_n8057;
  wire _abc_17692_n8058;
  wire _abc_17692_n8059;
  wire _abc_17692_n806;
  wire _abc_17692_n8060;
  wire _abc_17692_n8061;
  wire _abc_17692_n8062;
  wire _abc_17692_n8063;
  wire _abc_17692_n8064;
  wire _abc_17692_n8065;
  wire _abc_17692_n8066;
  wire _abc_17692_n8067;
  wire _abc_17692_n8068;
  wire _abc_17692_n8069;
  wire _abc_17692_n8070;
  wire _abc_17692_n8071;
  wire _abc_17692_n8072;
  wire _abc_17692_n8073;
  wire _abc_17692_n8074;
  wire _abc_17692_n8075;
  wire _abc_17692_n8076;
  wire _abc_17692_n8077;
  wire _abc_17692_n8078;
  wire _abc_17692_n8079;
  wire _abc_17692_n808;
  wire _abc_17692_n8080;
  wire _abc_17692_n8081;
  wire _abc_17692_n8082;
  wire _abc_17692_n8083;
  wire _abc_17692_n8084;
  wire _abc_17692_n8085;
  wire _abc_17692_n8086;
  wire _abc_17692_n8087;
  wire _abc_17692_n8088;
  wire _abc_17692_n8089;
  wire _abc_17692_n809;
  wire _abc_17692_n8090;
  wire _abc_17692_n8091;
  wire _abc_17692_n8092;
  wire _abc_17692_n8093;
  wire _abc_17692_n8094;
  wire _abc_17692_n8095;
  wire _abc_17692_n8096;
  wire _abc_17692_n8097;
  wire _abc_17692_n8098;
  wire _abc_17692_n8099;
  wire _abc_17692_n8100;
  wire _abc_17692_n8101;
  wire _abc_17692_n8102;
  wire _abc_17692_n8103;
  wire _abc_17692_n8104;
  wire _abc_17692_n8105;
  wire _abc_17692_n8106;
  wire _abc_17692_n8107;
  wire _abc_17692_n8108;
  wire _abc_17692_n8109;
  wire _abc_17692_n811;
  wire _abc_17692_n8110;
  wire _abc_17692_n8111;
  wire _abc_17692_n8112;
  wire _abc_17692_n8113;
  wire _abc_17692_n8114;
  wire _abc_17692_n8115;
  wire _abc_17692_n8116;
  wire _abc_17692_n8117;
  wire _abc_17692_n8118;
  wire _abc_17692_n8119;
  wire _abc_17692_n812;
  wire _abc_17692_n8120;
  wire _abc_17692_n8121;
  wire _abc_17692_n8122;
  wire _abc_17692_n8123;
  wire _abc_17692_n8124;
  wire _abc_17692_n8125;
  wire _abc_17692_n8126;
  wire _abc_17692_n8127;
  wire _abc_17692_n8128;
  wire _abc_17692_n8129;
  wire _abc_17692_n8130;
  wire _abc_17692_n8131;
  wire _abc_17692_n8132;
  wire _abc_17692_n8133;
  wire _abc_17692_n8134;
  wire _abc_17692_n8135;
  wire _abc_17692_n8136;
  wire _abc_17692_n8137;
  wire _abc_17692_n8138;
  wire _abc_17692_n8139;
  wire _abc_17692_n8140;
  wire _abc_17692_n8141;
  wire _abc_17692_n8142;
  wire _abc_17692_n8143;
  wire _abc_17692_n8144;
  wire _abc_17692_n8145;
  wire _abc_17692_n8146;
  wire _abc_17692_n8147;
  wire _abc_17692_n8148;
  wire _abc_17692_n8149;
  wire _abc_17692_n814_1;
  wire _abc_17692_n8150;
  wire _abc_17692_n8151;
  wire _abc_17692_n8152;
  wire _abc_17692_n8153;
  wire _abc_17692_n8154;
  wire _abc_17692_n8155;
  wire _abc_17692_n8156;
  wire _abc_17692_n8157;
  wire _abc_17692_n8158;
  wire _abc_17692_n8159;
  wire _abc_17692_n815_1;
  wire _abc_17692_n8160;
  wire _abc_17692_n8161;
  wire _abc_17692_n8162;
  wire _abc_17692_n8163;
  wire _abc_17692_n8164;
  wire _abc_17692_n8165;
  wire _abc_17692_n8166;
  wire _abc_17692_n8167;
  wire _abc_17692_n8168;
  wire _abc_17692_n8169;
  wire _abc_17692_n817;
  wire _abc_17692_n8170;
  wire _abc_17692_n8171;
  wire _abc_17692_n8172;
  wire _abc_17692_n8173;
  wire _abc_17692_n8174;
  wire _abc_17692_n8175;
  wire _abc_17692_n8176;
  wire _abc_17692_n8177;
  wire _abc_17692_n8178;
  wire _abc_17692_n8179;
  wire _abc_17692_n818;
  wire _abc_17692_n8180;
  wire _abc_17692_n8181;
  wire _abc_17692_n8182;
  wire _abc_17692_n8183;
  wire _abc_17692_n8184;
  wire _abc_17692_n8185;
  wire _abc_17692_n8186;
  wire _abc_17692_n8187;
  wire _abc_17692_n8189;
  wire _abc_17692_n8190;
  wire _abc_17692_n8191;
  wire _abc_17692_n8192;
  wire _abc_17692_n8193;
  wire _abc_17692_n8194;
  wire _abc_17692_n8195;
  wire _abc_17692_n8196;
  wire _abc_17692_n8197;
  wire _abc_17692_n8198;
  wire _abc_17692_n8199;
  wire _abc_17692_n820;
  wire _abc_17692_n8200;
  wire _abc_17692_n8201;
  wire _abc_17692_n8202;
  wire _abc_17692_n8203;
  wire _abc_17692_n8204;
  wire _abc_17692_n8205;
  wire _abc_17692_n8206;
  wire _abc_17692_n8207;
  wire _abc_17692_n8208;
  wire _abc_17692_n8209;
  wire _abc_17692_n821;
  wire _abc_17692_n8210;
  wire _abc_17692_n8211;
  wire _abc_17692_n8212;
  wire _abc_17692_n8213;
  wire _abc_17692_n8214;
  wire _abc_17692_n8215;
  wire _abc_17692_n8216;
  wire _abc_17692_n8217;
  wire _abc_17692_n8218;
  wire _abc_17692_n8219;
  wire _abc_17692_n8220;
  wire _abc_17692_n8221;
  wire _abc_17692_n8222;
  wire _abc_17692_n8223;
  wire _abc_17692_n8224;
  wire _abc_17692_n8225;
  wire _abc_17692_n8226;
  wire _abc_17692_n8227;
  wire _abc_17692_n8228;
  wire _abc_17692_n8229;
  wire _abc_17692_n823;
  wire _abc_17692_n8230;
  wire _abc_17692_n8231;
  wire _abc_17692_n8232;
  wire _abc_17692_n8233;
  wire _abc_17692_n8234;
  wire _abc_17692_n8235;
  wire _abc_17692_n8236;
  wire _abc_17692_n8237;
  wire _abc_17692_n8238;
  wire _abc_17692_n8239;
  wire _abc_17692_n824;
  wire _abc_17692_n8240;
  wire _abc_17692_n8241;
  wire _abc_17692_n8242;
  wire _abc_17692_n8243;
  wire _abc_17692_n8244;
  wire _abc_17692_n8245;
  wire _abc_17692_n8246;
  wire _abc_17692_n8247;
  wire _abc_17692_n8248;
  wire _abc_17692_n8249;
  wire _abc_17692_n8250;
  wire _abc_17692_n8251;
  wire _abc_17692_n8252;
  wire _abc_17692_n8253;
  wire _abc_17692_n8254;
  wire _abc_17692_n8255;
  wire _abc_17692_n8256;
  wire _abc_17692_n8257;
  wire _abc_17692_n8258;
  wire _abc_17692_n8259;
  wire _abc_17692_n826;
  wire _abc_17692_n8260;
  wire _abc_17692_n8261;
  wire _abc_17692_n8262;
  wire _abc_17692_n8263;
  wire _abc_17692_n8264;
  wire _abc_17692_n8265;
  wire _abc_17692_n8266;
  wire _abc_17692_n8267;
  wire _abc_17692_n8268;
  wire _abc_17692_n8269;
  wire _abc_17692_n827;
  wire _abc_17692_n8270;
  wire _abc_17692_n8271;
  wire _abc_17692_n8272;
  wire _abc_17692_n8273;
  wire _abc_17692_n8274;
  wire _abc_17692_n8275;
  wire _abc_17692_n8276;
  wire _abc_17692_n8277;
  wire _abc_17692_n8278;
  wire _abc_17692_n8279;
  wire _abc_17692_n8280;
  wire _abc_17692_n8281;
  wire _abc_17692_n8282;
  wire _abc_17692_n8283;
  wire _abc_17692_n8284;
  wire _abc_17692_n8285;
  wire _abc_17692_n8286;
  wire _abc_17692_n8287;
  wire _abc_17692_n8288;
  wire _abc_17692_n8289;
  wire _abc_17692_n829;
  wire _abc_17692_n8290;
  wire _abc_17692_n8291;
  wire _abc_17692_n8292;
  wire _abc_17692_n8293;
  wire _abc_17692_n8294;
  wire _abc_17692_n8295;
  wire _abc_17692_n8296;
  wire _abc_17692_n8297;
  wire _abc_17692_n8298;
  wire _abc_17692_n8299;
  wire _abc_17692_n830;
  wire _abc_17692_n8300;
  wire _abc_17692_n8301;
  wire _abc_17692_n8302;
  wire _abc_17692_n8303;
  wire _abc_17692_n8304;
  wire _abc_17692_n8305;
  wire _abc_17692_n8306;
  wire _abc_17692_n8307;
  wire _abc_17692_n8308;
  wire _abc_17692_n8309;
  wire _abc_17692_n8310;
  wire _abc_17692_n8311;
  wire _abc_17692_n8312;
  wire _abc_17692_n8313;
  wire _abc_17692_n8314;
  wire _abc_17692_n8315;
  wire _abc_17692_n8316;
  wire _abc_17692_n8317;
  wire _abc_17692_n8318;
  wire _abc_17692_n8319;
  wire _abc_17692_n832;
  wire _abc_17692_n8320;
  wire _abc_17692_n8321;
  wire _abc_17692_n8322;
  wire _abc_17692_n8323;
  wire _abc_17692_n8324;
  wire _abc_17692_n8325;
  wire _abc_17692_n8326;
  wire _abc_17692_n8327;
  wire _abc_17692_n8328;
  wire _abc_17692_n8329;
  wire _abc_17692_n833;
  wire _abc_17692_n8330;
  wire _abc_17692_n8331;
  wire _abc_17692_n8332;
  wire _abc_17692_n8333;
  wire _abc_17692_n8334;
  wire _abc_17692_n8335;
  wire _abc_17692_n8336;
  wire _abc_17692_n8338;
  wire _abc_17692_n8339;
  wire _abc_17692_n8340;
  wire _abc_17692_n8341;
  wire _abc_17692_n8342;
  wire _abc_17692_n8343;
  wire _abc_17692_n8344;
  wire _abc_17692_n8345;
  wire _abc_17692_n8346;
  wire _abc_17692_n8347;
  wire _abc_17692_n8348;
  wire _abc_17692_n8349;
  wire _abc_17692_n835;
  wire _abc_17692_n8350;
  wire _abc_17692_n8351;
  wire _abc_17692_n8352;
  wire _abc_17692_n8353;
  wire _abc_17692_n8354;
  wire _abc_17692_n8355;
  wire _abc_17692_n8356;
  wire _abc_17692_n8357;
  wire _abc_17692_n8358;
  wire _abc_17692_n8359;
  wire _abc_17692_n8360;
  wire _abc_17692_n8361;
  wire _abc_17692_n8362;
  wire _abc_17692_n8363;
  wire _abc_17692_n8364;
  wire _abc_17692_n8365;
  wire _abc_17692_n8366;
  wire _abc_17692_n8367;
  wire _abc_17692_n8368;
  wire _abc_17692_n8369;
  wire _abc_17692_n836_1;
  wire _abc_17692_n8370;
  wire _abc_17692_n8371;
  wire _abc_17692_n8372;
  wire _abc_17692_n8373;
  wire _abc_17692_n8374;
  wire _abc_17692_n8375;
  wire _abc_17692_n8376;
  wire _abc_17692_n8377;
  wire _abc_17692_n8378;
  wire _abc_17692_n8379;
  wire _abc_17692_n838;
  wire _abc_17692_n8380;
  wire _abc_17692_n8381;
  wire _abc_17692_n8382;
  wire _abc_17692_n8383;
  wire _abc_17692_n8383_bF_buf0;
  wire _abc_17692_n8383_bF_buf1;
  wire _abc_17692_n8383_bF_buf2;
  wire _abc_17692_n8383_bF_buf3;
  wire _abc_17692_n8383_bF_buf4;
  wire _abc_17692_n8384;
  wire _abc_17692_n8385;
  wire _abc_17692_n8386;
  wire _abc_17692_n8388;
  wire _abc_17692_n8389;
  wire _abc_17692_n839;
  wire _abc_17692_n8390;
  wire _abc_17692_n8391;
  wire _abc_17692_n8392;
  wire _abc_17692_n8393;
  wire _abc_17692_n8394;
  wire _abc_17692_n8395;
  wire _abc_17692_n8396;
  wire _abc_17692_n8397;
  wire _abc_17692_n8398;
  wire _abc_17692_n8399;
  wire _abc_17692_n8400;
  wire _abc_17692_n8401;
  wire _abc_17692_n8402;
  wire _abc_17692_n8403;
  wire _abc_17692_n8404;
  wire _abc_17692_n8405;
  wire _abc_17692_n8406;
  wire _abc_17692_n8407;
  wire _abc_17692_n8408;
  wire _abc_17692_n8409;
  wire _abc_17692_n841;
  wire _abc_17692_n8410;
  wire _abc_17692_n8411;
  wire _abc_17692_n8412;
  wire _abc_17692_n8413;
  wire _abc_17692_n8414;
  wire _abc_17692_n8415;
  wire _abc_17692_n8416;
  wire _abc_17692_n8417;
  wire _abc_17692_n8418;
  wire _abc_17692_n8419;
  wire _abc_17692_n842;
  wire _abc_17692_n8420;
  wire _abc_17692_n8421;
  wire _abc_17692_n8422;
  wire _abc_17692_n8423;
  wire _abc_17692_n8424;
  wire _abc_17692_n8425;
  wire _abc_17692_n8426;
  wire _abc_17692_n8427;
  wire _abc_17692_n8428;
  wire _abc_17692_n8429;
  wire _abc_17692_n8430;
  wire _abc_17692_n8431;
  wire _abc_17692_n8432;
  wire _abc_17692_n8433;
  wire _abc_17692_n8434;
  wire _abc_17692_n8435;
  wire _abc_17692_n8436;
  wire _abc_17692_n8437;
  wire _abc_17692_n8438;
  wire _abc_17692_n8439;
  wire _abc_17692_n844;
  wire _abc_17692_n8440;
  wire _abc_17692_n8441;
  wire _abc_17692_n8442;
  wire _abc_17692_n8443;
  wire _abc_17692_n8444;
  wire _abc_17692_n8445;
  wire _abc_17692_n8446;
  wire _abc_17692_n8447;
  wire _abc_17692_n8448;
  wire _abc_17692_n8449;
  wire _abc_17692_n845;
  wire _abc_17692_n8450;
  wire _abc_17692_n8451;
  wire _abc_17692_n8452;
  wire _abc_17692_n8453;
  wire _abc_17692_n8454;
  wire _abc_17692_n8455;
  wire _abc_17692_n8456;
  wire _abc_17692_n8457;
  wire _abc_17692_n8458;
  wire _abc_17692_n8459;
  wire _abc_17692_n8460;
  wire _abc_17692_n8461;
  wire _abc_17692_n8462;
  wire _abc_17692_n8463;
  wire _abc_17692_n8464;
  wire _abc_17692_n8465;
  wire _abc_17692_n8466;
  wire _abc_17692_n8467;
  wire _abc_17692_n8468;
  wire _abc_17692_n8469;
  wire _abc_17692_n847;
  wire _abc_17692_n8470;
  wire _abc_17692_n8471;
  wire _abc_17692_n8472;
  wire _abc_17692_n8473;
  wire _abc_17692_n8474;
  wire _abc_17692_n8475;
  wire _abc_17692_n8476;
  wire _abc_17692_n8477;
  wire _abc_17692_n8478;
  wire _abc_17692_n8479;
  wire _abc_17692_n848;
  wire _abc_17692_n8480;
  wire _abc_17692_n8481;
  wire _abc_17692_n8482;
  wire _abc_17692_n8483;
  wire _abc_17692_n8484;
  wire _abc_17692_n8485;
  wire _abc_17692_n8486;
  wire _abc_17692_n8487;
  wire _abc_17692_n8488;
  wire _abc_17692_n8489;
  wire _abc_17692_n8490;
  wire _abc_17692_n8491;
  wire _abc_17692_n8492;
  wire _abc_17692_n8493;
  wire _abc_17692_n8494;
  wire _abc_17692_n8496;
  wire _abc_17692_n8497;
  wire _abc_17692_n8498;
  wire _abc_17692_n8499;
  wire _abc_17692_n8500;
  wire _abc_17692_n8501;
  wire _abc_17692_n8502;
  wire _abc_17692_n8503;
  wire _abc_17692_n8504;
  wire _abc_17692_n8505;
  wire _abc_17692_n8506;
  wire _abc_17692_n8507;
  wire _abc_17692_n8508;
  wire _abc_17692_n8509;
  wire _abc_17692_n850_1;
  wire _abc_17692_n8510;
  wire _abc_17692_n8511;
  wire _abc_17692_n8512;
  wire _abc_17692_n8513;
  wire _abc_17692_n8514;
  wire _abc_17692_n8515;
  wire _abc_17692_n8516;
  wire _abc_17692_n8517;
  wire _abc_17692_n8518;
  wire _abc_17692_n8519;
  wire _abc_17692_n851_1;
  wire _abc_17692_n8520;
  wire _abc_17692_n8521;
  wire _abc_17692_n8522;
  wire _abc_17692_n8523;
  wire _abc_17692_n8524;
  wire _abc_17692_n8525;
  wire _abc_17692_n8526;
  wire _abc_17692_n8527;
  wire _abc_17692_n8528;
  wire _abc_17692_n8529;
  wire _abc_17692_n853;
  wire _abc_17692_n8530;
  wire _abc_17692_n8531;
  wire _abc_17692_n8532;
  wire _abc_17692_n8533;
  wire _abc_17692_n8534;
  wire _abc_17692_n8535;
  wire _abc_17692_n8536;
  wire _abc_17692_n8537;
  wire _abc_17692_n8538;
  wire _abc_17692_n8539;
  wire _abc_17692_n854;
  wire _abc_17692_n8540;
  wire _abc_17692_n8541;
  wire _abc_17692_n8542;
  wire _abc_17692_n8543;
  wire _abc_17692_n8544;
  wire _abc_17692_n8545;
  wire _abc_17692_n8546;
  wire _abc_17692_n8547;
  wire _abc_17692_n8548;
  wire _abc_17692_n8549;
  wire _abc_17692_n8550;
  wire _abc_17692_n8551;
  wire _abc_17692_n8552;
  wire _abc_17692_n8553;
  wire _abc_17692_n8554;
  wire _abc_17692_n8555;
  wire _abc_17692_n8556;
  wire _abc_17692_n8557;
  wire _abc_17692_n8558;
  wire _abc_17692_n8559;
  wire _abc_17692_n856;
  wire _abc_17692_n8560;
  wire _abc_17692_n8561;
  wire _abc_17692_n8562;
  wire _abc_17692_n8563;
  wire _abc_17692_n8564;
  wire _abc_17692_n8565;
  wire _abc_17692_n8566;
  wire _abc_17692_n8567;
  wire _abc_17692_n8568;
  wire _abc_17692_n8569;
  wire _abc_17692_n857;
  wire _abc_17692_n8570;
  wire _abc_17692_n8571;
  wire _abc_17692_n8572;
  wire _abc_17692_n8573;
  wire _abc_17692_n8574;
  wire _abc_17692_n8575;
  wire _abc_17692_n8576;
  wire _abc_17692_n8577;
  wire _abc_17692_n8578;
  wire _abc_17692_n8579;
  wire _abc_17692_n8580;
  wire _abc_17692_n8581;
  wire _abc_17692_n8582;
  wire _abc_17692_n8583;
  wire _abc_17692_n8584;
  wire _abc_17692_n8585;
  wire _abc_17692_n8586;
  wire _abc_17692_n8587;
  wire _abc_17692_n8588;
  wire _abc_17692_n8589;
  wire _abc_17692_n859;
  wire _abc_17692_n8590;
  wire _abc_17692_n8591;
  wire _abc_17692_n8592;
  wire _abc_17692_n8593;
  wire _abc_17692_n8594;
  wire _abc_17692_n8595;
  wire _abc_17692_n8596;
  wire _abc_17692_n8597;
  wire _abc_17692_n8598;
  wire _abc_17692_n8599;
  wire _abc_17692_n860;
  wire _abc_17692_n8600;
  wire _abc_17692_n8601;
  wire _abc_17692_n8602;
  wire _abc_17692_n8603;
  wire _abc_17692_n8604;
  wire _abc_17692_n8605;
  wire _abc_17692_n8606;
  wire _abc_17692_n8607;
  wire _abc_17692_n8608;
  wire _abc_17692_n8609;
  wire _abc_17692_n8610;
  wire _abc_17692_n8611;
  wire _abc_17692_n8612;
  wire _abc_17692_n8613;
  wire _abc_17692_n8614;
  wire _abc_17692_n8615;
  wire _abc_17692_n8616;
  wire _abc_17692_n8618;
  wire _abc_17692_n8619;
  wire _abc_17692_n862;
  wire _abc_17692_n8620;
  wire _abc_17692_n8621;
  wire _abc_17692_n8622;
  wire _abc_17692_n8623;
  wire _abc_17692_n8624;
  wire _abc_17692_n8625;
  wire _abc_17692_n8626;
  wire _abc_17692_n8627;
  wire _abc_17692_n8628;
  wire _abc_17692_n8629;
  wire _abc_17692_n863;
  wire _abc_17692_n8630;
  wire _abc_17692_n8631;
  wire _abc_17692_n8632;
  wire _abc_17692_n8633;
  wire _abc_17692_n8634;
  wire _abc_17692_n8635;
  wire _abc_17692_n8636;
  wire _abc_17692_n8637;
  wire _abc_17692_n8638;
  wire _abc_17692_n8639;
  wire _abc_17692_n8640;
  wire _abc_17692_n8641;
  wire _abc_17692_n8642;
  wire _abc_17692_n8643;
  wire _abc_17692_n8644;
  wire _abc_17692_n8645;
  wire _abc_17692_n8646;
  wire _abc_17692_n8647;
  wire _abc_17692_n8648;
  wire _abc_17692_n8649;
  wire _abc_17692_n865;
  wire _abc_17692_n8650;
  wire _abc_17692_n8651;
  wire _abc_17692_n8652;
  wire _abc_17692_n8653;
  wire _abc_17692_n8654;
  wire _abc_17692_n8655;
  wire _abc_17692_n8656;
  wire _abc_17692_n8657;
  wire _abc_17692_n8658;
  wire _abc_17692_n8659;
  wire _abc_17692_n866;
  wire _abc_17692_n8660;
  wire _abc_17692_n8661;
  wire _abc_17692_n8662;
  wire _abc_17692_n8663;
  wire _abc_17692_n8664;
  wire _abc_17692_n8665;
  wire _abc_17692_n8666;
  wire _abc_17692_n8667;
  wire _abc_17692_n8668;
  wire _abc_17692_n8669;
  wire _abc_17692_n8670;
  wire _abc_17692_n8671;
  wire _abc_17692_n8672;
  wire _abc_17692_n8673;
  wire _abc_17692_n8674;
  wire _abc_17692_n8675;
  wire _abc_17692_n8676;
  wire _abc_17692_n8677;
  wire _abc_17692_n8678;
  wire _abc_17692_n8679;
  wire _abc_17692_n868;
  wire _abc_17692_n8680;
  wire _abc_17692_n8681;
  wire _abc_17692_n8682;
  wire _abc_17692_n8683;
  wire _abc_17692_n8684;
  wire _abc_17692_n8685;
  wire _abc_17692_n8686;
  wire _abc_17692_n8687;
  wire _abc_17692_n8688;
  wire _abc_17692_n8689;
  wire _abc_17692_n869;
  wire _abc_17692_n8690;
  wire _abc_17692_n8691;
  wire _abc_17692_n8692;
  wire _abc_17692_n8693;
  wire _abc_17692_n8694;
  wire _abc_17692_n8695;
  wire _abc_17692_n8696;
  wire _abc_17692_n8697;
  wire _abc_17692_n8698;
  wire _abc_17692_n8699;
  wire _abc_17692_n8700;
  wire _abc_17692_n8701;
  wire _abc_17692_n8702;
  wire _abc_17692_n8703;
  wire _abc_17692_n8704;
  wire _abc_17692_n8705;
  wire _abc_17692_n8706;
  wire _abc_17692_n8707;
  wire _abc_17692_n8708;
  wire _abc_17692_n8709;
  wire _abc_17692_n871;
  wire _abc_17692_n8710;
  wire _abc_17692_n8711;
  wire _abc_17692_n8712;
  wire _abc_17692_n8713;
  wire _abc_17692_n8714;
  wire _abc_17692_n8715;
  wire _abc_17692_n8716;
  wire _abc_17692_n8717;
  wire _abc_17692_n8718;
  wire _abc_17692_n8719;
  wire _abc_17692_n872;
  wire _abc_17692_n8720;
  wire _abc_17692_n8721;
  wire _abc_17692_n8722;
  wire _abc_17692_n8723;
  wire _abc_17692_n8724;
  wire _abc_17692_n8725;
  wire _abc_17692_n8726;
  wire _abc_17692_n8727;
  wire _abc_17692_n8728;
  wire _abc_17692_n8729;
  wire _abc_17692_n8730;
  wire _abc_17692_n8731;
  wire _abc_17692_n8732;
  wire _abc_17692_n8733;
  wire _abc_17692_n8734;
  wire _abc_17692_n8735;
  wire _abc_17692_n8736;
  wire _abc_17692_n8737;
  wire _abc_17692_n8738;
  wire _abc_17692_n8739;
  wire _abc_17692_n874;
  wire _abc_17692_n8740;
  wire _abc_17692_n8742;
  wire _abc_17692_n8743;
  wire _abc_17692_n8744;
  wire _abc_17692_n8745;
  wire _abc_17692_n8746;
  wire _abc_17692_n8747;
  wire _abc_17692_n8748;
  wire _abc_17692_n8749;
  wire _abc_17692_n8750;
  wire _abc_17692_n8751;
  wire _abc_17692_n8752;
  wire _abc_17692_n8753;
  wire _abc_17692_n8754;
  wire _abc_17692_n8755;
  wire _abc_17692_n8756;
  wire _abc_17692_n8757;
  wire _abc_17692_n8758;
  wire _abc_17692_n8759;
  wire _abc_17692_n875_1;
  wire _abc_17692_n8760;
  wire _abc_17692_n8761;
  wire _abc_17692_n8762;
  wire _abc_17692_n8763;
  wire _abc_17692_n8764;
  wire _abc_17692_n8765;
  wire _abc_17692_n8766;
  wire _abc_17692_n8767;
  wire _abc_17692_n8768;
  wire _abc_17692_n8769;
  wire _abc_17692_n877;
  wire _abc_17692_n8770;
  wire _abc_17692_n8771;
  wire _abc_17692_n8772;
  wire _abc_17692_n8773;
  wire _abc_17692_n8774;
  wire _abc_17692_n8775;
  wire _abc_17692_n8776;
  wire _abc_17692_n8777;
  wire _abc_17692_n8778;
  wire _abc_17692_n8779;
  wire _abc_17692_n878;
  wire _abc_17692_n8780;
  wire _abc_17692_n8781;
  wire _abc_17692_n8782;
  wire _abc_17692_n8783;
  wire _abc_17692_n8784;
  wire _abc_17692_n8785;
  wire _abc_17692_n8786;
  wire _abc_17692_n8787;
  wire _abc_17692_n8788;
  wire _abc_17692_n8789;
  wire _abc_17692_n8790;
  wire _abc_17692_n8791;
  wire _abc_17692_n8792;
  wire _abc_17692_n8793;
  wire _abc_17692_n8794;
  wire _abc_17692_n8795;
  wire _abc_17692_n8796;
  wire _abc_17692_n8797;
  wire _abc_17692_n8798;
  wire _abc_17692_n8799;
  wire _abc_17692_n880;
  wire _abc_17692_n8800;
  wire _abc_17692_n8801;
  wire _abc_17692_n8802;
  wire _abc_17692_n8803;
  wire _abc_17692_n8804;
  wire _abc_17692_n8805;
  wire _abc_17692_n8806;
  wire _abc_17692_n8807;
  wire _abc_17692_n8808;
  wire _abc_17692_n8809;
  wire _abc_17692_n881;
  wire _abc_17692_n8810;
  wire _abc_17692_n8811;
  wire _abc_17692_n8812;
  wire _abc_17692_n8813;
  wire _abc_17692_n8814;
  wire _abc_17692_n8815;
  wire _abc_17692_n8816;
  wire _abc_17692_n8817;
  wire _abc_17692_n8818;
  wire _abc_17692_n8819;
  wire _abc_17692_n8820;
  wire _abc_17692_n8821;
  wire _abc_17692_n8822;
  wire _abc_17692_n8823;
  wire _abc_17692_n8824;
  wire _abc_17692_n8825;
  wire _abc_17692_n8826;
  wire _abc_17692_n8827;
  wire _abc_17692_n8828;
  wire _abc_17692_n8829;
  wire _abc_17692_n883;
  wire _abc_17692_n8830;
  wire _abc_17692_n8831;
  wire _abc_17692_n8832;
  wire _abc_17692_n8833;
  wire _abc_17692_n8834;
  wire _abc_17692_n8835;
  wire _abc_17692_n8836;
  wire _abc_17692_n8837;
  wire _abc_17692_n8838;
  wire _abc_17692_n8839;
  wire _abc_17692_n884;
  wire _abc_17692_n8840;
  wire _abc_17692_n8841;
  wire _abc_17692_n8842;
  wire _abc_17692_n8843;
  wire _abc_17692_n8844;
  wire _abc_17692_n8845;
  wire _abc_17692_n8846;
  wire _abc_17692_n8847;
  wire _abc_17692_n8848;
  wire _abc_17692_n8849;
  wire _abc_17692_n8850;
  wire _abc_17692_n8851;
  wire _abc_17692_n8852;
  wire _abc_17692_n8853;
  wire _abc_17692_n8854;
  wire _abc_17692_n8855;
  wire _abc_17692_n8856;
  wire _abc_17692_n8857;
  wire _abc_17692_n8858;
  wire _abc_17692_n8859;
  wire _abc_17692_n886;
  wire _abc_17692_n8860;
  wire _abc_17692_n8861;
  wire _abc_17692_n8862;
  wire _abc_17692_n8863;
  wire _abc_17692_n8864;
  wire _abc_17692_n8865;
  wire _abc_17692_n8866;
  wire _abc_17692_n8867;
  wire _abc_17692_n8868;
  wire _abc_17692_n8869;
  wire _abc_17692_n887;
  wire _abc_17692_n8870;
  wire _abc_17692_n8871;
  wire _abc_17692_n8873;
  wire _abc_17692_n8874;
  wire _abc_17692_n8875;
  wire _abc_17692_n8876;
  wire _abc_17692_n8877;
  wire _abc_17692_n8878;
  wire _abc_17692_n8879;
  wire _abc_17692_n8880;
  wire _abc_17692_n8881;
  wire _abc_17692_n8882;
  wire _abc_17692_n8883;
  wire _abc_17692_n8884;
  wire _abc_17692_n8885;
  wire _abc_17692_n8886;
  wire _abc_17692_n8887;
  wire _abc_17692_n8888;
  wire _abc_17692_n8889;
  wire _abc_17692_n8890;
  wire _abc_17692_n8891;
  wire _abc_17692_n8892;
  wire _abc_17692_n8893;
  wire _abc_17692_n8894;
  wire _abc_17692_n8895;
  wire _abc_17692_n8896;
  wire _abc_17692_n8897;
  wire _abc_17692_n8898;
  wire _abc_17692_n8899;
  wire _abc_17692_n889_1;
  wire _abc_17692_n8900;
  wire _abc_17692_n8901;
  wire _abc_17692_n8902;
  wire _abc_17692_n8903;
  wire _abc_17692_n8904;
  wire _abc_17692_n8905;
  wire _abc_17692_n8906;
  wire _abc_17692_n8907;
  wire _abc_17692_n8908;
  wire _abc_17692_n8909;
  wire _abc_17692_n890_1;
  wire _abc_17692_n8910;
  wire _abc_17692_n8911;
  wire _abc_17692_n8912;
  wire _abc_17692_n8913;
  wire _abc_17692_n8914;
  wire _abc_17692_n8915;
  wire _abc_17692_n8916;
  wire _abc_17692_n8917;
  wire _abc_17692_n8918;
  wire _abc_17692_n8919;
  wire _abc_17692_n892;
  wire _abc_17692_n8920;
  wire _abc_17692_n8921;
  wire _abc_17692_n8922;
  wire _abc_17692_n8923;
  wire _abc_17692_n8924;
  wire _abc_17692_n8925;
  wire _abc_17692_n8926;
  wire _abc_17692_n8927;
  wire _abc_17692_n8928;
  wire _abc_17692_n8929;
  wire _abc_17692_n893;
  wire _abc_17692_n8930;
  wire _abc_17692_n8931;
  wire _abc_17692_n8932;
  wire _abc_17692_n8933;
  wire _abc_17692_n8934;
  wire _abc_17692_n8935;
  wire _abc_17692_n8936;
  wire _abc_17692_n8937;
  wire _abc_17692_n8938;
  wire _abc_17692_n8939;
  wire _abc_17692_n8940;
  wire _abc_17692_n8941;
  wire _abc_17692_n8942;
  wire _abc_17692_n8943;
  wire _abc_17692_n8944;
  wire _abc_17692_n8945;
  wire _abc_17692_n8946;
  wire _abc_17692_n8947;
  wire _abc_17692_n8948;
  wire _abc_17692_n8949;
  wire _abc_17692_n895;
  wire _abc_17692_n8950;
  wire _abc_17692_n8951;
  wire _abc_17692_n8952;
  wire _abc_17692_n8953;
  wire _abc_17692_n8954;
  wire _abc_17692_n8955;
  wire _abc_17692_n8956;
  wire _abc_17692_n8957;
  wire _abc_17692_n8958;
  wire _abc_17692_n8959;
  wire _abc_17692_n896;
  wire _abc_17692_n8960;
  wire _abc_17692_n8961;
  wire _abc_17692_n8962;
  wire _abc_17692_n8963;
  wire _abc_17692_n8964;
  wire _abc_17692_n8965;
  wire _abc_17692_n8966;
  wire _abc_17692_n8967;
  wire _abc_17692_n8968;
  wire _abc_17692_n8969;
  wire _abc_17692_n8970;
  wire _abc_17692_n8971;
  wire _abc_17692_n8972;
  wire _abc_17692_n8973;
  wire _abc_17692_n8974;
  wire _abc_17692_n8975;
  wire _abc_17692_n8976;
  wire _abc_17692_n8977;
  wire _abc_17692_n8978;
  wire _abc_17692_n8979;
  wire _abc_17692_n898;
  wire _abc_17692_n8980;
  wire _abc_17692_n8981;
  wire _abc_17692_n8982;
  wire _abc_17692_n8983;
  wire _abc_17692_n8984;
  wire _abc_17692_n8985;
  wire _abc_17692_n8986;
  wire _abc_17692_n8987;
  wire _abc_17692_n8988;
  wire _abc_17692_n8989;
  wire _abc_17692_n899;
  wire _abc_17692_n8990;
  wire _abc_17692_n8991;
  wire _abc_17692_n8992;
  wire _abc_17692_n8993;
  wire _abc_17692_n8994;
  wire _abc_17692_n8995;
  wire _abc_17692_n8996;
  wire _abc_17692_n8997;
  wire _abc_17692_n8998;
  wire _abc_17692_n9000;
  wire _abc_17692_n9001;
  wire _abc_17692_n9002;
  wire _abc_17692_n9003;
  wire _abc_17692_n9004;
  wire _abc_17692_n9005;
  wire _abc_17692_n9006;
  wire _abc_17692_n9007;
  wire _abc_17692_n9008;
  wire _abc_17692_n9009;
  wire _abc_17692_n901;
  wire _abc_17692_n9010;
  wire _abc_17692_n9011;
  wire _abc_17692_n9012;
  wire _abc_17692_n9013;
  wire _abc_17692_n9014;
  wire _abc_17692_n9015;
  wire _abc_17692_n9016;
  wire _abc_17692_n9017;
  wire _abc_17692_n9018;
  wire _abc_17692_n9019;
  wire _abc_17692_n902;
  wire _abc_17692_n9020;
  wire _abc_17692_n9021;
  wire _abc_17692_n9022;
  wire _abc_17692_n9023;
  wire _abc_17692_n9024;
  wire _abc_17692_n9025;
  wire _abc_17692_n9026;
  wire _abc_17692_n9027;
  wire _abc_17692_n9028;
  wire _abc_17692_n9029;
  wire _abc_17692_n9030;
  wire _abc_17692_n9031;
  wire _abc_17692_n9032;
  wire _abc_17692_n9033;
  wire _abc_17692_n9034;
  wire _abc_17692_n9035;
  wire _abc_17692_n9036;
  wire _abc_17692_n9037;
  wire _abc_17692_n9038;
  wire _abc_17692_n9039;
  wire _abc_17692_n904;
  wire _abc_17692_n9040;
  wire _abc_17692_n9041;
  wire _abc_17692_n9042;
  wire _abc_17692_n9043;
  wire _abc_17692_n9044;
  wire _abc_17692_n9045;
  wire _abc_17692_n9046;
  wire _abc_17692_n9047;
  wire _abc_17692_n9048;
  wire _abc_17692_n9049;
  wire _abc_17692_n905;
  wire _abc_17692_n9050;
  wire _abc_17692_n9051;
  wire _abc_17692_n9052;
  wire _abc_17692_n9053;
  wire _abc_17692_n9054;
  wire _abc_17692_n9055;
  wire _abc_17692_n9056;
  wire _abc_17692_n9057;
  wire _abc_17692_n9058;
  wire _abc_17692_n9059;
  wire _abc_17692_n9060;
  wire _abc_17692_n9061;
  wire _abc_17692_n9062;
  wire _abc_17692_n9063;
  wire _abc_17692_n9064;
  wire _abc_17692_n9065;
  wire _abc_17692_n9066;
  wire _abc_17692_n9067;
  wire _abc_17692_n9068;
  wire _abc_17692_n9069;
  wire _abc_17692_n907;
  wire _abc_17692_n9070;
  wire _abc_17692_n9071;
  wire _abc_17692_n9072;
  wire _abc_17692_n9073;
  wire _abc_17692_n9074;
  wire _abc_17692_n9075;
  wire _abc_17692_n9076;
  wire _abc_17692_n9077;
  wire _abc_17692_n9078;
  wire _abc_17692_n9079;
  wire _abc_17692_n908;
  wire _abc_17692_n9080;
  wire _abc_17692_n9081;
  wire _abc_17692_n9082;
  wire _abc_17692_n9083;
  wire _abc_17692_n9084;
  wire _abc_17692_n9085;
  wire _abc_17692_n9086;
  wire _abc_17692_n9087;
  wire _abc_17692_n9088;
  wire _abc_17692_n9089;
  wire _abc_17692_n9090;
  wire _abc_17692_n9091;
  wire _abc_17692_n9092;
  wire _abc_17692_n9093;
  wire _abc_17692_n9094;
  wire _abc_17692_n9095;
  wire _abc_17692_n9096;
  wire _abc_17692_n9097;
  wire _abc_17692_n9098;
  wire _abc_17692_n9099;
  wire _abc_17692_n9100;
  wire _abc_17692_n9101;
  wire _abc_17692_n9102;
  wire _abc_17692_n9103;
  wire _abc_17692_n9104;
  wire _abc_17692_n9105;
  wire _abc_17692_n9106;
  wire _abc_17692_n9107;
  wire _abc_17692_n9108;
  wire _abc_17692_n9109;
  wire _abc_17692_n910_1;
  wire _abc_17692_n9110;
  wire _abc_17692_n9111;
  wire _abc_17692_n9112;
  wire _abc_17692_n9113;
  wire _abc_17692_n9114;
  wire _abc_17692_n9115;
  wire _abc_17692_n9116;
  wire _abc_17692_n9117;
  wire _abc_17692_n9118;
  wire _abc_17692_n9119;
  wire _abc_17692_n911_1;
  wire _abc_17692_n9120;
  wire _abc_17692_n9121;
  wire _abc_17692_n9122;
  wire _abc_17692_n9123;
  wire _abc_17692_n9124;
  wire _abc_17692_n9125;
  wire _abc_17692_n9126;
  wire _abc_17692_n9127;
  wire _abc_17692_n9128;
  wire _abc_17692_n9129;
  wire _abc_17692_n913;
  wire _abc_17692_n9130;
  wire _abc_17692_n9131;
  wire _abc_17692_n9132;
  wire _abc_17692_n9133;
  wire _abc_17692_n9134;
  wire _abc_17692_n9136;
  wire _abc_17692_n9137;
  wire _abc_17692_n9138;
  wire _abc_17692_n9139;
  wire _abc_17692_n914;
  wire _abc_17692_n9140;
  wire _abc_17692_n9141;
  wire _abc_17692_n9142;
  wire _abc_17692_n9143;
  wire _abc_17692_n9144;
  wire _abc_17692_n9145;
  wire _abc_17692_n9146;
  wire _abc_17692_n9147;
  wire _abc_17692_n9148;
  wire _abc_17692_n9149;
  wire _abc_17692_n9150;
  wire _abc_17692_n9151;
  wire _abc_17692_n9152;
  wire _abc_17692_n9153;
  wire _abc_17692_n9154;
  wire _abc_17692_n9155;
  wire _abc_17692_n9156;
  wire _abc_17692_n9157;
  wire _abc_17692_n9158;
  wire _abc_17692_n9159;
  wire _abc_17692_n916;
  wire _abc_17692_n9160;
  wire _abc_17692_n9161;
  wire _abc_17692_n9162;
  wire _abc_17692_n9163;
  wire _abc_17692_n9164;
  wire _abc_17692_n9165;
  wire _abc_17692_n9166;
  wire _abc_17692_n9167;
  wire _abc_17692_n9168;
  wire _abc_17692_n9169;
  wire _abc_17692_n917;
  wire _abc_17692_n9170;
  wire _abc_17692_n9171;
  wire _abc_17692_n9172;
  wire _abc_17692_n9173;
  wire _abc_17692_n9174;
  wire _abc_17692_n9175;
  wire _abc_17692_n9176;
  wire _abc_17692_n9177;
  wire _abc_17692_n9178;
  wire _abc_17692_n9179;
  wire _abc_17692_n9180;
  wire _abc_17692_n9181;
  wire _abc_17692_n9182;
  wire _abc_17692_n9183;
  wire _abc_17692_n9184;
  wire _abc_17692_n9185;
  wire _abc_17692_n9186;
  wire _abc_17692_n9187;
  wire _abc_17692_n9188;
  wire _abc_17692_n9189;
  wire _abc_17692_n919;
  wire _abc_17692_n9190;
  wire _abc_17692_n9191;
  wire _abc_17692_n9192;
  wire _abc_17692_n9193;
  wire _abc_17692_n9194;
  wire _abc_17692_n9195;
  wire _abc_17692_n9196;
  wire _abc_17692_n9197;
  wire _abc_17692_n9198;
  wire _abc_17692_n9199;
  wire _abc_17692_n920;
  wire _abc_17692_n9200;
  wire _abc_17692_n9201;
  wire _abc_17692_n9202;
  wire _abc_17692_n9203;
  wire _abc_17692_n9204;
  wire _abc_17692_n9205;
  wire _abc_17692_n9206;
  wire _abc_17692_n9207;
  wire _abc_17692_n9208;
  wire _abc_17692_n9209;
  wire _abc_17692_n921;
  wire _abc_17692_n9210;
  wire _abc_17692_n9211;
  wire _abc_17692_n9212;
  wire _abc_17692_n9213;
  wire _abc_17692_n9214;
  wire _abc_17692_n9215;
  wire _abc_17692_n9216;
  wire _abc_17692_n9217;
  wire _abc_17692_n9218;
  wire _abc_17692_n9219;
  wire _abc_17692_n922;
  wire _abc_17692_n9220;
  wire _abc_17692_n9221;
  wire _abc_17692_n9222;
  wire _abc_17692_n9223;
  wire _abc_17692_n9224;
  wire _abc_17692_n9225;
  wire _abc_17692_n9226;
  wire _abc_17692_n9227;
  wire _abc_17692_n9228;
  wire _abc_17692_n9229;
  wire _abc_17692_n9230;
  wire _abc_17692_n9231;
  wire _abc_17692_n9232;
  wire _abc_17692_n9233;
  wire _abc_17692_n9234;
  wire _abc_17692_n9235;
  wire _abc_17692_n9236;
  wire _abc_17692_n9237;
  wire _abc_17692_n9238;
  wire _abc_17692_n9239;
  wire _abc_17692_n923_1;
  wire _abc_17692_n924;
  wire _abc_17692_n9240;
  wire _abc_17692_n9241;
  wire _abc_17692_n9242;
  wire _abc_17692_n9243;
  wire _abc_17692_n9244;
  wire _abc_17692_n9245;
  wire _abc_17692_n9246;
  wire _abc_17692_n9247;
  wire _abc_17692_n9248;
  wire _abc_17692_n9249;
  wire _abc_17692_n9250;
  wire _abc_17692_n9251;
  wire _abc_17692_n9252;
  wire _abc_17692_n9253;
  wire _abc_17692_n9254;
  wire _abc_17692_n9255;
  wire _abc_17692_n9256;
  wire _abc_17692_n9257;
  wire _abc_17692_n9258;
  wire _abc_17692_n9259;
  wire _abc_17692_n9260;
  wire _abc_17692_n9261;
  wire _abc_17692_n9262;
  wire _abc_17692_n9263;
  wire _abc_17692_n9264;
  wire _abc_17692_n9265;
  wire _abc_17692_n9266;
  wire _abc_17692_n9267;
  wire _abc_17692_n9268;
  wire _abc_17692_n926_1;
  wire _abc_17692_n9270;
  wire _abc_17692_n9271;
  wire _abc_17692_n9272;
  wire _abc_17692_n9273;
  wire _abc_17692_n9274;
  wire _abc_17692_n9275;
  wire _abc_17692_n9276;
  wire _abc_17692_n9277;
  wire _abc_17692_n9278;
  wire _abc_17692_n9279;
  wire _abc_17692_n927_1;
  wire _abc_17692_n928;
  wire _abc_17692_n9280;
  wire _abc_17692_n9281;
  wire _abc_17692_n9282;
  wire _abc_17692_n9283;
  wire _abc_17692_n9284;
  wire _abc_17692_n9285;
  wire _abc_17692_n9286;
  wire _abc_17692_n9287;
  wire _abc_17692_n9288;
  wire _abc_17692_n9289;
  wire _abc_17692_n929;
  wire _abc_17692_n9290;
  wire _abc_17692_n9291;
  wire _abc_17692_n9292;
  wire _abc_17692_n9293;
  wire _abc_17692_n9294;
  wire _abc_17692_n9295;
  wire _abc_17692_n9296;
  wire _abc_17692_n9297;
  wire _abc_17692_n9298;
  wire _abc_17692_n9299;
  wire _abc_17692_n9300;
  wire _abc_17692_n9301;
  wire _abc_17692_n9302;
  wire _abc_17692_n9303;
  wire _abc_17692_n9304;
  wire _abc_17692_n9305;
  wire _abc_17692_n9306;
  wire _abc_17692_n9307;
  wire _abc_17692_n9308;
  wire _abc_17692_n9309;
  wire _abc_17692_n930_1;
  wire _abc_17692_n931;
  wire _abc_17692_n9310;
  wire _abc_17692_n9311;
  wire _abc_17692_n9312;
  wire _abc_17692_n9313;
  wire _abc_17692_n9314;
  wire _abc_17692_n9315;
  wire _abc_17692_n9316;
  wire _abc_17692_n9317;
  wire _abc_17692_n9318;
  wire _abc_17692_n9319;
  wire _abc_17692_n932;
  wire _abc_17692_n9320;
  wire _abc_17692_n9321;
  wire _abc_17692_n9322;
  wire _abc_17692_n9323;
  wire _abc_17692_n9324;
  wire _abc_17692_n9325;
  wire _abc_17692_n9326;
  wire _abc_17692_n9327;
  wire _abc_17692_n9328;
  wire _abc_17692_n9329;
  wire _abc_17692_n933;
  wire _abc_17692_n9330;
  wire _abc_17692_n9331;
  wire _abc_17692_n9332;
  wire _abc_17692_n9333;
  wire _abc_17692_n9334;
  wire _abc_17692_n9335;
  wire _abc_17692_n9336;
  wire _abc_17692_n9337;
  wire _abc_17692_n9338;
  wire _abc_17692_n9339;
  wire _abc_17692_n934;
  wire _abc_17692_n9340;
  wire _abc_17692_n9341;
  wire _abc_17692_n9342;
  wire _abc_17692_n9343;
  wire _abc_17692_n9344;
  wire _abc_17692_n9345;
  wire _abc_17692_n9346;
  wire _abc_17692_n9347;
  wire _abc_17692_n9348;
  wire _abc_17692_n9349;
  wire _abc_17692_n935;
  wire _abc_17692_n9350;
  wire _abc_17692_n9351;
  wire _abc_17692_n9352;
  wire _abc_17692_n9353;
  wire _abc_17692_n9354;
  wire _abc_17692_n9355;
  wire _abc_17692_n9356;
  wire _abc_17692_n9357;
  wire _abc_17692_n9358;
  wire _abc_17692_n9359;
  wire _abc_17692_n936;
  wire _abc_17692_n9360;
  wire _abc_17692_n9361;
  wire _abc_17692_n9362;
  wire _abc_17692_n9363;
  wire _abc_17692_n9364;
  wire _abc_17692_n9365;
  wire _abc_17692_n9366;
  wire _abc_17692_n9367;
  wire _abc_17692_n9368;
  wire _abc_17692_n9369;
  wire _abc_17692_n9370;
  wire _abc_17692_n9371;
  wire _abc_17692_n9372;
  wire _abc_17692_n9373;
  wire _abc_17692_n9374;
  wire _abc_17692_n9375;
  wire _abc_17692_n9376;
  wire _abc_17692_n9377;
  wire _abc_17692_n9378;
  wire _abc_17692_n9379;
  wire _abc_17692_n937_1;
  wire _abc_17692_n938;
  wire _abc_17692_n9380;
  wire _abc_17692_n9381;
  wire _abc_17692_n9382;
  wire _abc_17692_n9383;
  wire _abc_17692_n9384;
  wire _abc_17692_n9385;
  wire _abc_17692_n9386;
  wire _abc_17692_n9387;
  wire _abc_17692_n9388;
  wire _abc_17692_n9389;
  wire _abc_17692_n939;
  wire _abc_17692_n9390;
  wire _abc_17692_n9391;
  wire _abc_17692_n9392;
  wire _abc_17692_n9393;
  wire _abc_17692_n9394;
  wire _abc_17692_n9395;
  wire _abc_17692_n9396;
  wire _abc_17692_n9397;
  wire _abc_17692_n9398;
  wire _abc_17692_n9399;
  wire _abc_17692_n940;
  wire _abc_17692_n9400;
  wire _abc_17692_n9401;
  wire _abc_17692_n9402;
  wire _abc_17692_n9403;
  wire _abc_17692_n9404;
  wire _abc_17692_n9405;
  wire _abc_17692_n9406;
  wire _abc_17692_n9407;
  wire _abc_17692_n9408;
  wire _abc_17692_n9409;
  wire _abc_17692_n941;
  wire _abc_17692_n9410;
  wire _abc_17692_n9411;
  wire _abc_17692_n9412;
  wire _abc_17692_n9413;
  wire _abc_17692_n9414;
  wire _abc_17692_n9415;
  wire _abc_17692_n9417;
  wire _abc_17692_n9418;
  wire _abc_17692_n9419;
  wire _abc_17692_n942;
  wire _abc_17692_n9420;
  wire _abc_17692_n9421;
  wire _abc_17692_n9422;
  wire _abc_17692_n9423;
  wire _abc_17692_n9424;
  wire _abc_17692_n9425;
  wire _abc_17692_n9426;
  wire _abc_17692_n9427;
  wire _abc_17692_n9428;
  wire _abc_17692_n9429;
  wire _abc_17692_n943;
  wire _abc_17692_n9430;
  wire _abc_17692_n9431;
  wire _abc_17692_n9432;
  wire _abc_17692_n9433;
  wire _abc_17692_n9434;
  wire _abc_17692_n9435;
  wire _abc_17692_n9436;
  wire _abc_17692_n9437;
  wire _abc_17692_n9438;
  wire _abc_17692_n9439;
  wire _abc_17692_n944;
  wire _abc_17692_n9440;
  wire _abc_17692_n9441;
  wire _abc_17692_n9442;
  wire _abc_17692_n9443;
  wire _abc_17692_n9444;
  wire _abc_17692_n9445;
  wire _abc_17692_n9446;
  wire _abc_17692_n9447;
  wire _abc_17692_n9448;
  wire _abc_17692_n9449;
  wire _abc_17692_n9450;
  wire _abc_17692_n9451;
  wire _abc_17692_n9452;
  wire _abc_17692_n9453;
  wire _abc_17692_n9454;
  wire _abc_17692_n9455;
  wire _abc_17692_n9456;
  wire _abc_17692_n9457;
  wire _abc_17692_n9458;
  wire _abc_17692_n9459;
  wire _abc_17692_n946;
  wire _abc_17692_n9460;
  wire _abc_17692_n9461;
  wire _abc_17692_n9462;
  wire _abc_17692_n9463;
  wire _abc_17692_n9464;
  wire _abc_17692_n9465;
  wire _abc_17692_n9466;
  wire _abc_17692_n9467;
  wire _abc_17692_n9468;
  wire _abc_17692_n9469;
  wire _abc_17692_n947;
  wire _abc_17692_n9470;
  wire _abc_17692_n9471;
  wire _abc_17692_n9472;
  wire _abc_17692_n9473;
  wire _abc_17692_n9474;
  wire _abc_17692_n9475;
  wire _abc_17692_n9476;
  wire _abc_17692_n9477;
  wire _abc_17692_n9478;
  wire _abc_17692_n9479;
  wire _abc_17692_n948;
  wire _abc_17692_n9480;
  wire _abc_17692_n9481;
  wire _abc_17692_n9482;
  wire _abc_17692_n9483;
  wire _abc_17692_n9484;
  wire _abc_17692_n9485;
  wire _abc_17692_n9486;
  wire _abc_17692_n9487;
  wire _abc_17692_n9488;
  wire _abc_17692_n9489;
  wire _abc_17692_n9490;
  wire _abc_17692_n9491;
  wire _abc_17692_n9492;
  wire _abc_17692_n9493;
  wire _abc_17692_n9494;
  wire _abc_17692_n9495;
  wire _abc_17692_n9496;
  wire _abc_17692_n9497;
  wire _abc_17692_n9498;
  wire _abc_17692_n9499;
  wire _abc_17692_n949_1;
  wire _abc_17692_n950;
  wire _abc_17692_n9500;
  wire _abc_17692_n9501;
  wire _abc_17692_n9502;
  wire _abc_17692_n9503;
  wire _abc_17692_n9504;
  wire _abc_17692_n9505;
  wire _abc_17692_n9506;
  wire _abc_17692_n9507;
  wire _abc_17692_n9508;
  wire _abc_17692_n9509;
  wire _abc_17692_n951;
  wire _abc_17692_n9510;
  wire _abc_17692_n9511;
  wire _abc_17692_n9512;
  wire _abc_17692_n9513;
  wire _abc_17692_n9514;
  wire _abc_17692_n9515;
  wire _abc_17692_n9516;
  wire _abc_17692_n9517;
  wire _abc_17692_n9518;
  wire _abc_17692_n9519;
  wire _abc_17692_n952;
  wire _abc_17692_n9520;
  wire _abc_17692_n9521;
  wire _abc_17692_n9522;
  wire _abc_17692_n9523;
  wire _abc_17692_n9524;
  wire _abc_17692_n9525;
  wire _abc_17692_n9526;
  wire _abc_17692_n9527;
  wire _abc_17692_n9528;
  wire _abc_17692_n9529;
  wire _abc_17692_n953;
  wire _abc_17692_n9530;
  wire _abc_17692_n9531;
  wire _abc_17692_n9532;
  wire _abc_17692_n9533;
  wire _abc_17692_n9534;
  wire _abc_17692_n9535;
  wire _abc_17692_n9536;
  wire _abc_17692_n9537;
  wire _abc_17692_n9538;
  wire _abc_17692_n9539;
  wire _abc_17692_n954;
  wire _abc_17692_n9540;
  wire _abc_17692_n9542;
  wire _abc_17692_n9543;
  wire _abc_17692_n9544;
  wire _abc_17692_n9545;
  wire _abc_17692_n9546;
  wire _abc_17692_n9547;
  wire _abc_17692_n9548;
  wire _abc_17692_n9549;
  wire _abc_17692_n955;
  wire _abc_17692_n9550;
  wire _abc_17692_n9551;
  wire _abc_17692_n9552;
  wire _abc_17692_n9553;
  wire _abc_17692_n9554;
  wire _abc_17692_n9555;
  wire _abc_17692_n9556;
  wire _abc_17692_n9557;
  wire _abc_17692_n9558;
  wire _abc_17692_n9559;
  wire _abc_17692_n956;
  wire _abc_17692_n9560;
  wire _abc_17692_n9561;
  wire _abc_17692_n9562;
  wire _abc_17692_n9563;
  wire _abc_17692_n9564;
  wire _abc_17692_n9565;
  wire _abc_17692_n9566;
  wire _abc_17692_n9567;
  wire _abc_17692_n9568;
  wire _abc_17692_n9569;
  wire _abc_17692_n957;
  wire _abc_17692_n9570;
  wire _abc_17692_n9571;
  wire _abc_17692_n9572;
  wire _abc_17692_n9573;
  wire _abc_17692_n9574;
  wire _abc_17692_n9575;
  wire _abc_17692_n9576;
  wire _abc_17692_n9577;
  wire _abc_17692_n9578;
  wire _abc_17692_n9579;
  wire _abc_17692_n958;
  wire _abc_17692_n9580;
  wire _abc_17692_n9581;
  wire _abc_17692_n9582;
  wire _abc_17692_n9583;
  wire _abc_17692_n9584;
  wire _abc_17692_n9585;
  wire _abc_17692_n9586;
  wire _abc_17692_n9587;
  wire _abc_17692_n9588;
  wire _abc_17692_n9589;
  wire _abc_17692_n959;
  wire _abc_17692_n9590;
  wire _abc_17692_n9591;
  wire _abc_17692_n9592;
  wire _abc_17692_n9593;
  wire _abc_17692_n9594;
  wire _abc_17692_n9595;
  wire _abc_17692_n9596;
  wire _abc_17692_n9597;
  wire _abc_17692_n9598;
  wire _abc_17692_n9599;
  wire _abc_17692_n960;
  wire _abc_17692_n9600;
  wire _abc_17692_n9601;
  wire _abc_17692_n9602;
  wire _abc_17692_n9603;
  wire _abc_17692_n9604;
  wire _abc_17692_n9605;
  wire _abc_17692_n9606;
  wire _abc_17692_n9607;
  wire _abc_17692_n9608;
  wire _abc_17692_n9609;
  wire _abc_17692_n961;
  wire _abc_17692_n9610;
  wire _abc_17692_n9611;
  wire _abc_17692_n9612;
  wire _abc_17692_n9613;
  wire _abc_17692_n9614;
  wire _abc_17692_n9615;
  wire _abc_17692_n9616;
  wire _abc_17692_n9617;
  wire _abc_17692_n9618;
  wire _abc_17692_n9619;
  wire _abc_17692_n962;
  wire _abc_17692_n9620;
  wire _abc_17692_n9621;
  wire _abc_17692_n9622;
  wire _abc_17692_n9623;
  wire _abc_17692_n9624;
  wire _abc_17692_n9625;
  wire _abc_17692_n9626;
  wire _abc_17692_n9627;
  wire _abc_17692_n9628;
  wire _abc_17692_n9629;
  wire _abc_17692_n963;
  wire _abc_17692_n9630;
  wire _abc_17692_n9631;
  wire _abc_17692_n9632;
  wire _abc_17692_n9633;
  wire _abc_17692_n9634;
  wire _abc_17692_n9635;
  wire _abc_17692_n9636;
  wire _abc_17692_n9637;
  wire _abc_17692_n9638;
  wire _abc_17692_n9639;
  wire _abc_17692_n9640;
  wire _abc_17692_n9641;
  wire _abc_17692_n9642;
  wire _abc_17692_n9643;
  wire _abc_17692_n9644;
  wire _abc_17692_n9645;
  wire _abc_17692_n9646;
  wire _abc_17692_n9647;
  wire _abc_17692_n9648;
  wire _abc_17692_n9649;
  wire _abc_17692_n964_1;
  wire _abc_17692_n965;
  wire _abc_17692_n9650;
  wire _abc_17692_n9651;
  wire _abc_17692_n9652;
  wire _abc_17692_n9653;
  wire _abc_17692_n9654;
  wire _abc_17692_n9655;
  wire _abc_17692_n9656;
  wire _abc_17692_n9657;
  wire _abc_17692_n9658;
  wire _abc_17692_n9659;
  wire _abc_17692_n966;
  wire _abc_17692_n9660;
  wire _abc_17692_n9661;
  wire _abc_17692_n9662;
  wire _abc_17692_n9663;
  wire _abc_17692_n9664;
  wire _abc_17692_n9665;
  wire _abc_17692_n9666;
  wire _abc_17692_n9667;
  wire _abc_17692_n9668;
  wire _abc_17692_n9669;
  wire _abc_17692_n9670;
  wire _abc_17692_n9671;
  wire _abc_17692_n9672;
  wire _abc_17692_n9673;
  wire _abc_17692_n9674;
  wire _abc_17692_n9675;
  wire _abc_17692_n9676;
  wire _abc_17692_n9677;
  wire _abc_17692_n9678;
  wire _abc_17692_n9679;
  wire _abc_17692_n967_1;
  wire _abc_17692_n9680;
  wire _abc_17692_n9681;
  wire _abc_17692_n9682;
  wire _abc_17692_n9683;
  wire _abc_17692_n9684;
  wire _abc_17692_n9685;
  wire _abc_17692_n9686;
  wire _abc_17692_n9687;
  wire _abc_17692_n9688;
  wire _abc_17692_n9689;
  wire _abc_17692_n969;
  wire _abc_17692_n9690;
  wire _abc_17692_n9691;
  wire _abc_17692_n9692;
  wire _abc_17692_n9693;
  wire _abc_17692_n9694;
  wire _abc_17692_n9695;
  wire _abc_17692_n9696;
  wire _abc_17692_n9697;
  wire _abc_17692_n9698;
  wire _abc_17692_n9699;
  wire _abc_17692_n970;
  wire _abc_17692_n9700;
  wire _abc_17692_n9701;
  wire _abc_17692_n9702;
  wire _abc_17692_n9703;
  wire _abc_17692_n9704;
  wire _abc_17692_n9705;
  wire _abc_17692_n9706;
  wire _abc_17692_n9707;
  wire _abc_17692_n9708;
  wire _abc_17692_n9709;
  wire _abc_17692_n971;
  wire _abc_17692_n9710;
  wire _abc_17692_n9711;
  wire _abc_17692_n9712;
  wire _abc_17692_n9713;
  wire _abc_17692_n9715;
  wire _abc_17692_n9716;
  wire _abc_17692_n9717;
  wire _abc_17692_n9718;
  wire _abc_17692_n9719;
  wire _abc_17692_n9720;
  wire _abc_17692_n9721;
  wire _abc_17692_n9722;
  wire _abc_17692_n9723;
  wire _abc_17692_n9724;
  wire _abc_17692_n9725;
  wire _abc_17692_n9726;
  wire _abc_17692_n9727;
  wire _abc_17692_n9728;
  wire _abc_17692_n9729;
  wire _abc_17692_n972_1;
  wire _abc_17692_n973;
  wire _abc_17692_n9730;
  wire _abc_17692_n9731;
  wire _abc_17692_n9732;
  wire _abc_17692_n9733;
  wire _abc_17692_n9734;
  wire _abc_17692_n9735;
  wire _abc_17692_n9736;
  wire _abc_17692_n9737;
  wire _abc_17692_n9738;
  wire _abc_17692_n9739;
  wire _abc_17692_n974;
  wire _abc_17692_n9740;
  wire _abc_17692_n9741;
  wire _abc_17692_n9742;
  wire _abc_17692_n9743;
  wire _abc_17692_n9744;
  wire _abc_17692_n9745;
  wire _abc_17692_n9746;
  wire _abc_17692_n9747;
  wire _abc_17692_n9748;
  wire _abc_17692_n9749;
  wire _abc_17692_n975;
  wire _abc_17692_n9750;
  wire _abc_17692_n9751;
  wire _abc_17692_n9752;
  wire _abc_17692_n9753;
  wire _abc_17692_n9754;
  wire _abc_17692_n9755;
  wire _abc_17692_n9756;
  wire _abc_17692_n9757;
  wire _abc_17692_n9758;
  wire _abc_17692_n9759;
  wire _abc_17692_n976;
  wire _abc_17692_n9760;
  wire _abc_17692_n9761;
  wire _abc_17692_n9762;
  wire _abc_17692_n9763;
  wire _abc_17692_n9764;
  wire _abc_17692_n9765;
  wire _abc_17692_n9766;
  wire _abc_17692_n9767;
  wire _abc_17692_n9768;
  wire _abc_17692_n9769;
  wire _abc_17692_n977;
  wire _abc_17692_n9770;
  wire _abc_17692_n9771;
  wire _abc_17692_n9772;
  wire _abc_17692_n9773;
  wire _abc_17692_n9774;
  wire _abc_17692_n9775;
  wire _abc_17692_n9776;
  wire _abc_17692_n9777;
  wire _abc_17692_n9778;
  wire _abc_17692_n9779;
  wire _abc_17692_n978;
  wire _abc_17692_n9780;
  wire _abc_17692_n9781;
  wire _abc_17692_n9782;
  wire _abc_17692_n9783;
  wire _abc_17692_n9784;
  wire _abc_17692_n9785;
  wire _abc_17692_n9786;
  wire _abc_17692_n9787;
  wire _abc_17692_n9788;
  wire _abc_17692_n9789;
  wire _abc_17692_n979;
  wire _abc_17692_n9790;
  wire _abc_17692_n9791;
  wire _abc_17692_n9792;
  wire _abc_17692_n9793;
  wire _abc_17692_n9794;
  wire _abc_17692_n9795;
  wire _abc_17692_n9796;
  wire _abc_17692_n9797;
  wire _abc_17692_n9798;
  wire _abc_17692_n9799;
  wire _abc_17692_n9800;
  wire _abc_17692_n9801;
  wire _abc_17692_n9802;
  wire _abc_17692_n9803;
  wire _abc_17692_n9804;
  wire _abc_17692_n9805;
  wire _abc_17692_n9806;
  wire _abc_17692_n9807;
  wire _abc_17692_n9808;
  wire _abc_17692_n9809;
  wire _abc_17692_n980_1;
  wire _abc_17692_n981;
  wire _abc_17692_n9810;
  wire _abc_17692_n9811;
  wire _abc_17692_n9812;
  wire _abc_17692_n9813;
  wire _abc_17692_n9814;
  wire _abc_17692_n9815;
  wire _abc_17692_n9816;
  wire _abc_17692_n9817;
  wire _abc_17692_n9818;
  wire _abc_17692_n9819;
  wire _abc_17692_n982;
  wire _abc_17692_n9820;
  wire _abc_17692_n9821;
  wire _abc_17692_n9822;
  wire _abc_17692_n9823;
  wire _abc_17692_n9824;
  wire _abc_17692_n9825;
  wire _abc_17692_n9826;
  wire _abc_17692_n9827;
  wire _abc_17692_n9828;
  wire _abc_17692_n9829;
  wire _abc_17692_n983;
  wire _abc_17692_n9830;
  wire _abc_17692_n9831;
  wire _abc_17692_n9832;
  wire _abc_17692_n9833;
  wire _abc_17692_n9834;
  wire _abc_17692_n9835;
  wire _abc_17692_n9836;
  wire _abc_17692_n9837;
  wire _abc_17692_n9838;
  wire _abc_17692_n9839;
  wire _abc_17692_n984;
  wire _abc_17692_n9840;
  wire _abc_17692_n9841;
  wire _abc_17692_n9842;
  wire _abc_17692_n9843;
  wire _abc_17692_n9844;
  wire _abc_17692_n9845;
  wire _abc_17692_n9846;
  wire _abc_17692_n9847;
  wire _abc_17692_n9848;
  wire _abc_17692_n9849;
  wire _abc_17692_n985;
  wire _abc_17692_n9851;
  wire _abc_17692_n9852;
  wire _abc_17692_n9853;
  wire _abc_17692_n9854;
  wire _abc_17692_n9855;
  wire _abc_17692_n9856;
  wire _abc_17692_n9857;
  wire _abc_17692_n9858;
  wire _abc_17692_n9859;
  wire _abc_17692_n986;
  wire _abc_17692_n9860;
  wire _abc_17692_n9861;
  wire _abc_17692_n9862;
  wire _abc_17692_n9863;
  wire _abc_17692_n9864;
  wire _abc_17692_n9865;
  wire _abc_17692_n9866;
  wire _abc_17692_n9867;
  wire _abc_17692_n9868;
  wire _abc_17692_n9869;
  wire _abc_17692_n987;
  wire _abc_17692_n9870;
  wire _abc_17692_n9871;
  wire _abc_17692_n9872;
  wire _abc_17692_n9873;
  wire _abc_17692_n9874;
  wire _abc_17692_n9875;
  wire _abc_17692_n9876;
  wire _abc_17692_n9877;
  wire _abc_17692_n9878;
  wire _abc_17692_n9879;
  wire _abc_17692_n9880;
  wire _abc_17692_n9881;
  wire _abc_17692_n9882;
  wire _abc_17692_n9883;
  wire _abc_17692_n9884;
  wire _abc_17692_n9885;
  wire _abc_17692_n9886;
  wire _abc_17692_n9887;
  wire _abc_17692_n9888;
  wire _abc_17692_n9889;
  wire _abc_17692_n988_1;
  wire _abc_17692_n989;
  wire _abc_17692_n9890;
  wire _abc_17692_n9891;
  wire _abc_17692_n9892;
  wire _abc_17692_n9893;
  wire _abc_17692_n9894;
  wire _abc_17692_n9895;
  wire _abc_17692_n9896;
  wire _abc_17692_n9897;
  wire _abc_17692_n9898;
  wire _abc_17692_n9899;
  wire _abc_17692_n990;
  wire _abc_17692_n9900;
  wire _abc_17692_n9901;
  wire _abc_17692_n9902;
  wire _abc_17692_n9903;
  wire _abc_17692_n9904;
  wire _abc_17692_n9905;
  wire _abc_17692_n9906;
  wire _abc_17692_n9907;
  wire _abc_17692_n9908;
  wire _abc_17692_n9909;
  wire _abc_17692_n991;
  wire _abc_17692_n9910;
  wire _abc_17692_n9911;
  wire _abc_17692_n9912;
  wire _abc_17692_n9913;
  wire _abc_17692_n9914;
  wire _abc_17692_n9915;
  wire _abc_17692_n9916;
  wire _abc_17692_n9917;
  wire _abc_17692_n9918;
  wire _abc_17692_n9919;
  wire _abc_17692_n992;
  wire _abc_17692_n9920;
  wire _abc_17692_n9921;
  wire _abc_17692_n9922;
  wire _abc_17692_n9923;
  wire _abc_17692_n9924;
  wire _abc_17692_n9925;
  wire _abc_17692_n9926;
  wire _abc_17692_n9927;
  wire _abc_17692_n9928;
  wire _abc_17692_n9929;
  wire _abc_17692_n993;
  wire _abc_17692_n9930;
  wire _abc_17692_n9931;
  wire _abc_17692_n9932;
  wire _abc_17692_n9933;
  wire _abc_17692_n9934;
  wire _abc_17692_n9935;
  wire _abc_17692_n9936;
  wire _abc_17692_n9937;
  wire _abc_17692_n9938;
  wire _abc_17692_n9939;
  wire _abc_17692_n9940;
  wire _abc_17692_n9941;
  wire _abc_17692_n9942;
  wire _abc_17692_n9943;
  wire _abc_17692_n9944;
  wire _abc_17692_n9945;
  wire _abc_17692_n9946;
  wire _abc_17692_n9947;
  wire _abc_17692_n9948;
  wire _abc_17692_n9949;
  wire _abc_17692_n995;
  wire _abc_17692_n9950;
  wire _abc_17692_n9951;
  wire _abc_17692_n9952;
  wire _abc_17692_n9953;
  wire _abc_17692_n9954;
  wire _abc_17692_n9955;
  wire _abc_17692_n9956;
  wire _abc_17692_n9957;
  wire _abc_17692_n9958;
  wire _abc_17692_n9959;
  wire _abc_17692_n9960;
  wire _abc_17692_n9961;
  wire _abc_17692_n9962;
  wire _abc_17692_n9963;
  wire _abc_17692_n9964;
  wire _abc_17692_n9965;
  wire _abc_17692_n9966;
  wire _abc_17692_n9967;
  wire _abc_17692_n9968;
  wire _abc_17692_n9969;
  wire _abc_17692_n996_1;
  wire _abc_17692_n997;
  wire _abc_17692_n9970;
  wire _abc_17692_n9971;
  wire _abc_17692_n9972;
  wire _abc_17692_n9973;
  wire _abc_17692_n9974;
  wire _abc_17692_n9975;
  wire _abc_17692_n9976;
  wire _abc_17692_n9977;
  wire _abc_17692_n9978;
  wire _abc_17692_n9979;
  wire _abc_17692_n998;
  wire _abc_17692_n9980;
  wire _abc_17692_n9981;
  wire _abc_17692_n9982;
  wire _abc_17692_n9983;
  wire _abc_17692_n9984;
  wire _abc_17692_n9985;
  wire _abc_17692_n9986;
  wire _abc_17692_n9987;
  wire _abc_17692_n9988;
  wire _abc_17692_n9989;
  wire _abc_17692_n999;
  wire _abc_17692_n9990;
  wire _abc_17692_n9991;
  wire _abc_17692_n9992;
  wire _abc_17692_n9993;
  wire _abc_17692_n9994;
  wire _abc_17692_n9995;
  wire _abc_17692_n9996;
  wire _abc_17692_n9997;
  wire _abc_17692_n9998;
  wire _abc_17692_n9999;
  wire _auto_iopadmap_cc_313_execute_30032_0_;
  wire _auto_iopadmap_cc_313_execute_30032_10_;
  wire _auto_iopadmap_cc_313_execute_30032_11_;
  wire _auto_iopadmap_cc_313_execute_30032_12_;
  wire _auto_iopadmap_cc_313_execute_30032_13_;
  wire _auto_iopadmap_cc_313_execute_30032_14_;
  wire _auto_iopadmap_cc_313_execute_30032_15_;
  wire _auto_iopadmap_cc_313_execute_30032_16_;
  wire _auto_iopadmap_cc_313_execute_30032_17_;
  wire _auto_iopadmap_cc_313_execute_30032_18_;
  wire _auto_iopadmap_cc_313_execute_30032_19_;
  wire _auto_iopadmap_cc_313_execute_30032_1_;
  wire _auto_iopadmap_cc_313_execute_30032_20_;
  wire _auto_iopadmap_cc_313_execute_30032_21_;
  wire _auto_iopadmap_cc_313_execute_30032_22_;
  wire _auto_iopadmap_cc_313_execute_30032_23_;
  wire _auto_iopadmap_cc_313_execute_30032_24_;
  wire _auto_iopadmap_cc_313_execute_30032_25_;
  wire _auto_iopadmap_cc_313_execute_30032_26_;
  wire _auto_iopadmap_cc_313_execute_30032_27_;
  wire _auto_iopadmap_cc_313_execute_30032_28_;
  wire _auto_iopadmap_cc_313_execute_30032_29_;
  wire _auto_iopadmap_cc_313_execute_30032_2_;
  wire _auto_iopadmap_cc_313_execute_30032_30_;
  wire _auto_iopadmap_cc_313_execute_30032_31_;
  wire _auto_iopadmap_cc_313_execute_30032_3_;
  wire _auto_iopadmap_cc_313_execute_30032_4_;
  wire _auto_iopadmap_cc_313_execute_30032_5_;
  wire _auto_iopadmap_cc_313_execute_30032_6_;
  wire _auto_iopadmap_cc_313_execute_30032_7_;
  wire _auto_iopadmap_cc_313_execute_30032_8_;
  wire _auto_iopadmap_cc_313_execute_30032_9_;
  wire _auto_iopadmap_cc_313_execute_30065_0_;
  wire _auto_iopadmap_cc_313_execute_30065_10_;
  wire _auto_iopadmap_cc_313_execute_30065_11_;
  wire _auto_iopadmap_cc_313_execute_30065_12_;
  wire _auto_iopadmap_cc_313_execute_30065_13_;
  wire _auto_iopadmap_cc_313_execute_30065_14_;
  wire _auto_iopadmap_cc_313_execute_30065_15_;
  wire _auto_iopadmap_cc_313_execute_30065_16_;
  wire _auto_iopadmap_cc_313_execute_30065_17_;
  wire _auto_iopadmap_cc_313_execute_30065_18_;
  wire _auto_iopadmap_cc_313_execute_30065_19_;
  wire _auto_iopadmap_cc_313_execute_30065_1_;
  wire _auto_iopadmap_cc_313_execute_30065_20_;
  wire _auto_iopadmap_cc_313_execute_30065_21_;
  wire _auto_iopadmap_cc_313_execute_30065_22_;
  wire _auto_iopadmap_cc_313_execute_30065_23_;
  wire _auto_iopadmap_cc_313_execute_30065_24_;
  wire _auto_iopadmap_cc_313_execute_30065_25_;
  wire _auto_iopadmap_cc_313_execute_30065_26_;
  wire _auto_iopadmap_cc_313_execute_30065_27_;
  wire _auto_iopadmap_cc_313_execute_30065_28_;
  wire _auto_iopadmap_cc_313_execute_30065_29_;
  wire _auto_iopadmap_cc_313_execute_30065_2_;
  wire _auto_iopadmap_cc_313_execute_30065_30_;
  wire _auto_iopadmap_cc_313_execute_30065_31_;
  wire _auto_iopadmap_cc_313_execute_30065_3_;
  wire _auto_iopadmap_cc_313_execute_30065_4_;
  wire _auto_iopadmap_cc_313_execute_30065_5_;
  wire _auto_iopadmap_cc_313_execute_30065_6_;
  wire _auto_iopadmap_cc_313_execute_30065_7_;
  wire _auto_iopadmap_cc_313_execute_30065_8_;
  wire _auto_iopadmap_cc_313_execute_30065_9_;
  output all_done;
  input clock;
  wire clock_bF_buf0;
  wire clock_bF_buf1;
  wire clock_bF_buf10;
  wire clock_bF_buf11;
  wire clock_bF_buf12;
  wire clock_bF_buf13;
  wire clock_bF_buf2;
  wire clock_bF_buf3;
  wire clock_bF_buf4;
  wire clock_bF_buf5;
  wire clock_bF_buf6;
  wire clock_bF_buf7;
  wire clock_bF_buf8;
  wire clock_bF_buf9;
  input \data_in1[0] ;
  input \data_in1[10] ;
  input \data_in1[11] ;
  input \data_in1[12] ;
  input \data_in1[13] ;
  input \data_in1[14] ;
  input \data_in1[15] ;
  input \data_in1[16] ;
  input \data_in1[17] ;
  input \data_in1[18] ;
  input \data_in1[19] ;
  input \data_in1[1] ;
  input \data_in1[20] ;
  input \data_in1[21] ;
  input \data_in1[22] ;
  input \data_in1[23] ;
  input \data_in1[24] ;
  input \data_in1[25] ;
  input \data_in1[26] ;
  input \data_in1[27] ;
  input \data_in1[28] ;
  input \data_in1[29] ;
  input \data_in1[2] ;
  input \data_in1[30] ;
  input \data_in1[31] ;
  input \data_in1[3] ;
  input \data_in1[4] ;
  input \data_in1[5] ;
  input \data_in1[6] ;
  input \data_in1[7] ;
  input \data_in1[8] ;
  input \data_in1[9] ;
  input \data_in2[0] ;
  input \data_in2[10] ;
  input \data_in2[11] ;
  input \data_in2[12] ;
  input \data_in2[13] ;
  input \data_in2[14] ;
  input \data_in2[15] ;
  input \data_in2[16] ;
  input \data_in2[17] ;
  input \data_in2[18] ;
  input \data_in2[19] ;
  input \data_in2[1] ;
  input \data_in2[20] ;
  input \data_in2[21] ;
  input \data_in2[22] ;
  input \data_in2[23] ;
  input \data_in2[24] ;
  input \data_in2[25] ;
  input \data_in2[26] ;
  input \data_in2[27] ;
  input \data_in2[28] ;
  input \data_in2[29] ;
  input \data_in2[2] ;
  input \data_in2[30] ;
  input \data_in2[31] ;
  input \data_in2[3] ;
  input \data_in2[4] ;
  input \data_in2[5] ;
  input \data_in2[6] ;
  input \data_in2[7] ;
  input \data_in2[8] ;
  input \data_in2[9] ;
  output \data_out1[0] ;
  output \data_out1[10] ;
  output \data_out1[11] ;
  output \data_out1[12] ;
  output \data_out1[13] ;
  output \data_out1[14] ;
  output \data_out1[15] ;
  output \data_out1[16] ;
  output \data_out1[17] ;
  output \data_out1[18] ;
  output \data_out1[19] ;
  output \data_out1[1] ;
  output \data_out1[20] ;
  output \data_out1[21] ;
  output \data_out1[22] ;
  output \data_out1[23] ;
  output \data_out1[24] ;
  output \data_out1[25] ;
  output \data_out1[26] ;
  output \data_out1[27] ;
  output \data_out1[28] ;
  output \data_out1[29] ;
  output \data_out1[2] ;
  output \data_out1[30] ;
  output \data_out1[31] ;
  output \data_out1[3] ;
  output \data_out1[4] ;
  output \data_out1[5] ;
  output \data_out1[6] ;
  output \data_out1[7] ;
  output \data_out1[8] ;
  output \data_out1[9] ;
  wire data_out1_0__FF_INPUT;
  wire data_out1_10__FF_INPUT;
  wire data_out1_11__FF_INPUT;
  wire data_out1_12__FF_INPUT;
  wire data_out1_13__FF_INPUT;
  wire data_out1_14__FF_INPUT;
  wire data_out1_15__FF_INPUT;
  wire data_out1_16__FF_INPUT;
  wire data_out1_17__FF_INPUT;
  wire data_out1_18__FF_INPUT;
  wire data_out1_19__FF_INPUT;
  wire data_out1_1__FF_INPUT;
  wire data_out1_20__FF_INPUT;
  wire data_out1_21__FF_INPUT;
  wire data_out1_22__FF_INPUT;
  wire data_out1_23__FF_INPUT;
  wire data_out1_24__FF_INPUT;
  wire data_out1_25__FF_INPUT;
  wire data_out1_26__FF_INPUT;
  wire data_out1_27__FF_INPUT;
  wire data_out1_28__FF_INPUT;
  wire data_out1_29__FF_INPUT;
  wire data_out1_2__FF_INPUT;
  wire data_out1_30__FF_INPUT;
  wire data_out1_31__FF_INPUT;
  wire data_out1_3__FF_INPUT;
  wire data_out1_4__FF_INPUT;
  wire data_out1_5__FF_INPUT;
  wire data_out1_6__FF_INPUT;
  wire data_out1_7__FF_INPUT;
  wire data_out1_8__FF_INPUT;
  wire data_out1_9__FF_INPUT;
  output \data_out2[0] ;
  output \data_out2[10] ;
  output \data_out2[11] ;
  output \data_out2[12] ;
  output \data_out2[13] ;
  output \data_out2[14] ;
  output \data_out2[15] ;
  output \data_out2[16] ;
  output \data_out2[17] ;
  output \data_out2[18] ;
  output \data_out2[19] ;
  output \data_out2[1] ;
  output \data_out2[20] ;
  output \data_out2[21] ;
  output \data_out2[22] ;
  output \data_out2[23] ;
  output \data_out2[24] ;
  output \data_out2[25] ;
  output \data_out2[26] ;
  output \data_out2[27] ;
  output \data_out2[28] ;
  output \data_out2[29] ;
  output \data_out2[2] ;
  output \data_out2[30] ;
  output \data_out2[31] ;
  output \data_out2[3] ;
  output \data_out2[4] ;
  output \data_out2[5] ;
  output \data_out2[6] ;
  output \data_out2[7] ;
  output \data_out2[8] ;
  output \data_out2[9] ;
  wire data_out2_0__FF_INPUT;
  wire data_out2_10__FF_INPUT;
  wire data_out2_11__FF_INPUT;
  wire data_out2_12__FF_INPUT;
  wire data_out2_13__FF_INPUT;
  wire data_out2_14__FF_INPUT;
  wire data_out2_15__FF_INPUT;
  wire data_out2_16__FF_INPUT;
  wire data_out2_17__FF_INPUT;
  wire data_out2_18__FF_INPUT;
  wire data_out2_19__FF_INPUT;
  wire data_out2_1__FF_INPUT;
  wire data_out2_20__FF_INPUT;
  wire data_out2_21__FF_INPUT;
  wire data_out2_22__FF_INPUT;
  wire data_out2_23__FF_INPUT;
  wire data_out2_24__FF_INPUT;
  wire data_out2_25__FF_INPUT;
  wire data_out2_26__FF_INPUT;
  wire data_out2_27__FF_INPUT;
  wire data_out2_28__FF_INPUT;
  wire data_out2_29__FF_INPUT;
  wire data_out2_2__FF_INPUT;
  wire data_out2_30__FF_INPUT;
  wire data_out2_31__FF_INPUT;
  wire data_out2_3__FF_INPUT;
  wire data_out2_4__FF_INPUT;
  wire data_out2_5__FF_INPUT;
  wire data_out2_6__FF_INPUT;
  wire data_out2_7__FF_INPUT;
  wire data_out2_8__FF_INPUT;
  wire data_out2_9__FF_INPUT;
  wire delta_0_;
  wire delta_0__FF_INPUT;
  wire delta_10_;
  wire delta_10__FF_INPUT;
  wire delta_11_;
  wire delta_11__FF_INPUT;
  wire delta_12_;
  wire delta_12__FF_INPUT;
  wire delta_13_;
  wire delta_13__FF_INPUT;
  wire delta_14_;
  wire delta_14__FF_INPUT;
  wire delta_15_;
  wire delta_15__FF_INPUT;
  wire delta_16_;
  wire delta_16__FF_INPUT;
  wire delta_17_;
  wire delta_17__FF_INPUT;
  wire delta_18_;
  wire delta_18__FF_INPUT;
  wire delta_19_;
  wire delta_19__FF_INPUT;
  wire delta_1_;
  wire delta_1__FF_INPUT;
  wire delta_20_;
  wire delta_20__FF_INPUT;
  wire delta_21_;
  wire delta_21__FF_INPUT;
  wire delta_22_;
  wire delta_22__FF_INPUT;
  wire delta_23_;
  wire delta_23__FF_INPUT;
  wire delta_24_;
  wire delta_24__FF_INPUT;
  wire delta_25_;
  wire delta_25__FF_INPUT;
  wire delta_26_;
  wire delta_26__FF_INPUT;
  wire delta_27_;
  wire delta_27__FF_INPUT;
  wire delta_28_;
  wire delta_28__FF_INPUT;
  wire delta_29_;
  wire delta_29__FF_INPUT;
  wire delta_2_;
  wire delta_2__FF_INPUT;
  wire delta_30_;
  wire delta_30__FF_INPUT;
  wire delta_31_;
  wire delta_31__FF_INPUT;
  wire delta_3_;
  wire delta_3__FF_INPUT;
  wire delta_4_;
  wire delta_4__FF_INPUT;
  wire delta_5_;
  wire delta_5__FF_INPUT;
  wire delta_6_;
  wire delta_6__FF_INPUT;
  wire delta_7_;
  wire delta_7__FF_INPUT;
  wire delta_8_;
  wire delta_8__FF_INPUT;
  wire delta_9_;
  wire delta_9__FF_INPUT;
  input \key_in[0] ;
  input \key_in[100] ;
  input \key_in[101] ;
  input \key_in[102] ;
  input \key_in[103] ;
  input \key_in[104] ;
  input \key_in[105] ;
  input \key_in[106] ;
  input \key_in[107] ;
  input \key_in[108] ;
  input \key_in[109] ;
  input \key_in[10] ;
  input \key_in[110] ;
  input \key_in[111] ;
  input \key_in[112] ;
  input \key_in[113] ;
  input \key_in[114] ;
  input \key_in[115] ;
  input \key_in[116] ;
  input \key_in[117] ;
  input \key_in[118] ;
  input \key_in[119] ;
  input \key_in[11] ;
  input \key_in[120] ;
  input \key_in[121] ;
  input \key_in[122] ;
  input \key_in[123] ;
  input \key_in[124] ;
  input \key_in[125] ;
  input \key_in[126] ;
  input \key_in[127] ;
  input \key_in[12] ;
  input \key_in[13] ;
  input \key_in[14] ;
  input \key_in[15] ;
  input \key_in[16] ;
  input \key_in[17] ;
  input \key_in[18] ;
  input \key_in[19] ;
  input \key_in[1] ;
  input \key_in[20] ;
  input \key_in[21] ;
  input \key_in[22] ;
  input \key_in[23] ;
  input \key_in[24] ;
  input \key_in[25] ;
  input \key_in[26] ;
  input \key_in[27] ;
  input \key_in[28] ;
  input \key_in[29] ;
  input \key_in[2] ;
  input \key_in[30] ;
  input \key_in[31] ;
  input \key_in[32] ;
  input \key_in[33] ;
  input \key_in[34] ;
  input \key_in[35] ;
  input \key_in[36] ;
  input \key_in[37] ;
  input \key_in[38] ;
  input \key_in[39] ;
  input \key_in[3] ;
  input \key_in[40] ;
  input \key_in[41] ;
  input \key_in[42] ;
  input \key_in[43] ;
  input \key_in[44] ;
  input \key_in[45] ;
  input \key_in[46] ;
  input \key_in[47] ;
  input \key_in[48] ;
  input \key_in[49] ;
  input \key_in[4] ;
  input \key_in[50] ;
  input \key_in[51] ;
  input \key_in[52] ;
  input \key_in[53] ;
  input \key_in[54] ;
  input \key_in[55] ;
  input \key_in[56] ;
  input \key_in[57] ;
  input \key_in[58] ;
  input \key_in[59] ;
  input \key_in[5] ;
  input \key_in[60] ;
  input \key_in[61] ;
  input \key_in[62] ;
  input \key_in[63] ;
  input \key_in[64] ;
  input \key_in[65] ;
  input \key_in[66] ;
  input \key_in[67] ;
  input \key_in[68] ;
  input \key_in[69] ;
  input \key_in[6] ;
  input \key_in[70] ;
  input \key_in[71] ;
  input \key_in[72] ;
  input \key_in[73] ;
  input \key_in[74] ;
  input \key_in[75] ;
  input \key_in[76] ;
  input \key_in[77] ;
  input \key_in[78] ;
  input \key_in[79] ;
  input \key_in[7] ;
  input \key_in[80] ;
  input \key_in[81] ;
  input \key_in[82] ;
  input \key_in[83] ;
  input \key_in[84] ;
  input \key_in[85] ;
  input \key_in[86] ;
  input \key_in[87] ;
  input \key_in[88] ;
  input \key_in[89] ;
  input \key_in[8] ;
  input \key_in[90] ;
  input \key_in[91] ;
  input \key_in[92] ;
  input \key_in[93] ;
  input \key_in[94] ;
  input \key_in[95] ;
  input \key_in[96] ;
  input \key_in[97] ;
  input \key_in[98] ;
  input \key_in[99] ;
  input \key_in[9] ;
  input mode;
  wire modereg;
  wire modereg_FF_INPUT;
  input reset;
  wire selectslice_0_;
  wire selectslice_0__FF_INPUT;
  wire selectslice_1_;
  wire selectslice_1__FF_INPUT;
  wire state_0_;
  wire state_10_;
  wire state_10_bF_buf0;
  wire state_10_bF_buf1;
  wire state_10_bF_buf2;
  wire state_10_bF_buf3;
  wire state_10_bF_buf4;
  wire state_11_;
  wire state_12_;
  wire state_13_;
  wire state_14_;
  wire state_14_bF_buf0;
  wire state_14_bF_buf1;
  wire state_14_bF_buf2;
  wire state_14_bF_buf3;
  wire state_14_bF_buf4;
  wire state_15_;
  wire state_15_bF_buf0;
  wire state_15_bF_buf1;
  wire state_15_bF_buf2;
  wire state_15_bF_buf3;
  wire state_15_bF_buf4;
  wire state_1_;
  wire state_2_;
  wire state_3_;
  wire state_3_bF_buf0;
  wire state_3_bF_buf1;
  wire state_3_bF_buf2;
  wire state_3_bF_buf3;
  wire state_3_bF_buf4;
  wire state_4_;
  wire state_5_;
  wire state_6_;
  wire state_6_bF_buf0;
  wire state_6_bF_buf1;
  wire state_6_bF_buf2;
  wire state_6_bF_buf3;
  wire state_6_bF_buf4;
  wire state_7_;
  wire state_7_bF_buf0;
  wire state_7_bF_buf1;
  wire state_7_bF_buf2;
  wire state_7_bF_buf3;
  wire state_7_bF_buf4;
  wire state_8_;
  wire state_8_bF_buf0;
  wire state_8_bF_buf1;
  wire state_8_bF_buf2;
  wire state_8_bF_buf3;
  wire state_8_bF_buf4;
  wire state_8_bF_buf5;
  wire state_8_bF_buf6;
  wire state_8_bF_buf7;
  wire state_8_bF_buf8;
  wire state_8_bF_buf9;
  wire sum_0_;
  wire sum_0__FF_INPUT;
  wire sum_10_;
  wire sum_10__FF_INPUT;
  wire sum_11_;
  wire sum_11__FF_INPUT;
  wire sum_12_;
  wire sum_12__FF_INPUT;
  wire sum_13_;
  wire sum_13__FF_INPUT;
  wire sum_14_;
  wire sum_14__FF_INPUT;
  wire sum_15_;
  wire sum_15__FF_INPUT;
  wire sum_16_;
  wire sum_16__FF_INPUT;
  wire sum_17_;
  wire sum_17__FF_INPUT;
  wire sum_18_;
  wire sum_18__FF_INPUT;
  wire sum_19_;
  wire sum_19__FF_INPUT;
  wire sum_1_;
  wire sum_1__FF_INPUT;
  wire sum_20_;
  wire sum_20__FF_INPUT;
  wire sum_21_;
  wire sum_21__FF_INPUT;
  wire sum_22_;
  wire sum_22__FF_INPUT;
  wire sum_23_;
  wire sum_23__FF_INPUT;
  wire sum_24_;
  wire sum_24__FF_INPUT;
  wire sum_25_;
  wire sum_25__FF_INPUT;
  wire sum_26_;
  wire sum_26__FF_INPUT;
  wire sum_27_;
  wire sum_27__FF_INPUT;
  wire sum_28_;
  wire sum_28__FF_INPUT;
  wire sum_29_;
  wire sum_29__FF_INPUT;
  wire sum_2_;
  wire sum_2__FF_INPUT;
  wire sum_30_;
  wire sum_30__FF_INPUT;
  wire sum_31_;
  wire sum_31__FF_INPUT;
  wire sum_3_;
  wire sum_3__FF_INPUT;
  wire sum_4_;
  wire sum_4__FF_INPUT;
  wire sum_5_;
  wire sum_5__FF_INPUT;
  wire sum_6_;
  wire sum_6__FF_INPUT;
  wire sum_7_;
  wire sum_7__FF_INPUT;
  wire sum_8_;
  wire sum_8__FF_INPUT;
  wire sum_9_;
  wire sum_9__FF_INPUT;
  wire while_flag;
  wire while_flag_FF_INPUT;
  wire workunit1_0_;
  wire workunit1_0__FF_INPUT;
  wire workunit1_10_;
  wire workunit1_10__FF_INPUT;
  wire workunit1_11_;
  wire workunit1_11__FF_INPUT;
  wire workunit1_11_bF_buf0;
  wire workunit1_11_bF_buf1;
  wire workunit1_11_bF_buf2;
  wire workunit1_11_bF_buf3;
  wire workunit1_12_;
  wire workunit1_12__FF_INPUT;
  wire workunit1_12_bF_buf0;
  wire workunit1_12_bF_buf1;
  wire workunit1_12_bF_buf2;
  wire workunit1_12_bF_buf3;
  wire workunit1_13_;
  wire workunit1_13__FF_INPUT;
  wire workunit1_13_bF_buf0;
  wire workunit1_13_bF_buf1;
  wire workunit1_13_bF_buf2;
  wire workunit1_13_bF_buf3;
  wire workunit1_14_;
  wire workunit1_14__FF_INPUT;
  wire workunit1_14_bF_buf0;
  wire workunit1_14_bF_buf1;
  wire workunit1_14_bF_buf2;
  wire workunit1_14_bF_buf3;
  wire workunit1_15_;
  wire workunit1_15__FF_INPUT;
  wire workunit1_16_;
  wire workunit1_16__FF_INPUT;
  wire workunit1_16_bF_buf0;
  wire workunit1_16_bF_buf1;
  wire workunit1_16_bF_buf2;
  wire workunit1_16_bF_buf3;
  wire workunit1_17_;
  wire workunit1_17__FF_INPUT;
  wire workunit1_18_;
  wire workunit1_18__FF_INPUT;
  wire workunit1_19_;
  wire workunit1_19__FF_INPUT;
  wire workunit1_1_;
  wire workunit1_1__FF_INPUT;
  wire workunit1_1_bF_buf0;
  wire workunit1_1_bF_buf1;
  wire workunit1_1_bF_buf2;
  wire workunit1_1_bF_buf3;
  wire workunit1_20_;
  wire workunit1_20__FF_INPUT;
  wire workunit1_21_;
  wire workunit1_21__FF_INPUT;
  wire workunit1_22_;
  wire workunit1_22__FF_INPUT;
  wire workunit1_23_;
  wire workunit1_23__FF_INPUT;
  wire workunit1_24_;
  wire workunit1_24__FF_INPUT;
  wire workunit1_25_;
  wire workunit1_25__FF_INPUT;
  wire workunit1_26_;
  wire workunit1_26__FF_INPUT;
  wire workunit1_27_;
  wire workunit1_27__FF_INPUT;
  wire workunit1_28_;
  wire workunit1_28__FF_INPUT;
  wire workunit1_29_;
  wire workunit1_29__FF_INPUT;
  wire workunit1_2_;
  wire workunit1_2__FF_INPUT;
  wire workunit1_30_;
  wire workunit1_30__FF_INPUT;
  wire workunit1_31_;
  wire workunit1_31__FF_INPUT;
  wire workunit1_3_;
  wire workunit1_3__FF_INPUT;
  wire workunit1_4_;
  wire workunit1_4__FF_INPUT;
  wire workunit1_5_;
  wire workunit1_5__FF_INPUT;
  wire workunit1_6_;
  wire workunit1_6__FF_INPUT;
  wire workunit1_7_;
  wire workunit1_7__FF_INPUT;
  wire workunit1_8_;
  wire workunit1_8__FF_INPUT;
  wire workunit1_8_bF_buf0;
  wire workunit1_8_bF_buf1;
  wire workunit1_8_bF_buf2;
  wire workunit1_8_bF_buf3;
  wire workunit1_9_;
  wire workunit1_9__FF_INPUT;
  wire workunit2_0_;
  wire workunit2_0__FF_INPUT;
  wire workunit2_10_;
  wire workunit2_10__FF_INPUT;
  wire workunit2_10_bF_buf0;
  wire workunit2_10_bF_buf1;
  wire workunit2_10_bF_buf2;
  wire workunit2_10_bF_buf3;
  wire workunit2_11_;
  wire workunit2_11__FF_INPUT;
  wire workunit2_12_;
  wire workunit2_12__FF_INPUT;
  wire workunit2_12_bF_buf0;
  wire workunit2_12_bF_buf1;
  wire workunit2_12_bF_buf2;
  wire workunit2_12_bF_buf3;
  wire workunit2_13_;
  wire workunit2_13__FF_INPUT;
  wire workunit2_14_;
  wire workunit2_14__FF_INPUT;
  wire workunit2_14_bF_buf0;
  wire workunit2_14_bF_buf1;
  wire workunit2_14_bF_buf2;
  wire workunit2_14_bF_buf3;
  wire workunit2_15_;
  wire workunit2_15__FF_INPUT;
  wire workunit2_16_;
  wire workunit2_16__FF_INPUT;
  wire workunit2_16_bF_buf0;
  wire workunit2_16_bF_buf1;
  wire workunit2_16_bF_buf2;
  wire workunit2_16_bF_buf3;
  wire workunit2_17_;
  wire workunit2_17__FF_INPUT;
  wire workunit2_18_;
  wire workunit2_18__FF_INPUT;
  wire workunit2_19_;
  wire workunit2_19__FF_INPUT;
  wire workunit2_1_;
  wire workunit2_1__FF_INPUT;
  wire workunit2_1_bF_buf0;
  wire workunit2_1_bF_buf1;
  wire workunit2_1_bF_buf2;
  wire workunit2_1_bF_buf3;
  wire workunit2_20_;
  wire workunit2_20__FF_INPUT;
  wire workunit2_21_;
  wire workunit2_21__FF_INPUT;
  wire workunit2_22_;
  wire workunit2_22__FF_INPUT;
  wire workunit2_23_;
  wire workunit2_23__FF_INPUT;
  wire workunit2_24_;
  wire workunit2_24__FF_INPUT;
  wire workunit2_25_;
  wire workunit2_25__FF_INPUT;
  wire workunit2_26_;
  wire workunit2_26__FF_INPUT;
  wire workunit2_27_;
  wire workunit2_27__FF_INPUT;
  wire workunit2_28_;
  wire workunit2_28__FF_INPUT;
  wire workunit2_29_;
  wire workunit2_29__FF_INPUT;
  wire workunit2_2_;
  wire workunit2_2__FF_INPUT;
  wire workunit2_30_;
  wire workunit2_30__FF_INPUT;
  wire workunit2_31_;
  wire workunit2_31__FF_INPUT;
  wire workunit2_3_;
  wire workunit2_3__FF_INPUT;
  wire workunit2_4_;
  wire workunit2_4__FF_INPUT;
  wire workunit2_5_;
  wire workunit2_5__FF_INPUT;
  wire workunit2_6_;
  wire workunit2_6__FF_INPUT;
  wire workunit2_7_;
  wire workunit2_7__FF_INPUT;
  wire workunit2_8_;
  wire workunit2_8__FF_INPUT;
  wire workunit2_8_bF_buf0;
  wire workunit2_8_bF_buf1;
  wire workunit2_8_bF_buf2;
  wire workunit2_8_bF_buf3;
  wire workunit2_9_;
  wire workunit2_9__FF_INPUT;
  wire x_0_;
  wire x_0__FF_INPUT;
  wire x_1_;
  wire x_1__FF_INPUT;
  wire x_2_;
  wire x_2__FF_INPUT;
  wire x_3_;
  wire x_3__FF_INPUT;
  wire x_4_;
  wire x_4__FF_INPUT;
  wire x_5_;
  wire x_5__FF_INPUT;
  wire x_6_;
  wire x_6__FF_INPUT;
  wire x_7_;
  wire x_7__FF_INPUT;
  AND2X2 AND2X2_1 ( .A(_abc_17692_n623), .B(state_13_), .Y(_abc_17692_n624) );
  AND2X2 AND2X2_10 ( .A(_abc_17692_n632), .B(delta_19_), .Y(delta_19__FF_INPUT) );
  AND2X2 AND2X2_100 ( .A(_abc_17692_n905), .B(_abc_17692_n904), .Y(data_out1_27__FF_INPUT) );
  AND2X2 AND2X2_1000 ( .A(_abc_17692_n2969), .B(_abc_17692_n2967), .Y(_abc_17692_n2970) );
  AND2X2 AND2X2_1001 ( .A(_abc_17692_n2766), .B(_abc_17692_n2767), .Y(_abc_17692_n2971) );
  AND2X2 AND2X2_1002 ( .A(_abc_17692_n2975), .B(_abc_17692_n1863_bF_buf10), .Y(_abc_17692_n2976) );
  AND2X2 AND2X2_1003 ( .A(_abc_17692_n2976), .B(_abc_17692_n2973), .Y(_abc_17692_n2977) );
  AND2X2 AND2X2_1004 ( .A(_abc_17692_n2978), .B(state_6_bF_buf3), .Y(_abc_17692_n2979) );
  AND2X2 AND2X2_1005 ( .A(_abc_17692_n2982), .B(_abc_17692_n2896), .Y(_abc_17692_n2983) );
  AND2X2 AND2X2_1006 ( .A(_abc_17692_n2985), .B(_abc_17692_n1830_bF_buf9), .Y(_abc_17692_n2986) );
  AND2X2 AND2X2_1007 ( .A(_abc_17692_n2986), .B(_abc_17692_n2984), .Y(_abc_17692_n2987) );
  AND2X2 AND2X2_1008 ( .A(_abc_17692_n2804), .B(_abc_17692_n2732), .Y(_abc_17692_n2989) );
  AND2X2 AND2X2_1009 ( .A(_abc_17692_n2990), .B(_abc_17692_n2931), .Y(_abc_17692_n2992) );
  AND2X2 AND2X2_101 ( .A(_abc_17692_n908), .B(_abc_17692_n907), .Y(data_out1_28__FF_INPUT) );
  AND2X2 AND2X2_1010 ( .A(_abc_17692_n2993), .B(_abc_17692_n1846_bF_buf9), .Y(_abc_17692_n2994) );
  AND2X2 AND2X2_1011 ( .A(_abc_17692_n2994), .B(_abc_17692_n2991), .Y(_abc_17692_n2995_1) );
  AND2X2 AND2X2_1012 ( .A(_abc_17692_n2793), .B(_abc_17692_n2759), .Y(_abc_17692_n2997) );
  AND2X2 AND2X2_1013 ( .A(_abc_17692_n2796), .B(_abc_17692_n2764), .Y(_abc_17692_n3000) );
  AND2X2 AND2X2_1014 ( .A(_abc_17692_n3002), .B(_abc_17692_n1863_bF_buf9), .Y(_abc_17692_n3003) );
  AND2X2 AND2X2_1015 ( .A(_abc_17692_n3003), .B(_abc_17692_n2998_1), .Y(_abc_17692_n3004) );
  AND2X2 AND2X2_1016 ( .A(_abc_17692_n2782), .B(_abc_17692_n3005), .Y(_abc_17692_n3006) );
  AND2X2 AND2X2_1017 ( .A(_abc_17692_n2779), .B(_abc_17692_n2776), .Y(_abc_17692_n3010) );
  AND2X2 AND2X2_1018 ( .A(_abc_17692_n3012), .B(_abc_17692_n1877_bF_buf9), .Y(_abc_17692_n3013) );
  AND2X2 AND2X2_1019 ( .A(_abc_17692_n3013), .B(_abc_17692_n3007), .Y(_abc_17692_n3014) );
  AND2X2 AND2X2_102 ( .A(_abc_17692_n911_1), .B(_abc_17692_n910_1), .Y(data_out1_29__FF_INPUT) );
  AND2X2 AND2X2_1020 ( .A(_abc_17692_n3016), .B(state_7_bF_buf2), .Y(_abc_17692_n3017) );
  AND2X2 AND2X2_1021 ( .A(_abc_17692_n1885_bF_buf3), .B(workunit2_6_), .Y(_abc_17692_n3018) );
  AND2X2 AND2X2_1022 ( .A(state_8_bF_buf3), .B(\data_in2[6] ), .Y(_abc_17692_n3019) );
  AND2X2 AND2X2_1023 ( .A(_abc_17692_n3023), .B(_abc_17692_n2826), .Y(_abc_17692_n3024) );
  AND2X2 AND2X2_1024 ( .A(workunit1_3_), .B(workunit1_12_bF_buf2), .Y(_abc_17692_n3025) );
  AND2X2 AND2X2_1025 ( .A(_abc_17692_n2249), .B(_abc_17692_n3026), .Y(_abc_17692_n3027) );
  AND2X2 AND2X2_1026 ( .A(_abc_17692_n3030), .B(_abc_17692_n3031), .Y(_abc_17692_n3032) );
  AND2X2 AND2X2_1027 ( .A(_abc_17692_n3029), .B(_abc_17692_n3033), .Y(_abc_17692_n3034_1) );
  AND2X2 AND2X2_1028 ( .A(_abc_17692_n3024), .B(_abc_17692_n3034_1), .Y(_abc_17692_n3035) );
  AND2X2 AND2X2_1029 ( .A(_abc_17692_n3032), .B(workunit1_7_), .Y(_abc_17692_n3037) );
  AND2X2 AND2X2_103 ( .A(_abc_17692_n914), .B(_abc_17692_n913), .Y(data_out1_30__FF_INPUT) );
  AND2X2 AND2X2_1030 ( .A(_abc_17692_n3028), .B(_abc_17692_n2063), .Y(_abc_17692_n3038) );
  AND2X2 AND2X2_1031 ( .A(_abc_17692_n3036), .B(_abc_17692_n3039), .Y(_abc_17692_n3040) );
  AND2X2 AND2X2_1032 ( .A(sum_7_), .B(\key_in[7] ), .Y(_abc_17692_n3044) );
  AND2X2 AND2X2_1033 ( .A(_abc_17692_n3045), .B(_abc_17692_n3046), .Y(_abc_17692_n3047) );
  AND2X2 AND2X2_1034 ( .A(_abc_17692_n3043), .B(_abc_17692_n3047), .Y(_abc_17692_n3048) );
  AND2X2 AND2X2_1035 ( .A(_abc_17692_n3042), .B(_abc_17692_n3049), .Y(_abc_17692_n3050) );
  AND2X2 AND2X2_1036 ( .A(_abc_17692_n3051), .B(_abc_17692_n3041), .Y(_abc_17692_n3052) );
  AND2X2 AND2X2_1037 ( .A(_abc_17692_n3054), .B(_abc_17692_n3053), .Y(_abc_17692_n3055) );
  AND2X2 AND2X2_1038 ( .A(_abc_17692_n3056), .B(_abc_17692_n3055), .Y(_abc_17692_n3057) );
  AND2X2 AND2X2_1039 ( .A(_abc_17692_n3058_1), .B(workunit2_7_), .Y(_abc_17692_n3059) );
  AND2X2 AND2X2_104 ( .A(_abc_17692_n917), .B(_abc_17692_n916), .Y(data_out1_31__FF_INPUT) );
  AND2X2 AND2X2_1040 ( .A(_abc_17692_n3061), .B(_abc_17692_n3060), .Y(_abc_17692_n3062) );
  AND2X2 AND2X2_1041 ( .A(_abc_17692_n2898), .B(_abc_17692_n3065), .Y(_abc_17692_n3066) );
  AND2X2 AND2X2_1042 ( .A(_abc_17692_n3069), .B(_abc_17692_n1830_bF_buf8), .Y(_abc_17692_n3070) );
  AND2X2 AND2X2_1043 ( .A(_abc_17692_n3070), .B(_abc_17692_n3068), .Y(_abc_17692_n3071) );
  AND2X2 AND2X2_1044 ( .A(sum_7_), .B(\key_in[71] ), .Y(_abc_17692_n3073) );
  AND2X2 AND2X2_1045 ( .A(_abc_17692_n3074), .B(_abc_17692_n3075), .Y(_abc_17692_n3076) );
  AND2X2 AND2X2_1046 ( .A(_abc_17692_n3072), .B(_abc_17692_n3077), .Y(_abc_17692_n3079) );
  AND2X2 AND2X2_1047 ( .A(_abc_17692_n3080_1), .B(_abc_17692_n3078), .Y(_abc_17692_n3081) );
  AND2X2 AND2X2_1048 ( .A(_abc_17692_n3082), .B(_abc_17692_n3041), .Y(_abc_17692_n3083) );
  AND2X2 AND2X2_1049 ( .A(_abc_17692_n3081), .B(_abc_17692_n3055), .Y(_abc_17692_n3084) );
  AND2X2 AND2X2_105 ( .A(_abc_17692_n723), .B(sum_0_), .Y(_abc_17692_n919) );
  AND2X2 AND2X2_1050 ( .A(_abc_17692_n3087), .B(_abc_17692_n3088), .Y(_abc_17692_n3089) );
  AND2X2 AND2X2_1051 ( .A(_abc_17692_n2863), .B(workunit2_6_), .Y(_abc_17692_n3091) );
  AND2X2 AND2X2_1052 ( .A(_abc_17692_n3095), .B(_abc_17692_n1877_bF_buf8), .Y(_abc_17692_n3096) );
  AND2X2 AND2X2_1053 ( .A(_abc_17692_n3096), .B(_abc_17692_n3094), .Y(_abc_17692_n3097) );
  AND2X2 AND2X2_1054 ( .A(_abc_17692_n3098), .B(_abc_17692_n2913), .Y(_abc_17692_n3099) );
  AND2X2 AND2X2_1055 ( .A(sum_7_), .B(\key_in[39] ), .Y(_abc_17692_n3100) );
  AND2X2 AND2X2_1056 ( .A(_abc_17692_n3101), .B(_abc_17692_n3102), .Y(_abc_17692_n3103) );
  AND2X2 AND2X2_1057 ( .A(_abc_17692_n3099), .B(_abc_17692_n3103), .Y(_abc_17692_n3104) );
  AND2X2 AND2X2_1058 ( .A(_abc_17692_n3105), .B(_abc_17692_n3106), .Y(_abc_17692_n3107) );
  AND2X2 AND2X2_1059 ( .A(_abc_17692_n3111), .B(_abc_17692_n3110), .Y(_abc_17692_n3112) );
  AND2X2 AND2X2_106 ( .A(delta_0_), .B(sum_0_), .Y(_abc_17692_n921) );
  AND2X2 AND2X2_1060 ( .A(_abc_17692_n3109), .B(_abc_17692_n3113), .Y(_abc_17692_n3114) );
  AND2X2 AND2X2_1061 ( .A(_abc_17692_n3114), .B(workunit2_7_), .Y(_abc_17692_n3115) );
  AND2X2 AND2X2_1062 ( .A(_abc_17692_n3116), .B(_abc_17692_n3117), .Y(_abc_17692_n3118) );
  AND2X2 AND2X2_1063 ( .A(_abc_17692_n3118), .B(_abc_17692_n3060), .Y(_abc_17692_n3119) );
  AND2X2 AND2X2_1064 ( .A(_abc_17692_n2928), .B(workunit2_6_), .Y(_abc_17692_n3122) );
  AND2X2 AND2X2_1065 ( .A(_abc_17692_n2944), .B(_abc_17692_n3123), .Y(_abc_17692_n3124) );
  AND2X2 AND2X2_1066 ( .A(_abc_17692_n3127), .B(_abc_17692_n1846_bF_buf8), .Y(_abc_17692_n3128) );
  AND2X2 AND2X2_1067 ( .A(_abc_17692_n3128), .B(_abc_17692_n3126), .Y(_abc_17692_n3129) );
  AND2X2 AND2X2_1068 ( .A(sum_7_), .B(\key_in[103] ), .Y(_abc_17692_n3133) );
  AND2X2 AND2X2_1069 ( .A(_abc_17692_n3134), .B(_abc_17692_n3135), .Y(_abc_17692_n3136) );
  AND2X2 AND2X2_107 ( .A(_abc_17692_n922), .B(_abc_17692_n920), .Y(_abc_17692_n923_1) );
  AND2X2 AND2X2_1070 ( .A(_abc_17692_n3132), .B(_abc_17692_n3137), .Y(_abc_17692_n3139) );
  AND2X2 AND2X2_1071 ( .A(_abc_17692_n3140), .B(_abc_17692_n3138), .Y(_abc_17692_n3141_1) );
  AND2X2 AND2X2_1072 ( .A(_abc_17692_n3142), .B(_abc_17692_n3041), .Y(_abc_17692_n3143) );
  AND2X2 AND2X2_1073 ( .A(_abc_17692_n3141_1), .B(_abc_17692_n3055), .Y(_abc_17692_n3144_1) );
  AND2X2 AND2X2_1074 ( .A(_abc_17692_n3147), .B(_abc_17692_n3148), .Y(_abc_17692_n3149) );
  AND2X2 AND2X2_1075 ( .A(_abc_17692_n2975), .B(_abc_17692_n2967), .Y(_abc_17692_n3150) );
  AND2X2 AND2X2_1076 ( .A(_abc_17692_n3154), .B(_abc_17692_n1863_bF_buf8), .Y(_abc_17692_n3155) );
  AND2X2 AND2X2_1077 ( .A(_abc_17692_n3155), .B(_abc_17692_n3152), .Y(_abc_17692_n3156) );
  AND2X2 AND2X2_1078 ( .A(_abc_17692_n3157), .B(state_6_bF_buf2), .Y(_abc_17692_n3158) );
  AND2X2 AND2X2_1079 ( .A(_abc_17692_n2984), .B(_abc_17692_n2894), .Y(_abc_17692_n3159) );
  AND2X2 AND2X2_108 ( .A(_abc_17692_n923_1), .B(_abc_17692_n721), .Y(_abc_17692_n924) );
  AND2X2 AND2X2_1080 ( .A(_abc_17692_n3162), .B(_abc_17692_n1830_bF_buf7), .Y(_abc_17692_n3163) );
  AND2X2 AND2X2_1081 ( .A(_abc_17692_n3163), .B(_abc_17692_n3160), .Y(_abc_17692_n3164) );
  AND2X2 AND2X2_1082 ( .A(_abc_17692_n2993), .B(_abc_17692_n2929), .Y(_abc_17692_n3165) );
  AND2X2 AND2X2_1083 ( .A(_abc_17692_n3168), .B(_abc_17692_n1846_bF_buf7), .Y(_abc_17692_n3169) );
  AND2X2 AND2X2_1084 ( .A(_abc_17692_n3169), .B(_abc_17692_n3167), .Y(_abc_17692_n3170) );
  AND2X2 AND2X2_1085 ( .A(_abc_17692_n3001), .B(_abc_17692_n2974), .Y(_abc_17692_n3174) );
  AND2X2 AND2X2_1086 ( .A(_abc_17692_n2998_1), .B(_abc_17692_n3172), .Y(_abc_17692_n3177) );
  AND2X2 AND2X2_1087 ( .A(_abc_17692_n3178_1), .B(_abc_17692_n1863_bF_buf7), .Y(_abc_17692_n3179) );
  AND2X2 AND2X2_1088 ( .A(_abc_17692_n3179), .B(_abc_17692_n3176), .Y(_abc_17692_n3180) );
  AND2X2 AND2X2_1089 ( .A(_abc_17692_n3011), .B(_abc_17692_n3008), .Y(_abc_17692_n3181) );
  AND2X2 AND2X2_109 ( .A(_abc_17692_n926_1), .B(sum_1_), .Y(_abc_17692_n928) );
  AND2X2 AND2X2_1090 ( .A(_abc_17692_n3185), .B(_abc_17692_n1877_bF_buf7), .Y(_abc_17692_n3186) );
  AND2X2 AND2X2_1091 ( .A(_abc_17692_n3187), .B(_abc_17692_n3186), .Y(_abc_17692_n3188) );
  AND2X2 AND2X2_1092 ( .A(_abc_17692_n3188), .B(_abc_17692_n3183), .Y(_abc_17692_n3189_1) );
  AND2X2 AND2X2_1093 ( .A(_abc_17692_n3191), .B(state_7_bF_buf1), .Y(_abc_17692_n3192) );
  AND2X2 AND2X2_1094 ( .A(_abc_17692_n1885_bF_buf2), .B(workunit2_7_), .Y(_abc_17692_n3193) );
  AND2X2 AND2X2_1095 ( .A(state_8_bF_buf2), .B(\data_in2[7] ), .Y(_abc_17692_n3194) );
  AND2X2 AND2X2_1096 ( .A(_abc_17692_n2831), .B(_abc_17692_n3034_1), .Y(_abc_17692_n3199) );
  AND2X2 AND2X2_1097 ( .A(_abc_17692_n2816), .B(_abc_17692_n3199), .Y(_abc_17692_n3200) );
  AND2X2 AND2X2_1098 ( .A(_abc_17692_n3200), .B(_abc_17692_n2448), .Y(_abc_17692_n3201) );
  AND2X2 AND2X2_1099 ( .A(_abc_17692_n2819), .B(_abc_17692_n3199), .Y(_abc_17692_n3202) );
  AND2X2 AND2X2_11 ( .A(_abc_17692_n632), .B(delta_22_), .Y(delta_22__FF_INPUT) );
  AND2X2 AND2X2_110 ( .A(_abc_17692_n929), .B(_abc_17692_n927_1), .Y(_abc_17692_n930_1) );
  AND2X2 AND2X2_1100 ( .A(_abc_17692_n2826), .B(_abc_17692_n3029), .Y(_abc_17692_n3203) );
  AND2X2 AND2X2_1101 ( .A(_abc_17692_n3208), .B(workunit1_4_), .Y(_abc_17692_n3209) );
  AND2X2 AND2X2_1102 ( .A(_abc_17692_n2433), .B(workunit1_13_bF_buf1), .Y(_abc_17692_n3210) );
  AND2X2 AND2X2_1103 ( .A(_abc_17692_n3211), .B(workunit1_8_bF_buf0), .Y(_abc_17692_n3212) );
  AND2X2 AND2X2_1104 ( .A(_abc_17692_n3213), .B(_abc_17692_n3214), .Y(_abc_17692_n3215) );
  AND2X2 AND2X2_1105 ( .A(_abc_17692_n3215), .B(_abc_17692_n2250), .Y(_abc_17692_n3216) );
  AND2X2 AND2X2_1106 ( .A(_abc_17692_n3207), .B(_abc_17692_n3218), .Y(_abc_17692_n3219) );
  AND2X2 AND2X2_1107 ( .A(_abc_17692_n3224_1), .B(_abc_17692_n3204), .Y(_abc_17692_n3225) );
  AND2X2 AND2X2_1108 ( .A(_abc_17692_n3223), .B(_abc_17692_n3225), .Y(_abc_17692_n3226) );
  AND2X2 AND2X2_1109 ( .A(_abc_17692_n3226), .B(_abc_17692_n3217), .Y(_abc_17692_n3227_1) );
  AND2X2 AND2X2_111 ( .A(_abc_17692_n930_1), .B(_abc_17692_n932), .Y(_abc_17692_n933) );
  AND2X2 AND2X2_1110 ( .A(_abc_17692_n2852), .B(_abc_17692_n3076), .Y(_abc_17692_n3229) );
  AND2X2 AND2X2_1111 ( .A(_abc_17692_n2843), .B(_abc_17692_n3229), .Y(_abc_17692_n3230) );
  AND2X2 AND2X2_1112 ( .A(_abc_17692_n2503), .B(_abc_17692_n3230), .Y(_abc_17692_n3231) );
  AND2X2 AND2X2_1113 ( .A(_abc_17692_n2847), .B(_abc_17692_n3229), .Y(_abc_17692_n3232) );
  AND2X2 AND2X2_1114 ( .A(_abc_17692_n3075), .B(_abc_17692_n2849_1), .Y(_abc_17692_n3233) );
  AND2X2 AND2X2_1115 ( .A(sum_8_), .B(\key_in[72] ), .Y(_abc_17692_n3237) );
  AND2X2 AND2X2_1116 ( .A(_abc_17692_n3238), .B(_abc_17692_n3239), .Y(_abc_17692_n3240_1) );
  AND2X2 AND2X2_1117 ( .A(_abc_17692_n3236), .B(_abc_17692_n3240_1), .Y(_abc_17692_n3241) );
  AND2X2 AND2X2_1118 ( .A(_abc_17692_n3242), .B(_abc_17692_n3243), .Y(_abc_17692_n3244) );
  AND2X2 AND2X2_1119 ( .A(_abc_17692_n3247), .B(_abc_17692_n3249), .Y(_abc_17692_n3250) );
  AND2X2 AND2X2_112 ( .A(_abc_17692_n935), .B(state_15_bF_buf3), .Y(_abc_17692_n936) );
  AND2X2 AND2X2_1120 ( .A(_abc_17692_n3251), .B(_abc_17692_n3198), .Y(_abc_17692_n3252) );
  AND2X2 AND2X2_1121 ( .A(_abc_17692_n3250), .B(workunit2_8_bF_buf1), .Y(_abc_17692_n3253) );
  AND2X2 AND2X2_1122 ( .A(_abc_17692_n3257), .B(_abc_17692_n3088), .Y(_abc_17692_n3258_1) );
  AND2X2 AND2X2_1123 ( .A(_abc_17692_n3258_1), .B(_abc_17692_n3255), .Y(_abc_17692_n3260) );
  AND2X2 AND2X2_1124 ( .A(_abc_17692_n3261), .B(_abc_17692_n1877_bF_buf6), .Y(_abc_17692_n3262) );
  AND2X2 AND2X2_1125 ( .A(_abc_17692_n3262), .B(_abc_17692_n3259), .Y(_abc_17692_n3263) );
  AND2X2 AND2X2_1126 ( .A(_abc_17692_n3265), .B(_abc_17692_n3264), .Y(_abc_17692_n3266) );
  AND2X2 AND2X2_1127 ( .A(_abc_17692_n3268), .B(_abc_17692_n3266), .Y(_abc_17692_n3269) );
  AND2X2 AND2X2_1128 ( .A(_abc_17692_n2915), .B(_abc_17692_n3103), .Y(_abc_17692_n3271) );
  AND2X2 AND2X2_1129 ( .A(_abc_17692_n2906), .B(_abc_17692_n3271), .Y(_abc_17692_n3272) );
  AND2X2 AND2X2_113 ( .A(_abc_17692_n936), .B(_abc_17692_n934), .Y(_abc_17692_n937_1) );
  AND2X2 AND2X2_1130 ( .A(_abc_17692_n2529), .B(_abc_17692_n3272), .Y(_abc_17692_n3273) );
  AND2X2 AND2X2_1131 ( .A(_abc_17692_n3271), .B(_abc_17692_n2910), .Y(_abc_17692_n3274) );
  AND2X2 AND2X2_1132 ( .A(_abc_17692_n3102), .B(_abc_17692_n2912), .Y(_abc_17692_n3275) );
  AND2X2 AND2X2_1133 ( .A(sum_8_), .B(\key_in[40] ), .Y(_abc_17692_n3279) );
  AND2X2 AND2X2_1134 ( .A(_abc_17692_n3280), .B(_abc_17692_n3281), .Y(_abc_17692_n3282) );
  AND2X2 AND2X2_1135 ( .A(_abc_17692_n3278_1), .B(_abc_17692_n3282), .Y(_abc_17692_n3283) );
  AND2X2 AND2X2_1136 ( .A(_abc_17692_n3285), .B(_abc_17692_n3286), .Y(_abc_17692_n3287) );
  AND2X2 AND2X2_1137 ( .A(_abc_17692_n3287), .B(_abc_17692_n3288), .Y(_abc_17692_n3289) );
  AND2X2 AND2X2_1138 ( .A(_abc_17692_n3293), .B(_abc_17692_n3292), .Y(_abc_17692_n3294) );
  AND2X2 AND2X2_1139 ( .A(_abc_17692_n3294), .B(workunit2_8_bF_buf0), .Y(_abc_17692_n3295_1) );
  AND2X2 AND2X2_114 ( .A(_abc_17692_n723), .B(sum_1_), .Y(_abc_17692_n938) );
  AND2X2 AND2X2_1140 ( .A(_abc_17692_n3296), .B(_abc_17692_n3297), .Y(_abc_17692_n3298) );
  AND2X2 AND2X2_1141 ( .A(_abc_17692_n3270), .B(_abc_17692_n3298), .Y(_abc_17692_n3300) );
  AND2X2 AND2X2_1142 ( .A(_abc_17692_n3301), .B(_abc_17692_n1846_bF_buf6), .Y(_abc_17692_n3302) );
  AND2X2 AND2X2_1143 ( .A(_abc_17692_n3302), .B(_abc_17692_n3299), .Y(_abc_17692_n3303) );
  AND2X2 AND2X2_1144 ( .A(_abc_17692_n2883), .B(_abc_17692_n3047), .Y(_abc_17692_n3304) );
  AND2X2 AND2X2_1145 ( .A(_abc_17692_n2874), .B(_abc_17692_n3304), .Y(_abc_17692_n3305) );
  AND2X2 AND2X2_1146 ( .A(_abc_17692_n2464), .B(_abc_17692_n3305), .Y(_abc_17692_n3306) );
  AND2X2 AND2X2_1147 ( .A(_abc_17692_n3304), .B(_abc_17692_n2878), .Y(_abc_17692_n3307) );
  AND2X2 AND2X2_1148 ( .A(_abc_17692_n3046), .B(_abc_17692_n2880), .Y(_abc_17692_n3308) );
  AND2X2 AND2X2_1149 ( .A(sum_8_), .B(\key_in[8] ), .Y(_abc_17692_n3312) );
  AND2X2 AND2X2_115 ( .A(_abc_17692_n941), .B(state_3_bF_buf3), .Y(_abc_17692_n942) );
  AND2X2 AND2X2_1150 ( .A(_abc_17692_n3313), .B(_abc_17692_n3314), .Y(_abc_17692_n3315) );
  AND2X2 AND2X2_1151 ( .A(_abc_17692_n3311), .B(_abc_17692_n3315), .Y(_abc_17692_n3316) );
  AND2X2 AND2X2_1152 ( .A(_abc_17692_n3318), .B(_abc_17692_n3319), .Y(_abc_17692_n3320) );
  AND2X2 AND2X2_1153 ( .A(_abc_17692_n3320), .B(_abc_17692_n3321), .Y(_abc_17692_n3322) );
  AND2X2 AND2X2_1154 ( .A(_abc_17692_n3326), .B(_abc_17692_n3325), .Y(_abc_17692_n3327) );
  AND2X2 AND2X2_1155 ( .A(_abc_17692_n3327), .B(workunit2_8_bF_buf2), .Y(_abc_17692_n3328) );
  AND2X2 AND2X2_1156 ( .A(_abc_17692_n3329), .B(_abc_17692_n3330), .Y(_abc_17692_n3331) );
  AND2X2 AND2X2_1157 ( .A(_abc_17692_n2902), .B(_abc_17692_n2899), .Y(_abc_17692_n3333) );
  AND2X2 AND2X2_1158 ( .A(_abc_17692_n3334), .B(_abc_17692_n3065), .Y(_abc_17692_n3335) );
  AND2X2 AND2X2_1159 ( .A(_abc_17692_n3337), .B(_abc_17692_n3332), .Y(_abc_17692_n3338) );
  AND2X2 AND2X2_116 ( .A(_abc_17692_n942), .B(_abc_17692_n939), .Y(_abc_17692_n943) );
  AND2X2 AND2X2_1160 ( .A(_abc_17692_n3338), .B(_abc_17692_n3331), .Y(_abc_17692_n3340) );
  AND2X2 AND2X2_1161 ( .A(_abc_17692_n3341), .B(_abc_17692_n1830_bF_buf6), .Y(_abc_17692_n3342) );
  AND2X2 AND2X2_1162 ( .A(_abc_17692_n3342), .B(_abc_17692_n3339), .Y(_abc_17692_n3343) );
  AND2X2 AND2X2_1163 ( .A(_abc_17692_n3154), .B(_abc_17692_n3147), .Y(_abc_17692_n3346_1) );
  AND2X2 AND2X2_1164 ( .A(sum_8_), .B(\key_in[104] ), .Y(_abc_17692_n3348) );
  AND2X2 AND2X2_1165 ( .A(_abc_17692_n3349_1), .B(_abc_17692_n3350), .Y(_abc_17692_n3351) );
  AND2X2 AND2X2_1166 ( .A(_abc_17692_n3135), .B(_abc_17692_n2955), .Y(_abc_17692_n3352) );
  AND2X2 AND2X2_1167 ( .A(_abc_17692_n2958), .B(_abc_17692_n3136), .Y(_abc_17692_n3354) );
  AND2X2 AND2X2_1168 ( .A(_abc_17692_n2953), .B(_abc_17692_n3354), .Y(_abc_17692_n3355_1) );
  AND2X2 AND2X2_1169 ( .A(_abc_17692_n2949_1), .B(_abc_17692_n3354), .Y(_abc_17692_n3357) );
  AND2X2 AND2X2_117 ( .A(_abc_17692_n946), .B(delta_2_), .Y(_abc_17692_n947) );
  AND2X2 AND2X2_1170 ( .A(_abc_17692_n2559), .B(_abc_17692_n3357), .Y(_abc_17692_n3358) );
  AND2X2 AND2X2_1171 ( .A(_abc_17692_n3359), .B(_abc_17692_n3351), .Y(_abc_17692_n3360) );
  AND2X2 AND2X2_1172 ( .A(_abc_17692_n3363), .B(_abc_17692_n3362), .Y(_abc_17692_n3364) );
  AND2X2 AND2X2_1173 ( .A(_abc_17692_n3364), .B(_abc_17692_n3361), .Y(_abc_17692_n3365) );
  AND2X2 AND2X2_1174 ( .A(_abc_17692_n3366_1), .B(_abc_17692_n3228), .Y(_abc_17692_n3367) );
  AND2X2 AND2X2_1175 ( .A(_abc_17692_n3368), .B(_abc_17692_n3248), .Y(_abc_17692_n3369) );
  AND2X2 AND2X2_1176 ( .A(_abc_17692_n3370), .B(workunit2_8_bF_buf0), .Y(_abc_17692_n3371) );
  AND2X2 AND2X2_1177 ( .A(_abc_17692_n3372), .B(_abc_17692_n3373), .Y(_abc_17692_n3374) );
  AND2X2 AND2X2_1178 ( .A(_abc_17692_n3347), .B(_abc_17692_n3374), .Y(_abc_17692_n3376_1) );
  AND2X2 AND2X2_1179 ( .A(_abc_17692_n3377), .B(_abc_17692_n1863_bF_buf6), .Y(_abc_17692_n3378) );
  AND2X2 AND2X2_118 ( .A(_abc_17692_n948), .B(_abc_17692_n949_1), .Y(_abc_17692_n950) );
  AND2X2 AND2X2_1180 ( .A(_abc_17692_n3378), .B(_abc_17692_n3375), .Y(_abc_17692_n3379) );
  AND2X2 AND2X2_1181 ( .A(_abc_17692_n3380), .B(state_6_bF_buf1), .Y(_abc_17692_n3381) );
  AND2X2 AND2X2_1182 ( .A(_abc_17692_n3175), .B(_abc_17692_n3153_1), .Y(_abc_17692_n3385) );
  AND2X2 AND2X2_1183 ( .A(_abc_17692_n3386), .B(_abc_17692_n3382), .Y(_abc_17692_n3388_1) );
  AND2X2 AND2X2_1184 ( .A(_abc_17692_n3389), .B(_abc_17692_n1863_bF_buf5), .Y(_abc_17692_n3390) );
  AND2X2 AND2X2_1185 ( .A(_abc_17692_n3390), .B(_abc_17692_n3387), .Y(_abc_17692_n3391) );
  AND2X2 AND2X2_1186 ( .A(_abc_17692_n3181), .B(_abc_17692_n3090), .Y(_abc_17692_n3392) );
  AND2X2 AND2X2_1187 ( .A(_abc_17692_n3086), .B(workunit2_7_), .Y(_abc_17692_n3393) );
  AND2X2 AND2X2_1188 ( .A(_abc_17692_n3185), .B(_abc_17692_n3394), .Y(_abc_17692_n3395) );
  AND2X2 AND2X2_1189 ( .A(_abc_17692_n3397), .B(_abc_17692_n3254), .Y(_abc_17692_n3398) );
  AND2X2 AND2X2_119 ( .A(delta_1_), .B(sum_1_), .Y(_abc_17692_n952) );
  AND2X2 AND2X2_1190 ( .A(_abc_17692_n3400), .B(_abc_17692_n1877_bF_buf5), .Y(_abc_17692_n3401) );
  AND2X2 AND2X2_1191 ( .A(_abc_17692_n3401), .B(_abc_17692_n3399), .Y(_abc_17692_n3402) );
  AND2X2 AND2X2_1192 ( .A(_abc_17692_n3118), .B(workunit2_7_), .Y(_abc_17692_n3404) );
  AND2X2 AND2X2_1193 ( .A(_abc_17692_n3120), .B(_abc_17692_n3405), .Y(_abc_17692_n3406) );
  AND2X2 AND2X2_1194 ( .A(_abc_17692_n3120), .B(_abc_17692_n2931), .Y(_abc_17692_n3408) );
  AND2X2 AND2X2_1195 ( .A(_abc_17692_n2990), .B(_abc_17692_n3408), .Y(_abc_17692_n3409) );
  AND2X2 AND2X2_1196 ( .A(_abc_17692_n3410), .B(_abc_17692_n3403), .Y(_abc_17692_n3412) );
  AND2X2 AND2X2_1197 ( .A(_abc_17692_n3413), .B(_abc_17692_n1846_bF_buf5), .Y(_abc_17692_n3414) );
  AND2X2 AND2X2_1198 ( .A(_abc_17692_n3414), .B(_abc_17692_n3411), .Y(_abc_17692_n3415) );
  AND2X2 AND2X2_1199 ( .A(_abc_17692_n3061), .B(workunit2_7_), .Y(_abc_17692_n3417) );
  AND2X2 AND2X2_12 ( .A(_abc_17692_n632), .B(delta_23_), .Y(delta_23__FF_INPUT) );
  AND2X2 AND2X2_120 ( .A(_abc_17692_n939), .B(_abc_17692_n953), .Y(_abc_17692_n954) );
  AND2X2 AND2X2_1200 ( .A(_abc_17692_n3063), .B(_abc_17692_n2893), .Y(_abc_17692_n3418) );
  AND2X2 AND2X2_1201 ( .A(_abc_17692_n3063), .B(_abc_17692_n2896), .Y(_abc_17692_n3420) );
  AND2X2 AND2X2_1202 ( .A(_abc_17692_n3420), .B(_abc_17692_n2982), .Y(_abc_17692_n3421) );
  AND2X2 AND2X2_1203 ( .A(_abc_17692_n3422), .B(_abc_17692_n3416), .Y(_abc_17692_n3423) );
  AND2X2 AND2X2_1204 ( .A(_abc_17692_n3425), .B(_abc_17692_n1830_bF_buf5), .Y(_abc_17692_n3426) );
  AND2X2 AND2X2_1205 ( .A(_abc_17692_n3426), .B(_abc_17692_n3424_1), .Y(_abc_17692_n3427_1) );
  AND2X2 AND2X2_1206 ( .A(_abc_17692_n3430), .B(state_7_bF_buf0), .Y(_abc_17692_n3431) );
  AND2X2 AND2X2_1207 ( .A(_abc_17692_n1885_bF_buf1), .B(workunit2_8_bF_buf2), .Y(_abc_17692_n3432) );
  AND2X2 AND2X2_1208 ( .A(state_8_bF_buf1), .B(\data_in2[8] ), .Y(_abc_17692_n3433) );
  AND2X2 AND2X2_1209 ( .A(_abc_17692_n3261), .B(_abc_17692_n3437), .Y(_abc_17692_n3438) );
  AND2X2 AND2X2_121 ( .A(_abc_17692_n957), .B(state_3_bF_buf2), .Y(_abc_17692_n958) );
  AND2X2 AND2X2_1210 ( .A(workunit1_5_), .B(workunit1_14_bF_buf2), .Y(_abc_17692_n3441) );
  AND2X2 AND2X2_1211 ( .A(_abc_17692_n3442), .B(_abc_17692_n3443), .Y(_abc_17692_n3444_1) );
  AND2X2 AND2X2_1212 ( .A(_abc_17692_n3444_1), .B(workunit1_9_), .Y(_abc_17692_n3445) );
  AND2X2 AND2X2_1213 ( .A(_abc_17692_n3447), .B(_abc_17692_n2435), .Y(_abc_17692_n3448) );
  AND2X2 AND2X2_1214 ( .A(_abc_17692_n3440), .B(_abc_17692_n3450), .Y(_abc_17692_n3451) );
  AND2X2 AND2X2_1215 ( .A(_abc_17692_n3439), .B(_abc_17692_n3449), .Y(_abc_17692_n3452) );
  AND2X2 AND2X2_1216 ( .A(sum_9_), .B(\key_in[73] ), .Y(_abc_17692_n3456) );
  AND2X2 AND2X2_1217 ( .A(_abc_17692_n3457), .B(_abc_17692_n3458), .Y(_abc_17692_n3459) );
  AND2X2 AND2X2_1218 ( .A(_abc_17692_n3455), .B(_abc_17692_n3459), .Y(_abc_17692_n3460) );
  AND2X2 AND2X2_1219 ( .A(_abc_17692_n3454), .B(_abc_17692_n3461), .Y(_abc_17692_n3462) );
  AND2X2 AND2X2_122 ( .A(_abc_17692_n958), .B(_abc_17692_n956), .Y(_abc_17692_n959) );
  AND2X2 AND2X2_1220 ( .A(_abc_17692_n3453), .B(_abc_17692_n3463), .Y(_abc_17692_n3464) );
  AND2X2 AND2X2_1221 ( .A(_abc_17692_n3465), .B(_abc_17692_n3466), .Y(_abc_17692_n3467) );
  AND2X2 AND2X2_1222 ( .A(_abc_17692_n3469), .B(workunit2_9_), .Y(_abc_17692_n3470) );
  AND2X2 AND2X2_1223 ( .A(_abc_17692_n3468), .B(_abc_17692_n3471), .Y(_abc_17692_n3472_1) );
  AND2X2 AND2X2_1224 ( .A(_abc_17692_n3438), .B(_abc_17692_n3473), .Y(_abc_17692_n3474) );
  AND2X2 AND2X2_1225 ( .A(_abc_17692_n3475), .B(_abc_17692_n3476), .Y(_abc_17692_n3477) );
  AND2X2 AND2X2_1226 ( .A(_abc_17692_n3478), .B(_abc_17692_n1877_bF_buf4), .Y(_abc_17692_n3479) );
  AND2X2 AND2X2_1227 ( .A(_abc_17692_n3301), .B(_abc_17692_n3296), .Y(_abc_17692_n3480) );
  AND2X2 AND2X2_1228 ( .A(sum_9_), .B(\key_in[41] ), .Y(_abc_17692_n3484) );
  AND2X2 AND2X2_1229 ( .A(_abc_17692_n3485), .B(_abc_17692_n3486), .Y(_abc_17692_n3487) );
  AND2X2 AND2X2_123 ( .A(_abc_17692_n723), .B(sum_2_), .Y(_abc_17692_n960) );
  AND2X2 AND2X2_1230 ( .A(_abc_17692_n3483), .B(_abc_17692_n3487), .Y(_abc_17692_n3488) );
  AND2X2 AND2X2_1231 ( .A(_abc_17692_n3493), .B(_abc_17692_n3489), .Y(_abc_17692_n3494) );
  AND2X2 AND2X2_1232 ( .A(_abc_17692_n3492), .B(_abc_17692_n3495), .Y(_abc_17692_n3496) );
  AND2X2 AND2X2_1233 ( .A(_abc_17692_n3498), .B(_abc_17692_n3499), .Y(_abc_17692_n3500) );
  AND2X2 AND2X2_1234 ( .A(_abc_17692_n3497), .B(_abc_17692_n3501), .Y(_abc_17692_n3502) );
  AND2X2 AND2X2_1235 ( .A(_abc_17692_n3505), .B(_abc_17692_n1846_bF_buf4), .Y(_abc_17692_n3506) );
  AND2X2 AND2X2_1236 ( .A(_abc_17692_n3506), .B(_abc_17692_n3504), .Y(_abc_17692_n3507) );
  AND2X2 AND2X2_1237 ( .A(_abc_17692_n3341), .B(_abc_17692_n3329), .Y(_abc_17692_n3508) );
  AND2X2 AND2X2_1238 ( .A(sum_9_), .B(\key_in[9] ), .Y(_abc_17692_n3511) );
  AND2X2 AND2X2_1239 ( .A(_abc_17692_n3512), .B(_abc_17692_n3513), .Y(_abc_17692_n3514) );
  AND2X2 AND2X2_124 ( .A(_abc_17692_n961), .B(_abc_17692_n950), .Y(_abc_17692_n962) );
  AND2X2 AND2X2_1240 ( .A(_abc_17692_n3510), .B(_abc_17692_n3515), .Y(_abc_17692_n3517) );
  AND2X2 AND2X2_1241 ( .A(_abc_17692_n3518), .B(_abc_17692_n3516), .Y(_abc_17692_n3519) );
  AND2X2 AND2X2_1242 ( .A(_abc_17692_n3520), .B(_abc_17692_n3522), .Y(_abc_17692_n3523) );
  AND2X2 AND2X2_1243 ( .A(_abc_17692_n3525), .B(_abc_17692_n3526), .Y(_abc_17692_n3527) );
  AND2X2 AND2X2_1244 ( .A(_abc_17692_n3530), .B(_abc_17692_n1830_bF_buf4), .Y(_abc_17692_n3531) );
  AND2X2 AND2X2_1245 ( .A(_abc_17692_n3531), .B(_abc_17692_n3529), .Y(_abc_17692_n3532) );
  AND2X2 AND2X2_1246 ( .A(_abc_17692_n3377), .B(_abc_17692_n3372), .Y(_abc_17692_n3535) );
  AND2X2 AND2X2_1247 ( .A(sum_9_), .B(\key_in[105] ), .Y(_abc_17692_n3537) );
  AND2X2 AND2X2_1248 ( .A(_abc_17692_n3538), .B(_abc_17692_n3539), .Y(_abc_17692_n3540) );
  AND2X2 AND2X2_1249 ( .A(_abc_17692_n3536), .B(_abc_17692_n3541), .Y(_abc_17692_n3543) );
  AND2X2 AND2X2_125 ( .A(_abc_17692_n964_1), .B(state_15_bF_buf2), .Y(_abc_17692_n965) );
  AND2X2 AND2X2_1250 ( .A(_abc_17692_n3544), .B(_abc_17692_n3542), .Y(_abc_17692_n3545) );
  AND2X2 AND2X2_1251 ( .A(_abc_17692_n3548), .B(_abc_17692_n3546), .Y(_abc_17692_n3549) );
  AND2X2 AND2X2_1252 ( .A(_abc_17692_n3551), .B(_abc_17692_n3552), .Y(_abc_17692_n3553) );
  AND2X2 AND2X2_1253 ( .A(_abc_17692_n3535), .B(_abc_17692_n3554), .Y(_abc_17692_n3555) );
  AND2X2 AND2X2_1254 ( .A(_abc_17692_n3556), .B(_abc_17692_n3553), .Y(_abc_17692_n3557) );
  AND2X2 AND2X2_1255 ( .A(_abc_17692_n3558), .B(_abc_17692_n1863_bF_buf4), .Y(_abc_17692_n3559) );
  AND2X2 AND2X2_1256 ( .A(_abc_17692_n3560), .B(state_6_bF_buf0), .Y(_abc_17692_n3561) );
  AND2X2 AND2X2_1257 ( .A(_abc_17692_n3562), .B(workunit2_8_bF_buf1), .Y(_abc_17692_n3563) );
  AND2X2 AND2X2_1258 ( .A(_abc_17692_n3389), .B(_abc_17692_n3564), .Y(_abc_17692_n3565) );
  AND2X2 AND2X2_1259 ( .A(_abc_17692_n3566), .B(_abc_17692_n3554), .Y(_abc_17692_n3567) );
  AND2X2 AND2X2_126 ( .A(_abc_17692_n965), .B(_abc_17692_n963), .Y(_abc_17692_n966) );
  AND2X2 AND2X2_1260 ( .A(_abc_17692_n3565), .B(_abc_17692_n3553), .Y(_abc_17692_n3568) );
  AND2X2 AND2X2_1261 ( .A(_abc_17692_n3569), .B(_abc_17692_n1863_bF_buf3), .Y(_abc_17692_n3570) );
  AND2X2 AND2X2_1262 ( .A(_abc_17692_n3251), .B(workunit2_8_bF_buf0), .Y(_abc_17692_n3571) );
  AND2X2 AND2X2_1263 ( .A(_abc_17692_n3399), .B(_abc_17692_n3572), .Y(_abc_17692_n3573) );
  AND2X2 AND2X2_1264 ( .A(_abc_17692_n3576), .B(_abc_17692_n1877_bF_buf3), .Y(_abc_17692_n3577) );
  AND2X2 AND2X2_1265 ( .A(_abc_17692_n3577), .B(_abc_17692_n3575), .Y(_abc_17692_n3578) );
  AND2X2 AND2X2_1266 ( .A(_abc_17692_n3579), .B(workunit2_8_bF_buf3), .Y(_abc_17692_n3580) );
  AND2X2 AND2X2_1267 ( .A(_abc_17692_n3424_1), .B(_abc_17692_n3581), .Y(_abc_17692_n3582) );
  AND2X2 AND2X2_1268 ( .A(_abc_17692_n3585), .B(_abc_17692_n1830_bF_buf3), .Y(_abc_17692_n3586) );
  AND2X2 AND2X2_1269 ( .A(_abc_17692_n3586), .B(_abc_17692_n3583), .Y(_abc_17692_n3587) );
  AND2X2 AND2X2_127 ( .A(_abc_17692_n969), .B(delta_3_), .Y(_abc_17692_n970) );
  AND2X2 AND2X2_1270 ( .A(_abc_17692_n3588), .B(workunit2_8_bF_buf2), .Y(_abc_17692_n3589) );
  AND2X2 AND2X2_1271 ( .A(_abc_17692_n3413), .B(_abc_17692_n3590), .Y(_abc_17692_n3591) );
  AND2X2 AND2X2_1272 ( .A(_abc_17692_n3594), .B(_abc_17692_n1846_bF_buf3), .Y(_abc_17692_n3595) );
  AND2X2 AND2X2_1273 ( .A(_abc_17692_n3595), .B(_abc_17692_n3593), .Y(_abc_17692_n3596) );
  AND2X2 AND2X2_1274 ( .A(_abc_17692_n3599), .B(state_7_bF_buf4), .Y(_abc_17692_n3600) );
  AND2X2 AND2X2_1275 ( .A(_abc_17692_n1885_bF_buf0), .B(workunit2_9_), .Y(_abc_17692_n3601) );
  AND2X2 AND2X2_1276 ( .A(state_8_bF_buf0), .B(\data_in2[9] ), .Y(_abc_17692_n3602) );
  AND2X2 AND2X2_1277 ( .A(_abc_17692_n3207), .B(_abc_17692_n3607), .Y(_abc_17692_n3608) );
  AND2X2 AND2X2_1278 ( .A(_abc_17692_n3610), .B(_abc_17692_n3609), .Y(_abc_17692_n3611) );
  AND2X2 AND2X2_1279 ( .A(_abc_17692_n3613), .B(_abc_17692_n3615), .Y(_abc_17692_n3616) );
  AND2X2 AND2X2_128 ( .A(_abc_17692_n972_1), .B(sum_3_), .Y(_abc_17692_n973) );
  AND2X2 AND2X2_1280 ( .A(_abc_17692_n3614), .B(workunit1_6_), .Y(_abc_17692_n3618_1) );
  AND2X2 AND2X2_1281 ( .A(_abc_17692_n2821), .B(workunit1_15_), .Y(_abc_17692_n3619) );
  AND2X2 AND2X2_1282 ( .A(_abc_17692_n3621_1), .B(_abc_17692_n3617), .Y(_abc_17692_n3622) );
  AND2X2 AND2X2_1283 ( .A(_abc_17692_n3612), .B(_abc_17692_n3622), .Y(_abc_17692_n3623) );
  AND2X2 AND2X2_1284 ( .A(_abc_17692_n3627), .B(_abc_17692_n3625), .Y(_abc_17692_n3628) );
  AND2X2 AND2X2_1285 ( .A(_abc_17692_n3624), .B(_abc_17692_n3628), .Y(_abc_17692_n3629) );
  AND2X2 AND2X2_1286 ( .A(_abc_17692_n3620), .B(workunit1_10_), .Y(_abc_17692_n3630_1) );
  AND2X2 AND2X2_1287 ( .A(_abc_17692_n3616), .B(_abc_17692_n2638), .Y(_abc_17692_n3631) );
  AND2X2 AND2X2_1288 ( .A(_abc_17692_n3629), .B(_abc_17692_n3632), .Y(_abc_17692_n3633) );
  AND2X2 AND2X2_1289 ( .A(_abc_17692_n3240_1), .B(_abc_17692_n3459), .Y(_abc_17692_n3635) );
  AND2X2 AND2X2_129 ( .A(_abc_17692_n971), .B(_abc_17692_n974), .Y(_abc_17692_n975) );
  AND2X2 AND2X2_1290 ( .A(_abc_17692_n3236), .B(_abc_17692_n3635), .Y(_abc_17692_n3636) );
  AND2X2 AND2X2_1291 ( .A(_abc_17692_n3238), .B(_abc_17692_n3457), .Y(_abc_17692_n3638) );
  AND2X2 AND2X2_1292 ( .A(sum_10_), .B(\key_in[74] ), .Y(_abc_17692_n3642) );
  AND2X2 AND2X2_1293 ( .A(_abc_17692_n3643), .B(_abc_17692_n3644), .Y(_abc_17692_n3645) );
  AND2X2 AND2X2_1294 ( .A(_abc_17692_n3641), .B(_abc_17692_n3645), .Y(_abc_17692_n3646) );
  AND2X2 AND2X2_1295 ( .A(_abc_17692_n3647), .B(_abc_17692_n3648), .Y(_abc_17692_n3649) );
  AND2X2 AND2X2_1296 ( .A(_abc_17692_n3652), .B(_abc_17692_n3654), .Y(_abc_17692_n3655) );
  AND2X2 AND2X2_1297 ( .A(_abc_17692_n3655), .B(workunit2_10_bF_buf2), .Y(_abc_17692_n3656) );
  AND2X2 AND2X2_1298 ( .A(_abc_17692_n3657), .B(_abc_17692_n3658), .Y(_abc_17692_n3659) );
  AND2X2 AND2X2_1299 ( .A(_abc_17692_n3473), .B(_abc_17692_n3255), .Y(_abc_17692_n3661_1) );
  AND2X2 AND2X2_13 ( .A(_abc_17692_n632), .B(delta_24_), .Y(delta_24__FF_INPUT) );
  AND2X2 AND2X2_130 ( .A(_abc_17692_n981), .B(state_15_bF_buf1), .Y(_abc_17692_n982) );
  AND2X2 AND2X2_1300 ( .A(_abc_17692_n3468), .B(workunit2_9_), .Y(_abc_17692_n3664) );
  AND2X2 AND2X2_1301 ( .A(_abc_17692_n3473), .B(_abc_17692_n3253), .Y(_abc_17692_n3665) );
  AND2X2 AND2X2_1302 ( .A(_abc_17692_n3663), .B(_abc_17692_n3667), .Y(_abc_17692_n3668) );
  AND2X2 AND2X2_1303 ( .A(_abc_17692_n3669), .B(_abc_17692_n3659), .Y(_abc_17692_n3671) );
  AND2X2 AND2X2_1304 ( .A(_abc_17692_n3672), .B(_abc_17692_n1877_bF_buf2), .Y(_abc_17692_n3673) );
  AND2X2 AND2X2_1305 ( .A(_abc_17692_n3673), .B(_abc_17692_n3670), .Y(_abc_17692_n3674) );
  AND2X2 AND2X2_1306 ( .A(_abc_17692_n3282), .B(_abc_17692_n3487), .Y(_abc_17692_n3675) );
  AND2X2 AND2X2_1307 ( .A(_abc_17692_n3278_1), .B(_abc_17692_n3675), .Y(_abc_17692_n3676) );
  AND2X2 AND2X2_1308 ( .A(_abc_17692_n3677), .B(_abc_17692_n3486), .Y(_abc_17692_n3678) );
  AND2X2 AND2X2_1309 ( .A(sum_10_), .B(\key_in[42] ), .Y(_abc_17692_n3680) );
  AND2X2 AND2X2_131 ( .A(_abc_17692_n982), .B(_abc_17692_n978), .Y(_abc_17692_n983) );
  AND2X2 AND2X2_1310 ( .A(_abc_17692_n3681), .B(_abc_17692_n3682), .Y(_abc_17692_n3683) );
  AND2X2 AND2X2_1311 ( .A(_abc_17692_n3679), .B(_abc_17692_n3683), .Y(_abc_17692_n3684) );
  AND2X2 AND2X2_1312 ( .A(_abc_17692_n3685), .B(_abc_17692_n3686), .Y(_abc_17692_n3687) );
  AND2X2 AND2X2_1313 ( .A(_abc_17692_n3687), .B(_abc_17692_n3688), .Y(_abc_17692_n3689) );
  AND2X2 AND2X2_1314 ( .A(_abc_17692_n3653), .B(_abc_17692_n3690), .Y(_abc_17692_n3691) );
  AND2X2 AND2X2_1315 ( .A(_abc_17692_n3692), .B(_abc_17692_n3634), .Y(_abc_17692_n3693) );
  AND2X2 AND2X2_1316 ( .A(_abc_17692_n3694), .B(workunit2_10_bF_buf0), .Y(_abc_17692_n3695) );
  AND2X2 AND2X2_1317 ( .A(_abc_17692_n3696_1), .B(_abc_17692_n3697), .Y(_abc_17692_n3698) );
  AND2X2 AND2X2_1318 ( .A(_abc_17692_n3496), .B(workunit2_9_), .Y(_abc_17692_n3702) );
  AND2X2 AND2X2_1319 ( .A(_abc_17692_n3704), .B(_abc_17692_n3703), .Y(_abc_17692_n3705) );
  AND2X2 AND2X2_132 ( .A(_abc_17692_n723), .B(sum_3_), .Y(_abc_17692_n984) );
  AND2X2 AND2X2_1320 ( .A(_abc_17692_n3701), .B(_abc_17692_n3705), .Y(_abc_17692_n3706) );
  AND2X2 AND2X2_1321 ( .A(_abc_17692_n3707), .B(_abc_17692_n3699_1), .Y(_abc_17692_n3708) );
  AND2X2 AND2X2_1322 ( .A(_abc_17692_n3710), .B(_abc_17692_n1846_bF_buf2), .Y(_abc_17692_n3711) );
  AND2X2 AND2X2_1323 ( .A(_abc_17692_n3711), .B(_abc_17692_n3709), .Y(_abc_17692_n3712_1) );
  AND2X2 AND2X2_1324 ( .A(_abc_17692_n3315), .B(_abc_17692_n3514), .Y(_abc_17692_n3713) );
  AND2X2 AND2X2_1325 ( .A(_abc_17692_n3311), .B(_abc_17692_n3713), .Y(_abc_17692_n3714) );
  AND2X2 AND2X2_1326 ( .A(_abc_17692_n3715), .B(_abc_17692_n3513), .Y(_abc_17692_n3716) );
  AND2X2 AND2X2_1327 ( .A(sum_10_), .B(\key_in[10] ), .Y(_abc_17692_n3718) );
  AND2X2 AND2X2_1328 ( .A(_abc_17692_n3719), .B(_abc_17692_n3720), .Y(_abc_17692_n3721) );
  AND2X2 AND2X2_1329 ( .A(_abc_17692_n3717), .B(_abc_17692_n3721), .Y(_abc_17692_n3722) );
  AND2X2 AND2X2_133 ( .A(delta_2_), .B(sum_2_), .Y(_abc_17692_n985) );
  AND2X2 AND2X2_1330 ( .A(_abc_17692_n3723), .B(_abc_17692_n3724), .Y(_abc_17692_n3725) );
  AND2X2 AND2X2_1331 ( .A(_abc_17692_n3728), .B(_abc_17692_n3729), .Y(_abc_17692_n3730) );
  AND2X2 AND2X2_1332 ( .A(_abc_17692_n3730), .B(workunit2_10_bF_buf1), .Y(_abc_17692_n3732) );
  AND2X2 AND2X2_1333 ( .A(_abc_17692_n3733_1), .B(_abc_17692_n3731), .Y(_abc_17692_n3734) );
  AND2X2 AND2X2_1334 ( .A(_abc_17692_n3338), .B(_abc_17692_n3736), .Y(_abc_17692_n3737) );
  AND2X2 AND2X2_1335 ( .A(_abc_17692_n3524), .B(workunit2_9_), .Y(_abc_17692_n3738) );
  AND2X2 AND2X2_1336 ( .A(_abc_17692_n3740), .B(_abc_17692_n3739), .Y(_abc_17692_n3741) );
  AND2X2 AND2X2_1337 ( .A(_abc_17692_n3743), .B(_abc_17692_n3734), .Y(_abc_17692_n3744) );
  AND2X2 AND2X2_1338 ( .A(_abc_17692_n3746), .B(_abc_17692_n1830_bF_buf2), .Y(_abc_17692_n3747) );
  AND2X2 AND2X2_1339 ( .A(_abc_17692_n3747), .B(_abc_17692_n3745), .Y(_abc_17692_n3748) );
  AND2X2 AND2X2_134 ( .A(_abc_17692_n957), .B(_abc_17692_n986), .Y(_abc_17692_n987) );
  AND2X2 AND2X2_1340 ( .A(_abc_17692_n3351), .B(_abc_17692_n3540), .Y(_abc_17692_n3752) );
  AND2X2 AND2X2_1341 ( .A(_abc_17692_n3359), .B(_abc_17692_n3752), .Y(_abc_17692_n3753) );
  AND2X2 AND2X2_1342 ( .A(_abc_17692_n3349_1), .B(_abc_17692_n3538), .Y(_abc_17692_n3755) );
  AND2X2 AND2X2_1343 ( .A(sum_10_), .B(\key_in[106] ), .Y(_abc_17692_n3759) );
  AND2X2 AND2X2_1344 ( .A(_abc_17692_n3760), .B(_abc_17692_n3761), .Y(_abc_17692_n3762) );
  AND2X2 AND2X2_1345 ( .A(_abc_17692_n3758), .B(_abc_17692_n3762), .Y(_abc_17692_n3763) );
  AND2X2 AND2X2_1346 ( .A(_abc_17692_n3764), .B(_abc_17692_n3765), .Y(_abc_17692_n3766) );
  AND2X2 AND2X2_1347 ( .A(_abc_17692_n3769), .B(_abc_17692_n3770), .Y(_abc_17692_n3771) );
  AND2X2 AND2X2_1348 ( .A(_abc_17692_n3774), .B(_abc_17692_n3772), .Y(_abc_17692_n3775) );
  AND2X2 AND2X2_1349 ( .A(_abc_17692_n3550), .B(workunit2_9_), .Y(_abc_17692_n3777) );
  AND2X2 AND2X2_135 ( .A(_abc_17692_n989), .B(_abc_17692_n990), .Y(_abc_17692_n991) );
  AND2X2 AND2X2_1350 ( .A(_abc_17692_n3779), .B(_abc_17692_n3778), .Y(_abc_17692_n3780) );
  AND2X2 AND2X2_1351 ( .A(_abc_17692_n3554), .B(_abc_17692_n3374), .Y(_abc_17692_n3782) );
  AND2X2 AND2X2_1352 ( .A(_abc_17692_n3347), .B(_abc_17692_n3782), .Y(_abc_17692_n3783) );
  AND2X2 AND2X2_1353 ( .A(_abc_17692_n3784), .B(_abc_17692_n3776_1), .Y(_abc_17692_n3786) );
  AND2X2 AND2X2_1354 ( .A(_abc_17692_n3787), .B(_abc_17692_n1863_bF_buf2), .Y(_abc_17692_n3788) );
  AND2X2 AND2X2_1355 ( .A(_abc_17692_n3788), .B(_abc_17692_n3785), .Y(_abc_17692_n3789) );
  AND2X2 AND2X2_1356 ( .A(_abc_17692_n3790), .B(state_6_bF_buf4), .Y(_abc_17692_n3791) );
  AND2X2 AND2X2_1357 ( .A(_abc_17692_n3178_1), .B(_abc_17692_n3383), .Y(_abc_17692_n3792) );
  AND2X2 AND2X2_1358 ( .A(_abc_17692_n3553), .B(_abc_17692_n3382), .Y(_abc_17692_n3793) );
  AND2X2 AND2X2_1359 ( .A(_abc_17692_n3552), .B(_abc_17692_n3563), .Y(_abc_17692_n3797) );
  AND2X2 AND2X2_136 ( .A(_abc_17692_n991), .B(state_3_bF_buf1), .Y(_abc_17692_n992) );
  AND2X2 AND2X2_1360 ( .A(_abc_17692_n3795), .B(_abc_17692_n3799), .Y(_abc_17692_n3800) );
  AND2X2 AND2X2_1361 ( .A(_abc_17692_n3801), .B(_abc_17692_n3775), .Y(_abc_17692_n3803) );
  AND2X2 AND2X2_1362 ( .A(_abc_17692_n3804), .B(_abc_17692_n1863_bF_buf1), .Y(_abc_17692_n3805) );
  AND2X2 AND2X2_1363 ( .A(_abc_17692_n3805), .B(_abc_17692_n3802), .Y(_abc_17692_n3806) );
  AND2X2 AND2X2_1364 ( .A(_abc_17692_n3397), .B(_abc_17692_n3809), .Y(_abc_17692_n3810) );
  AND2X2 AND2X2_1365 ( .A(_abc_17692_n3811), .B(_abc_17692_n3812), .Y(_abc_17692_n3813) );
  AND2X2 AND2X2_1366 ( .A(_abc_17692_n3815), .B(_abc_17692_n3807), .Y(_abc_17692_n3816) );
  AND2X2 AND2X2_1367 ( .A(_abc_17692_n3818), .B(_abc_17692_n1877_bF_buf1), .Y(_abc_17692_n3819) );
  AND2X2 AND2X2_1368 ( .A(_abc_17692_n3819), .B(_abc_17692_n3817), .Y(_abc_17692_n3820) );
  AND2X2 AND2X2_1369 ( .A(_abc_17692_n2802), .B(_abc_17692_n2727), .Y(_abc_17692_n3822) );
  AND2X2 AND2X2_137 ( .A(_abc_17692_n995), .B(delta_4_), .Y(_abc_17692_n996_1) );
  AND2X2 AND2X2_1370 ( .A(_abc_17692_n3824), .B(_abc_17692_n3821), .Y(_abc_17692_n3825) );
  AND2X2 AND2X2_1371 ( .A(_abc_17692_n3502), .B(_abc_17692_n3403), .Y(_abc_17692_n3826) );
  AND2X2 AND2X2_1372 ( .A(_abc_17692_n3830), .B(_abc_17692_n3501), .Y(_abc_17692_n3831) );
  AND2X2 AND2X2_1373 ( .A(_abc_17692_n3828), .B(_abc_17692_n3832), .Y(_abc_17692_n3833) );
  AND2X2 AND2X2_1374 ( .A(_abc_17692_n3834_1), .B(_abc_17692_n3698), .Y(_abc_17692_n3836) );
  AND2X2 AND2X2_1375 ( .A(_abc_17692_n3837_1), .B(_abc_17692_n1846_bF_buf1), .Y(_abc_17692_n3838) );
  AND2X2 AND2X2_1376 ( .A(_abc_17692_n3838), .B(_abc_17692_n3835), .Y(_abc_17692_n3839) );
  AND2X2 AND2X2_1377 ( .A(_abc_17692_n3527), .B(_abc_17692_n3416), .Y(_abc_17692_n3842) );
  AND2X2 AND2X2_1378 ( .A(_abc_17692_n3526), .B(_abc_17692_n3580), .Y(_abc_17692_n3846) );
  AND2X2 AND2X2_1379 ( .A(_abc_17692_n3844), .B(_abc_17692_n3848), .Y(_abc_17692_n3849) );
  AND2X2 AND2X2_138 ( .A(delta_3_), .B(sum_3_), .Y(_abc_17692_n1000) );
  AND2X2 AND2X2_1380 ( .A(_abc_17692_n3850), .B(_abc_17692_n3840), .Y(_abc_17692_n3851) );
  AND2X2 AND2X2_1381 ( .A(_abc_17692_n3853), .B(_abc_17692_n1830_bF_buf1), .Y(_abc_17692_n3854) );
  AND2X2 AND2X2_1382 ( .A(_abc_17692_n3854), .B(_abc_17692_n3852), .Y(_abc_17692_n3855_1) );
  AND2X2 AND2X2_1383 ( .A(_abc_17692_n3858), .B(state_7_bF_buf3), .Y(_abc_17692_n3859) );
  AND2X2 AND2X2_1384 ( .A(_abc_17692_n1885_bF_buf4), .B(workunit2_10_bF_buf2), .Y(_abc_17692_n3860) );
  AND2X2 AND2X2_1385 ( .A(state_8_bF_buf9), .B(\data_in2[10] ), .Y(_abc_17692_n3861) );
  AND2X2 AND2X2_1386 ( .A(_abc_17692_n3672), .B(_abc_17692_n3657), .Y(_abc_17692_n3865) );
  AND2X2 AND2X2_1387 ( .A(_abc_17692_n3867), .B(workunit1_7_), .Y(_abc_17692_n3868) );
  AND2X2 AND2X2_1388 ( .A(_abc_17692_n2063), .B(workunit1_16_bF_buf1), .Y(_abc_17692_n3869) );
  AND2X2 AND2X2_1389 ( .A(_abc_17692_n3870), .B(workunit1_11_bF_buf3), .Y(_abc_17692_n3871) );
  AND2X2 AND2X2_139 ( .A(_abc_17692_n972_1), .B(_abc_17692_n969), .Y(_abc_17692_n1002) );
  AND2X2 AND2X2_1390 ( .A(_abc_17692_n3872), .B(_abc_17692_n3873), .Y(_abc_17692_n3874) );
  AND2X2 AND2X2_1391 ( .A(_abc_17692_n3874), .B(_abc_17692_n2823), .Y(_abc_17692_n3875) );
  AND2X2 AND2X2_1392 ( .A(_abc_17692_n3878), .B(_abc_17692_n3617), .Y(_abc_17692_n3879) );
  AND2X2 AND2X2_1393 ( .A(_abc_17692_n3881), .B(_abc_17692_n3880), .Y(_abc_17692_n3882) );
  AND2X2 AND2X2_1394 ( .A(_abc_17692_n3883), .B(_abc_17692_n3877_1), .Y(_abc_17692_n3884) );
  AND2X2 AND2X2_1395 ( .A(sum_11_), .B(\key_in[75] ), .Y(_abc_17692_n3887) );
  AND2X2 AND2X2_1396 ( .A(_abc_17692_n3888), .B(_abc_17692_n3889), .Y(_abc_17692_n3890) );
  AND2X2 AND2X2_1397 ( .A(_abc_17692_n3886), .B(_abc_17692_n3890), .Y(_abc_17692_n3891) );
  AND2X2 AND2X2_1398 ( .A(_abc_17692_n3885), .B(_abc_17692_n3893), .Y(_abc_17692_n3894) );
  AND2X2 AND2X2_1399 ( .A(_abc_17692_n3892), .B(_abc_17692_n3895), .Y(_abc_17692_n3896) );
  AND2X2 AND2X2_14 ( .A(_abc_17692_n632), .B(delta_29_), .Y(delta_29__FF_INPUT) );
  AND2X2 AND2X2_140 ( .A(_abc_17692_n1003), .B(_abc_17692_n1001), .Y(_abc_17692_n1004) );
  AND2X2 AND2X2_1400 ( .A(_abc_17692_n3879), .B(_abc_17692_n3882), .Y(_abc_17692_n3898) );
  AND2X2 AND2X2_1401 ( .A(_abc_17692_n3866_1), .B(_abc_17692_n3876), .Y(_abc_17692_n3899) );
  AND2X2 AND2X2_1402 ( .A(_abc_17692_n3897), .B(_abc_17692_n3902), .Y(_abc_17692_n3903) );
  AND2X2 AND2X2_1403 ( .A(_abc_17692_n3903), .B(workunit2_11_), .Y(_abc_17692_n3904) );
  AND2X2 AND2X2_1404 ( .A(_abc_17692_n3907), .B(_abc_17692_n3906), .Y(_abc_17692_n3908) );
  AND2X2 AND2X2_1405 ( .A(_abc_17692_n3908), .B(_abc_17692_n3905), .Y(_abc_17692_n3909) );
  AND2X2 AND2X2_1406 ( .A(_abc_17692_n3914), .B(_abc_17692_n1877_bF_buf0), .Y(_abc_17692_n3915_1) );
  AND2X2 AND2X2_1407 ( .A(_abc_17692_n3915_1), .B(_abc_17692_n3912_1), .Y(_abc_17692_n3916) );
  AND2X2 AND2X2_1408 ( .A(_abc_17692_n3709), .B(_abc_17692_n3917), .Y(_abc_17692_n3918) );
  AND2X2 AND2X2_1409 ( .A(_abc_17692_n3920), .B(_abc_17692_n3681), .Y(_abc_17692_n3921) );
  AND2X2 AND2X2_141 ( .A(_abc_17692_n1008), .B(state_3_bF_buf0), .Y(_abc_17692_n1009) );
  AND2X2 AND2X2_1410 ( .A(sum_11_), .B(\key_in[43] ), .Y(_abc_17692_n3922) );
  AND2X2 AND2X2_1411 ( .A(_abc_17692_n3923), .B(_abc_17692_n3924), .Y(_abc_17692_n3925) );
  AND2X2 AND2X2_1412 ( .A(_abc_17692_n3921), .B(_abc_17692_n3925), .Y(_abc_17692_n3926) );
  AND2X2 AND2X2_1413 ( .A(_abc_17692_n3927), .B(_abc_17692_n3928), .Y(_abc_17692_n3929) );
  AND2X2 AND2X2_1414 ( .A(_abc_17692_n3933), .B(_abc_17692_n3932), .Y(_abc_17692_n3934) );
  AND2X2 AND2X2_1415 ( .A(_abc_17692_n3931), .B(_abc_17692_n3935), .Y(_abc_17692_n3936) );
  AND2X2 AND2X2_1416 ( .A(_abc_17692_n3936), .B(workunit2_11_), .Y(_abc_17692_n3937) );
  AND2X2 AND2X2_1417 ( .A(_abc_17692_n3938), .B(_abc_17692_n3939), .Y(_abc_17692_n3940) );
  AND2X2 AND2X2_1418 ( .A(_abc_17692_n3940), .B(_abc_17692_n3905), .Y(_abc_17692_n3941) );
  AND2X2 AND2X2_1419 ( .A(_abc_17692_n3945), .B(_abc_17692_n1846_bF_buf0), .Y(_abc_17692_n3946) );
  AND2X2 AND2X2_142 ( .A(_abc_17692_n1009), .B(_abc_17692_n1006), .Y(_abc_17692_n1010) );
  AND2X2 AND2X2_1420 ( .A(_abc_17692_n3946), .B(_abc_17692_n3944), .Y(_abc_17692_n3947) );
  AND2X2 AND2X2_1421 ( .A(_abc_17692_n3745), .B(_abc_17692_n3733_1), .Y(_abc_17692_n3948) );
  AND2X2 AND2X2_1422 ( .A(sum_11_), .B(\key_in[11] ), .Y(_abc_17692_n3952) );
  AND2X2 AND2X2_1423 ( .A(_abc_17692_n3953), .B(_abc_17692_n3954_1), .Y(_abc_17692_n3955) );
  AND2X2 AND2X2_1424 ( .A(_abc_17692_n3951), .B(_abc_17692_n3955), .Y(_abc_17692_n3956) );
  AND2X2 AND2X2_1425 ( .A(_abc_17692_n3950), .B(_abc_17692_n3957), .Y(_abc_17692_n3958) );
  AND2X2 AND2X2_1426 ( .A(_abc_17692_n3962), .B(_abc_17692_n3960), .Y(_abc_17692_n3963) );
  AND2X2 AND2X2_1427 ( .A(_abc_17692_n3963), .B(workunit2_11_), .Y(_abc_17692_n3964) );
  AND2X2 AND2X2_1428 ( .A(_abc_17692_n3965), .B(_abc_17692_n3966), .Y(_abc_17692_n3967) );
  AND2X2 AND2X2_1429 ( .A(_abc_17692_n3967), .B(_abc_17692_n3905), .Y(_abc_17692_n3968) );
  AND2X2 AND2X2_143 ( .A(_abc_17692_n723), .B(sum_4_), .Y(_abc_17692_n1011) );
  AND2X2 AND2X2_1430 ( .A(_abc_17692_n3972), .B(_abc_17692_n1830_bF_buf0), .Y(_abc_17692_n3973) );
  AND2X2 AND2X2_1431 ( .A(_abc_17692_n3973), .B(_abc_17692_n3971), .Y(_abc_17692_n3974) );
  AND2X2 AND2X2_1432 ( .A(_abc_17692_n3771), .B(workunit2_10_bF_buf1), .Y(_abc_17692_n3977) );
  AND2X2 AND2X2_1433 ( .A(_abc_17692_n3787), .B(_abc_17692_n3978_1), .Y(_abc_17692_n3979) );
  AND2X2 AND2X2_1434 ( .A(sum_11_), .B(\key_in[107] ), .Y(_abc_17692_n3982) );
  AND2X2 AND2X2_1435 ( .A(_abc_17692_n3983), .B(_abc_17692_n3984), .Y(_abc_17692_n3985) );
  AND2X2 AND2X2_1436 ( .A(_abc_17692_n3981), .B(_abc_17692_n3985), .Y(_abc_17692_n3986) );
  AND2X2 AND2X2_1437 ( .A(_abc_17692_n3980), .B(_abc_17692_n3987), .Y(_abc_17692_n3988) );
  AND2X2 AND2X2_1438 ( .A(_abc_17692_n3992), .B(_abc_17692_n3991), .Y(_abc_17692_n3993) );
  AND2X2 AND2X2_1439 ( .A(_abc_17692_n3990), .B(_abc_17692_n3994), .Y(_abc_17692_n3995) );
  AND2X2 AND2X2_144 ( .A(_abc_17692_n977), .B(_abc_17692_n971), .Y(_abc_17692_n1012) );
  AND2X2 AND2X2_1440 ( .A(_abc_17692_n3995), .B(workunit2_11_), .Y(_abc_17692_n3996) );
  AND2X2 AND2X2_1441 ( .A(_abc_17692_n3998), .B(_abc_17692_n3997), .Y(_abc_17692_n3999) );
  AND2X2 AND2X2_1442 ( .A(_abc_17692_n3999), .B(_abc_17692_n3905), .Y(_abc_17692_n4000) );
  AND2X2 AND2X2_1443 ( .A(_abc_17692_n3979), .B(_abc_17692_n4002_1), .Y(_abc_17692_n4003) );
  AND2X2 AND2X2_1444 ( .A(_abc_17692_n4004), .B(_abc_17692_n4001), .Y(_abc_17692_n4005) );
  AND2X2 AND2X2_1445 ( .A(_abc_17692_n4006), .B(_abc_17692_n1863_bF_buf0), .Y(_abc_17692_n4007) );
  AND2X2 AND2X2_1446 ( .A(_abc_17692_n4008), .B(state_6_bF_buf3), .Y(_abc_17692_n4009) );
  AND2X2 AND2X2_1447 ( .A(_abc_17692_n3804), .B(_abc_17692_n3772), .Y(_abc_17692_n4010) );
  AND2X2 AND2X2_1448 ( .A(_abc_17692_n4011), .B(_abc_17692_n4002_1), .Y(_abc_17692_n4012) );
  AND2X2 AND2X2_1449 ( .A(_abc_17692_n4010), .B(_abc_17692_n4001), .Y(_abc_17692_n4013) );
  AND2X2 AND2X2_145 ( .A(_abc_17692_n1013), .B(_abc_17692_n1007), .Y(_abc_17692_n1014) );
  AND2X2 AND2X2_1450 ( .A(_abc_17692_n4014), .B(_abc_17692_n1863_bF_buf10), .Y(_abc_17692_n4015) );
  AND2X2 AND2X2_1451 ( .A(_abc_17692_n4016), .B(workunit2_10_bF_buf0), .Y(_abc_17692_n4017) );
  AND2X2 AND2X2_1452 ( .A(_abc_17692_n3817), .B(_abc_17692_n4018), .Y(_abc_17692_n4019) );
  AND2X2 AND2X2_1453 ( .A(_abc_17692_n4022), .B(_abc_17692_n1877_bF_buf10), .Y(_abc_17692_n4023) );
  AND2X2 AND2X2_1454 ( .A(_abc_17692_n4023), .B(_abc_17692_n4021), .Y(_abc_17692_n4024) );
  AND2X2 AND2X2_1455 ( .A(_abc_17692_n3837_1), .B(_abc_17692_n3696_1), .Y(_abc_17692_n4025) );
  AND2X2 AND2X2_1456 ( .A(_abc_17692_n4028), .B(_abc_17692_n1846_bF_buf10), .Y(_abc_17692_n4029) );
  AND2X2 AND2X2_1457 ( .A(_abc_17692_n4029), .B(_abc_17692_n4027), .Y(_abc_17692_n4030) );
  AND2X2 AND2X2_1458 ( .A(_abc_17692_n3852), .B(_abc_17692_n4031), .Y(_abc_17692_n4032) );
  AND2X2 AND2X2_1459 ( .A(_abc_17692_n4035), .B(_abc_17692_n1830_bF_buf10), .Y(_abc_17692_n4036) );
  AND2X2 AND2X2_146 ( .A(_abc_17692_n1016), .B(state_15_bF_buf0), .Y(_abc_17692_n1017) );
  AND2X2 AND2X2_1460 ( .A(_abc_17692_n4036), .B(_abc_17692_n4034), .Y(_abc_17692_n4037) );
  AND2X2 AND2X2_1461 ( .A(_abc_17692_n4040), .B(state_7_bF_buf2), .Y(_abc_17692_n4041) );
  AND2X2 AND2X2_1462 ( .A(_abc_17692_n1885_bF_buf3), .B(workunit2_11_), .Y(_abc_17692_n4042) );
  AND2X2 AND2X2_1463 ( .A(state_8_bF_buf8), .B(\data_in2[11] ), .Y(_abc_17692_n4043) );
  AND2X2 AND2X2_1464 ( .A(_abc_17692_n3622), .B(_abc_17692_n3882), .Y(_abc_17692_n4048) );
  AND2X2 AND2X2_1465 ( .A(_abc_17692_n4048), .B(_abc_17692_n3611), .Y(_abc_17692_n4049) );
  AND2X2 AND2X2_1466 ( .A(_abc_17692_n3617), .B(_abc_17692_n3880), .Y(_abc_17692_n4050) );
  AND2X2 AND2X2_1467 ( .A(_abc_17692_n3207), .B(_abc_17692_n4056), .Y(_abc_17692_n4057) );
  AND2X2 AND2X2_1468 ( .A(_abc_17692_n4059), .B(workunit1_8_bF_buf3), .Y(_abc_17692_n4060) );
  AND2X2 AND2X2_1469 ( .A(_abc_17692_n2250), .B(workunit1_17_), .Y(_abc_17692_n4061) );
  AND2X2 AND2X2_147 ( .A(_abc_17692_n1017), .B(_abc_17692_n1015), .Y(_abc_17692_n1018) );
  AND2X2 AND2X2_1470 ( .A(_abc_17692_n4062), .B(workunit1_12_bF_buf3), .Y(_abc_17692_n4063) );
  AND2X2 AND2X2_1471 ( .A(_abc_17692_n4064_1), .B(_abc_17692_n4065), .Y(_abc_17692_n4066) );
  AND2X2 AND2X2_1472 ( .A(_abc_17692_n4058), .B(_abc_17692_n4066), .Y(_abc_17692_n4067_1) );
  AND2X2 AND2X2_1473 ( .A(_abc_17692_n4068), .B(_abc_17692_n4051), .Y(_abc_17692_n4069) );
  AND2X2 AND2X2_1474 ( .A(_abc_17692_n4070), .B(_abc_17692_n4069), .Y(_abc_17692_n4071) );
  AND2X2 AND2X2_1475 ( .A(_abc_17692_n4071), .B(_abc_17692_n4072), .Y(_abc_17692_n4073_1) );
  AND2X2 AND2X2_1476 ( .A(_abc_17692_n3762), .B(_abc_17692_n3985), .Y(_abc_17692_n4075) );
  AND2X2 AND2X2_1477 ( .A(_abc_17692_n3757), .B(_abc_17692_n4075), .Y(_abc_17692_n4076) );
  AND2X2 AND2X2_1478 ( .A(_abc_17692_n3984), .B(_abc_17692_n3759), .Y(_abc_17692_n4077) );
  AND2X2 AND2X2_1479 ( .A(_abc_17692_n3752), .B(_abc_17692_n4075), .Y(_abc_17692_n4080) );
  AND2X2 AND2X2_148 ( .A(delta_5_), .B(sum_5_), .Y(_abc_17692_n1021) );
  AND2X2 AND2X2_1480 ( .A(_abc_17692_n3359), .B(_abc_17692_n4080), .Y(_abc_17692_n4081) );
  AND2X2 AND2X2_1481 ( .A(sum_12_), .B(\key_in[108] ), .Y(_abc_17692_n4083) );
  AND2X2 AND2X2_1482 ( .A(_abc_17692_n4084_1), .B(_abc_17692_n4085), .Y(_abc_17692_n4086) );
  AND2X2 AND2X2_1483 ( .A(_abc_17692_n4082), .B(_abc_17692_n4086), .Y(_abc_17692_n4087) );
  AND2X2 AND2X2_1484 ( .A(_abc_17692_n4089), .B(_abc_17692_n4088), .Y(_abc_17692_n4090) );
  AND2X2 AND2X2_1485 ( .A(_abc_17692_n4090), .B(_abc_17692_n4091), .Y(_abc_17692_n4092) );
  AND2X2 AND2X2_1486 ( .A(_abc_17692_n4095), .B(_abc_17692_n4097), .Y(_abc_17692_n4098) );
  AND2X2 AND2X2_1487 ( .A(_abc_17692_n4098), .B(workunit2_12_bF_buf2), .Y(_abc_17692_n4099) );
  AND2X2 AND2X2_1488 ( .A(_abc_17692_n4100), .B(_abc_17692_n4101), .Y(_abc_17692_n4102) );
  AND2X2 AND2X2_1489 ( .A(_abc_17692_n4002_1), .B(_abc_17692_n3776_1), .Y(_abc_17692_n4104) );
  AND2X2 AND2X2_149 ( .A(_abc_17692_n1023), .B(_abc_17692_n1024), .Y(_abc_17692_n1025_1) );
  AND2X2 AND2X2_1490 ( .A(_abc_17692_n4108), .B(_abc_17692_n3978_1), .Y(_abc_17692_n4109) );
  AND2X2 AND2X2_1491 ( .A(_abc_17692_n4111), .B(_abc_17692_n4110), .Y(_abc_17692_n4112) );
  AND2X2 AND2X2_1492 ( .A(_abc_17692_n4107_1), .B(_abc_17692_n4112), .Y(_abc_17692_n4113) );
  AND2X2 AND2X2_1493 ( .A(_abc_17692_n4114), .B(_abc_17692_n4102), .Y(_abc_17692_n4115) );
  AND2X2 AND2X2_1494 ( .A(_abc_17692_n4116), .B(_abc_17692_n4117), .Y(_abc_17692_n4118) );
  AND2X2 AND2X2_1495 ( .A(_abc_17692_n3645), .B(_abc_17692_n3890), .Y(_abc_17692_n4121) );
  AND2X2 AND2X2_1496 ( .A(_abc_17692_n3640_1), .B(_abc_17692_n4121), .Y(_abc_17692_n4122) );
  AND2X2 AND2X2_1497 ( .A(_abc_17692_n3889), .B(_abc_17692_n3642), .Y(_abc_17692_n4123) );
  AND2X2 AND2X2_1498 ( .A(_abc_17692_n3635), .B(_abc_17692_n4121), .Y(_abc_17692_n4126) );
  AND2X2 AND2X2_1499 ( .A(_abc_17692_n3236), .B(_abc_17692_n4126), .Y(_abc_17692_n4127) );
  AND2X2 AND2X2_15 ( .A(_abc_17692_n632), .B(delta_30_), .Y(delta_30__FF_INPUT) );
  AND2X2 AND2X2_150 ( .A(_abc_17692_n1026), .B(_abc_17692_n1022), .Y(_abc_17692_n1027) );
  AND2X2 AND2X2_1500 ( .A(sum_12_), .B(\key_in[76] ), .Y(_abc_17692_n4129) );
  AND2X2 AND2X2_1501 ( .A(_abc_17692_n4130), .B(_abc_17692_n4131), .Y(_abc_17692_n4132) );
  AND2X2 AND2X2_1502 ( .A(_abc_17692_n4128), .B(_abc_17692_n4132), .Y(_abc_17692_n4133) );
  AND2X2 AND2X2_1503 ( .A(_abc_17692_n4134), .B(_abc_17692_n4135), .Y(_abc_17692_n4136) );
  AND2X2 AND2X2_1504 ( .A(_abc_17692_n4139), .B(_abc_17692_n4140_1), .Y(_abc_17692_n4141) );
  AND2X2 AND2X2_1505 ( .A(_abc_17692_n4142), .B(_abc_17692_n4120), .Y(_abc_17692_n4143_1) );
  AND2X2 AND2X2_1506 ( .A(_abc_17692_n4141), .B(workunit2_12_bF_buf3), .Y(_abc_17692_n4144) );
  AND2X2 AND2X2_1507 ( .A(_abc_17692_n3910), .B(_abc_17692_n3659), .Y(_abc_17692_n4147) );
  AND2X2 AND2X2_1508 ( .A(_abc_17692_n4147), .B(_abc_17692_n3661_1), .Y(_abc_17692_n4148) );
  AND2X2 AND2X2_1509 ( .A(_abc_17692_n3258_1), .B(_abc_17692_n4148), .Y(_abc_17692_n4149) );
  AND2X2 AND2X2_151 ( .A(delta_4_), .B(sum_4_), .Y(_abc_17692_n1029) );
  AND2X2 AND2X2_1510 ( .A(_abc_17692_n4147), .B(_abc_17692_n3666), .Y(_abc_17692_n4150) );
  AND2X2 AND2X2_1511 ( .A(_abc_17692_n3908), .B(workunit2_11_), .Y(_abc_17692_n4151) );
  AND2X2 AND2X2_1512 ( .A(_abc_17692_n3910), .B(_abc_17692_n3656), .Y(_abc_17692_n4152_1) );
  AND2X2 AND2X2_1513 ( .A(_abc_17692_n4155), .B(_abc_17692_n4146), .Y(_abc_17692_n4157) );
  AND2X2 AND2X2_1514 ( .A(_abc_17692_n4158), .B(_abc_17692_n1877_bF_buf9), .Y(_abc_17692_n4159) );
  AND2X2 AND2X2_1515 ( .A(_abc_17692_n4159), .B(_abc_17692_n4156), .Y(_abc_17692_n4160) );
  AND2X2 AND2X2_1516 ( .A(_abc_17692_n3721), .B(_abc_17692_n3955), .Y(_abc_17692_n4161) );
  AND2X2 AND2X2_1517 ( .A(_abc_17692_n4161), .B(_abc_17692_n3716), .Y(_abc_17692_n4162) );
  AND2X2 AND2X2_1518 ( .A(_abc_17692_n3954_1), .B(_abc_17692_n3718), .Y(_abc_17692_n4163) );
  AND2X2 AND2X2_1519 ( .A(_abc_17692_n3713), .B(_abc_17692_n4161), .Y(_abc_17692_n4166) );
  AND2X2 AND2X2_152 ( .A(_abc_17692_n1008), .B(_abc_17692_n1030), .Y(_abc_17692_n1031) );
  AND2X2 AND2X2_1520 ( .A(_abc_17692_n3311), .B(_abc_17692_n4166), .Y(_abc_17692_n4167) );
  AND2X2 AND2X2_1521 ( .A(sum_12_), .B(\key_in[12] ), .Y(_abc_17692_n4169_1) );
  AND2X2 AND2X2_1522 ( .A(_abc_17692_n4170), .B(_abc_17692_n4171), .Y(_abc_17692_n4172) );
  AND2X2 AND2X2_1523 ( .A(_abc_17692_n4168), .B(_abc_17692_n4172), .Y(_abc_17692_n4173) );
  AND2X2 AND2X2_1524 ( .A(_abc_17692_n4174), .B(_abc_17692_n4175), .Y(_abc_17692_n4176) );
  AND2X2 AND2X2_1525 ( .A(_abc_17692_n4179), .B(_abc_17692_n4180), .Y(_abc_17692_n4181) );
  AND2X2 AND2X2_1526 ( .A(_abc_17692_n4181), .B(workunit2_12_bF_buf2), .Y(_abc_17692_n4182) );
  AND2X2 AND2X2_1527 ( .A(_abc_17692_n4183), .B(_abc_17692_n4184), .Y(_abc_17692_n4185) );
  AND2X2 AND2X2_1528 ( .A(_abc_17692_n2898), .B(_abc_17692_n3335), .Y(_abc_17692_n4186_1) );
  AND2X2 AND2X2_1529 ( .A(_abc_17692_n4192), .B(_abc_17692_n4191), .Y(_abc_17692_n4193) );
  AND2X2 AND2X2_153 ( .A(_abc_17692_n1034), .B(state_3_bF_buf4), .Y(_abc_17692_n1035_1) );
  AND2X2 AND2X2_1530 ( .A(_abc_17692_n4194), .B(_abc_17692_n4193), .Y(_abc_17692_n4195) );
  AND2X2 AND2X2_1531 ( .A(_abc_17692_n4190), .B(_abc_17692_n4195), .Y(_abc_17692_n4196) );
  AND2X2 AND2X2_1532 ( .A(_abc_17692_n4197), .B(_abc_17692_n4185), .Y(_abc_17692_n4199) );
  AND2X2 AND2X2_1533 ( .A(_abc_17692_n4200), .B(_abc_17692_n1830_bF_buf9), .Y(_abc_17692_n4201) );
  AND2X2 AND2X2_1534 ( .A(_abc_17692_n4201), .B(_abc_17692_n4198), .Y(_abc_17692_n4202_1) );
  AND2X2 AND2X2_1535 ( .A(_abc_17692_n3683), .B(_abc_17692_n3925), .Y(_abc_17692_n4203) );
  AND2X2 AND2X2_1536 ( .A(_abc_17692_n4203), .B(_abc_17692_n3678), .Y(_abc_17692_n4204) );
  AND2X2 AND2X2_1537 ( .A(_abc_17692_n3924), .B(_abc_17692_n3680), .Y(_abc_17692_n4205) );
  AND2X2 AND2X2_1538 ( .A(_abc_17692_n3675), .B(_abc_17692_n4203), .Y(_abc_17692_n4208) );
  AND2X2 AND2X2_1539 ( .A(_abc_17692_n3278_1), .B(_abc_17692_n4208), .Y(_abc_17692_n4209) );
  AND2X2 AND2X2_154 ( .A(_abc_17692_n1035_1), .B(_abc_17692_n1032), .Y(_abc_17692_n1036) );
  AND2X2 AND2X2_1540 ( .A(sum_12_), .B(\key_in[44] ), .Y(_abc_17692_n4211) );
  AND2X2 AND2X2_1541 ( .A(_abc_17692_n4212), .B(_abc_17692_n4213), .Y(_abc_17692_n4214) );
  AND2X2 AND2X2_1542 ( .A(_abc_17692_n4210), .B(_abc_17692_n4214), .Y(_abc_17692_n4215) );
  AND2X2 AND2X2_1543 ( .A(_abc_17692_n4217), .B(_abc_17692_n4216), .Y(_abc_17692_n4218) );
  AND2X2 AND2X2_1544 ( .A(_abc_17692_n4218), .B(_abc_17692_n4219), .Y(_abc_17692_n4220) );
  AND2X2 AND2X2_1545 ( .A(_abc_17692_n4224), .B(_abc_17692_n4223), .Y(_abc_17692_n4225) );
  AND2X2 AND2X2_1546 ( .A(_abc_17692_n4225), .B(workunit2_12_bF_buf0), .Y(_abc_17692_n4226) );
  AND2X2 AND2X2_1547 ( .A(_abc_17692_n4227), .B(_abc_17692_n4228), .Y(_abc_17692_n4229) );
  AND2X2 AND2X2_1548 ( .A(_abc_17692_n4232), .B(_abc_17692_n4231), .Y(_abc_17692_n4233) );
  AND2X2 AND2X2_1549 ( .A(_abc_17692_n4230), .B(_abc_17692_n4233), .Y(_abc_17692_n4234) );
  AND2X2 AND2X2_155 ( .A(_abc_17692_n1037), .B(_abc_17692_n1028_1), .Y(_abc_17692_n1039) );
  AND2X2 AND2X2_1550 ( .A(_abc_17692_n4233), .B(_abc_17692_n3705), .Y(_abc_17692_n4235) );
  AND2X2 AND2X2_1551 ( .A(_abc_17692_n3701), .B(_abc_17692_n4235), .Y(_abc_17692_n4236) );
  AND2X2 AND2X2_1552 ( .A(_abc_17692_n4238), .B(_abc_17692_n4229), .Y(_abc_17692_n4240) );
  AND2X2 AND2X2_1553 ( .A(_abc_17692_n4241), .B(_abc_17692_n1846_bF_buf9), .Y(_abc_17692_n4242) );
  AND2X2 AND2X2_1554 ( .A(_abc_17692_n4242), .B(_abc_17692_n4239), .Y(_abc_17692_n4243) );
  AND2X2 AND2X2_1555 ( .A(_abc_17692_n4246), .B(state_6_bF_buf2), .Y(_abc_17692_n4247) );
  AND2X2 AND2X2_1556 ( .A(_abc_17692_n4247), .B(_abc_17692_n4119), .Y(_abc_17692_n4248) );
  AND2X2 AND2X2_1557 ( .A(_abc_17692_n4001), .B(_abc_17692_n3775), .Y(_abc_17692_n4250_1) );
  AND2X2 AND2X2_1558 ( .A(_abc_17692_n4250_1), .B(_abc_17692_n3793), .Y(_abc_17692_n4251) );
  AND2X2 AND2X2_1559 ( .A(_abc_17692_n3386), .B(_abc_17692_n4251), .Y(_abc_17692_n4252) );
  AND2X2 AND2X2_156 ( .A(_abc_17692_n1040), .B(state_15_bF_buf4), .Y(_abc_17692_n1041) );
  AND2X2 AND2X2_1560 ( .A(_abc_17692_n4250_1), .B(_abc_17692_n3798), .Y(_abc_17692_n4253_1) );
  AND2X2 AND2X2_1561 ( .A(_abc_17692_n3999), .B(workunit2_11_), .Y(_abc_17692_n4254) );
  AND2X2 AND2X2_1562 ( .A(_abc_17692_n4001), .B(_abc_17692_n4255), .Y(_abc_17692_n4256) );
  AND2X2 AND2X2_1563 ( .A(_abc_17692_n4259), .B(_abc_17692_n4249), .Y(_abc_17692_n4261) );
  AND2X2 AND2X2_1564 ( .A(_abc_17692_n4262), .B(_abc_17692_n1863_bF_buf7), .Y(_abc_17692_n4263) );
  AND2X2 AND2X2_1565 ( .A(_abc_17692_n4263), .B(_abc_17692_n4260), .Y(_abc_17692_n4264) );
  AND2X2 AND2X2_1566 ( .A(_abc_17692_n3187), .B(_abc_17692_n3395), .Y(_abc_17692_n4265) );
  AND2X2 AND2X2_1567 ( .A(_abc_17692_n4270), .B(_abc_17692_n4269_1), .Y(_abc_17692_n4271) );
  AND2X2 AND2X2_1568 ( .A(_abc_17692_n4272), .B(_abc_17692_n4271), .Y(_abc_17692_n4273) );
  AND2X2 AND2X2_1569 ( .A(_abc_17692_n4268), .B(_abc_17692_n4273), .Y(_abc_17692_n4274) );
  AND2X2 AND2X2_157 ( .A(_abc_17692_n1041), .B(_abc_17692_n1038), .Y(_abc_17692_n1042) );
  AND2X2 AND2X2_1570 ( .A(_abc_17692_n4275), .B(_abc_17692_n4145), .Y(_abc_17692_n4277) );
  AND2X2 AND2X2_1571 ( .A(_abc_17692_n4278), .B(_abc_17692_n1877_bF_buf8), .Y(_abc_17692_n4279_1) );
  AND2X2 AND2X2_1572 ( .A(_abc_17692_n4279_1), .B(_abc_17692_n4276), .Y(_abc_17692_n4280) );
  AND2X2 AND2X2_1573 ( .A(_abc_17692_n3942), .B(_abc_17692_n3698), .Y(_abc_17692_n4282) );
  AND2X2 AND2X2_1574 ( .A(_abc_17692_n4282), .B(_abc_17692_n3826), .Y(_abc_17692_n4283) );
  AND2X2 AND2X2_1575 ( .A(_abc_17692_n4283), .B(_abc_17692_n3410), .Y(_abc_17692_n4284) );
  AND2X2 AND2X2_1576 ( .A(_abc_17692_n4282), .B(_abc_17692_n3831), .Y(_abc_17692_n4285) );
  AND2X2 AND2X2_1577 ( .A(_abc_17692_n3940), .B(workunit2_11_), .Y(_abc_17692_n4286) );
  AND2X2 AND2X2_1578 ( .A(_abc_17692_n3942), .B(_abc_17692_n3695), .Y(_abc_17692_n4287) );
  AND2X2 AND2X2_1579 ( .A(_abc_17692_n4290), .B(_abc_17692_n4281), .Y(_abc_17692_n4292) );
  AND2X2 AND2X2_158 ( .A(_abc_17692_n722_bF_buf2), .B(sum_5_), .Y(_abc_17692_n1043) );
  AND2X2 AND2X2_1580 ( .A(_abc_17692_n4293), .B(_abc_17692_n1846_bF_buf8), .Y(_abc_17692_n4294) );
  AND2X2 AND2X2_1581 ( .A(_abc_17692_n4294), .B(_abc_17692_n4291), .Y(_abc_17692_n4295) );
  AND2X2 AND2X2_1582 ( .A(_abc_17692_n3969), .B(_abc_17692_n3840), .Y(_abc_17692_n4297) );
  AND2X2 AND2X2_1583 ( .A(_abc_17692_n4297), .B(_abc_17692_n3842), .Y(_abc_17692_n4298) );
  AND2X2 AND2X2_1584 ( .A(_abc_17692_n4298), .B(_abc_17692_n3422), .Y(_abc_17692_n4299) );
  AND2X2 AND2X2_1585 ( .A(_abc_17692_n4297), .B(_abc_17692_n3847), .Y(_abc_17692_n4300) );
  AND2X2 AND2X2_1586 ( .A(_abc_17692_n3967), .B(workunit2_11_), .Y(_abc_17692_n4301) );
  AND2X2 AND2X2_1587 ( .A(_abc_17692_n3969), .B(_abc_17692_n4302), .Y(_abc_17692_n4303) );
  AND2X2 AND2X2_1588 ( .A(_abc_17692_n4306), .B(_abc_17692_n4296), .Y(_abc_17692_n4307) );
  AND2X2 AND2X2_1589 ( .A(_abc_17692_n4309), .B(_abc_17692_n1830_bF_buf8), .Y(_abc_17692_n4310) );
  AND2X2 AND2X2_159 ( .A(_abc_17692_n1047), .B(delta_6_), .Y(_abc_17692_n1048) );
  AND2X2 AND2X2_1590 ( .A(_abc_17692_n4310), .B(_abc_17692_n4308), .Y(_abc_17692_n4311) );
  AND2X2 AND2X2_1591 ( .A(_abc_17692_n4314), .B(state_7_bF_buf1), .Y(_abc_17692_n4315) );
  AND2X2 AND2X2_1592 ( .A(_abc_17692_n1885_bF_buf2), .B(workunit2_12_bF_buf2), .Y(_abc_17692_n4316) );
  AND2X2 AND2X2_1593 ( .A(state_8_bF_buf7), .B(\data_in2[12] ), .Y(_abc_17692_n4317_1) );
  AND2X2 AND2X2_1594 ( .A(_abc_17692_n4322), .B(workunit1_9_), .Y(_abc_17692_n4323) );
  AND2X2 AND2X2_1595 ( .A(_abc_17692_n2435), .B(workunit1_18_), .Y(_abc_17692_n4324) );
  AND2X2 AND2X2_1596 ( .A(_abc_17692_n4325), .B(workunit1_13_bF_buf3), .Y(_abc_17692_n4326) );
  AND2X2 AND2X2_1597 ( .A(_abc_17692_n4321), .B(_abc_17692_n4329), .Y(_abc_17692_n4330) );
  AND2X2 AND2X2_1598 ( .A(_abc_17692_n4331), .B(_abc_17692_n4332), .Y(_abc_17692_n4333) );
  AND2X2 AND2X2_1599 ( .A(sum_13_), .B(\key_in[77] ), .Y(_abc_17692_n4337) );
  AND2X2 AND2X2_16 ( .A(_abc_17692_n629), .B(x_0_), .Y(_abc_17692_n667) );
  AND2X2 AND2X2_160 ( .A(_abc_17692_n1023), .B(sum_5_), .Y(_abc_17692_n1053) );
  AND2X2 AND2X2_1600 ( .A(_abc_17692_n4338), .B(_abc_17692_n4339), .Y(_abc_17692_n4340) );
  AND2X2 AND2X2_1601 ( .A(_abc_17692_n4336), .B(_abc_17692_n4340), .Y(_abc_17692_n4341) );
  AND2X2 AND2X2_1602 ( .A(_abc_17692_n4335), .B(_abc_17692_n4342), .Y(_abc_17692_n4343) );
  AND2X2 AND2X2_1603 ( .A(_abc_17692_n4334), .B(_abc_17692_n4344_1), .Y(_abc_17692_n4345) );
  AND2X2 AND2X2_1604 ( .A(_abc_17692_n4346), .B(_abc_17692_n4333), .Y(_abc_17692_n4347_1) );
  AND2X2 AND2X2_1605 ( .A(_abc_17692_n4349), .B(workunit2_13_), .Y(_abc_17692_n4350) );
  AND2X2 AND2X2_1606 ( .A(_abc_17692_n4348), .B(_abc_17692_n4351), .Y(_abc_17692_n4352) );
  AND2X2 AND2X2_1607 ( .A(_abc_17692_n4158), .B(_abc_17692_n4355), .Y(_abc_17692_n4356) );
  AND2X2 AND2X2_1608 ( .A(_abc_17692_n4359), .B(_abc_17692_n1877_bF_buf7), .Y(_abc_17692_n4360) );
  AND2X2 AND2X2_1609 ( .A(_abc_17692_n4360), .B(_abc_17692_n4357), .Y(_abc_17692_n4361) );
  AND2X2 AND2X2_161 ( .A(_abc_17692_n1054), .B(_abc_17692_n1052), .Y(_abc_17692_n1056) );
  AND2X2 AND2X2_1610 ( .A(sum_13_), .B(\key_in[45] ), .Y(_abc_17692_n4364) );
  AND2X2 AND2X2_1611 ( .A(_abc_17692_n4365), .B(_abc_17692_n4366), .Y(_abc_17692_n4367) );
  AND2X2 AND2X2_1612 ( .A(_abc_17692_n4363), .B(_abc_17692_n4367), .Y(_abc_17692_n4368) );
  AND2X2 AND2X2_1613 ( .A(_abc_17692_n4373), .B(_abc_17692_n4369), .Y(_abc_17692_n4374) );
  AND2X2 AND2X2_1614 ( .A(_abc_17692_n4372), .B(_abc_17692_n4375), .Y(_abc_17692_n4376) );
  AND2X2 AND2X2_1615 ( .A(_abc_17692_n4379), .B(_abc_17692_n4378), .Y(_abc_17692_n4380) );
  AND2X2 AND2X2_1616 ( .A(_abc_17692_n4381), .B(_abc_17692_n4377), .Y(_abc_17692_n4382) );
  AND2X2 AND2X2_1617 ( .A(_abc_17692_n4241), .B(_abc_17692_n4227), .Y(_abc_17692_n4384) );
  AND2X2 AND2X2_1618 ( .A(_abc_17692_n4387), .B(_abc_17692_n1846_bF_buf7), .Y(_abc_17692_n4388) );
  AND2X2 AND2X2_1619 ( .A(_abc_17692_n4388), .B(_abc_17692_n4386), .Y(_abc_17692_n4389_1) );
  AND2X2 AND2X2_162 ( .A(_abc_17692_n1057_1), .B(state_15_bF_buf3), .Y(_abc_17692_n1058) );
  AND2X2 AND2X2_1620 ( .A(sum_13_), .B(\key_in[13] ), .Y(_abc_17692_n4391) );
  AND2X2 AND2X2_1621 ( .A(_abc_17692_n4392_1), .B(_abc_17692_n4393), .Y(_abc_17692_n4394) );
  AND2X2 AND2X2_1622 ( .A(_abc_17692_n4390), .B(_abc_17692_n4395), .Y(_abc_17692_n4397) );
  AND2X2 AND2X2_1623 ( .A(_abc_17692_n4398), .B(_abc_17692_n4396), .Y(_abc_17692_n4399) );
  AND2X2 AND2X2_1624 ( .A(_abc_17692_n4402), .B(_abc_17692_n4400), .Y(_abc_17692_n4403) );
  AND2X2 AND2X2_1625 ( .A(_abc_17692_n4405), .B(_abc_17692_n4406), .Y(_abc_17692_n4407) );
  AND2X2 AND2X2_1626 ( .A(_abc_17692_n4200), .B(_abc_17692_n4183), .Y(_abc_17692_n4409) );
  AND2X2 AND2X2_1627 ( .A(_abc_17692_n4412), .B(_abc_17692_n1830_bF_buf7), .Y(_abc_17692_n4413) );
  AND2X2 AND2X2_1628 ( .A(_abc_17692_n4413), .B(_abc_17692_n4411), .Y(_abc_17692_n4414) );
  AND2X2 AND2X2_1629 ( .A(sum_13_), .B(\key_in[109] ), .Y(_abc_17692_n4418) );
  AND2X2 AND2X2_163 ( .A(_abc_17692_n1058), .B(_abc_17692_n1055), .Y(_abc_17692_n1059) );
  AND2X2 AND2X2_1630 ( .A(_abc_17692_n4419), .B(_abc_17692_n4420), .Y(_abc_17692_n4421) );
  AND2X2 AND2X2_1631 ( .A(_abc_17692_n4417), .B(_abc_17692_n4422), .Y(_abc_17692_n4424) );
  AND2X2 AND2X2_1632 ( .A(_abc_17692_n4425), .B(_abc_17692_n4423), .Y(_abc_17692_n4426) );
  AND2X2 AND2X2_1633 ( .A(_abc_17692_n4429), .B(_abc_17692_n4427), .Y(_abc_17692_n4430) );
  AND2X2 AND2X2_1634 ( .A(_abc_17692_n4432), .B(_abc_17692_n4433), .Y(_abc_17692_n4434) );
  AND2X2 AND2X2_1635 ( .A(_abc_17692_n4116), .B(_abc_17692_n4100), .Y(_abc_17692_n4436) );
  AND2X2 AND2X2_1636 ( .A(_abc_17692_n4439), .B(_abc_17692_n1863_bF_buf6), .Y(_abc_17692_n4440) );
  AND2X2 AND2X2_1637 ( .A(_abc_17692_n4440), .B(_abc_17692_n4438), .Y(_abc_17692_n4441) );
  AND2X2 AND2X2_1638 ( .A(_abc_17692_n4442), .B(state_6_bF_buf1), .Y(_abc_17692_n4443) );
  AND2X2 AND2X2_1639 ( .A(_abc_17692_n4444_1), .B(workunit2_12_bF_buf1), .Y(_abc_17692_n4445) );
  AND2X2 AND2X2_164 ( .A(_abc_17692_n723), .B(sum_6_), .Y(_abc_17692_n1060) );
  AND2X2 AND2X2_1640 ( .A(_abc_17692_n4262), .B(_abc_17692_n4446), .Y(_abc_17692_n4447_1) );
  AND2X2 AND2X2_1641 ( .A(_abc_17692_n4450), .B(_abc_17692_n1863_bF_buf5), .Y(_abc_17692_n4451) );
  AND2X2 AND2X2_1642 ( .A(_abc_17692_n4451), .B(_abc_17692_n4448), .Y(_abc_17692_n4452) );
  AND2X2 AND2X2_1643 ( .A(_abc_17692_n4142), .B(workunit2_12_bF_buf0), .Y(_abc_17692_n4453) );
  AND2X2 AND2X2_1644 ( .A(_abc_17692_n4278), .B(_abc_17692_n4454), .Y(_abc_17692_n4455) );
  AND2X2 AND2X2_1645 ( .A(_abc_17692_n4456), .B(_abc_17692_n4353), .Y(_abc_17692_n4457) );
  AND2X2 AND2X2_1646 ( .A(_abc_17692_n4455), .B(_abc_17692_n4354), .Y(_abc_17692_n4458) );
  AND2X2 AND2X2_1647 ( .A(_abc_17692_n4459), .B(_abc_17692_n1877_bF_buf6), .Y(_abc_17692_n4460) );
  AND2X2 AND2X2_1648 ( .A(_abc_17692_n4461), .B(workunit2_12_bF_buf3), .Y(_abc_17692_n4462) );
  AND2X2 AND2X2_1649 ( .A(_abc_17692_n4293), .B(_abc_17692_n4463), .Y(_abc_17692_n4464) );
  AND2X2 AND2X2_165 ( .A(_abc_17692_n1061), .B(_abc_17692_n1022), .Y(_abc_17692_n1062) );
  AND2X2 AND2X2_1650 ( .A(_abc_17692_n4467), .B(_abc_17692_n1846_bF_buf6), .Y(_abc_17692_n4468) );
  AND2X2 AND2X2_1651 ( .A(_abc_17692_n4468), .B(_abc_17692_n4466), .Y(_abc_17692_n4469) );
  AND2X2 AND2X2_1652 ( .A(_abc_17692_n4470), .B(workunit2_12_bF_buf2), .Y(_abc_17692_n4471) );
  AND2X2 AND2X2_1653 ( .A(_abc_17692_n4308), .B(_abc_17692_n4472), .Y(_abc_17692_n4473) );
  AND2X2 AND2X2_1654 ( .A(_abc_17692_n4476), .B(_abc_17692_n1830_bF_buf6), .Y(_abc_17692_n4477) );
  AND2X2 AND2X2_1655 ( .A(_abc_17692_n4477), .B(_abc_17692_n4474), .Y(_abc_17692_n4478) );
  AND2X2 AND2X2_1656 ( .A(_abc_17692_n4481), .B(state_7_bF_buf0), .Y(_abc_17692_n4482) );
  AND2X2 AND2X2_1657 ( .A(_abc_17692_n1885_bF_buf1), .B(workunit2_13_), .Y(_abc_17692_n4483) );
  AND2X2 AND2X2_1658 ( .A(state_8_bF_buf6), .B(\data_in2[13] ), .Y(_abc_17692_n4484) );
  AND2X2 AND2X2_1659 ( .A(_abc_17692_n4488), .B(_abc_17692_n4066), .Y(_abc_17692_n4489) );
  AND2X2 AND2X2_166 ( .A(_abc_17692_n1065), .B(state_3_bF_buf3), .Y(_abc_17692_n1066) );
  AND2X2 AND2X2_1660 ( .A(_abc_17692_n4058), .B(_abc_17692_n4489), .Y(_abc_17692_n4490) );
  AND2X2 AND2X2_1661 ( .A(_abc_17692_n4491), .B(_abc_17692_n4327), .Y(_abc_17692_n4492) );
  AND2X2 AND2X2_1662 ( .A(_abc_17692_n4494), .B(workunit1_10_), .Y(_abc_17692_n4495) );
  AND2X2 AND2X2_1663 ( .A(_abc_17692_n2638), .B(workunit1_19_), .Y(_abc_17692_n4496) );
  AND2X2 AND2X2_1664 ( .A(_abc_17692_n4497), .B(workunit1_14_bF_buf0), .Y(_abc_17692_n4498) );
  AND2X2 AND2X2_1665 ( .A(_abc_17692_n4499), .B(_abc_17692_n4500), .Y(_abc_17692_n4501) );
  AND2X2 AND2X2_1666 ( .A(_abc_17692_n4493), .B(_abc_17692_n4501), .Y(_abc_17692_n4502) );
  AND2X2 AND2X2_1667 ( .A(_abc_17692_n4504), .B(_abc_17692_n4505), .Y(_abc_17692_n4506) );
  AND2X2 AND2X2_1668 ( .A(_abc_17692_n4506), .B(_abc_17692_n4508), .Y(_abc_17692_n4509) );
  AND2X2 AND2X2_1669 ( .A(_abc_17692_n4086), .B(_abc_17692_n4421), .Y(_abc_17692_n4511) );
  AND2X2 AND2X2_167 ( .A(_abc_17692_n1066), .B(_abc_17692_n1063), .Y(_abc_17692_n1067) );
  AND2X2 AND2X2_1670 ( .A(_abc_17692_n4082), .B(_abc_17692_n4511), .Y(_abc_17692_n4512) );
  AND2X2 AND2X2_1671 ( .A(_abc_17692_n4084_1), .B(_abc_17692_n4419), .Y(_abc_17692_n4514) );
  AND2X2 AND2X2_1672 ( .A(sum_14_), .B(\key_in[110] ), .Y(_abc_17692_n4518) );
  AND2X2 AND2X2_1673 ( .A(_abc_17692_n4519), .B(_abc_17692_n4520), .Y(_abc_17692_n4521) );
  AND2X2 AND2X2_1674 ( .A(_abc_17692_n4517), .B(_abc_17692_n4521), .Y(_abc_17692_n4522) );
  AND2X2 AND2X2_1675 ( .A(_abc_17692_n4523), .B(_abc_17692_n4515), .Y(_abc_17692_n4524) );
  AND2X2 AND2X2_1676 ( .A(_abc_17692_n4524), .B(_abc_17692_n4525), .Y(_abc_17692_n4526) );
  AND2X2 AND2X2_1677 ( .A(_abc_17692_n4529), .B(_abc_17692_n4531), .Y(_abc_17692_n4532) );
  AND2X2 AND2X2_1678 ( .A(_abc_17692_n4532), .B(workunit2_14_bF_buf1), .Y(_abc_17692_n4534) );
  AND2X2 AND2X2_1679 ( .A(_abc_17692_n4535), .B(_abc_17692_n4533), .Y(_abc_17692_n4536) );
  AND2X2 AND2X2_168 ( .A(_abc_17692_n1070), .B(delta_7_), .Y(_abc_17692_n1071) );
  AND2X2 AND2X2_1680 ( .A(_abc_17692_n4431), .B(workunit2_13_), .Y(_abc_17692_n4537) );
  AND2X2 AND2X2_1681 ( .A(_abc_17692_n4539), .B(_abc_17692_n4538), .Y(_abc_17692_n4540) );
  AND2X2 AND2X2_1682 ( .A(_abc_17692_n4435), .B(_abc_17692_n4102), .Y(_abc_17692_n4542) );
  AND2X2 AND2X2_1683 ( .A(_abc_17692_n4114), .B(_abc_17692_n4542), .Y(_abc_17692_n4543) );
  AND2X2 AND2X2_1684 ( .A(_abc_17692_n4544), .B(_abc_17692_n4536), .Y(_abc_17692_n4546) );
  AND2X2 AND2X2_1685 ( .A(_abc_17692_n4547), .B(_abc_17692_n4545), .Y(_abc_17692_n4548) );
  AND2X2 AND2X2_1686 ( .A(_abc_17692_n4132), .B(_abc_17692_n4340), .Y(_abc_17692_n4550) );
  AND2X2 AND2X2_1687 ( .A(_abc_17692_n4128), .B(_abc_17692_n4550), .Y(_abc_17692_n4551) );
  AND2X2 AND2X2_1688 ( .A(_abc_17692_n4130), .B(_abc_17692_n4338), .Y(_abc_17692_n4553) );
  AND2X2 AND2X2_1689 ( .A(sum_14_), .B(\key_in[78] ), .Y(_abc_17692_n4557) );
  AND2X2 AND2X2_169 ( .A(delta_6_), .B(sum_6_), .Y(_abc_17692_n1076) );
  AND2X2 AND2X2_1690 ( .A(_abc_17692_n4558), .B(_abc_17692_n4559), .Y(_abc_17692_n4560) );
  AND2X2 AND2X2_1691 ( .A(_abc_17692_n4556), .B(_abc_17692_n4560), .Y(_abc_17692_n4561) );
  AND2X2 AND2X2_1692 ( .A(_abc_17692_n4562), .B(_abc_17692_n4563), .Y(_abc_17692_n4564) );
  AND2X2 AND2X2_1693 ( .A(_abc_17692_n4567), .B(_abc_17692_n4568), .Y(_abc_17692_n4569) );
  AND2X2 AND2X2_1694 ( .A(_abc_17692_n4569), .B(workunit2_14_bF_buf0), .Y(_abc_17692_n4570) );
  AND2X2 AND2X2_1695 ( .A(_abc_17692_n4571), .B(_abc_17692_n4572), .Y(_abc_17692_n4573) );
  AND2X2 AND2X2_1696 ( .A(_abc_17692_n4348), .B(workunit2_13_), .Y(_abc_17692_n4574) );
  AND2X2 AND2X2_1697 ( .A(_abc_17692_n4353), .B(_abc_17692_n4144), .Y(_abc_17692_n4575) );
  AND2X2 AND2X2_1698 ( .A(_abc_17692_n4353), .B(_abc_17692_n4146), .Y(_abc_17692_n4577) );
  AND2X2 AND2X2_1699 ( .A(_abc_17692_n4155), .B(_abc_17692_n4577), .Y(_abc_17692_n4578) );
  AND2X2 AND2X2_17 ( .A(_abc_17692_n668), .B(_abc_17692_n669), .Y(x_0__FF_INPUT) );
  AND2X2 AND2X2_170 ( .A(_abc_17692_n1063), .B(_abc_17692_n1077), .Y(_abc_17692_n1078) );
  AND2X2 AND2X2_1700 ( .A(_abc_17692_n4579), .B(_abc_17692_n4573), .Y(_abc_17692_n4580) );
  AND2X2 AND2X2_1701 ( .A(_abc_17692_n4582), .B(_abc_17692_n1877_bF_buf5), .Y(_abc_17692_n4583) );
  AND2X2 AND2X2_1702 ( .A(_abc_17692_n4583), .B(_abc_17692_n4581), .Y(_abc_17692_n4584_1) );
  AND2X2 AND2X2_1703 ( .A(_abc_17692_n4172), .B(_abc_17692_n4394), .Y(_abc_17692_n4585) );
  AND2X2 AND2X2_1704 ( .A(_abc_17692_n4168), .B(_abc_17692_n4585), .Y(_abc_17692_n4586) );
  AND2X2 AND2X2_1705 ( .A(_abc_17692_n4170), .B(_abc_17692_n4392_1), .Y(_abc_17692_n4588) );
  AND2X2 AND2X2_1706 ( .A(sum_14_), .B(\key_in[14] ), .Y(_abc_17692_n4592) );
  AND2X2 AND2X2_1707 ( .A(_abc_17692_n4593), .B(_abc_17692_n4594), .Y(_abc_17692_n4595) );
  AND2X2 AND2X2_1708 ( .A(_abc_17692_n4591), .B(_abc_17692_n4595), .Y(_abc_17692_n4596) );
  AND2X2 AND2X2_1709 ( .A(_abc_17692_n4597), .B(_abc_17692_n4598), .Y(_abc_17692_n4599) );
  AND2X2 AND2X2_171 ( .A(_abc_17692_n1081), .B(state_3_bF_buf2), .Y(_abc_17692_n1082) );
  AND2X2 AND2X2_1710 ( .A(_abc_17692_n4602), .B(_abc_17692_n4603), .Y(_abc_17692_n4604) );
  AND2X2 AND2X2_1711 ( .A(_abc_17692_n4604), .B(workunit2_14_bF_buf1), .Y(_abc_17692_n4606) );
  AND2X2 AND2X2_1712 ( .A(_abc_17692_n4607), .B(_abc_17692_n4605), .Y(_abc_17692_n4608) );
  AND2X2 AND2X2_1713 ( .A(_abc_17692_n4404), .B(workunit2_13_), .Y(_abc_17692_n4609) );
  AND2X2 AND2X2_1714 ( .A(_abc_17692_n4611), .B(_abc_17692_n4610), .Y(_abc_17692_n4612) );
  AND2X2 AND2X2_1715 ( .A(_abc_17692_n4197), .B(_abc_17692_n4615), .Y(_abc_17692_n4616) );
  AND2X2 AND2X2_1716 ( .A(_abc_17692_n4617), .B(_abc_17692_n4608), .Y(_abc_17692_n4618) );
  AND2X2 AND2X2_1717 ( .A(_abc_17692_n4620), .B(_abc_17692_n1830_bF_buf5), .Y(_abc_17692_n4621) );
  AND2X2 AND2X2_1718 ( .A(_abc_17692_n4621), .B(_abc_17692_n4619), .Y(_abc_17692_n4622) );
  AND2X2 AND2X2_1719 ( .A(_abc_17692_n4214), .B(_abc_17692_n4367), .Y(_abc_17692_n4624) );
  AND2X2 AND2X2_172 ( .A(_abc_17692_n1082), .B(_abc_17692_n1079), .Y(_abc_17692_n1083) );
  AND2X2 AND2X2_1720 ( .A(_abc_17692_n4210), .B(_abc_17692_n4624), .Y(_abc_17692_n4625) );
  AND2X2 AND2X2_1721 ( .A(_abc_17692_n4212), .B(_abc_17692_n4365), .Y(_abc_17692_n4627) );
  AND2X2 AND2X2_1722 ( .A(sum_14_), .B(\key_in[46] ), .Y(_abc_17692_n4631) );
  AND2X2 AND2X2_1723 ( .A(_abc_17692_n4632), .B(_abc_17692_n4633), .Y(_abc_17692_n4634) );
  AND2X2 AND2X2_1724 ( .A(_abc_17692_n4630), .B(_abc_17692_n4634), .Y(_abc_17692_n4635) );
  AND2X2 AND2X2_1725 ( .A(_abc_17692_n4636), .B(_abc_17692_n4628), .Y(_abc_17692_n4637) );
  AND2X2 AND2X2_1726 ( .A(_abc_17692_n4637), .B(_abc_17692_n4638), .Y(_abc_17692_n4639) );
  AND2X2 AND2X2_1727 ( .A(_abc_17692_n4530), .B(_abc_17692_n4640), .Y(_abc_17692_n4641) );
  AND2X2 AND2X2_1728 ( .A(_abc_17692_n4642), .B(_abc_17692_n4510_1), .Y(_abc_17692_n4643_1) );
  AND2X2 AND2X2_1729 ( .A(_abc_17692_n4646_1), .B(_abc_17692_n4647), .Y(_abc_17692_n4648) );
  AND2X2 AND2X2_173 ( .A(_abc_17692_n723), .B(sum_7_), .Y(_abc_17692_n1084) );
  AND2X2 AND2X2_1730 ( .A(_abc_17692_n4376), .B(workunit2_13_), .Y(_abc_17692_n4650) );
  AND2X2 AND2X2_1731 ( .A(_abc_17692_n4652), .B(_abc_17692_n4651), .Y(_abc_17692_n4653) );
  AND2X2 AND2X2_1732 ( .A(_abc_17692_n4238), .B(_abc_17692_n4656), .Y(_abc_17692_n4657) );
  AND2X2 AND2X2_1733 ( .A(_abc_17692_n4658), .B(_abc_17692_n4649), .Y(_abc_17692_n4659) );
  AND2X2 AND2X2_1734 ( .A(_abc_17692_n4661), .B(_abc_17692_n1846_bF_buf5), .Y(_abc_17692_n4662) );
  AND2X2 AND2X2_1735 ( .A(_abc_17692_n4662), .B(_abc_17692_n4660), .Y(_abc_17692_n4663) );
  AND2X2 AND2X2_1736 ( .A(_abc_17692_n4666), .B(state_6_bF_buf0), .Y(_abc_17692_n4667) );
  AND2X2 AND2X2_1737 ( .A(_abc_17692_n4667), .B(_abc_17692_n4549), .Y(_abc_17692_n4668) );
  AND2X2 AND2X2_1738 ( .A(_abc_17692_n4433), .B(_abc_17692_n4445), .Y(_abc_17692_n4671) );
  AND2X2 AND2X2_1739 ( .A(_abc_17692_n4434), .B(_abc_17692_n4249), .Y(_abc_17692_n4673) );
  AND2X2 AND2X2_174 ( .A(_abc_17692_n1056), .B(_abc_17692_n1075), .Y(_abc_17692_n1087) );
  AND2X2 AND2X2_1740 ( .A(_abc_17692_n4259), .B(_abc_17692_n4673), .Y(_abc_17692_n4674) );
  AND2X2 AND2X2_1741 ( .A(_abc_17692_n4675), .B(_abc_17692_n4669), .Y(_abc_17692_n4676) );
  AND2X2 AND2X2_1742 ( .A(_abc_17692_n4678), .B(_abc_17692_n1863_bF_buf3), .Y(_abc_17692_n4679) );
  AND2X2 AND2X2_1743 ( .A(_abc_17692_n4679), .B(_abc_17692_n4677), .Y(_abc_17692_n4680) );
  AND2X2 AND2X2_1744 ( .A(_abc_17692_n4682), .B(_abc_17692_n4683), .Y(_abc_17692_n4684) );
  AND2X2 AND2X2_1745 ( .A(_abc_17692_n4275), .B(_abc_17692_n4687), .Y(_abc_17692_n4688) );
  AND2X2 AND2X2_1746 ( .A(_abc_17692_n4689), .B(_abc_17692_n4681), .Y(_abc_17692_n4690) );
  AND2X2 AND2X2_1747 ( .A(_abc_17692_n4692), .B(_abc_17692_n1877_bF_buf4), .Y(_abc_17692_n4693) );
  AND2X2 AND2X2_1748 ( .A(_abc_17692_n4693), .B(_abc_17692_n4691), .Y(_abc_17692_n4694) );
  AND2X2 AND2X2_1749 ( .A(_abc_17692_n4377), .B(_abc_17692_n4463), .Y(_abc_17692_n4696) );
  AND2X2 AND2X2_175 ( .A(_abc_17692_n1075), .B(_abc_17692_n1050), .Y(_abc_17692_n1089) );
  AND2X2 AND2X2_1750 ( .A(_abc_17692_n4382), .B(_abc_17692_n4281), .Y(_abc_17692_n4699) );
  AND2X2 AND2X2_1751 ( .A(_abc_17692_n4290), .B(_abc_17692_n4699), .Y(_abc_17692_n4700) );
  AND2X2 AND2X2_1752 ( .A(_abc_17692_n4701), .B(_abc_17692_n4648), .Y(_abc_17692_n4702) );
  AND2X2 AND2X2_1753 ( .A(_abc_17692_n4704), .B(_abc_17692_n1846_bF_buf4), .Y(_abc_17692_n4705) );
  AND2X2 AND2X2_1754 ( .A(_abc_17692_n4705), .B(_abc_17692_n4703), .Y(_abc_17692_n4706) );
  AND2X2 AND2X2_1755 ( .A(_abc_17692_n4405), .B(_abc_17692_n4472), .Y(_abc_17692_n4709) );
  AND2X2 AND2X2_1756 ( .A(_abc_17692_n4407), .B(_abc_17692_n4296), .Y(_abc_17692_n4712) );
  AND2X2 AND2X2_1757 ( .A(_abc_17692_n4306), .B(_abc_17692_n4712), .Y(_abc_17692_n4713) );
  AND2X2 AND2X2_1758 ( .A(_abc_17692_n4714), .B(_abc_17692_n4707), .Y(_abc_17692_n4715) );
  AND2X2 AND2X2_1759 ( .A(_abc_17692_n4717), .B(_abc_17692_n1830_bF_buf4), .Y(_abc_17692_n4718) );
  AND2X2 AND2X2_176 ( .A(_abc_17692_n1090), .B(state_15_bF_buf2), .Y(_abc_17692_n1091) );
  AND2X2 AND2X2_1760 ( .A(_abc_17692_n4718), .B(_abc_17692_n4716), .Y(_abc_17692_n4719) );
  AND2X2 AND2X2_1761 ( .A(_abc_17692_n4722), .B(state_7_bF_buf4), .Y(_abc_17692_n4723) );
  AND2X2 AND2X2_1762 ( .A(_abc_17692_n1885_bF_buf0), .B(workunit2_14_bF_buf2), .Y(_abc_17692_n4724) );
  AND2X2 AND2X2_1763 ( .A(state_8_bF_buf5), .B(\data_in2[14] ), .Y(_abc_17692_n4725) );
  AND2X2 AND2X2_1764 ( .A(_abc_17692_n4730), .B(workunit1_11_bF_buf1), .Y(_abc_17692_n4731) );
  AND2X2 AND2X2_1765 ( .A(_abc_17692_n2823), .B(workunit1_20_), .Y(_abc_17692_n4732) );
  AND2X2 AND2X2_1766 ( .A(_abc_17692_n4733), .B(workunit1_15_), .Y(_abc_17692_n4734) );
  AND2X2 AND2X2_1767 ( .A(_abc_17692_n4739), .B(_abc_17692_n4499), .Y(_abc_17692_n4740) );
  AND2X2 AND2X2_1768 ( .A(_abc_17692_n4741), .B(_abc_17692_n4735_1), .Y(_abc_17692_n4742) );
  AND2X2 AND2X2_1769 ( .A(_abc_17692_n4743), .B(_abc_17692_n4738_1), .Y(_abc_17692_n4744) );
  AND2X2 AND2X2_177 ( .A(_abc_17692_n1088), .B(_abc_17692_n1091), .Y(_abc_17692_n1092) );
  AND2X2 AND2X2_1770 ( .A(sum_15_), .B(\key_in[79] ), .Y(_abc_17692_n4747) );
  AND2X2 AND2X2_1771 ( .A(_abc_17692_n4748), .B(_abc_17692_n4749), .Y(_abc_17692_n4750) );
  AND2X2 AND2X2_1772 ( .A(_abc_17692_n4746), .B(_abc_17692_n4750), .Y(_abc_17692_n4751) );
  AND2X2 AND2X2_1773 ( .A(_abc_17692_n4745), .B(_abc_17692_n4753), .Y(_abc_17692_n4754) );
  AND2X2 AND2X2_1774 ( .A(_abc_17692_n4752), .B(_abc_17692_n4755), .Y(_abc_17692_n4756) );
  AND2X2 AND2X2_1775 ( .A(_abc_17692_n4740), .B(_abc_17692_n4742), .Y(_abc_17692_n4758) );
  AND2X2 AND2X2_1776 ( .A(_abc_17692_n4729), .B(_abc_17692_n4737), .Y(_abc_17692_n4759) );
  AND2X2 AND2X2_1777 ( .A(_abc_17692_n4757), .B(_abc_17692_n4762), .Y(_abc_17692_n4763) );
  AND2X2 AND2X2_1778 ( .A(_abc_17692_n4763), .B(workunit2_15_), .Y(_abc_17692_n4764) );
  AND2X2 AND2X2_1779 ( .A(_abc_17692_n4767), .B(_abc_17692_n4766), .Y(_abc_17692_n4768) );
  AND2X2 AND2X2_178 ( .A(_abc_17692_n1092), .B(_abc_17692_n1086), .Y(_abc_17692_n1093) );
  AND2X2 AND2X2_1780 ( .A(_abc_17692_n4768), .B(_abc_17692_n4765), .Y(_abc_17692_n4769) );
  AND2X2 AND2X2_1781 ( .A(_abc_17692_n4581), .B(_abc_17692_n4571), .Y(_abc_17692_n4771) );
  AND2X2 AND2X2_1782 ( .A(_abc_17692_n4775), .B(_abc_17692_n1877_bF_buf3), .Y(_abc_17692_n4776) );
  AND2X2 AND2X2_1783 ( .A(_abc_17692_n4776), .B(_abc_17692_n4773), .Y(_abc_17692_n4777) );
  AND2X2 AND2X2_1784 ( .A(sum_15_), .B(\key_in[15] ), .Y(_abc_17692_n4780) );
  AND2X2 AND2X2_1785 ( .A(_abc_17692_n4781), .B(_abc_17692_n4782), .Y(_abc_17692_n4783) );
  AND2X2 AND2X2_1786 ( .A(_abc_17692_n4779), .B(_abc_17692_n4783), .Y(_abc_17692_n4784) );
  AND2X2 AND2X2_1787 ( .A(_abc_17692_n4778), .B(_abc_17692_n4785), .Y(_abc_17692_n4786) );
  AND2X2 AND2X2_1788 ( .A(_abc_17692_n4790), .B(_abc_17692_n4788), .Y(_abc_17692_n4791) );
  AND2X2 AND2X2_1789 ( .A(_abc_17692_n4791), .B(workunit2_15_), .Y(_abc_17692_n4792_1) );
  AND2X2 AND2X2_179 ( .A(delta_8_), .B(sum_8_), .Y(_abc_17692_n1096) );
  AND2X2 AND2X2_1790 ( .A(_abc_17692_n4793), .B(_abc_17692_n4794), .Y(_abc_17692_n4795) );
  AND2X2 AND2X2_1791 ( .A(_abc_17692_n4795), .B(_abc_17692_n4765), .Y(_abc_17692_n4796) );
  AND2X2 AND2X2_1792 ( .A(_abc_17692_n4619), .B(_abc_17692_n4607), .Y(_abc_17692_n4798) );
  AND2X2 AND2X2_1793 ( .A(_abc_17692_n4802), .B(_abc_17692_n1830_bF_buf3), .Y(_abc_17692_n4803) );
  AND2X2 AND2X2_1794 ( .A(_abc_17692_n4803), .B(_abc_17692_n4799), .Y(_abc_17692_n4804) );
  AND2X2 AND2X2_1795 ( .A(_abc_17692_n4805), .B(_abc_17692_n4632), .Y(_abc_17692_n4806) );
  AND2X2 AND2X2_1796 ( .A(sum_15_), .B(\key_in[47] ), .Y(_abc_17692_n4807) );
  AND2X2 AND2X2_1797 ( .A(_abc_17692_n4808), .B(_abc_17692_n4809), .Y(_abc_17692_n4810) );
  AND2X2 AND2X2_1798 ( .A(_abc_17692_n4806), .B(_abc_17692_n4810), .Y(_abc_17692_n4811) );
  AND2X2 AND2X2_1799 ( .A(_abc_17692_n4812), .B(_abc_17692_n4813), .Y(_abc_17692_n4814) );
  AND2X2 AND2X2_18 ( .A(_abc_17692_n667), .B(x_1_), .Y(_abc_17692_n671) );
  AND2X2 AND2X2_180 ( .A(_abc_17692_n1097), .B(_abc_17692_n1098), .Y(_abc_17692_n1099) );
  AND2X2 AND2X2_1800 ( .A(_abc_17692_n4818), .B(_abc_17692_n4817), .Y(_abc_17692_n4819) );
  AND2X2 AND2X2_1801 ( .A(_abc_17692_n4816), .B(_abc_17692_n4820), .Y(_abc_17692_n4821) );
  AND2X2 AND2X2_1802 ( .A(_abc_17692_n4821), .B(workunit2_15_), .Y(_abc_17692_n4822) );
  AND2X2 AND2X2_1803 ( .A(_abc_17692_n4823), .B(_abc_17692_n4824), .Y(_abc_17692_n4825) );
  AND2X2 AND2X2_1804 ( .A(_abc_17692_n4825), .B(_abc_17692_n4765), .Y(_abc_17692_n4826) );
  AND2X2 AND2X2_1805 ( .A(_abc_17692_n4645), .B(workunit2_14_bF_buf1), .Y(_abc_17692_n4829) );
  AND2X2 AND2X2_1806 ( .A(_abc_17692_n4660), .B(_abc_17692_n4830), .Y(_abc_17692_n4831) );
  AND2X2 AND2X2_1807 ( .A(_abc_17692_n4834), .B(_abc_17692_n1846_bF_buf3), .Y(_abc_17692_n4835) );
  AND2X2 AND2X2_1808 ( .A(_abc_17692_n4835), .B(_abc_17692_n4833), .Y(_abc_17692_n4836) );
  AND2X2 AND2X2_1809 ( .A(_abc_17692_n4840), .B(_abc_17692_n4519), .Y(_abc_17692_n4841) );
  AND2X2 AND2X2_181 ( .A(delta_7_), .B(sum_7_), .Y(_abc_17692_n1102) );
  AND2X2 AND2X2_1810 ( .A(sum_15_), .B(\key_in[111] ), .Y(_abc_17692_n4842) );
  AND2X2 AND2X2_1811 ( .A(_abc_17692_n4843), .B(_abc_17692_n4844), .Y(_abc_17692_n4845) );
  AND2X2 AND2X2_1812 ( .A(_abc_17692_n4841), .B(_abc_17692_n4845), .Y(_abc_17692_n4846) );
  AND2X2 AND2X2_1813 ( .A(_abc_17692_n4847), .B(_abc_17692_n4848), .Y(_abc_17692_n4849) );
  AND2X2 AND2X2_1814 ( .A(_abc_17692_n4853), .B(_abc_17692_n4852), .Y(_abc_17692_n4854) );
  AND2X2 AND2X2_1815 ( .A(_abc_17692_n4851), .B(_abc_17692_n4855), .Y(_abc_17692_n4856) );
  AND2X2 AND2X2_1816 ( .A(_abc_17692_n4856), .B(workunit2_15_), .Y(_abc_17692_n4857) );
  AND2X2 AND2X2_1817 ( .A(_abc_17692_n4858), .B(_abc_17692_n4859), .Y(_abc_17692_n4860) );
  AND2X2 AND2X2_1818 ( .A(_abc_17692_n4860), .B(_abc_17692_n4765), .Y(_abc_17692_n4861) );
  AND2X2 AND2X2_1819 ( .A(_abc_17692_n4547), .B(_abc_17692_n4535), .Y(_abc_17692_n4863) );
  AND2X2 AND2X2_182 ( .A(_abc_17692_n1079), .B(_abc_17692_n1103), .Y(_abc_17692_n1104_1) );
  AND2X2 AND2X2_1820 ( .A(_abc_17692_n4864), .B(_abc_17692_n4862), .Y(_abc_17692_n4865) );
  AND2X2 AND2X2_1821 ( .A(_abc_17692_n4863), .B(_abc_17692_n4866), .Y(_abc_17692_n4867) );
  AND2X2 AND2X2_1822 ( .A(_abc_17692_n4869), .B(state_6_bF_buf4), .Y(_abc_17692_n4870) );
  AND2X2 AND2X2_1823 ( .A(_abc_17692_n4870), .B(_abc_17692_n4839), .Y(_abc_17692_n4871) );
  AND2X2 AND2X2_1824 ( .A(_abc_17692_n4872), .B(workunit2_14_bF_buf0), .Y(_abc_17692_n4873) );
  AND2X2 AND2X2_1825 ( .A(_abc_17692_n4677), .B(_abc_17692_n4874), .Y(_abc_17692_n4875) );
  AND2X2 AND2X2_1826 ( .A(_abc_17692_n4878), .B(_abc_17692_n1863_bF_buf1), .Y(_abc_17692_n4879) );
  AND2X2 AND2X2_1827 ( .A(_abc_17692_n4879), .B(_abc_17692_n4877), .Y(_abc_17692_n4880) );
  AND2X2 AND2X2_1828 ( .A(_abc_17692_n4881), .B(workunit2_14_bF_buf3), .Y(_abc_17692_n4882) );
  AND2X2 AND2X2_1829 ( .A(_abc_17692_n4691), .B(_abc_17692_n4883), .Y(_abc_17692_n4884) );
  AND2X2 AND2X2_183 ( .A(_abc_17692_n1107_1), .B(state_3_bF_buf1), .Y(_abc_17692_n1108) );
  AND2X2 AND2X2_1830 ( .A(_abc_17692_n4887), .B(_abc_17692_n1877_bF_buf2), .Y(_abc_17692_n4888) );
  AND2X2 AND2X2_1831 ( .A(_abc_17692_n4888), .B(_abc_17692_n4886), .Y(_abc_17692_n4889) );
  AND2X2 AND2X2_1832 ( .A(_abc_17692_n4703), .B(_abc_17692_n4646_1), .Y(_abc_17692_n4890) );
  AND2X2 AND2X2_1833 ( .A(_abc_17692_n4893_1), .B(_abc_17692_n1846_bF_buf2), .Y(_abc_17692_n4894) );
  AND2X2 AND2X2_1834 ( .A(_abc_17692_n4894), .B(_abc_17692_n4892), .Y(_abc_17692_n4895) );
  AND2X2 AND2X2_1835 ( .A(_abc_17692_n4896_1), .B(workunit2_14_bF_buf2), .Y(_abc_17692_n4897) );
  AND2X2 AND2X2_1836 ( .A(_abc_17692_n4716), .B(_abc_17692_n4898), .Y(_abc_17692_n4899) );
  AND2X2 AND2X2_1837 ( .A(_abc_17692_n4902), .B(_abc_17692_n1830_bF_buf2), .Y(_abc_17692_n4903) );
  AND2X2 AND2X2_1838 ( .A(_abc_17692_n4903), .B(_abc_17692_n4900), .Y(_abc_17692_n4904) );
  AND2X2 AND2X2_1839 ( .A(_abc_17692_n4907), .B(state_7_bF_buf3), .Y(_abc_17692_n4908) );
  AND2X2 AND2X2_184 ( .A(_abc_17692_n1108), .B(_abc_17692_n1106), .Y(_abc_17692_n1109) );
  AND2X2 AND2X2_1840 ( .A(_abc_17692_n1885_bF_buf4), .B(workunit2_15_), .Y(_abc_17692_n4909) );
  AND2X2 AND2X2_1841 ( .A(state_8_bF_buf4), .B(\data_in2[15] ), .Y(_abc_17692_n4910) );
  AND2X2 AND2X2_1842 ( .A(_abc_17692_n4501), .B(_abc_17692_n4742), .Y(_abc_17692_n4914) );
  AND2X2 AND2X2_1843 ( .A(_abc_17692_n4489), .B(_abc_17692_n4914), .Y(_abc_17692_n4915) );
  AND2X2 AND2X2_1844 ( .A(_abc_17692_n4915), .B(_abc_17692_n4056), .Y(_abc_17692_n4916) );
  AND2X2 AND2X2_1845 ( .A(_abc_17692_n4916), .B(_abc_17692_n3207), .Y(_abc_17692_n4917) );
  AND2X2 AND2X2_1846 ( .A(_abc_17692_n4915), .B(_abc_17692_n4053), .Y(_abc_17692_n4918) );
  AND2X2 AND2X2_1847 ( .A(_abc_17692_n4914), .B(_abc_17692_n4492), .Y(_abc_17692_n4919) );
  AND2X2 AND2X2_1848 ( .A(_abc_17692_n4735_1), .B(_abc_17692_n4498), .Y(_abc_17692_n4920) );
  AND2X2 AND2X2_1849 ( .A(_abc_17692_n4925), .B(_abc_17692_n4927), .Y(_abc_17692_n4928) );
  AND2X2 AND2X2_185 ( .A(_abc_17692_n1111), .B(_abc_17692_n1100), .Y(_abc_17692_n1113) );
  AND2X2 AND2X2_1850 ( .A(_abc_17692_n4929), .B(workunit1_16_bF_buf3), .Y(_abc_17692_n4930) );
  AND2X2 AND2X2_1851 ( .A(_abc_17692_n4928), .B(_abc_17692_n3867), .Y(_abc_17692_n4931) );
  AND2X2 AND2X2_1852 ( .A(_abc_17692_n4924), .B(_abc_17692_n4933), .Y(_abc_17692_n4934) );
  AND2X2 AND2X2_1853 ( .A(_abc_17692_n4939), .B(_abc_17692_n4940), .Y(_abc_17692_n4941) );
  AND2X2 AND2X2_1854 ( .A(_abc_17692_n4938), .B(_abc_17692_n4941), .Y(_abc_17692_n4942) );
  AND2X2 AND2X2_1855 ( .A(_abc_17692_n4942), .B(_abc_17692_n4932), .Y(_abc_17692_n4943) );
  AND2X2 AND2X2_1856 ( .A(_abc_17692_n4560), .B(_abc_17692_n4750), .Y(_abc_17692_n4945) );
  AND2X2 AND2X2_1857 ( .A(_abc_17692_n4550), .B(_abc_17692_n4945), .Y(_abc_17692_n4946) );
  AND2X2 AND2X2_1858 ( .A(_abc_17692_n4126), .B(_abc_17692_n4946), .Y(_abc_17692_n4947) );
  AND2X2 AND2X2_1859 ( .A(_abc_17692_n3236), .B(_abc_17692_n4947), .Y(_abc_17692_n4948) );
  AND2X2 AND2X2_186 ( .A(_abc_17692_n1114), .B(state_15_bF_buf1), .Y(_abc_17692_n1115_1) );
  AND2X2 AND2X2_1860 ( .A(_abc_17692_n4125), .B(_abc_17692_n4946), .Y(_abc_17692_n4949) );
  AND2X2 AND2X2_1861 ( .A(_abc_17692_n4555), .B(_abc_17692_n4945), .Y(_abc_17692_n4950) );
  AND2X2 AND2X2_1862 ( .A(_abc_17692_n4749), .B(_abc_17692_n4557), .Y(_abc_17692_n4951) );
  AND2X2 AND2X2_1863 ( .A(sum_16_), .B(\key_in[80] ), .Y(_abc_17692_n4956) );
  AND2X2 AND2X2_1864 ( .A(_abc_17692_n4957), .B(_abc_17692_n4958), .Y(_abc_17692_n4959) );
  AND2X2 AND2X2_1865 ( .A(_abc_17692_n4955), .B(_abc_17692_n4959), .Y(_abc_17692_n4960) );
  AND2X2 AND2X2_1866 ( .A(_abc_17692_n4961), .B(_abc_17692_n4962), .Y(_abc_17692_n4963_1) );
  AND2X2 AND2X2_1867 ( .A(_abc_17692_n4966_1), .B(_abc_17692_n4968), .Y(_abc_17692_n4969) );
  AND2X2 AND2X2_1868 ( .A(_abc_17692_n4969), .B(workunit2_16_bF_buf2), .Y(_abc_17692_n4970) );
  AND2X2 AND2X2_1869 ( .A(_abc_17692_n4971), .B(_abc_17692_n4972), .Y(_abc_17692_n4973) );
  AND2X2 AND2X2_187 ( .A(_abc_17692_n1115_1), .B(_abc_17692_n1112), .Y(_abc_17692_n1116) );
  AND2X2 AND2X2_1870 ( .A(_abc_17692_n4770), .B(_abc_17692_n4573), .Y(_abc_17692_n4974) );
  AND2X2 AND2X2_1871 ( .A(_abc_17692_n4974), .B(_abc_17692_n4576), .Y(_abc_17692_n4975) );
  AND2X2 AND2X2_1872 ( .A(_abc_17692_n4768), .B(workunit2_15_), .Y(_abc_17692_n4976) );
  AND2X2 AND2X2_1873 ( .A(_abc_17692_n4770), .B(_abc_17692_n4570), .Y(_abc_17692_n4977) );
  AND2X2 AND2X2_1874 ( .A(_abc_17692_n4974), .B(_abc_17692_n4577), .Y(_abc_17692_n4980) );
  AND2X2 AND2X2_1875 ( .A(_abc_17692_n4155), .B(_abc_17692_n4980), .Y(_abc_17692_n4981) );
  AND2X2 AND2X2_1876 ( .A(_abc_17692_n4982), .B(_abc_17692_n4973), .Y(_abc_17692_n4983) );
  AND2X2 AND2X2_1877 ( .A(_abc_17692_n4985), .B(_abc_17692_n1877_bF_buf1), .Y(_abc_17692_n4986) );
  AND2X2 AND2X2_1878 ( .A(_abc_17692_n4986), .B(_abc_17692_n4984), .Y(_abc_17692_n4987) );
  AND2X2 AND2X2_1879 ( .A(_abc_17692_n4634), .B(_abc_17692_n4810), .Y(_abc_17692_n4988) );
  AND2X2 AND2X2_188 ( .A(_abc_17692_n722_bF_buf1), .B(sum_8_), .Y(_abc_17692_n1117) );
  AND2X2 AND2X2_1880 ( .A(_abc_17692_n4624), .B(_abc_17692_n4988), .Y(_abc_17692_n4989) );
  AND2X2 AND2X2_1881 ( .A(_abc_17692_n4208), .B(_abc_17692_n4989), .Y(_abc_17692_n4990) );
  AND2X2 AND2X2_1882 ( .A(_abc_17692_n3278_1), .B(_abc_17692_n4990), .Y(_abc_17692_n4991) );
  AND2X2 AND2X2_1883 ( .A(_abc_17692_n4207), .B(_abc_17692_n4989), .Y(_abc_17692_n4992) );
  AND2X2 AND2X2_1884 ( .A(_abc_17692_n4629), .B(_abc_17692_n4988), .Y(_abc_17692_n4993) );
  AND2X2 AND2X2_1885 ( .A(_abc_17692_n4809), .B(_abc_17692_n4631), .Y(_abc_17692_n4994) );
  AND2X2 AND2X2_1886 ( .A(sum_16_), .B(\key_in[48] ), .Y(_abc_17692_n4999) );
  AND2X2 AND2X2_1887 ( .A(_abc_17692_n5000), .B(_abc_17692_n5001), .Y(_abc_17692_n5002) );
  AND2X2 AND2X2_1888 ( .A(_abc_17692_n4998), .B(_abc_17692_n5002), .Y(_abc_17692_n5003) );
  AND2X2 AND2X2_1889 ( .A(_abc_17692_n5005), .B(_abc_17692_n5006), .Y(_abc_17692_n5007) );
  AND2X2 AND2X2_189 ( .A(delta_9_), .B(sum_9_), .Y(_abc_17692_n1121) );
  AND2X2 AND2X2_1890 ( .A(_abc_17692_n5007), .B(_abc_17692_n5008), .Y(_abc_17692_n5009) );
  AND2X2 AND2X2_1891 ( .A(_abc_17692_n5013), .B(_abc_17692_n5012), .Y(_abc_17692_n5014) );
  AND2X2 AND2X2_1892 ( .A(_abc_17692_n5014), .B(workunit2_16_bF_buf0), .Y(_abc_17692_n5015) );
  AND2X2 AND2X2_1893 ( .A(_abc_17692_n5016), .B(_abc_17692_n5017), .Y(_abc_17692_n5018) );
  AND2X2 AND2X2_1894 ( .A(_abc_17692_n5022), .B(_abc_17692_n5021), .Y(_abc_17692_n5023) );
  AND2X2 AND2X2_1895 ( .A(_abc_17692_n5020), .B(_abc_17692_n5023), .Y(_abc_17692_n5024) );
  AND2X2 AND2X2_1896 ( .A(_abc_17692_n5026), .B(_abc_17692_n5024), .Y(_abc_17692_n5027) );
  AND2X2 AND2X2_1897 ( .A(_abc_17692_n5028), .B(_abc_17692_n5018), .Y(_abc_17692_n5029) );
  AND2X2 AND2X2_1898 ( .A(_abc_17692_n5031), .B(_abc_17692_n1846_bF_buf1), .Y(_abc_17692_n5032) );
  AND2X2 AND2X2_1899 ( .A(_abc_17692_n5032), .B(_abc_17692_n5030), .Y(_abc_17692_n5033) );
  AND2X2 AND2X2_19 ( .A(_abc_17692_n672), .B(_abc_17692_n673), .Y(x_1__FF_INPUT) );
  AND2X2 AND2X2_190 ( .A(_abc_17692_n1123), .B(_abc_17692_n1124), .Y(_abc_17692_n1125) );
  AND2X2 AND2X2_1900 ( .A(_abc_17692_n4595), .B(_abc_17692_n4783), .Y(_abc_17692_n5034) );
  AND2X2 AND2X2_1901 ( .A(_abc_17692_n4585), .B(_abc_17692_n5034), .Y(_abc_17692_n5035) );
  AND2X2 AND2X2_1902 ( .A(_abc_17692_n4166), .B(_abc_17692_n5035), .Y(_abc_17692_n5036) );
  AND2X2 AND2X2_1903 ( .A(_abc_17692_n3311), .B(_abc_17692_n5036), .Y(_abc_17692_n5037) );
  AND2X2 AND2X2_1904 ( .A(_abc_17692_n4165), .B(_abc_17692_n5035), .Y(_abc_17692_n5038) );
  AND2X2 AND2X2_1905 ( .A(_abc_17692_n4590), .B(_abc_17692_n5034), .Y(_abc_17692_n5039) );
  AND2X2 AND2X2_1906 ( .A(_abc_17692_n4782), .B(_abc_17692_n4592), .Y(_abc_17692_n5040) );
  AND2X2 AND2X2_1907 ( .A(sum_16_), .B(\key_in[16] ), .Y(_abc_17692_n5045) );
  AND2X2 AND2X2_1908 ( .A(_abc_17692_n5046), .B(_abc_17692_n5047_1), .Y(_abc_17692_n5048) );
  AND2X2 AND2X2_1909 ( .A(_abc_17692_n5044_1), .B(_abc_17692_n5048), .Y(_abc_17692_n5049) );
  AND2X2 AND2X2_191 ( .A(_abc_17692_n1126), .B(_abc_17692_n1122), .Y(_abc_17692_n1127_1) );
  AND2X2 AND2X2_1910 ( .A(_abc_17692_n5051), .B(_abc_17692_n5052), .Y(_abc_17692_n5053) );
  AND2X2 AND2X2_1911 ( .A(_abc_17692_n5053), .B(_abc_17692_n5054), .Y(_abc_17692_n5055) );
  AND2X2 AND2X2_1912 ( .A(_abc_17692_n5059), .B(_abc_17692_n5058), .Y(_abc_17692_n5060) );
  AND2X2 AND2X2_1913 ( .A(_abc_17692_n5060), .B(workunit2_16_bF_buf2), .Y(_abc_17692_n5061) );
  AND2X2 AND2X2_1914 ( .A(_abc_17692_n5062), .B(_abc_17692_n5063), .Y(_abc_17692_n5064) );
  AND2X2 AND2X2_1915 ( .A(_abc_17692_n5068), .B(_abc_17692_n5067), .Y(_abc_17692_n5069) );
  AND2X2 AND2X2_1916 ( .A(_abc_17692_n5066), .B(_abc_17692_n5069), .Y(_abc_17692_n5070) );
  AND2X2 AND2X2_1917 ( .A(_abc_17692_n5072), .B(_abc_17692_n5070), .Y(_abc_17692_n5073) );
  AND2X2 AND2X2_1918 ( .A(_abc_17692_n5074), .B(_abc_17692_n5064), .Y(_abc_17692_n5075) );
  AND2X2 AND2X2_1919 ( .A(_abc_17692_n5077), .B(_abc_17692_n1830_bF_buf1), .Y(_abc_17692_n5078) );
  AND2X2 AND2X2_192 ( .A(_abc_17692_n1107_1), .B(_abc_17692_n1128), .Y(_abc_17692_n1129) );
  AND2X2 AND2X2_1920 ( .A(_abc_17692_n5078), .B(_abc_17692_n5076), .Y(_abc_17692_n5079) );
  AND2X2 AND2X2_1921 ( .A(_abc_17692_n4521), .B(_abc_17692_n4845), .Y(_abc_17692_n5082) );
  AND2X2 AND2X2_1922 ( .A(_abc_17692_n4511), .B(_abc_17692_n5082), .Y(_abc_17692_n5083) );
  AND2X2 AND2X2_1923 ( .A(_abc_17692_n4080), .B(_abc_17692_n5083), .Y(_abc_17692_n5084) );
  AND2X2 AND2X2_1924 ( .A(_abc_17692_n3359), .B(_abc_17692_n5084), .Y(_abc_17692_n5085) );
  AND2X2 AND2X2_1925 ( .A(_abc_17692_n4079), .B(_abc_17692_n5083), .Y(_abc_17692_n5086) );
  AND2X2 AND2X2_1926 ( .A(_abc_17692_n4516), .B(_abc_17692_n5082), .Y(_abc_17692_n5087) );
  AND2X2 AND2X2_1927 ( .A(_abc_17692_n4844), .B(_abc_17692_n4518), .Y(_abc_17692_n5088) );
  AND2X2 AND2X2_1928 ( .A(sum_16_), .B(\key_in[112] ), .Y(_abc_17692_n5093) );
  AND2X2 AND2X2_1929 ( .A(_abc_17692_n5094), .B(_abc_17692_n5095), .Y(_abc_17692_n5096) );
  AND2X2 AND2X2_193 ( .A(_abc_17692_n1133), .B(state_3_bF_buf0), .Y(_abc_17692_n1134) );
  AND2X2 AND2X2_1930 ( .A(_abc_17692_n5092), .B(_abc_17692_n5096), .Y(_abc_17692_n5097_1) );
  AND2X2 AND2X2_1931 ( .A(_abc_17692_n5098), .B(_abc_17692_n5099), .Y(_abc_17692_n5100_1) );
  AND2X2 AND2X2_1932 ( .A(_abc_17692_n5100_1), .B(_abc_17692_n5101), .Y(_abc_17692_n5102) );
  AND2X2 AND2X2_1933 ( .A(_abc_17692_n5105), .B(_abc_17692_n5106), .Y(_abc_17692_n5107) );
  AND2X2 AND2X2_1934 ( .A(_abc_17692_n5107), .B(workunit2_16_bF_buf0), .Y(_abc_17692_n5108) );
  AND2X2 AND2X2_1935 ( .A(_abc_17692_n5109), .B(_abc_17692_n5110), .Y(_abc_17692_n5111) );
  AND2X2 AND2X2_1936 ( .A(_abc_17692_n5114), .B(_abc_17692_n4535), .Y(_abc_17692_n5115) );
  AND2X2 AND2X2_1937 ( .A(_abc_17692_n5113), .B(_abc_17692_n5116), .Y(_abc_17692_n5117) );
  AND2X2 AND2X2_1938 ( .A(_abc_17692_n5120), .B(_abc_17692_n5117), .Y(_abc_17692_n5121) );
  AND2X2 AND2X2_1939 ( .A(_abc_17692_n5122), .B(_abc_17692_n5111), .Y(_abc_17692_n5124) );
  AND2X2 AND2X2_194 ( .A(_abc_17692_n1134), .B(_abc_17692_n1131), .Y(_abc_17692_n1135) );
  AND2X2 AND2X2_1940 ( .A(_abc_17692_n5125), .B(_abc_17692_n1863_bF_buf0), .Y(_abc_17692_n5126) );
  AND2X2 AND2X2_1941 ( .A(_abc_17692_n5126), .B(_abc_17692_n5123), .Y(_abc_17692_n5127) );
  AND2X2 AND2X2_1942 ( .A(_abc_17692_n5128), .B(state_6_bF_buf3), .Y(_abc_17692_n5129) );
  AND2X2 AND2X2_1943 ( .A(_abc_17692_n4862), .B(_abc_17692_n4669), .Y(_abc_17692_n5131) );
  AND2X2 AND2X2_1944 ( .A(_abc_17692_n5131), .B(_abc_17692_n4672), .Y(_abc_17692_n5132) );
  AND2X2 AND2X2_1945 ( .A(_abc_17692_n4860), .B(workunit2_15_), .Y(_abc_17692_n5133) );
  AND2X2 AND2X2_1946 ( .A(_abc_17692_n4862), .B(_abc_17692_n4873), .Y(_abc_17692_n5134) );
  AND2X2 AND2X2_1947 ( .A(_abc_17692_n5131), .B(_abc_17692_n4673), .Y(_abc_17692_n5137) );
  AND2X2 AND2X2_1948 ( .A(_abc_17692_n4259), .B(_abc_17692_n5137), .Y(_abc_17692_n5138) );
  AND2X2 AND2X2_1949 ( .A(_abc_17692_n5139), .B(_abc_17692_n5130), .Y(_abc_17692_n5141) );
  AND2X2 AND2X2_195 ( .A(_abc_17692_n1113), .B(_abc_17692_n1132), .Y(_abc_17692_n1136) );
  AND2X2 AND2X2_1950 ( .A(_abc_17692_n5142), .B(_abc_17692_n1863_bF_buf10), .Y(_abc_17692_n5143) );
  AND2X2 AND2X2_1951 ( .A(_abc_17692_n5143), .B(_abc_17692_n5140), .Y(_abc_17692_n5144) );
  AND2X2 AND2X2_1952 ( .A(_abc_17692_n5149), .B(_abc_17692_n5148), .Y(_abc_17692_n5150) );
  AND2X2 AND2X2_1953 ( .A(_abc_17692_n5147), .B(_abc_17692_n5151), .Y(_abc_17692_n5152) );
  AND2X2 AND2X2_1954 ( .A(_abc_17692_n5154), .B(_abc_17692_n5152), .Y(_abc_17692_n5155) );
  AND2X2 AND2X2_1955 ( .A(_abc_17692_n5156), .B(_abc_17692_n5145), .Y(_abc_17692_n5157) );
  AND2X2 AND2X2_1956 ( .A(_abc_17692_n5159), .B(_abc_17692_n1877_bF_buf0), .Y(_abc_17692_n5160) );
  AND2X2 AND2X2_1957 ( .A(_abc_17692_n5160), .B(_abc_17692_n5158), .Y(_abc_17692_n5161) );
  AND2X2 AND2X2_1958 ( .A(_abc_17692_n4827), .B(_abc_17692_n4648), .Y(_abc_17692_n5163) );
  AND2X2 AND2X2_1959 ( .A(_abc_17692_n5163), .B(_abc_17692_n4698), .Y(_abc_17692_n5164) );
  AND2X2 AND2X2_196 ( .A(_abc_17692_n1097), .B(sum_8_), .Y(_abc_17692_n1138_1) );
  AND2X2 AND2X2_1960 ( .A(_abc_17692_n4825), .B(workunit2_15_), .Y(_abc_17692_n5165) );
  AND2X2 AND2X2_1961 ( .A(_abc_17692_n4827), .B(_abc_17692_n5166), .Y(_abc_17692_n5167) );
  AND2X2 AND2X2_1962 ( .A(_abc_17692_n5163), .B(_abc_17692_n4699), .Y(_abc_17692_n5170) );
  AND2X2 AND2X2_1963 ( .A(_abc_17692_n4290), .B(_abc_17692_n5170), .Y(_abc_17692_n5171) );
  AND2X2 AND2X2_1964 ( .A(_abc_17692_n5172), .B(_abc_17692_n5162), .Y(_abc_17692_n5174) );
  AND2X2 AND2X2_1965 ( .A(_abc_17692_n5175), .B(_abc_17692_n1846_bF_buf0), .Y(_abc_17692_n5176) );
  AND2X2 AND2X2_1966 ( .A(_abc_17692_n5176), .B(_abc_17692_n5173), .Y(_abc_17692_n5177) );
  AND2X2 AND2X2_1967 ( .A(_abc_17692_n4797), .B(_abc_17692_n4707), .Y(_abc_17692_n5179) );
  AND2X2 AND2X2_1968 ( .A(_abc_17692_n5179), .B(_abc_17692_n4711), .Y(_abc_17692_n5180) );
  AND2X2 AND2X2_1969 ( .A(_abc_17692_n4795), .B(workunit2_15_), .Y(_abc_17692_n5181) );
  AND2X2 AND2X2_197 ( .A(_abc_17692_n1132), .B(_abc_17692_n1138_1), .Y(_abc_17692_n1141) );
  AND2X2 AND2X2_1970 ( .A(_abc_17692_n4797), .B(_abc_17692_n4897), .Y(_abc_17692_n5182) );
  AND2X2 AND2X2_1971 ( .A(_abc_17692_n5179), .B(_abc_17692_n4712), .Y(_abc_17692_n5185) );
  AND2X2 AND2X2_1972 ( .A(_abc_17692_n4306), .B(_abc_17692_n5185), .Y(_abc_17692_n5186) );
  AND2X2 AND2X2_1973 ( .A(_abc_17692_n5187), .B(_abc_17692_n5178), .Y(_abc_17692_n5188) );
  AND2X2 AND2X2_1974 ( .A(_abc_17692_n5190), .B(_abc_17692_n1830_bF_buf0), .Y(_abc_17692_n5191) );
  AND2X2 AND2X2_1975 ( .A(_abc_17692_n5191), .B(_abc_17692_n5189), .Y(_abc_17692_n5192) );
  AND2X2 AND2X2_1976 ( .A(_abc_17692_n5195), .B(state_7_bF_buf2), .Y(_abc_17692_n5196) );
  AND2X2 AND2X2_1977 ( .A(_abc_17692_n1885_bF_buf3), .B(workunit2_16_bF_buf2), .Y(_abc_17692_n5197) );
  AND2X2 AND2X2_1978 ( .A(state_8_bF_buf3), .B(\data_in2[16] ), .Y(_abc_17692_n5198) );
  AND2X2 AND2X2_1979 ( .A(_abc_17692_n5076), .B(_abc_17692_n5062), .Y(_abc_17692_n5202) );
  AND2X2 AND2X2_198 ( .A(_abc_17692_n1142), .B(state_15_bF_buf0), .Y(_abc_17692_n1143) );
  AND2X2 AND2X2_1980 ( .A(_abc_17692_n5204), .B(_abc_17692_n5206), .Y(_abc_17692_n5207) );
  AND2X2 AND2X2_1981 ( .A(_abc_17692_n5208), .B(workunit1_17_), .Y(_abc_17692_n5209) );
  AND2X2 AND2X2_1982 ( .A(_abc_17692_n5207), .B(_abc_17692_n4059), .Y(_abc_17692_n5211) );
  AND2X2 AND2X2_1983 ( .A(_abc_17692_n5210), .B(_abc_17692_n5212_1), .Y(_abc_17692_n5213) );
  AND2X2 AND2X2_1984 ( .A(_abc_17692_n5203), .B(_abc_17692_n5214), .Y(_abc_17692_n5216) );
  AND2X2 AND2X2_1985 ( .A(_abc_17692_n5217), .B(_abc_17692_n5215_1), .Y(_abc_17692_n5218) );
  AND2X2 AND2X2_1986 ( .A(_abc_17692_n5219), .B(_abc_17692_n5046), .Y(_abc_17692_n5220) );
  AND2X2 AND2X2_1987 ( .A(sum_17_), .B(\key_in[17] ), .Y(_abc_17692_n5221) );
  AND2X2 AND2X2_1988 ( .A(_abc_17692_n5222), .B(_abc_17692_n5223), .Y(_abc_17692_n5224) );
  AND2X2 AND2X2_1989 ( .A(_abc_17692_n5220), .B(_abc_17692_n5224), .Y(_abc_17692_n5225) );
  AND2X2 AND2X2_199 ( .A(_abc_17692_n1140), .B(_abc_17692_n1143), .Y(_abc_17692_n1144) );
  AND2X2 AND2X2_1990 ( .A(_abc_17692_n5226), .B(_abc_17692_n5227), .Y(_abc_17692_n5228) );
  AND2X2 AND2X2_1991 ( .A(_abc_17692_n5232), .B(_abc_17692_n5229), .Y(_abc_17692_n5233) );
  AND2X2 AND2X2_1992 ( .A(_abc_17692_n5233), .B(workunit2_17_), .Y(_abc_17692_n5234) );
  AND2X2 AND2X2_1993 ( .A(_abc_17692_n5235), .B(_abc_17692_n5236), .Y(_abc_17692_n5237) );
  AND2X2 AND2X2_1994 ( .A(_abc_17692_n5202), .B(_abc_17692_n5238), .Y(_abc_17692_n5239) );
  AND2X2 AND2X2_1995 ( .A(_abc_17692_n5240), .B(_abc_17692_n5237), .Y(_abc_17692_n5241) );
  AND2X2 AND2X2_1996 ( .A(_abc_17692_n5242), .B(_abc_17692_n1830_bF_buf10), .Y(_abc_17692_n5243) );
  AND2X2 AND2X2_1997 ( .A(_abc_17692_n5244), .B(_abc_17692_n4957), .Y(_abc_17692_n5245) );
  AND2X2 AND2X2_1998 ( .A(sum_17_), .B(\key_in[81] ), .Y(_abc_17692_n5246) );
  AND2X2 AND2X2_1999 ( .A(_abc_17692_n5247), .B(_abc_17692_n5248), .Y(_abc_17692_n5249) );
  AND2X2 AND2X2_2 ( .A(_abc_17692_n626), .B(_abc_17692_n627), .Y(_abc_17692_n628) );
  AND2X2 AND2X2_20 ( .A(_abc_17692_n671), .B(x_2_), .Y(_abc_17692_n675) );
  AND2X2 AND2X2_200 ( .A(_abc_17692_n1144), .B(_abc_17692_n1137), .Y(_abc_17692_n1145) );
  AND2X2 AND2X2_2000 ( .A(_abc_17692_n5245), .B(_abc_17692_n5249), .Y(_abc_17692_n5250) );
  AND2X2 AND2X2_2001 ( .A(_abc_17692_n5251), .B(_abc_17692_n5252), .Y(_abc_17692_n5253) );
  AND2X2 AND2X2_2002 ( .A(_abc_17692_n5256), .B(_abc_17692_n5254), .Y(_abc_17692_n5257) );
  AND2X2 AND2X2_2003 ( .A(_abc_17692_n5257), .B(workunit2_17_), .Y(_abc_17692_n5258) );
  AND2X2 AND2X2_2004 ( .A(_abc_17692_n5261), .B(_abc_17692_n5260), .Y(_abc_17692_n5262) );
  AND2X2 AND2X2_2005 ( .A(_abc_17692_n5263), .B(_abc_17692_n5259), .Y(_abc_17692_n5264) );
  AND2X2 AND2X2_2006 ( .A(_abc_17692_n5265), .B(_abc_17692_n4973), .Y(_abc_17692_n5268) );
  AND2X2 AND2X2_2007 ( .A(_abc_17692_n4982), .B(_abc_17692_n5268), .Y(_abc_17692_n5269) );
  AND2X2 AND2X2_2008 ( .A(_abc_17692_n5271), .B(_abc_17692_n1877_bF_buf10), .Y(_abc_17692_n5272) );
  AND2X2 AND2X2_2009 ( .A(_abc_17692_n5270), .B(_abc_17692_n5272), .Y(_abc_17692_n5273) );
  AND2X2 AND2X2_201 ( .A(_abc_17692_n722_bF_buf0), .B(sum_9_), .Y(_abc_17692_n1146) );
  AND2X2 AND2X2_2010 ( .A(_abc_17692_n5273), .B(_abc_17692_n5267), .Y(_abc_17692_n5274) );
  AND2X2 AND2X2_2011 ( .A(_abc_17692_n5030), .B(_abc_17692_n5016), .Y(_abc_17692_n5275_1) );
  AND2X2 AND2X2_2012 ( .A(_abc_17692_n5277), .B(_abc_17692_n5000), .Y(_abc_17692_n5278_1) );
  AND2X2 AND2X2_2013 ( .A(sum_17_), .B(\key_in[49] ), .Y(_abc_17692_n5279) );
  AND2X2 AND2X2_2014 ( .A(_abc_17692_n5280), .B(_abc_17692_n5281), .Y(_abc_17692_n5282) );
  AND2X2 AND2X2_2015 ( .A(_abc_17692_n5278_1), .B(_abc_17692_n5282), .Y(_abc_17692_n5283) );
  AND2X2 AND2X2_2016 ( .A(_abc_17692_n5284), .B(_abc_17692_n5285), .Y(_abc_17692_n5286) );
  AND2X2 AND2X2_2017 ( .A(_abc_17692_n5287), .B(_abc_17692_n5230), .Y(_abc_17692_n5288) );
  AND2X2 AND2X2_2018 ( .A(_abc_17692_n5286), .B(_abc_17692_n5218), .Y(_abc_17692_n5289) );
  AND2X2 AND2X2_2019 ( .A(_abc_17692_n5293), .B(_abc_17692_n5291), .Y(_abc_17692_n5294) );
  AND2X2 AND2X2_202 ( .A(delta_10_), .B(sum_10_), .Y(_abc_17692_n1150) );
  AND2X2 AND2X2_2020 ( .A(_abc_17692_n5297), .B(_abc_17692_n1846_bF_buf10), .Y(_abc_17692_n5298) );
  AND2X2 AND2X2_2021 ( .A(_abc_17692_n5298), .B(_abc_17692_n5296), .Y(_abc_17692_n5299) );
  AND2X2 AND2X2_2022 ( .A(_abc_17692_n5125), .B(_abc_17692_n5109), .Y(_abc_17692_n5302) );
  AND2X2 AND2X2_2023 ( .A(_abc_17692_n5303), .B(_abc_17692_n5094), .Y(_abc_17692_n5304) );
  AND2X2 AND2X2_2024 ( .A(sum_17_), .B(\key_in[113] ), .Y(_abc_17692_n5305) );
  AND2X2 AND2X2_2025 ( .A(_abc_17692_n5306), .B(_abc_17692_n5307), .Y(_abc_17692_n5308) );
  AND2X2 AND2X2_2026 ( .A(_abc_17692_n5304), .B(_abc_17692_n5308), .Y(_abc_17692_n5309) );
  AND2X2 AND2X2_2027 ( .A(_abc_17692_n5310), .B(_abc_17692_n5311), .Y(_abc_17692_n5312) );
  AND2X2 AND2X2_2028 ( .A(_abc_17692_n5315), .B(_abc_17692_n5313), .Y(_abc_17692_n5316) );
  AND2X2 AND2X2_2029 ( .A(_abc_17692_n5316), .B(workunit2_17_), .Y(_abc_17692_n5317) );
  AND2X2 AND2X2_203 ( .A(_abc_17692_n1151), .B(_abc_17692_n1152_1), .Y(_abc_17692_n1153) );
  AND2X2 AND2X2_2030 ( .A(_abc_17692_n5319), .B(_abc_17692_n5260), .Y(_abc_17692_n5320) );
  AND2X2 AND2X2_2031 ( .A(_abc_17692_n5321), .B(_abc_17692_n5318), .Y(_abc_17692_n5322) );
  AND2X2 AND2X2_2032 ( .A(_abc_17692_n5302), .B(_abc_17692_n5323), .Y(_abc_17692_n5324) );
  AND2X2 AND2X2_2033 ( .A(_abc_17692_n5325), .B(_abc_17692_n5322), .Y(_abc_17692_n5326) );
  AND2X2 AND2X2_2034 ( .A(_abc_17692_n5327), .B(_abc_17692_n1863_bF_buf9), .Y(_abc_17692_n5328) );
  AND2X2 AND2X2_2035 ( .A(_abc_17692_n5329), .B(state_6_bF_buf2), .Y(_abc_17692_n5330) );
  AND2X2 AND2X2_2036 ( .A(_abc_17692_n5331), .B(workunit2_16_bF_buf1), .Y(_abc_17692_n5332) );
  AND2X2 AND2X2_2037 ( .A(_abc_17692_n5142), .B(_abc_17692_n5333), .Y(_abc_17692_n5334) );
  AND2X2 AND2X2_2038 ( .A(_abc_17692_n5335), .B(_abc_17692_n5323), .Y(_abc_17692_n5336) );
  AND2X2 AND2X2_2039 ( .A(_abc_17692_n5334), .B(_abc_17692_n5322), .Y(_abc_17692_n5337) );
  AND2X2 AND2X2_204 ( .A(_abc_17692_n1128), .B(_abc_17692_n1122), .Y(_abc_17692_n1157) );
  AND2X2 AND2X2_2040 ( .A(_abc_17692_n5338), .B(_abc_17692_n1863_bF_buf8), .Y(_abc_17692_n5339) );
  AND2X2 AND2X2_2041 ( .A(_abc_17692_n5340), .B(workunit2_16_bF_buf0), .Y(_abc_17692_n5341) );
  AND2X2 AND2X2_2042 ( .A(_abc_17692_n5158), .B(_abc_17692_n5342), .Y(_abc_17692_n5343) );
  AND2X2 AND2X2_2043 ( .A(_abc_17692_n5346), .B(_abc_17692_n1877_bF_buf9), .Y(_abc_17692_n5347) );
  AND2X2 AND2X2_2044 ( .A(_abc_17692_n5347), .B(_abc_17692_n5345), .Y(_abc_17692_n5348) );
  AND2X2 AND2X2_2045 ( .A(_abc_17692_n5349), .B(workunit2_16_bF_buf3), .Y(_abc_17692_n5350) );
  AND2X2 AND2X2_2046 ( .A(_abc_17692_n5175), .B(_abc_17692_n5351), .Y(_abc_17692_n5352) );
  AND2X2 AND2X2_2047 ( .A(_abc_17692_n5355), .B(_abc_17692_n1846_bF_buf9), .Y(_abc_17692_n5356) );
  AND2X2 AND2X2_2048 ( .A(_abc_17692_n5356), .B(_abc_17692_n5354), .Y(_abc_17692_n5357) );
  AND2X2 AND2X2_2049 ( .A(_abc_17692_n5358), .B(workunit2_16_bF_buf2), .Y(_abc_17692_n5359) );
  AND2X2 AND2X2_205 ( .A(_abc_17692_n1156), .B(_abc_17692_n1158), .Y(_abc_17692_n1159) );
  AND2X2 AND2X2_2050 ( .A(_abc_17692_n5189), .B(_abc_17692_n5360), .Y(_abc_17692_n5361) );
  AND2X2 AND2X2_2051 ( .A(_abc_17692_n5364), .B(_abc_17692_n1830_bF_buf9), .Y(_abc_17692_n5365) );
  AND2X2 AND2X2_2052 ( .A(_abc_17692_n5365), .B(_abc_17692_n5363), .Y(_abc_17692_n5366_1) );
  AND2X2 AND2X2_2053 ( .A(_abc_17692_n5369_1), .B(state_7_bF_buf1), .Y(_abc_17692_n5370) );
  AND2X2 AND2X2_2054 ( .A(_abc_17692_n1885_bF_buf2), .B(workunit2_17_), .Y(_abc_17692_n5371) );
  AND2X2 AND2X2_2055 ( .A(state_8_bF_buf2), .B(\data_in2[17] ), .Y(_abc_17692_n5372) );
  AND2X2 AND2X2_2056 ( .A(_abc_17692_n5377), .B(_abc_17692_n5379), .Y(_abc_17692_n5380) );
  AND2X2 AND2X2_2057 ( .A(_abc_17692_n5381), .B(workunit1_18_), .Y(_abc_17692_n5382) );
  AND2X2 AND2X2_2058 ( .A(_abc_17692_n5380), .B(_abc_17692_n4322), .Y(_abc_17692_n5383) );
  AND2X2 AND2X2_2059 ( .A(_abc_17692_n5212_1), .B(_abc_17692_n4930), .Y(_abc_17692_n5386) );
  AND2X2 AND2X2_206 ( .A(_abc_17692_n1160), .B(_abc_17692_n1155), .Y(_abc_17692_n1161) );
  AND2X2 AND2X2_2060 ( .A(_abc_17692_n4933), .B(_abc_17692_n5213), .Y(_abc_17692_n5388) );
  AND2X2 AND2X2_2061 ( .A(_abc_17692_n4924), .B(_abc_17692_n5388), .Y(_abc_17692_n5389) );
  AND2X2 AND2X2_2062 ( .A(_abc_17692_n5390), .B(_abc_17692_n5385), .Y(_abc_17692_n5391) );
  AND2X2 AND2X2_2063 ( .A(_abc_17692_n5392), .B(_abc_17692_n5384), .Y(_abc_17692_n5393) );
  AND2X2 AND2X2_2064 ( .A(sum_18_), .B(\key_in[82] ), .Y(_abc_17692_n5395) );
  AND2X2 AND2X2_2065 ( .A(_abc_17692_n5396), .B(_abc_17692_n5397), .Y(_abc_17692_n5398) );
  AND2X2 AND2X2_2066 ( .A(_abc_17692_n5248), .B(_abc_17692_n4956), .Y(_abc_17692_n5400) );
  AND2X2 AND2X2_2067 ( .A(_abc_17692_n4959), .B(_abc_17692_n5249), .Y(_abc_17692_n5403) );
  AND2X2 AND2X2_2068 ( .A(_abc_17692_n5405), .B(_abc_17692_n5402), .Y(_abc_17692_n5406) );
  AND2X2 AND2X2_2069 ( .A(_abc_17692_n5406), .B(_abc_17692_n5399), .Y(_abc_17692_n5409) );
  AND2X2 AND2X2_207 ( .A(_abc_17692_n1163), .B(state_3_bF_buf4), .Y(_abc_17692_n1164) );
  AND2X2 AND2X2_2070 ( .A(_abc_17692_n5410), .B(_abc_17692_n5394), .Y(_abc_17692_n5411) );
  AND2X2 AND2X2_2071 ( .A(_abc_17692_n5413), .B(_abc_17692_n5412), .Y(_abc_17692_n5414) );
  AND2X2 AND2X2_2072 ( .A(_abc_17692_n5415), .B(workunit2_18_), .Y(_abc_17692_n5416) );
  AND2X2 AND2X2_2073 ( .A(_abc_17692_n5417), .B(_abc_17692_n5418), .Y(_abc_17692_n5419) );
  AND2X2 AND2X2_2074 ( .A(_abc_17692_n5261), .B(workunit2_17_), .Y(_abc_17692_n5420_1) );
  AND2X2 AND2X2_2075 ( .A(_abc_17692_n5271), .B(_abc_17692_n5421), .Y(_abc_17692_n5422) );
  AND2X2 AND2X2_2076 ( .A(_abc_17692_n5270), .B(_abc_17692_n5422), .Y(_abc_17692_n5423_1) );
  AND2X2 AND2X2_2077 ( .A(_abc_17692_n5424), .B(_abc_17692_n5419), .Y(_abc_17692_n5425) );
  AND2X2 AND2X2_2078 ( .A(_abc_17692_n5427), .B(_abc_17692_n1877_bF_buf8), .Y(_abc_17692_n5428) );
  AND2X2 AND2X2_2079 ( .A(_abc_17692_n5428), .B(_abc_17692_n5426), .Y(_abc_17692_n5429) );
  AND2X2 AND2X2_208 ( .A(_abc_17692_n1164), .B(_abc_17692_n1162), .Y(_abc_17692_n1165) );
  AND2X2 AND2X2_2080 ( .A(sum_18_), .B(\key_in[50] ), .Y(_abc_17692_n5431) );
  AND2X2 AND2X2_2081 ( .A(_abc_17692_n5432), .B(_abc_17692_n5433), .Y(_abc_17692_n5434) );
  AND2X2 AND2X2_2082 ( .A(_abc_17692_n5281), .B(_abc_17692_n4999), .Y(_abc_17692_n5435) );
  AND2X2 AND2X2_2083 ( .A(_abc_17692_n5002), .B(_abc_17692_n5282), .Y(_abc_17692_n5437) );
  AND2X2 AND2X2_2084 ( .A(_abc_17692_n4998), .B(_abc_17692_n5437), .Y(_abc_17692_n5438) );
  AND2X2 AND2X2_2085 ( .A(_abc_17692_n5439), .B(_abc_17692_n5434), .Y(_abc_17692_n5440) );
  AND2X2 AND2X2_2086 ( .A(_abc_17692_n5442), .B(_abc_17692_n5441), .Y(_abc_17692_n5443) );
  AND2X2 AND2X2_2087 ( .A(_abc_17692_n5394), .B(_abc_17692_n5444), .Y(_abc_17692_n5445) );
  AND2X2 AND2X2_2088 ( .A(_abc_17692_n5412), .B(_abc_17692_n5446), .Y(_abc_17692_n5447) );
  AND2X2 AND2X2_2089 ( .A(_abc_17692_n5451), .B(_abc_17692_n5449), .Y(_abc_17692_n5452) );
  AND2X2 AND2X2_209 ( .A(_abc_17692_n1123), .B(sum_9_), .Y(_abc_17692_n1166) );
  AND2X2 AND2X2_2090 ( .A(_abc_17692_n5290), .B(workunit2_17_), .Y(_abc_17692_n5454) );
  AND2X2 AND2X2_2091 ( .A(_abc_17692_n5456), .B(_abc_17692_n5455), .Y(_abc_17692_n5457) );
  AND2X2 AND2X2_2092 ( .A(_abc_17692_n5295), .B(_abc_17692_n5018), .Y(_abc_17692_n5459) );
  AND2X2 AND2X2_2093 ( .A(_abc_17692_n5028), .B(_abc_17692_n5459), .Y(_abc_17692_n5460) );
  AND2X2 AND2X2_2094 ( .A(_abc_17692_n5461), .B(_abc_17692_n5453), .Y(_abc_17692_n5462) );
  AND2X2 AND2X2_2095 ( .A(_abc_17692_n5464), .B(_abc_17692_n1846_bF_buf8), .Y(_abc_17692_n5465) );
  AND2X2 AND2X2_2096 ( .A(_abc_17692_n5465), .B(_abc_17692_n5463), .Y(_abc_17692_n5466) );
  AND2X2 AND2X2_2097 ( .A(_abc_17692_n5048), .B(_abc_17692_n5224), .Y(_abc_17692_n5467) );
  AND2X2 AND2X2_2098 ( .A(_abc_17692_n5044_1), .B(_abc_17692_n5467), .Y(_abc_17692_n5468) );
  AND2X2 AND2X2_2099 ( .A(_abc_17692_n5046), .B(_abc_17692_n5222), .Y(_abc_17692_n5470) );
  AND2X2 AND2X2_21 ( .A(_abc_17692_n676_1), .B(_abc_17692_n677_1), .Y(x_2__FF_INPUT) );
  AND2X2 AND2X2_210 ( .A(_abc_17692_n1137), .B(_abc_17692_n1168), .Y(_abc_17692_n1169) );
  AND2X2 AND2X2_2100 ( .A(sum_18_), .B(\key_in[18] ), .Y(_abc_17692_n5474) );
  AND2X2 AND2X2_2101 ( .A(_abc_17692_n5475), .B(_abc_17692_n5476), .Y(_abc_17692_n5477) );
  AND2X2 AND2X2_2102 ( .A(_abc_17692_n5473), .B(_abc_17692_n5477), .Y(_abc_17692_n5478) );
  AND2X2 AND2X2_2103 ( .A(_abc_17692_n5479), .B(_abc_17692_n5480), .Y(_abc_17692_n5481) );
  AND2X2 AND2X2_2104 ( .A(_abc_17692_n5485), .B(_abc_17692_n5484), .Y(_abc_17692_n5486) );
  AND2X2 AND2X2_2105 ( .A(_abc_17692_n5489), .B(_abc_17692_n5487), .Y(_abc_17692_n5490) );
  AND2X2 AND2X2_2106 ( .A(_abc_17692_n5493), .B(_abc_17692_n5492), .Y(_abc_17692_n5494) );
  AND2X2 AND2X2_2107 ( .A(_abc_17692_n5238), .B(_abc_17692_n5064), .Y(_abc_17692_n5496) );
  AND2X2 AND2X2_2108 ( .A(_abc_17692_n5074), .B(_abc_17692_n5496), .Y(_abc_17692_n5497) );
  AND2X2 AND2X2_2109 ( .A(_abc_17692_n5498), .B(_abc_17692_n5491), .Y(_abc_17692_n5500) );
  AND2X2 AND2X2_211 ( .A(_abc_17692_n1170), .B(_abc_17692_n1154), .Y(_abc_17692_n1171) );
  AND2X2 AND2X2_2110 ( .A(_abc_17692_n5501), .B(_abc_17692_n1830_bF_buf8), .Y(_abc_17692_n5502) );
  AND2X2 AND2X2_2111 ( .A(_abc_17692_n5502), .B(_abc_17692_n5499), .Y(_abc_17692_n5503) );
  AND2X2 AND2X2_2112 ( .A(_abc_17692_n5096), .B(_abc_17692_n5308), .Y(_abc_17692_n5506) );
  AND2X2 AND2X2_2113 ( .A(_abc_17692_n5092), .B(_abc_17692_n5506), .Y(_abc_17692_n5507) );
  AND2X2 AND2X2_2114 ( .A(_abc_17692_n5094), .B(_abc_17692_n5306), .Y(_abc_17692_n5509) );
  AND2X2 AND2X2_2115 ( .A(sum_18_), .B(\key_in[114] ), .Y(_abc_17692_n5513) );
  AND2X2 AND2X2_2116 ( .A(_abc_17692_n5514), .B(_abc_17692_n5515), .Y(_abc_17692_n5516) );
  AND2X2 AND2X2_2117 ( .A(_abc_17692_n5512), .B(_abc_17692_n5516), .Y(_abc_17692_n5517) );
  AND2X2 AND2X2_2118 ( .A(_abc_17692_n5518), .B(_abc_17692_n5519), .Y(_abc_17692_n5520) );
  AND2X2 AND2X2_2119 ( .A(_abc_17692_n5523), .B(_abc_17692_n5524), .Y(_abc_17692_n5525) );
  AND2X2 AND2X2_212 ( .A(_abc_17692_n1173), .B(state_15_bF_buf4), .Y(_abc_17692_n1174) );
  AND2X2 AND2X2_2120 ( .A(_abc_17692_n5526), .B(_abc_17692_n5430), .Y(_abc_17692_n5527) );
  AND2X2 AND2X2_2121 ( .A(_abc_17692_n5525), .B(workunit2_18_), .Y(_abc_17692_n5528) );
  AND2X2 AND2X2_2122 ( .A(_abc_17692_n5319), .B(workunit2_17_), .Y(_abc_17692_n5531) );
  AND2X2 AND2X2_2123 ( .A(_abc_17692_n5533), .B(_abc_17692_n5532), .Y(_abc_17692_n5534) );
  AND2X2 AND2X2_2124 ( .A(_abc_17692_n5323), .B(_abc_17692_n5111), .Y(_abc_17692_n5536) );
  AND2X2 AND2X2_2125 ( .A(_abc_17692_n5122), .B(_abc_17692_n5536), .Y(_abc_17692_n5537) );
  AND2X2 AND2X2_2126 ( .A(_abc_17692_n5538), .B(_abc_17692_n5530), .Y(_abc_17692_n5539) );
  AND2X2 AND2X2_2127 ( .A(_abc_17692_n5541), .B(_abc_17692_n1863_bF_buf7), .Y(_abc_17692_n5542) );
  AND2X2 AND2X2_2128 ( .A(_abc_17692_n5542), .B(_abc_17692_n5540), .Y(_abc_17692_n5543) );
  AND2X2 AND2X2_2129 ( .A(_abc_17692_n5544), .B(state_6_bF_buf1), .Y(_abc_17692_n5545_1) );
  AND2X2 AND2X2_213 ( .A(_abc_17692_n1174), .B(_abc_17692_n1172), .Y(_abc_17692_n1175) );
  AND2X2 AND2X2_2130 ( .A(_abc_17692_n5321), .B(_abc_17692_n5546), .Y(_abc_17692_n5547) );
  AND2X2 AND2X2_2131 ( .A(_abc_17692_n5322), .B(_abc_17692_n5130), .Y(_abc_17692_n5548_1) );
  AND2X2 AND2X2_2132 ( .A(_abc_17692_n5139), .B(_abc_17692_n5548_1), .Y(_abc_17692_n5549) );
  AND2X2 AND2X2_2133 ( .A(_abc_17692_n5550), .B(_abc_17692_n5529), .Y(_abc_17692_n5551) );
  AND2X2 AND2X2_2134 ( .A(_abc_17692_n5553), .B(_abc_17692_n1863_bF_buf6), .Y(_abc_17692_n5554) );
  AND2X2 AND2X2_2135 ( .A(_abc_17692_n5554), .B(_abc_17692_n5552), .Y(_abc_17692_n5555) );
  AND2X2 AND2X2_2136 ( .A(_abc_17692_n5344), .B(_abc_17692_n5263), .Y(_abc_17692_n5557) );
  AND2X2 AND2X2_2137 ( .A(_abc_17692_n5558), .B(_abc_17692_n5556), .Y(_abc_17692_n5559) );
  AND2X2 AND2X2_2138 ( .A(_abc_17692_n5561), .B(_abc_17692_n1877_bF_buf7), .Y(_abc_17692_n5562) );
  AND2X2 AND2X2_2139 ( .A(_abc_17692_n5562), .B(_abc_17692_n5560), .Y(_abc_17692_n5563) );
  AND2X2 AND2X2_214 ( .A(_abc_17692_n722_bF_buf3), .B(sum_10_), .Y(_abc_17692_n1176) );
  AND2X2 AND2X2_2140 ( .A(_abc_17692_n5564), .B(_abc_17692_n5236), .Y(_abc_17692_n5565) );
  AND2X2 AND2X2_2141 ( .A(_abc_17692_n5237), .B(_abc_17692_n5178), .Y(_abc_17692_n5566) );
  AND2X2 AND2X2_2142 ( .A(_abc_17692_n5187), .B(_abc_17692_n5566), .Y(_abc_17692_n5567) );
  AND2X2 AND2X2_2143 ( .A(_abc_17692_n5568), .B(_abc_17692_n5490), .Y(_abc_17692_n5569) );
  AND2X2 AND2X2_2144 ( .A(_abc_17692_n5571), .B(_abc_17692_n1830_bF_buf7), .Y(_abc_17692_n5572) );
  AND2X2 AND2X2_2145 ( .A(_abc_17692_n5572), .B(_abc_17692_n5570), .Y(_abc_17692_n5573) );
  AND2X2 AND2X2_2146 ( .A(_abc_17692_n5291), .B(_abc_17692_n5351), .Y(_abc_17692_n5575) );
  AND2X2 AND2X2_2147 ( .A(_abc_17692_n5294), .B(_abc_17692_n5162), .Y(_abc_17692_n5578) );
  AND2X2 AND2X2_2148 ( .A(_abc_17692_n5172), .B(_abc_17692_n5578), .Y(_abc_17692_n5579) );
  AND2X2 AND2X2_2149 ( .A(_abc_17692_n5580), .B(_abc_17692_n5452), .Y(_abc_17692_n5581) );
  AND2X2 AND2X2_215 ( .A(_abc_17692_n1180), .B(delta_11_), .Y(_abc_17692_n1181) );
  AND2X2 AND2X2_2150 ( .A(_abc_17692_n5583), .B(_abc_17692_n1846_bF_buf7), .Y(_abc_17692_n5584) );
  AND2X2 AND2X2_2151 ( .A(_abc_17692_n5584), .B(_abc_17692_n5582), .Y(_abc_17692_n5585) );
  AND2X2 AND2X2_2152 ( .A(_abc_17692_n5588), .B(state_7_bF_buf0), .Y(_abc_17692_n5589) );
  AND2X2 AND2X2_2153 ( .A(_abc_17692_n1885_bF_buf1), .B(workunit2_18_), .Y(_abc_17692_n5590) );
  AND2X2 AND2X2_2154 ( .A(state_8_bF_buf1), .B(\data_in2[18] ), .Y(_abc_17692_n5591) );
  AND2X2 AND2X2_2155 ( .A(_abc_17692_n5597), .B(_abc_17692_n5599), .Y(_abc_17692_n5600) );
  AND2X2 AND2X2_2156 ( .A(_abc_17692_n5601), .B(workunit1_19_), .Y(_abc_17692_n5602) );
  AND2X2 AND2X2_2157 ( .A(_abc_17692_n5600), .B(_abc_17692_n4494), .Y(_abc_17692_n5604) );
  AND2X2 AND2X2_2158 ( .A(_abc_17692_n5603), .B(_abc_17692_n5605), .Y(_abc_17692_n5606) );
  AND2X2 AND2X2_2159 ( .A(_abc_17692_n5596), .B(_abc_17692_n5606), .Y(_abc_17692_n5607) );
  AND2X2 AND2X2_216 ( .A(_abc_17692_n1182), .B(_abc_17692_n1183), .Y(_abc_17692_n1184) );
  AND2X2 AND2X2_2160 ( .A(_abc_17692_n5595), .B(_abc_17692_n5608_1), .Y(_abc_17692_n5609) );
  AND2X2 AND2X2_2161 ( .A(_abc_17692_n5407), .B(_abc_17692_n5396), .Y(_abc_17692_n5612) );
  AND2X2 AND2X2_2162 ( .A(sum_19_), .B(\key_in[83] ), .Y(_abc_17692_n5613) );
  AND2X2 AND2X2_2163 ( .A(_abc_17692_n5614), .B(_abc_17692_n5615), .Y(_abc_17692_n5616) );
  AND2X2 AND2X2_2164 ( .A(_abc_17692_n5612), .B(_abc_17692_n5616), .Y(_abc_17692_n5617) );
  AND2X2 AND2X2_2165 ( .A(_abc_17692_n5618), .B(_abc_17692_n5619), .Y(_abc_17692_n5620) );
  AND2X2 AND2X2_2166 ( .A(_abc_17692_n5623), .B(_abc_17692_n5621), .Y(_abc_17692_n5624) );
  AND2X2 AND2X2_2167 ( .A(_abc_17692_n5624), .B(workunit2_19_), .Y(_abc_17692_n5625) );
  AND2X2 AND2X2_2168 ( .A(_abc_17692_n5627), .B(_abc_17692_n5626), .Y(_abc_17692_n5628) );
  AND2X2 AND2X2_2169 ( .A(_abc_17692_n5630), .B(workunit2_18_), .Y(_abc_17692_n5631) );
  AND2X2 AND2X2_217 ( .A(_abc_17692_n1162), .B(_abc_17692_n1186), .Y(_abc_17692_n1187) );
  AND2X2 AND2X2_2170 ( .A(_abc_17692_n5632), .B(_abc_17692_n5629), .Y(_abc_17692_n5633) );
  AND2X2 AND2X2_2171 ( .A(_abc_17692_n5635), .B(_abc_17692_n5634), .Y(_abc_17692_n5636) );
  AND2X2 AND2X2_2172 ( .A(_abc_17692_n5637), .B(_abc_17692_n1877_bF_buf6), .Y(_abc_17692_n5638) );
  AND2X2 AND2X2_2173 ( .A(sum_19_), .B(\key_in[115] ), .Y(_abc_17692_n5641) );
  AND2X2 AND2X2_2174 ( .A(_abc_17692_n5642), .B(_abc_17692_n5643), .Y(_abc_17692_n5644) );
  AND2X2 AND2X2_2175 ( .A(_abc_17692_n5640), .B(_abc_17692_n5644), .Y(_abc_17692_n5645) );
  AND2X2 AND2X2_2176 ( .A(_abc_17692_n5646), .B(_abc_17692_n5647), .Y(_abc_17692_n5648) );
  AND2X2 AND2X2_2177 ( .A(_abc_17692_n5652), .B(_abc_17692_n5649), .Y(_abc_17692_n5653) );
  AND2X2 AND2X2_2178 ( .A(_abc_17692_n5653), .B(workunit2_19_), .Y(_abc_17692_n5654) );
  AND2X2 AND2X2_2179 ( .A(_abc_17692_n5655), .B(_abc_17692_n5656), .Y(_abc_17692_n5657) );
  AND2X2 AND2X2_218 ( .A(_abc_17692_n1190), .B(state_3_bF_buf3), .Y(_abc_17692_n1191) );
  AND2X2 AND2X2_2180 ( .A(_abc_17692_n5657), .B(_abc_17692_n5626), .Y(_abc_17692_n5658) );
  AND2X2 AND2X2_2181 ( .A(_abc_17692_n5526), .B(workunit2_18_), .Y(_abc_17692_n5660) );
  AND2X2 AND2X2_2182 ( .A(_abc_17692_n5552), .B(_abc_17692_n5661), .Y(_abc_17692_n5662) );
  AND2X2 AND2X2_2183 ( .A(_abc_17692_n5664), .B(_abc_17692_n5665), .Y(_abc_17692_n5666) );
  AND2X2 AND2X2_2184 ( .A(_abc_17692_n5668), .B(_abc_17692_n1863_bF_buf5), .Y(_abc_17692_n5669) );
  AND2X2 AND2X2_2185 ( .A(_abc_17692_n5669), .B(_abc_17692_n5663), .Y(_abc_17692_n5670) );
  AND2X2 AND2X2_2186 ( .A(sum_19_), .B(\key_in[51] ), .Y(_abc_17692_n5673) );
  AND2X2 AND2X2_2187 ( .A(_abc_17692_n5674), .B(_abc_17692_n5675), .Y(_abc_17692_n5676) );
  AND2X2 AND2X2_2188 ( .A(_abc_17692_n5672), .B(_abc_17692_n5676), .Y(_abc_17692_n5677) );
  AND2X2 AND2X2_2189 ( .A(_abc_17692_n5682), .B(_abc_17692_n5678), .Y(_abc_17692_n5683) );
  AND2X2 AND2X2_219 ( .A(_abc_17692_n1191), .B(_abc_17692_n1189), .Y(_abc_17692_n1192_1) );
  AND2X2 AND2X2_2190 ( .A(_abc_17692_n5681), .B(_abc_17692_n5684), .Y(_abc_17692_n5685) );
  AND2X2 AND2X2_2191 ( .A(_abc_17692_n5687), .B(_abc_17692_n5688), .Y(_abc_17692_n5689) );
  AND2X2 AND2X2_2192 ( .A(_abc_17692_n5686), .B(_abc_17692_n5690), .Y(_abc_17692_n5691) );
  AND2X2 AND2X2_2193 ( .A(_abc_17692_n5582), .B(_abc_17692_n5449), .Y(_abc_17692_n5692_1) );
  AND2X2 AND2X2_2194 ( .A(_abc_17692_n5696), .B(_abc_17692_n1846_bF_buf6), .Y(_abc_17692_n5697) );
  AND2X2 AND2X2_2195 ( .A(_abc_17692_n5697), .B(_abc_17692_n5694), .Y(_abc_17692_n5698) );
  AND2X2 AND2X2_2196 ( .A(sum_19_), .B(\key_in[19] ), .Y(_abc_17692_n5701) );
  AND2X2 AND2X2_2197 ( .A(_abc_17692_n5702), .B(_abc_17692_n5703), .Y(_abc_17692_n5704) );
  AND2X2 AND2X2_2198 ( .A(_abc_17692_n5700), .B(_abc_17692_n5704), .Y(_abc_17692_n5705) );
  AND2X2 AND2X2_2199 ( .A(_abc_17692_n5710), .B(_abc_17692_n5706), .Y(_abc_17692_n5711) );
  AND2X2 AND2X2_22 ( .A(_abc_17692_n675), .B(x_3_), .Y(_abc_17692_n679) );
  AND2X2 AND2X2_220 ( .A(_abc_17692_n723), .B(sum_11_), .Y(_abc_17692_n1193) );
  AND2X2 AND2X2_2200 ( .A(_abc_17692_n5709), .B(_abc_17692_n5712), .Y(_abc_17692_n5713) );
  AND2X2 AND2X2_2201 ( .A(_abc_17692_n5715), .B(_abc_17692_n5716), .Y(_abc_17692_n5717) );
  AND2X2 AND2X2_2202 ( .A(_abc_17692_n5714), .B(_abc_17692_n5718), .Y(_abc_17692_n5719) );
  AND2X2 AND2X2_2203 ( .A(_abc_17692_n5570), .B(_abc_17692_n5487), .Y(_abc_17692_n5721) );
  AND2X2 AND2X2_2204 ( .A(_abc_17692_n5724), .B(_abc_17692_n1830_bF_buf6), .Y(_abc_17692_n5725) );
  AND2X2 AND2X2_2205 ( .A(_abc_17692_n5725), .B(_abc_17692_n5722), .Y(_abc_17692_n5726) );
  AND2X2 AND2X2_2206 ( .A(_abc_17692_n5729), .B(state_7_bF_buf4), .Y(_abc_17692_n5730) );
  AND2X2 AND2X2_2207 ( .A(_abc_17692_n5540), .B(_abc_17692_n5731), .Y(_abc_17692_n5732) );
  AND2X2 AND2X2_2208 ( .A(_abc_17692_n5733), .B(_abc_17692_n5666), .Y(_abc_17692_n5734) );
  AND2X2 AND2X2_2209 ( .A(_abc_17692_n5732), .B(_abc_17692_n5659), .Y(_abc_17692_n5735) );
  AND2X2 AND2X2_221 ( .A(_abc_17692_n1151), .B(sum_10_), .Y(_abc_17692_n1194) );
  AND2X2 AND2X2_2210 ( .A(_abc_17692_n5426), .B(_abc_17692_n5417), .Y(_abc_17692_n5738) );
  AND2X2 AND2X2_2211 ( .A(_abc_17692_n5741), .B(_abc_17692_n1877_bF_buf5), .Y(_abc_17692_n5742) );
  AND2X2 AND2X2_2212 ( .A(_abc_17692_n5742), .B(_abc_17692_n5740), .Y(_abc_17692_n5743) );
  AND2X2 AND2X2_2213 ( .A(_abc_17692_n5486), .B(workunit2_18_), .Y(_abc_17692_n5744) );
  AND2X2 AND2X2_2214 ( .A(_abc_17692_n5748_1), .B(_abc_17692_n1830_bF_buf5), .Y(_abc_17692_n5749) );
  AND2X2 AND2X2_2215 ( .A(_abc_17692_n5749), .B(_abc_17692_n5747), .Y(_abc_17692_n5750) );
  AND2X2 AND2X2_2216 ( .A(_abc_17692_n5448), .B(workunit2_18_), .Y(_abc_17692_n5751) );
  AND2X2 AND2X2_2217 ( .A(_abc_17692_n5463), .B(_abc_17692_n5752), .Y(_abc_17692_n5753) );
  AND2X2 AND2X2_2218 ( .A(_abc_17692_n5756), .B(_abc_17692_n1846_bF_buf5), .Y(_abc_17692_n5757) );
  AND2X2 AND2X2_2219 ( .A(_abc_17692_n5757), .B(_abc_17692_n5755), .Y(_abc_17692_n5758) );
  AND2X2 AND2X2_222 ( .A(_abc_17692_n1172), .B(_abc_17692_n1195_1), .Y(_abc_17692_n1196) );
  AND2X2 AND2X2_2220 ( .A(_abc_17692_n5761), .B(state_6_bF_buf0), .Y(_abc_17692_n5762) );
  AND2X2 AND2X2_2221 ( .A(_abc_17692_n5762), .B(_abc_17692_n5737), .Y(_abc_17692_n5763) );
  AND2X2 AND2X2_2222 ( .A(_abc_17692_n1885_bF_buf0), .B(workunit2_19_), .Y(_abc_17692_n5764) );
  AND2X2 AND2X2_2223 ( .A(state_8_bF_buf0), .B(\data_in2[19] ), .Y(_abc_17692_n5765) );
  AND2X2 AND2X2_2224 ( .A(_abc_17692_n5385), .B(_abc_17692_n5606), .Y(_abc_17692_n5770) );
  AND2X2 AND2X2_2225 ( .A(_abc_17692_n5388), .B(_abc_17692_n5770), .Y(_abc_17692_n5771) );
  AND2X2 AND2X2_2226 ( .A(_abc_17692_n4924), .B(_abc_17692_n5771), .Y(_abc_17692_n5772) );
  AND2X2 AND2X2_2227 ( .A(_abc_17692_n5770), .B(_abc_17692_n5387), .Y(_abc_17692_n5773) );
  AND2X2 AND2X2_2228 ( .A(_abc_17692_n5775), .B(_abc_17692_n5603), .Y(_abc_17692_n5776) );
  AND2X2 AND2X2_2229 ( .A(_abc_17692_n5774), .B(_abc_17692_n5777), .Y(_abc_17692_n5778) );
  AND2X2 AND2X2_223 ( .A(_abc_17692_n1199), .B(state_15_bF_buf3), .Y(_abc_17692_n1200) );
  AND2X2 AND2X2_2230 ( .A(_abc_17692_n5781), .B(_abc_17692_n5783), .Y(_abc_17692_n5784) );
  AND2X2 AND2X2_2231 ( .A(_abc_17692_n5785), .B(workunit1_20_), .Y(_abc_17692_n5786) );
  AND2X2 AND2X2_2232 ( .A(_abc_17692_n5784), .B(_abc_17692_n4730), .Y(_abc_17692_n5787) );
  AND2X2 AND2X2_2233 ( .A(_abc_17692_n5780), .B(_abc_17692_n5789), .Y(_abc_17692_n5790) );
  AND2X2 AND2X2_2234 ( .A(_abc_17692_n5792), .B(_abc_17692_n5778), .Y(_abc_17692_n5793) );
  AND2X2 AND2X2_2235 ( .A(_abc_17692_n5793), .B(_abc_17692_n5788), .Y(_abc_17692_n5794) );
  AND2X2 AND2X2_2236 ( .A(_abc_17692_n5516), .B(_abc_17692_n5644), .Y(_abc_17692_n5796) );
  AND2X2 AND2X2_2237 ( .A(_abc_17692_n5506), .B(_abc_17692_n5796), .Y(_abc_17692_n5797) );
  AND2X2 AND2X2_2238 ( .A(_abc_17692_n5092), .B(_abc_17692_n5797), .Y(_abc_17692_n5798) );
  AND2X2 AND2X2_2239 ( .A(_abc_17692_n5511), .B(_abc_17692_n5796), .Y(_abc_17692_n5799) );
  AND2X2 AND2X2_224 ( .A(_abc_17692_n1200), .B(_abc_17692_n1197), .Y(_abc_17692_n1201) );
  AND2X2 AND2X2_2240 ( .A(_abc_17692_n5643), .B(_abc_17692_n5513), .Y(_abc_17692_n5800) );
  AND2X2 AND2X2_2241 ( .A(sum_20_), .B(\key_in[116] ), .Y(_abc_17692_n5804) );
  AND2X2 AND2X2_2242 ( .A(_abc_17692_n5805), .B(_abc_17692_n5806), .Y(_abc_17692_n5807) );
  AND2X2 AND2X2_2243 ( .A(_abc_17692_n5803), .B(_abc_17692_n5807), .Y(_abc_17692_n5808) );
  AND2X2 AND2X2_2244 ( .A(_abc_17692_n5809), .B(_abc_17692_n5810), .Y(_abc_17692_n5811) );
  AND2X2 AND2X2_2245 ( .A(_abc_17692_n5811), .B(_abc_17692_n5812), .Y(_abc_17692_n5813) );
  AND2X2 AND2X2_2246 ( .A(_abc_17692_n5816), .B(_abc_17692_n5818), .Y(_abc_17692_n5819) );
  AND2X2 AND2X2_2247 ( .A(_abc_17692_n5820), .B(_abc_17692_n5769), .Y(_abc_17692_n5821) );
  AND2X2 AND2X2_2248 ( .A(_abc_17692_n5819), .B(workunit2_20_), .Y(_abc_17692_n5822) );
  AND2X2 AND2X2_2249 ( .A(_abc_17692_n5659), .B(_abc_17692_n5530), .Y(_abc_17692_n5825) );
  AND2X2 AND2X2_225 ( .A(delta_12_), .B(sum_12_), .Y(_abc_17692_n1204) );
  AND2X2 AND2X2_2250 ( .A(_abc_17692_n5825), .B(_abc_17692_n5536), .Y(_abc_17692_n5826) );
  AND2X2 AND2X2_2251 ( .A(_abc_17692_n5535), .B(_abc_17692_n5825), .Y(_abc_17692_n5829) );
  AND2X2 AND2X2_2252 ( .A(_abc_17692_n5657), .B(workunit2_19_), .Y(_abc_17692_n5831) );
  AND2X2 AND2X2_2253 ( .A(_abc_17692_n5659), .B(_abc_17692_n5528), .Y(_abc_17692_n5832) );
  AND2X2 AND2X2_2254 ( .A(_abc_17692_n5830), .B(_abc_17692_n5834), .Y(_abc_17692_n5835) );
  AND2X2 AND2X2_2255 ( .A(_abc_17692_n5828), .B(_abc_17692_n5835), .Y(_abc_17692_n5836) );
  AND2X2 AND2X2_2256 ( .A(_abc_17692_n5837), .B(_abc_17692_n5824), .Y(_abc_17692_n5838) );
  AND2X2 AND2X2_2257 ( .A(_abc_17692_n5839), .B(_abc_17692_n5840), .Y(_abc_17692_n5841) );
  AND2X2 AND2X2_2258 ( .A(_abc_17692_n5398), .B(_abc_17692_n5616), .Y(_abc_17692_n5843_1) );
  AND2X2 AND2X2_2259 ( .A(_abc_17692_n5403), .B(_abc_17692_n5843_1), .Y(_abc_17692_n5844) );
  AND2X2 AND2X2_226 ( .A(_abc_17692_n1205), .B(_abc_17692_n1206_1), .Y(_abc_17692_n1207) );
  AND2X2 AND2X2_2260 ( .A(_abc_17692_n4955), .B(_abc_17692_n5844), .Y(_abc_17692_n5845) );
  AND2X2 AND2X2_2261 ( .A(_abc_17692_n5843_1), .B(_abc_17692_n5401), .Y(_abc_17692_n5846_1) );
  AND2X2 AND2X2_2262 ( .A(_abc_17692_n5615), .B(_abc_17692_n5395), .Y(_abc_17692_n5847) );
  AND2X2 AND2X2_2263 ( .A(sum_20_), .B(\key_in[84] ), .Y(_abc_17692_n5851) );
  AND2X2 AND2X2_2264 ( .A(_abc_17692_n5852), .B(_abc_17692_n5853), .Y(_abc_17692_n5854) );
  AND2X2 AND2X2_2265 ( .A(_abc_17692_n5850), .B(_abc_17692_n5854), .Y(_abc_17692_n5855) );
  AND2X2 AND2X2_2266 ( .A(_abc_17692_n5856), .B(_abc_17692_n5857), .Y(_abc_17692_n5858) );
  AND2X2 AND2X2_2267 ( .A(_abc_17692_n5861), .B(_abc_17692_n5862), .Y(_abc_17692_n5863) );
  AND2X2 AND2X2_2268 ( .A(_abc_17692_n5863), .B(workunit2_20_), .Y(_abc_17692_n5864) );
  AND2X2 AND2X2_2269 ( .A(_abc_17692_n5865), .B(_abc_17692_n5866), .Y(_abc_17692_n5867) );
  AND2X2 AND2X2_227 ( .A(_abc_17692_n1185), .B(_abc_17692_n1155), .Y(_abc_17692_n1210) );
  AND2X2 AND2X2_2270 ( .A(_abc_17692_n5629), .B(_abc_17692_n5419), .Y(_abc_17692_n5868) );
  AND2X2 AND2X2_2271 ( .A(_abc_17692_n5627), .B(workunit2_19_), .Y(_abc_17692_n5871) );
  AND2X2 AND2X2_2272 ( .A(_abc_17692_n5629), .B(_abc_17692_n5416), .Y(_abc_17692_n5872) );
  AND2X2 AND2X2_2273 ( .A(_abc_17692_n5870), .B(_abc_17692_n5874), .Y(_abc_17692_n5875) );
  AND2X2 AND2X2_2274 ( .A(_abc_17692_n5868), .B(_abc_17692_n5268), .Y(_abc_17692_n5876) );
  AND2X2 AND2X2_2275 ( .A(_abc_17692_n4982), .B(_abc_17692_n5876), .Y(_abc_17692_n5877) );
  AND2X2 AND2X2_2276 ( .A(_abc_17692_n5878), .B(_abc_17692_n5875), .Y(_abc_17692_n5879) );
  AND2X2 AND2X2_2277 ( .A(_abc_17692_n5880), .B(_abc_17692_n5867), .Y(_abc_17692_n5881) );
  AND2X2 AND2X2_2278 ( .A(_abc_17692_n5883), .B(_abc_17692_n1877_bF_buf4), .Y(_abc_17692_n5884) );
  AND2X2 AND2X2_2279 ( .A(_abc_17692_n5884), .B(_abc_17692_n5882), .Y(_abc_17692_n5885) );
  AND2X2 AND2X2_228 ( .A(_abc_17692_n1185), .B(_abc_17692_n1150), .Y(_abc_17692_n1214) );
  AND2X2 AND2X2_2280 ( .A(_abc_17692_n5477), .B(_abc_17692_n5704), .Y(_abc_17692_n5886) );
  AND2X2 AND2X2_2281 ( .A(_abc_17692_n5467), .B(_abc_17692_n5886), .Y(_abc_17692_n5887) );
  AND2X2 AND2X2_2282 ( .A(_abc_17692_n5044_1), .B(_abc_17692_n5887), .Y(_abc_17692_n5888) );
  AND2X2 AND2X2_2283 ( .A(_abc_17692_n5472), .B(_abc_17692_n5886), .Y(_abc_17692_n5889) );
  AND2X2 AND2X2_2284 ( .A(_abc_17692_n5703), .B(_abc_17692_n5474), .Y(_abc_17692_n5890) );
  AND2X2 AND2X2_2285 ( .A(sum_20_), .B(\key_in[20] ), .Y(_abc_17692_n5894) );
  AND2X2 AND2X2_2286 ( .A(_abc_17692_n5895), .B(_abc_17692_n5896), .Y(_abc_17692_n5897) );
  AND2X2 AND2X2_2287 ( .A(_abc_17692_n5893), .B(_abc_17692_n5897), .Y(_abc_17692_n5898) );
  AND2X2 AND2X2_2288 ( .A(_abc_17692_n5900_1), .B(_abc_17692_n5901), .Y(_abc_17692_n5902) );
  AND2X2 AND2X2_2289 ( .A(_abc_17692_n5902), .B(_abc_17692_n5903_1), .Y(_abc_17692_n5904) );
  AND2X2 AND2X2_229 ( .A(delta_11_), .B(sum_11_), .Y(_abc_17692_n1215) );
  AND2X2 AND2X2_2290 ( .A(_abc_17692_n5908), .B(_abc_17692_n5907), .Y(_abc_17692_n5909) );
  AND2X2 AND2X2_2291 ( .A(_abc_17692_n5910), .B(_abc_17692_n5769), .Y(_abc_17692_n5911) );
  AND2X2 AND2X2_2292 ( .A(_abc_17692_n5909), .B(workunit2_20_), .Y(_abc_17692_n5912) );
  AND2X2 AND2X2_2293 ( .A(_abc_17692_n5720), .B(_abc_17692_n5491), .Y(_abc_17692_n5914) );
  AND2X2 AND2X2_2294 ( .A(_abc_17692_n5713), .B(workunit2_19_), .Y(_abc_17692_n5917) );
  AND2X2 AND2X2_2295 ( .A(_abc_17692_n5720), .B(_abc_17692_n5744), .Y(_abc_17692_n5919) );
  AND2X2 AND2X2_2296 ( .A(_abc_17692_n5920), .B(_abc_17692_n5918), .Y(_abc_17692_n5921) );
  AND2X2 AND2X2_2297 ( .A(_abc_17692_n5916), .B(_abc_17692_n5921), .Y(_abc_17692_n5922) );
  AND2X2 AND2X2_2298 ( .A(_abc_17692_n5914), .B(_abc_17692_n5496), .Y(_abc_17692_n5923) );
  AND2X2 AND2X2_2299 ( .A(_abc_17692_n5925), .B(_abc_17692_n5922), .Y(_abc_17692_n5926) );
  AND2X2 AND2X2_23 ( .A(_abc_17692_n680), .B(_abc_17692_n681), .Y(x_3__FF_INPUT) );
  AND2X2 AND2X2_230 ( .A(_abc_17692_n1213), .B(_abc_17692_n1217), .Y(_abc_17692_n1218) );
  AND2X2 AND2X2_2300 ( .A(_abc_17692_n5930), .B(_abc_17692_n1830_bF_buf4), .Y(_abc_17692_n5931) );
  AND2X2 AND2X2_2301 ( .A(_abc_17692_n5931), .B(_abc_17692_n5927), .Y(_abc_17692_n5932) );
  AND2X2 AND2X2_2302 ( .A(_abc_17692_n5434), .B(_abc_17692_n5676), .Y(_abc_17692_n5933) );
  AND2X2 AND2X2_2303 ( .A(_abc_17692_n5437), .B(_abc_17692_n5933), .Y(_abc_17692_n5934) );
  AND2X2 AND2X2_2304 ( .A(_abc_17692_n4998), .B(_abc_17692_n5934), .Y(_abc_17692_n5935) );
  AND2X2 AND2X2_2305 ( .A(_abc_17692_n5933), .B(_abc_17692_n5436), .Y(_abc_17692_n5936) );
  AND2X2 AND2X2_2306 ( .A(_abc_17692_n5675), .B(_abc_17692_n5431), .Y(_abc_17692_n5937) );
  AND2X2 AND2X2_2307 ( .A(sum_20_), .B(\key_in[52] ), .Y(_abc_17692_n5941) );
  AND2X2 AND2X2_2308 ( .A(_abc_17692_n5942), .B(_abc_17692_n5943), .Y(_abc_17692_n5944) );
  AND2X2 AND2X2_2309 ( .A(_abc_17692_n5940), .B(_abc_17692_n5944), .Y(_abc_17692_n5945) );
  AND2X2 AND2X2_231 ( .A(_abc_17692_n1212), .B(_abc_17692_n1218), .Y(_abc_17692_n1219) );
  AND2X2 AND2X2_2310 ( .A(_abc_17692_n5947), .B(_abc_17692_n5948), .Y(_abc_17692_n5949) );
  AND2X2 AND2X2_2311 ( .A(_abc_17692_n5949), .B(_abc_17692_n5950), .Y(_abc_17692_n5951) );
  AND2X2 AND2X2_2312 ( .A(_abc_17692_n5955), .B(_abc_17692_n5954), .Y(_abc_17692_n5956) );
  AND2X2 AND2X2_2313 ( .A(_abc_17692_n5957), .B(_abc_17692_n5769), .Y(_abc_17692_n5958) );
  AND2X2 AND2X2_2314 ( .A(_abc_17692_n5956), .B(workunit2_20_), .Y(_abc_17692_n5959) );
  AND2X2 AND2X2_2315 ( .A(_abc_17692_n5685), .B(workunit2_19_), .Y(_abc_17692_n5963) );
  AND2X2 AND2X2_2316 ( .A(_abc_17692_n5965), .B(_abc_17692_n5964), .Y(_abc_17692_n5966) );
  AND2X2 AND2X2_2317 ( .A(_abc_17692_n5962), .B(_abc_17692_n5966), .Y(_abc_17692_n5967) );
  AND2X2 AND2X2_2318 ( .A(_abc_17692_n5968), .B(_abc_17692_n5459), .Y(_abc_17692_n5969) );
  AND2X2 AND2X2_2319 ( .A(_abc_17692_n5971), .B(_abc_17692_n5967), .Y(_abc_17692_n5972) );
  AND2X2 AND2X2_232 ( .A(_abc_17692_n1222), .B(state_3_bF_buf2), .Y(_abc_17692_n1223_1) );
  AND2X2 AND2X2_2320 ( .A(_abc_17692_n5976), .B(_abc_17692_n1846_bF_buf4), .Y(_abc_17692_n5977) );
  AND2X2 AND2X2_2321 ( .A(_abc_17692_n5977), .B(_abc_17692_n5973), .Y(_abc_17692_n5978) );
  AND2X2 AND2X2_2322 ( .A(_abc_17692_n5981_1), .B(state_6_bF_buf4), .Y(_abc_17692_n5982) );
  AND2X2 AND2X2_2323 ( .A(_abc_17692_n5982), .B(_abc_17692_n5842), .Y(_abc_17692_n5983) );
  AND2X2 AND2X2_2324 ( .A(_abc_17692_n5666), .B(_abc_17692_n5529), .Y(_abc_17692_n5984_1) );
  AND2X2 AND2X2_2325 ( .A(_abc_17692_n5984_1), .B(_abc_17692_n5547), .Y(_abc_17692_n5985) );
  AND2X2 AND2X2_2326 ( .A(_abc_17692_n5986), .B(_abc_17692_n5664), .Y(_abc_17692_n5987) );
  AND2X2 AND2X2_2327 ( .A(_abc_17692_n5984_1), .B(_abc_17692_n5548_1), .Y(_abc_17692_n5990) );
  AND2X2 AND2X2_2328 ( .A(_abc_17692_n5139), .B(_abc_17692_n5990), .Y(_abc_17692_n5991) );
  AND2X2 AND2X2_2329 ( .A(_abc_17692_n5992), .B(_abc_17692_n5823), .Y(_abc_17692_n5994) );
  AND2X2 AND2X2_233 ( .A(_abc_17692_n1223_1), .B(_abc_17692_n1221), .Y(_abc_17692_n1224) );
  AND2X2 AND2X2_2330 ( .A(_abc_17692_n5995), .B(_abc_17692_n1863_bF_buf2), .Y(_abc_17692_n5996) );
  AND2X2 AND2X2_2331 ( .A(_abc_17692_n5996), .B(_abc_17692_n5993), .Y(_abc_17692_n5997) );
  AND2X2 AND2X2_2332 ( .A(_abc_17692_n5259), .B(_abc_17692_n5342), .Y(_abc_17692_n5999) );
  AND2X2 AND2X2_2333 ( .A(_abc_17692_n6005), .B(_abc_17692_n6003), .Y(_abc_17692_n6006) );
  AND2X2 AND2X2_2334 ( .A(_abc_17692_n6002), .B(_abc_17692_n6006), .Y(_abc_17692_n6007) );
  AND2X2 AND2X2_2335 ( .A(_abc_17692_n5264), .B(_abc_17692_n5145), .Y(_abc_17692_n6008) );
  AND2X2 AND2X2_2336 ( .A(_abc_17692_n6009), .B(_abc_17692_n6008), .Y(_abc_17692_n6010) );
  AND2X2 AND2X2_2337 ( .A(_abc_17692_n6012), .B(_abc_17692_n6007), .Y(_abc_17692_n6013) );
  AND2X2 AND2X2_2338 ( .A(_abc_17692_n6014), .B(_abc_17692_n5998), .Y(_abc_17692_n6015) );
  AND2X2 AND2X2_2339 ( .A(_abc_17692_n6017), .B(_abc_17692_n1877_bF_buf3), .Y(_abc_17692_n6018) );
  AND2X2 AND2X2_234 ( .A(_abc_17692_n1184), .B(_abc_17692_n1154), .Y(_abc_17692_n1225) );
  AND2X2 AND2X2_2340 ( .A(_abc_17692_n6018), .B(_abc_17692_n6016), .Y(_abc_17692_n6019) );
  AND2X2 AND2X2_2341 ( .A(_abc_17692_n5691), .B(_abc_17692_n5452), .Y(_abc_17692_n6020) );
  AND2X2 AND2X2_2342 ( .A(_abc_17692_n6020), .B(_abc_17692_n5577), .Y(_abc_17692_n6021) );
  AND2X2 AND2X2_2343 ( .A(_abc_17692_n5690), .B(_abc_17692_n6023), .Y(_abc_17692_n6024) );
  AND2X2 AND2X2_2344 ( .A(_abc_17692_n6020), .B(_abc_17692_n5578), .Y(_abc_17692_n6028) );
  AND2X2 AND2X2_2345 ( .A(_abc_17692_n5172), .B(_abc_17692_n6028), .Y(_abc_17692_n6029) );
  AND2X2 AND2X2_2346 ( .A(_abc_17692_n6030), .B(_abc_17692_n6027), .Y(_abc_17692_n6031) );
  AND2X2 AND2X2_2347 ( .A(_abc_17692_n6032), .B(_abc_17692_n5960), .Y(_abc_17692_n6034) );
  AND2X2 AND2X2_2348 ( .A(_abc_17692_n6035), .B(_abc_17692_n1846_bF_buf3), .Y(_abc_17692_n6036) );
  AND2X2 AND2X2_2349 ( .A(_abc_17692_n6036), .B(_abc_17692_n6033), .Y(_abc_17692_n6037) );
  AND2X2 AND2X2_235 ( .A(_abc_17692_n1167), .B(_abc_17692_n1225), .Y(_abc_17692_n1226) );
  AND2X2 AND2X2_2350 ( .A(_abc_17692_n5719), .B(_abc_17692_n5490), .Y(_abc_17692_n6038_1) );
  AND2X2 AND2X2_2351 ( .A(_abc_17692_n6038_1), .B(_abc_17692_n5565), .Y(_abc_17692_n6039) );
  AND2X2 AND2X2_2352 ( .A(_abc_17692_n5718), .B(_abc_17692_n6041_1), .Y(_abc_17692_n6042) );
  AND2X2 AND2X2_2353 ( .A(_abc_17692_n6038_1), .B(_abc_17692_n5566), .Y(_abc_17692_n6045) );
  AND2X2 AND2X2_2354 ( .A(_abc_17692_n5187), .B(_abc_17692_n6045), .Y(_abc_17692_n6046) );
  AND2X2 AND2X2_2355 ( .A(_abc_17692_n6047), .B(_abc_17692_n5913), .Y(_abc_17692_n6048) );
  AND2X2 AND2X2_2356 ( .A(_abc_17692_n6050), .B(_abc_17692_n1830_bF_buf3), .Y(_abc_17692_n6051) );
  AND2X2 AND2X2_2357 ( .A(_abc_17692_n6051), .B(_abc_17692_n6049), .Y(_abc_17692_n6052) );
  AND2X2 AND2X2_2358 ( .A(_abc_17692_n6055), .B(state_7_bF_buf3), .Y(_abc_17692_n6056) );
  AND2X2 AND2X2_2359 ( .A(_abc_17692_n1885_bF_buf4), .B(workunit2_20_), .Y(_abc_17692_n6057) );
  AND2X2 AND2X2_236 ( .A(_abc_17692_n1228), .B(_abc_17692_n1183), .Y(_abc_17692_n1229) );
  AND2X2 AND2X2_2360 ( .A(state_8_bF_buf9), .B(\data_in2[20] ), .Y(_abc_17692_n6058) );
  AND2X2 AND2X2_2361 ( .A(_abc_17692_n6064), .B(_abc_17692_n6066), .Y(_abc_17692_n6067) );
  AND2X2 AND2X2_2362 ( .A(_abc_17692_n6068), .B(workunit1_21_), .Y(_abc_17692_n6069) );
  AND2X2 AND2X2_2363 ( .A(_abc_17692_n6067), .B(_abc_17692_n4926), .Y(_abc_17692_n6071) );
  AND2X2 AND2X2_2364 ( .A(_abc_17692_n6070), .B(_abc_17692_n6072), .Y(_abc_17692_n6073) );
  AND2X2 AND2X2_2365 ( .A(_abc_17692_n6063), .B(_abc_17692_n6073), .Y(_abc_17692_n6074) );
  AND2X2 AND2X2_2366 ( .A(_abc_17692_n6075), .B(_abc_17692_n6076), .Y(_abc_17692_n6077) );
  AND2X2 AND2X2_2367 ( .A(sum_21_), .B(\key_in[85] ), .Y(_abc_17692_n6080) );
  AND2X2 AND2X2_2368 ( .A(_abc_17692_n6081), .B(_abc_17692_n6082), .Y(_abc_17692_n6083) );
  AND2X2 AND2X2_2369 ( .A(_abc_17692_n6079), .B(_abc_17692_n6083), .Y(_abc_17692_n6084) );
  AND2X2 AND2X2_237 ( .A(_abc_17692_n1227), .B(_abc_17692_n1229), .Y(_abc_17692_n1230) );
  AND2X2 AND2X2_2370 ( .A(_abc_17692_n6078), .B(_abc_17692_n6085), .Y(_abc_17692_n6086) );
  AND2X2 AND2X2_2371 ( .A(_abc_17692_n6092), .B(_abc_17692_n6089), .Y(_abc_17692_n6093) );
  AND2X2 AND2X2_2372 ( .A(_abc_17692_n6093), .B(workunit2_21_), .Y(_abc_17692_n6094) );
  AND2X2 AND2X2_2373 ( .A(_abc_17692_n6096), .B(_abc_17692_n6095), .Y(_abc_17692_n6097) );
  AND2X2 AND2X2_2374 ( .A(_abc_17692_n5882), .B(_abc_17692_n5865), .Y(_abc_17692_n6099) );
  AND2X2 AND2X2_2375 ( .A(_abc_17692_n6103), .B(_abc_17692_n1877_bF_buf2), .Y(_abc_17692_n6104) );
  AND2X2 AND2X2_2376 ( .A(_abc_17692_n6104), .B(_abc_17692_n6101), .Y(_abc_17692_n6105) );
  AND2X2 AND2X2_2377 ( .A(sum_21_), .B(\key_in[21] ), .Y(_abc_17692_n6107) );
  AND2X2 AND2X2_2378 ( .A(_abc_17692_n6108), .B(_abc_17692_n6109), .Y(_abc_17692_n6110) );
  AND2X2 AND2X2_2379 ( .A(_abc_17692_n6106), .B(_abc_17692_n6111), .Y(_abc_17692_n6113) );
  AND2X2 AND2X2_238 ( .A(_abc_17692_n1136), .B(_abc_17692_n1225), .Y(_abc_17692_n1231) );
  AND2X2 AND2X2_2380 ( .A(_abc_17692_n6114), .B(_abc_17692_n6112), .Y(_abc_17692_n6115) );
  AND2X2 AND2X2_2381 ( .A(_abc_17692_n6091), .B(_abc_17692_n6116), .Y(_abc_17692_n6117) );
  AND2X2 AND2X2_2382 ( .A(_abc_17692_n6077), .B(_abc_17692_n6115), .Y(_abc_17692_n6118) );
  AND2X2 AND2X2_2383 ( .A(_abc_17692_n6120), .B(workunit2_21_), .Y(_abc_17692_n6121) );
  AND2X2 AND2X2_2384 ( .A(_abc_17692_n6119), .B(_abc_17692_n6095), .Y(_abc_17692_n6122) );
  AND2X2 AND2X2_2385 ( .A(_abc_17692_n5927), .B(_abc_17692_n6124), .Y(_abc_17692_n6125) );
  AND2X2 AND2X2_2386 ( .A(_abc_17692_n6128), .B(_abc_17692_n6129), .Y(_abc_17692_n6130) );
  AND2X2 AND2X2_2387 ( .A(_abc_17692_n6131), .B(_abc_17692_n1830_bF_buf2), .Y(_abc_17692_n6132) );
  AND2X2 AND2X2_2388 ( .A(_abc_17692_n6132), .B(_abc_17692_n6127), .Y(_abc_17692_n6133) );
  AND2X2 AND2X2_2389 ( .A(sum_21_), .B(\key_in[53] ), .Y(_abc_17692_n6136) );
  AND2X2 AND2X2_239 ( .A(_abc_17692_n1232), .B(_abc_17692_n1230), .Y(_abc_17692_n1233) );
  AND2X2 AND2X2_2390 ( .A(_abc_17692_n6137), .B(_abc_17692_n6138), .Y(_abc_17692_n6139) );
  AND2X2 AND2X2_2391 ( .A(_abc_17692_n6135), .B(_abc_17692_n6139), .Y(_abc_17692_n6140) );
  AND2X2 AND2X2_2392 ( .A(_abc_17692_n6141), .B(_abc_17692_n6142), .Y(_abc_17692_n6143) );
  AND2X2 AND2X2_2393 ( .A(_abc_17692_n6091), .B(_abc_17692_n6144), .Y(_abc_17692_n6145) );
  AND2X2 AND2X2_2394 ( .A(_abc_17692_n6077), .B(_abc_17692_n6143), .Y(_abc_17692_n6146) );
  AND2X2 AND2X2_2395 ( .A(_abc_17692_n6150), .B(_abc_17692_n6149), .Y(_abc_17692_n6151) );
  AND2X2 AND2X2_2396 ( .A(_abc_17692_n6152), .B(_abc_17692_n6148), .Y(_abc_17692_n6153) );
  AND2X2 AND2X2_2397 ( .A(_abc_17692_n5973), .B(_abc_17692_n6155), .Y(_abc_17692_n6156) );
  AND2X2 AND2X2_2398 ( .A(_abc_17692_n6159), .B(_abc_17692_n1846_bF_buf2), .Y(_abc_17692_n6160) );
  AND2X2 AND2X2_2399 ( .A(_abc_17692_n6160), .B(_abc_17692_n6158), .Y(_abc_17692_n6161) );
  AND2X2 AND2X2_24 ( .A(_abc_17692_n679), .B(x_4_), .Y(_abc_17692_n683) );
  AND2X2 AND2X2_240 ( .A(_abc_17692_n1234), .B(_abc_17692_n1208), .Y(_abc_17692_n1235) );
  AND2X2 AND2X2_2400 ( .A(sum_21_), .B(\key_in[117] ), .Y(_abc_17692_n6166_1) );
  AND2X2 AND2X2_2401 ( .A(_abc_17692_n6167), .B(_abc_17692_n6168), .Y(_abc_17692_n6169_1) );
  AND2X2 AND2X2_2402 ( .A(_abc_17692_n6165), .B(_abc_17692_n6170), .Y(_abc_17692_n6172) );
  AND2X2 AND2X2_2403 ( .A(_abc_17692_n6173), .B(_abc_17692_n6171), .Y(_abc_17692_n6174) );
  AND2X2 AND2X2_2404 ( .A(_abc_17692_n6177), .B(_abc_17692_n6175), .Y(_abc_17692_n6178) );
  AND2X2 AND2X2_2405 ( .A(_abc_17692_n6178), .B(workunit2_21_), .Y(_abc_17692_n6179) );
  AND2X2 AND2X2_2406 ( .A(_abc_17692_n6181), .B(_abc_17692_n6095), .Y(_abc_17692_n6182) );
  AND2X2 AND2X2_2407 ( .A(_abc_17692_n6183), .B(_abc_17692_n6180), .Y(_abc_17692_n6184) );
  AND2X2 AND2X2_2408 ( .A(_abc_17692_n5839), .B(_abc_17692_n6185), .Y(_abc_17692_n6186) );
  AND2X2 AND2X2_2409 ( .A(_abc_17692_n6187), .B(_abc_17692_n6184), .Y(_abc_17692_n6188) );
  AND2X2 AND2X2_241 ( .A(_abc_17692_n1237), .B(state_15_bF_buf2), .Y(_abc_17692_n1238) );
  AND2X2 AND2X2_2410 ( .A(_abc_17692_n6186), .B(_abc_17692_n6189), .Y(_abc_17692_n6190) );
  AND2X2 AND2X2_2411 ( .A(_abc_17692_n6192), .B(state_6_bF_buf3), .Y(_abc_17692_n6193) );
  AND2X2 AND2X2_2412 ( .A(_abc_17692_n6193), .B(_abc_17692_n6164), .Y(_abc_17692_n6194) );
  AND2X2 AND2X2_2413 ( .A(_abc_17692_n5820), .B(workunit2_20_), .Y(_abc_17692_n6195) );
  AND2X2 AND2X2_2414 ( .A(_abc_17692_n5995), .B(_abc_17692_n6196), .Y(_abc_17692_n6197) );
  AND2X2 AND2X2_2415 ( .A(_abc_17692_n6200), .B(_abc_17692_n1863_bF_buf0), .Y(_abc_17692_n6201) );
  AND2X2 AND2X2_2416 ( .A(_abc_17692_n6201), .B(_abc_17692_n6198), .Y(_abc_17692_n6202) );
  AND2X2 AND2X2_2417 ( .A(_abc_17692_n6203), .B(workunit2_20_), .Y(_abc_17692_n6204) );
  AND2X2 AND2X2_2418 ( .A(_abc_17692_n6016), .B(_abc_17692_n6205), .Y(_abc_17692_n6206) );
  AND2X2 AND2X2_2419 ( .A(_abc_17692_n6209), .B(_abc_17692_n1877_bF_buf1), .Y(_abc_17692_n6210) );
  AND2X2 AND2X2_242 ( .A(_abc_17692_n1238), .B(_abc_17692_n1236), .Y(_abc_17692_n1239) );
  AND2X2 AND2X2_2420 ( .A(_abc_17692_n6210), .B(_abc_17692_n6207), .Y(_abc_17692_n6211) );
  AND2X2 AND2X2_2421 ( .A(_abc_17692_n5910), .B(workunit2_20_), .Y(_abc_17692_n6212) );
  AND2X2 AND2X2_2422 ( .A(_abc_17692_n6049), .B(_abc_17692_n6213), .Y(_abc_17692_n6214) );
  AND2X2 AND2X2_2423 ( .A(_abc_17692_n6217), .B(_abc_17692_n1830_bF_buf1), .Y(_abc_17692_n6218) );
  AND2X2 AND2X2_2424 ( .A(_abc_17692_n6218), .B(_abc_17692_n6215), .Y(_abc_17692_n6219) );
  AND2X2 AND2X2_2425 ( .A(_abc_17692_n5957), .B(workunit2_20_), .Y(_abc_17692_n6220) );
  AND2X2 AND2X2_2426 ( .A(_abc_17692_n6224), .B(_abc_17692_n1846_bF_buf1), .Y(_abc_17692_n6225_1) );
  AND2X2 AND2X2_2427 ( .A(_abc_17692_n6225_1), .B(_abc_17692_n6222_1), .Y(_abc_17692_n6226) );
  AND2X2 AND2X2_2428 ( .A(_abc_17692_n6229), .B(state_7_bF_buf2), .Y(_abc_17692_n6230) );
  AND2X2 AND2X2_2429 ( .A(_abc_17692_n1885_bF_buf3), .B(workunit2_21_), .Y(_abc_17692_n6231) );
  AND2X2 AND2X2_243 ( .A(_abc_17692_n722_bF_buf2), .B(sum_12_), .Y(_abc_17692_n1240) );
  AND2X2 AND2X2_2430 ( .A(state_8_bF_buf8), .B(\data_in2[21] ), .Y(_abc_17692_n6232) );
  AND2X2 AND2X2_2431 ( .A(_abc_17692_n5789), .B(_abc_17692_n6073), .Y(_abc_17692_n6236) );
  AND2X2 AND2X2_2432 ( .A(_abc_17692_n5780), .B(_abc_17692_n6236), .Y(_abc_17692_n6237) );
  AND2X2 AND2X2_2433 ( .A(_abc_17692_n6072), .B(_abc_17692_n5786), .Y(_abc_17692_n6238) );
  AND2X2 AND2X2_2434 ( .A(_abc_17692_n6241), .B(_abc_17692_n6243), .Y(_abc_17692_n6244) );
  AND2X2 AND2X2_2435 ( .A(_abc_17692_n6245), .B(workunit1_22_), .Y(_abc_17692_n6246) );
  AND2X2 AND2X2_2436 ( .A(_abc_17692_n6244), .B(_abc_17692_n5205), .Y(_abc_17692_n6247) );
  AND2X2 AND2X2_2437 ( .A(_abc_17692_n6240), .B(_abc_17692_n6249), .Y(_abc_17692_n6250) );
  AND2X2 AND2X2_2438 ( .A(_abc_17692_n6252), .B(_abc_17692_n6253), .Y(_abc_17692_n6254) );
  AND2X2 AND2X2_2439 ( .A(_abc_17692_n6254), .B(_abc_17692_n6248), .Y(_abc_17692_n6255) );
  AND2X2 AND2X2_244 ( .A(delta_13_), .B(sum_13_), .Y(_abc_17692_n1244) );
  AND2X2 AND2X2_2440 ( .A(_abc_17692_n5854), .B(_abc_17692_n6083), .Y(_abc_17692_n6257) );
  AND2X2 AND2X2_2441 ( .A(_abc_17692_n5850), .B(_abc_17692_n6257), .Y(_abc_17692_n6258) );
  AND2X2 AND2X2_2442 ( .A(_abc_17692_n5852), .B(_abc_17692_n6081), .Y(_abc_17692_n6261) );
  AND2X2 AND2X2_2443 ( .A(_abc_17692_n6259), .B(_abc_17692_n6262), .Y(_abc_17692_n6263) );
  AND2X2 AND2X2_2444 ( .A(sum_22_), .B(\key_in[86] ), .Y(_abc_17692_n6265) );
  AND2X2 AND2X2_2445 ( .A(_abc_17692_n6266), .B(_abc_17692_n6267), .Y(_abc_17692_n6268) );
  AND2X2 AND2X2_2446 ( .A(_abc_17692_n6264), .B(_abc_17692_n6268), .Y(_abc_17692_n6269) );
  AND2X2 AND2X2_2447 ( .A(_abc_17692_n6263), .B(_abc_17692_n6270), .Y(_abc_17692_n6271) );
  AND2X2 AND2X2_2448 ( .A(_abc_17692_n6274), .B(_abc_17692_n6276), .Y(_abc_17692_n6277) );
  AND2X2 AND2X2_2449 ( .A(_abc_17692_n6277), .B(workunit2_22_), .Y(_abc_17692_n6278) );
  AND2X2 AND2X2_245 ( .A(_abc_17692_n1246), .B(_abc_17692_n1247), .Y(_abc_17692_n1248) );
  AND2X2 AND2X2_2450 ( .A(_abc_17692_n6279), .B(_abc_17692_n6280), .Y(_abc_17692_n6281) );
  AND2X2 AND2X2_2451 ( .A(_abc_17692_n6096), .B(workunit2_21_), .Y(_abc_17692_n6282) );
  AND2X2 AND2X2_2452 ( .A(_abc_17692_n6098), .B(_abc_17692_n5864), .Y(_abc_17692_n6283) );
  AND2X2 AND2X2_2453 ( .A(_abc_17692_n6098), .B(_abc_17692_n5867), .Y(_abc_17692_n6285) );
  AND2X2 AND2X2_2454 ( .A(_abc_17692_n5880), .B(_abc_17692_n6285), .Y(_abc_17692_n6286) );
  AND2X2 AND2X2_2455 ( .A(_abc_17692_n6287), .B(_abc_17692_n6281), .Y(_abc_17692_n6288) );
  AND2X2 AND2X2_2456 ( .A(_abc_17692_n6290), .B(_abc_17692_n1877_bF_buf0), .Y(_abc_17692_n6291) );
  AND2X2 AND2X2_2457 ( .A(_abc_17692_n6291), .B(_abc_17692_n6289), .Y(_abc_17692_n6292) );
  AND2X2 AND2X2_2458 ( .A(_abc_17692_n5897), .B(_abc_17692_n6110), .Y(_abc_17692_n6294) );
  AND2X2 AND2X2_2459 ( .A(_abc_17692_n5893), .B(_abc_17692_n6294), .Y(_abc_17692_n6295) );
  AND2X2 AND2X2_246 ( .A(_abc_17692_n1249), .B(_abc_17692_n1245), .Y(_abc_17692_n1250) );
  AND2X2 AND2X2_2460 ( .A(_abc_17692_n5895), .B(_abc_17692_n6108), .Y(_abc_17692_n6297) );
  AND2X2 AND2X2_2461 ( .A(sum_22_), .B(\key_in[22] ), .Y(_abc_17692_n6301) );
  AND2X2 AND2X2_2462 ( .A(_abc_17692_n6302), .B(_abc_17692_n6303), .Y(_abc_17692_n6304) );
  AND2X2 AND2X2_2463 ( .A(_abc_17692_n6300), .B(_abc_17692_n6304), .Y(_abc_17692_n6305) );
  AND2X2 AND2X2_2464 ( .A(_abc_17692_n6307), .B(_abc_17692_n6298), .Y(_abc_17692_n6308) );
  AND2X2 AND2X2_2465 ( .A(_abc_17692_n6308), .B(_abc_17692_n6309), .Y(_abc_17692_n6310) );
  AND2X2 AND2X2_2466 ( .A(_abc_17692_n6275), .B(_abc_17692_n6311), .Y(_abc_17692_n6312) );
  AND2X2 AND2X2_2467 ( .A(_abc_17692_n6313), .B(_abc_17692_n6256), .Y(_abc_17692_n6314) );
  AND2X2 AND2X2_2468 ( .A(_abc_17692_n6317), .B(_abc_17692_n6318), .Y(_abc_17692_n6319_1) );
  AND2X2 AND2X2_2469 ( .A(_abc_17692_n6119), .B(workunit2_21_), .Y(_abc_17692_n6321) );
  AND2X2 AND2X2_247 ( .A(_abc_17692_n1222), .B(_abc_17692_n1252), .Y(_abc_17692_n1253) );
  AND2X2 AND2X2_2470 ( .A(_abc_17692_n6123), .B(_abc_17692_n5912), .Y(_abc_17692_n6322) );
  AND2X2 AND2X2_2471 ( .A(_abc_17692_n6123), .B(_abc_17692_n5928), .Y(_abc_17692_n6324) );
  AND2X2 AND2X2_2472 ( .A(_abc_17692_n5929), .B(_abc_17692_n6324), .Y(_abc_17692_n6325) );
  AND2X2 AND2X2_2473 ( .A(_abc_17692_n6326), .B(_abc_17692_n6320), .Y(_abc_17692_n6327) );
  AND2X2 AND2X2_2474 ( .A(_abc_17692_n6329), .B(_abc_17692_n1830_bF_buf0), .Y(_abc_17692_n6330) );
  AND2X2 AND2X2_2475 ( .A(_abc_17692_n6330), .B(_abc_17692_n6328), .Y(_abc_17692_n6331) );
  AND2X2 AND2X2_2476 ( .A(_abc_17692_n5944), .B(_abc_17692_n6139), .Y(_abc_17692_n6332) );
  AND2X2 AND2X2_2477 ( .A(_abc_17692_n5940), .B(_abc_17692_n6332), .Y(_abc_17692_n6333) );
  AND2X2 AND2X2_2478 ( .A(_abc_17692_n5942), .B(_abc_17692_n6137), .Y(_abc_17692_n6335) );
  AND2X2 AND2X2_2479 ( .A(sum_22_), .B(\key_in[54] ), .Y(_abc_17692_n6339) );
  AND2X2 AND2X2_248 ( .A(_abc_17692_n1256), .B(state_3_bF_buf1), .Y(_abc_17692_n1257) );
  AND2X2 AND2X2_2480 ( .A(_abc_17692_n6340), .B(_abc_17692_n6341), .Y(_abc_17692_n6342) );
  AND2X2 AND2X2_2481 ( .A(_abc_17692_n6338), .B(_abc_17692_n6342), .Y(_abc_17692_n6343) );
  AND2X2 AND2X2_2482 ( .A(_abc_17692_n6345), .B(_abc_17692_n6336), .Y(_abc_17692_n6346) );
  AND2X2 AND2X2_2483 ( .A(_abc_17692_n6346), .B(_abc_17692_n6347), .Y(_abc_17692_n6348) );
  AND2X2 AND2X2_2484 ( .A(_abc_17692_n6352), .B(_abc_17692_n6351), .Y(_abc_17692_n6353) );
  AND2X2 AND2X2_2485 ( .A(_abc_17692_n6354), .B(_abc_17692_n6293), .Y(_abc_17692_n6355) );
  AND2X2 AND2X2_2486 ( .A(_abc_17692_n6353), .B(workunit2_22_), .Y(_abc_17692_n6356) );
  AND2X2 AND2X2_2487 ( .A(_abc_17692_n6147), .B(workunit2_21_), .Y(_abc_17692_n6359) );
  AND2X2 AND2X2_2488 ( .A(_abc_17692_n6361), .B(_abc_17692_n6360), .Y(_abc_17692_n6362) );
  AND2X2 AND2X2_2489 ( .A(_abc_17692_n6364), .B(_abc_17692_n6362), .Y(_abc_17692_n6365) );
  AND2X2 AND2X2_249 ( .A(_abc_17692_n1257), .B(_abc_17692_n1254), .Y(_abc_17692_n1258_1) );
  AND2X2 AND2X2_2490 ( .A(_abc_17692_n6368), .B(_abc_17692_n1846_bF_buf0), .Y(_abc_17692_n6369) );
  AND2X2 AND2X2_2491 ( .A(_abc_17692_n6369), .B(_abc_17692_n6367), .Y(_abc_17692_n6370) );
  AND2X2 AND2X2_2492 ( .A(_abc_17692_n5807), .B(_abc_17692_n6169_1), .Y(_abc_17692_n6373) );
  AND2X2 AND2X2_2493 ( .A(_abc_17692_n5803), .B(_abc_17692_n6373), .Y(_abc_17692_n6374_1) );
  AND2X2 AND2X2_2494 ( .A(_abc_17692_n5805), .B(_abc_17692_n6167), .Y(_abc_17692_n6376) );
  AND2X2 AND2X2_2495 ( .A(sum_22_), .B(\key_in[118] ), .Y(_abc_17692_n6380) );
  AND2X2 AND2X2_2496 ( .A(_abc_17692_n6381), .B(_abc_17692_n6382), .Y(_abc_17692_n6383) );
  AND2X2 AND2X2_2497 ( .A(_abc_17692_n6379), .B(_abc_17692_n6383), .Y(_abc_17692_n6384) );
  AND2X2 AND2X2_2498 ( .A(_abc_17692_n6385), .B(_abc_17692_n6377), .Y(_abc_17692_n6386) );
  AND2X2 AND2X2_2499 ( .A(_abc_17692_n6386), .B(_abc_17692_n6387), .Y(_abc_17692_n6388) );
  AND2X2 AND2X2_25 ( .A(_abc_17692_n684), .B(_abc_17692_n685), .Y(x_4__FF_INPUT) );
  AND2X2 AND2X2_250 ( .A(_abc_17692_n1205), .B(sum_12_), .Y(_abc_17692_n1259) );
  AND2X2 AND2X2_2500 ( .A(_abc_17692_n6389), .B(_abc_17692_n6275), .Y(_abc_17692_n6390) );
  AND2X2 AND2X2_2501 ( .A(_abc_17692_n6391), .B(_abc_17692_n6256), .Y(_abc_17692_n6392) );
  AND2X2 AND2X2_2502 ( .A(_abc_17692_n6395), .B(_abc_17692_n6396), .Y(_abc_17692_n6397) );
  AND2X2 AND2X2_2503 ( .A(_abc_17692_n6181), .B(workunit2_21_), .Y(_abc_17692_n6399) );
  AND2X2 AND2X2_2504 ( .A(_abc_17692_n6189), .B(_abc_17692_n5822), .Y(_abc_17692_n6400) );
  AND2X2 AND2X2_2505 ( .A(_abc_17692_n6189), .B(_abc_17692_n5824), .Y(_abc_17692_n6402) );
  AND2X2 AND2X2_2506 ( .A(_abc_17692_n5837), .B(_abc_17692_n6402), .Y(_abc_17692_n6403) );
  AND2X2 AND2X2_2507 ( .A(_abc_17692_n6404), .B(_abc_17692_n6398), .Y(_abc_17692_n6405) );
  AND2X2 AND2X2_2508 ( .A(_abc_17692_n6407), .B(_abc_17692_n1863_bF_buf10), .Y(_abc_17692_n6408) );
  AND2X2 AND2X2_2509 ( .A(_abc_17692_n6408), .B(_abc_17692_n6406), .Y(_abc_17692_n6409) );
  AND2X2 AND2X2_251 ( .A(_abc_17692_n1251), .B(_abc_17692_n1208), .Y(_abc_17692_n1262) );
  AND2X2 AND2X2_2510 ( .A(_abc_17692_n6410), .B(state_6_bF_buf2), .Y(_abc_17692_n6411) );
  AND2X2 AND2X2_2511 ( .A(_abc_17692_n6180), .B(_abc_17692_n6196), .Y(_abc_17692_n6412) );
  AND2X2 AND2X2_2512 ( .A(_abc_17692_n5995), .B(_abc_17692_n6412), .Y(_abc_17692_n6413) );
  AND2X2 AND2X2_2513 ( .A(_abc_17692_n6417), .B(_abc_17692_n1863_bF_buf9), .Y(_abc_17692_n6418) );
  AND2X2 AND2X2_2514 ( .A(_abc_17692_n6418), .B(_abc_17692_n6415), .Y(_abc_17692_n6419) );
  AND2X2 AND2X2_2515 ( .A(_abc_17692_n6014), .B(_abc_17692_n6422), .Y(_abc_17692_n6423) );
  AND2X2 AND2X2_2516 ( .A(_abc_17692_n6424), .B(_abc_17692_n6205), .Y(_abc_17692_n6425) );
  AND2X2 AND2X2_2517 ( .A(_abc_17692_n6428), .B(_abc_17692_n6420), .Y(_abc_17692_n6429) );
  AND2X2 AND2X2_2518 ( .A(_abc_17692_n6431), .B(_abc_17692_n1877_bF_buf10), .Y(_abc_17692_n6432) );
  AND2X2 AND2X2_2519 ( .A(_abc_17692_n6432), .B(_abc_17692_n6430), .Y(_abc_17692_n6433) );
  AND2X2 AND2X2_252 ( .A(_abc_17692_n1234), .B(_abc_17692_n1262), .Y(_abc_17692_n1263) );
  AND2X2 AND2X2_2520 ( .A(_abc_17692_n6435), .B(_abc_17692_n6152), .Y(_abc_17692_n6436) );
  AND2X2 AND2X2_2521 ( .A(_abc_17692_n6153), .B(_abc_17692_n5960), .Y(_abc_17692_n6438) );
  AND2X2 AND2X2_2522 ( .A(_abc_17692_n6440), .B(_abc_17692_n6437), .Y(_abc_17692_n6441) );
  AND2X2 AND2X2_2523 ( .A(_abc_17692_n6444), .B(_abc_17692_n1846_bF_buf10), .Y(_abc_17692_n6445) );
  AND2X2 AND2X2_2524 ( .A(_abc_17692_n6445), .B(_abc_17692_n6442), .Y(_abc_17692_n6446) );
  AND2X2 AND2X2_2525 ( .A(_abc_17692_n6447), .B(_abc_17692_n6129), .Y(_abc_17692_n6448) );
  AND2X2 AND2X2_2526 ( .A(_abc_17692_n6130), .B(_abc_17692_n5913), .Y(_abc_17692_n6449) );
  AND2X2 AND2X2_2527 ( .A(_abc_17692_n6047), .B(_abc_17692_n6449), .Y(_abc_17692_n6450) );
  AND2X2 AND2X2_2528 ( .A(_abc_17692_n6451), .B(_abc_17692_n6319_1), .Y(_abc_17692_n6452) );
  AND2X2 AND2X2_2529 ( .A(_abc_17692_n6454), .B(_abc_17692_n1830_bF_buf10), .Y(_abc_17692_n6455) );
  AND2X2 AND2X2_253 ( .A(_abc_17692_n1251), .B(_abc_17692_n1259), .Y(_abc_17692_n1265) );
  AND2X2 AND2X2_2530 ( .A(_abc_17692_n6455), .B(_abc_17692_n6453), .Y(_abc_17692_n6456) );
  AND2X2 AND2X2_2531 ( .A(_abc_17692_n6459), .B(state_7_bF_buf1), .Y(_abc_17692_n6460) );
  AND2X2 AND2X2_2532 ( .A(_abc_17692_n1885_bF_buf2), .B(workunit2_22_), .Y(_abc_17692_n6461) );
  AND2X2 AND2X2_2533 ( .A(state_8_bF_buf7), .B(\data_in2[22] ), .Y(_abc_17692_n6462) );
  AND2X2 AND2X2_2534 ( .A(_abc_17692_n6467), .B(_abc_17692_n6469), .Y(_abc_17692_n6470) );
  AND2X2 AND2X2_2535 ( .A(_abc_17692_n6471), .B(workunit1_23_), .Y(_abc_17692_n6472) );
  AND2X2 AND2X2_2536 ( .A(_abc_17692_n6470), .B(_abc_17692_n5378), .Y(_abc_17692_n6474) );
  AND2X2 AND2X2_2537 ( .A(_abc_17692_n6473), .B(_abc_17692_n6475), .Y(_abc_17692_n6476) );
  AND2X2 AND2X2_2538 ( .A(_abc_17692_n6480), .B(_abc_17692_n6479), .Y(_abc_17692_n6481) );
  AND2X2 AND2X2_2539 ( .A(_abc_17692_n6482), .B(_abc_17692_n6478), .Y(_abc_17692_n6483) );
  AND2X2 AND2X2_254 ( .A(_abc_17692_n1266), .B(state_15_bF_buf1), .Y(_abc_17692_n1267) );
  AND2X2 AND2X2_2540 ( .A(_abc_17692_n6484), .B(_abc_17692_n6266), .Y(_abc_17692_n6485) );
  AND2X2 AND2X2_2541 ( .A(sum_23_), .B(\key_in[87] ), .Y(_abc_17692_n6486) );
  AND2X2 AND2X2_2542 ( .A(_abc_17692_n6487), .B(_abc_17692_n6488), .Y(_abc_17692_n6489) );
  AND2X2 AND2X2_2543 ( .A(_abc_17692_n6485), .B(_abc_17692_n6489), .Y(_abc_17692_n6490) );
  AND2X2 AND2X2_2544 ( .A(_abc_17692_n6491), .B(_abc_17692_n6492), .Y(_abc_17692_n6493) );
  AND2X2 AND2X2_2545 ( .A(_abc_17692_n6481), .B(_abc_17692_n6476), .Y(_abc_17692_n6495) );
  AND2X2 AND2X2_2546 ( .A(_abc_17692_n6466), .B(_abc_17692_n6477), .Y(_abc_17692_n6496) );
  AND2X2 AND2X2_2547 ( .A(_abc_17692_n6498), .B(_abc_17692_n6499), .Y(_abc_17692_n6500) );
  AND2X2 AND2X2_2548 ( .A(_abc_17692_n6502), .B(_abc_17692_n6494), .Y(_abc_17692_n6503) );
  AND2X2 AND2X2_2549 ( .A(_abc_17692_n6503), .B(workunit2_23_), .Y(_abc_17692_n6504) );
  AND2X2 AND2X2_255 ( .A(_abc_17692_n1264), .B(_abc_17692_n1267), .Y(_abc_17692_n1268) );
  AND2X2 AND2X2_2550 ( .A(_abc_17692_n6506), .B(_abc_17692_n6507), .Y(_abc_17692_n6508) );
  AND2X2 AND2X2_2551 ( .A(_abc_17692_n6508), .B(_abc_17692_n6505), .Y(_abc_17692_n6509) );
  AND2X2 AND2X2_2552 ( .A(_abc_17692_n6289), .B(_abc_17692_n6279), .Y(_abc_17692_n6511) );
  AND2X2 AND2X2_2553 ( .A(_abc_17692_n6515), .B(_abc_17692_n1877_bF_buf9), .Y(_abc_17692_n6516) );
  AND2X2 AND2X2_2554 ( .A(_abc_17692_n6516), .B(_abc_17692_n6513), .Y(_abc_17692_n6517) );
  AND2X2 AND2X2_2555 ( .A(_abc_17692_n6518), .B(_abc_17692_n6340), .Y(_abc_17692_n6519) );
  AND2X2 AND2X2_2556 ( .A(sum_23_), .B(\key_in[55] ), .Y(_abc_17692_n6520) );
  AND2X2 AND2X2_2557 ( .A(_abc_17692_n6521), .B(_abc_17692_n6522), .Y(_abc_17692_n6523_1) );
  AND2X2 AND2X2_2558 ( .A(_abc_17692_n6519), .B(_abc_17692_n6523_1), .Y(_abc_17692_n6524) );
  AND2X2 AND2X2_2559 ( .A(_abc_17692_n6525), .B(_abc_17692_n6526_1), .Y(_abc_17692_n6527) );
  AND2X2 AND2X2_256 ( .A(_abc_17692_n1268), .B(_abc_17692_n1261), .Y(_abc_17692_n1269) );
  AND2X2 AND2X2_2560 ( .A(_abc_17692_n6531), .B(_abc_17692_n6530), .Y(_abc_17692_n6532) );
  AND2X2 AND2X2_2561 ( .A(_abc_17692_n6529), .B(_abc_17692_n6533), .Y(_abc_17692_n6534) );
  AND2X2 AND2X2_2562 ( .A(_abc_17692_n6536), .B(_abc_17692_n6537), .Y(_abc_17692_n6538) );
  AND2X2 AND2X2_2563 ( .A(_abc_17692_n6535), .B(_abc_17692_n6539), .Y(_abc_17692_n6540) );
  AND2X2 AND2X2_2564 ( .A(_abc_17692_n6368), .B(_abc_17692_n6542), .Y(_abc_17692_n6543) );
  AND2X2 AND2X2_2565 ( .A(_abc_17692_n6546), .B(_abc_17692_n1846_bF_buf9), .Y(_abc_17692_n6547) );
  AND2X2 AND2X2_2566 ( .A(_abc_17692_n6547), .B(_abc_17692_n6545), .Y(_abc_17692_n6548) );
  AND2X2 AND2X2_2567 ( .A(_abc_17692_n6549), .B(_abc_17692_n6302), .Y(_abc_17692_n6550) );
  AND2X2 AND2X2_2568 ( .A(sum_23_), .B(\key_in[23] ), .Y(_abc_17692_n6551) );
  AND2X2 AND2X2_2569 ( .A(_abc_17692_n6552), .B(_abc_17692_n6553), .Y(_abc_17692_n6554) );
  AND2X2 AND2X2_257 ( .A(_abc_17692_n722_bF_buf1), .B(sum_13_), .Y(_abc_17692_n1270) );
  AND2X2 AND2X2_2570 ( .A(_abc_17692_n6550), .B(_abc_17692_n6554), .Y(_abc_17692_n6555) );
  AND2X2 AND2X2_2571 ( .A(_abc_17692_n6556), .B(_abc_17692_n6557), .Y(_abc_17692_n6558) );
  AND2X2 AND2X2_2572 ( .A(_abc_17692_n6562), .B(_abc_17692_n6561), .Y(_abc_17692_n6563) );
  AND2X2 AND2X2_2573 ( .A(_abc_17692_n6560), .B(_abc_17692_n6564), .Y(_abc_17692_n6565) );
  AND2X2 AND2X2_2574 ( .A(_abc_17692_n6567), .B(_abc_17692_n6568), .Y(_abc_17692_n6569) );
  AND2X2 AND2X2_2575 ( .A(_abc_17692_n6566), .B(_abc_17692_n6570), .Y(_abc_17692_n6571) );
  AND2X2 AND2X2_2576 ( .A(_abc_17692_n6316_1), .B(workunit2_22_), .Y(_abc_17692_n6573) );
  AND2X2 AND2X2_2577 ( .A(_abc_17692_n6328), .B(_abc_17692_n6574), .Y(_abc_17692_n6575) );
  AND2X2 AND2X2_2578 ( .A(_abc_17692_n6578), .B(_abc_17692_n1830_bF_buf9), .Y(_abc_17692_n6579) );
  AND2X2 AND2X2_2579 ( .A(_abc_17692_n6579), .B(_abc_17692_n6577), .Y(_abc_17692_n6580) );
  AND2X2 AND2X2_258 ( .A(_abc_17692_n1274), .B(delta_14_), .Y(_abc_17692_n1275) );
  AND2X2 AND2X2_2580 ( .A(sum_23_), .B(\key_in[119] ), .Y(_abc_17692_n6584) );
  AND2X2 AND2X2_2581 ( .A(_abc_17692_n6585), .B(_abc_17692_n6586), .Y(_abc_17692_n6587) );
  AND2X2 AND2X2_2582 ( .A(_abc_17692_n6583), .B(_abc_17692_n6588), .Y(_abc_17692_n6590) );
  AND2X2 AND2X2_2583 ( .A(_abc_17692_n6591), .B(_abc_17692_n6589), .Y(_abc_17692_n6592) );
  AND2X2 AND2X2_2584 ( .A(_abc_17692_n6594), .B(_abc_17692_n6381), .Y(_abc_17692_n6595) );
  AND2X2 AND2X2_2585 ( .A(_abc_17692_n6595), .B(_abc_17692_n6587), .Y(_abc_17692_n6596) );
  AND2X2 AND2X2_2586 ( .A(_abc_17692_n6593), .B(_abc_17692_n6598), .Y(_abc_17692_n6599) );
  AND2X2 AND2X2_2587 ( .A(_abc_17692_n6599), .B(workunit2_23_), .Y(_abc_17692_n6600_1) );
  AND2X2 AND2X2_2588 ( .A(_abc_17692_n6601), .B(_abc_17692_n6602), .Y(_abc_17692_n6603) );
  AND2X2 AND2X2_2589 ( .A(_abc_17692_n6603), .B(_abc_17692_n6505), .Y(_abc_17692_n6604) );
  AND2X2 AND2X2_259 ( .A(_abc_17692_n1252), .B(_abc_17692_n1245), .Y(_abc_17692_n1280) );
  AND2X2 AND2X2_2590 ( .A(_abc_17692_n6609), .B(_abc_17692_n6605), .Y(_abc_17692_n6610) );
  AND2X2 AND2X2_2591 ( .A(_abc_17692_n6611), .B(_abc_17692_n6612), .Y(_abc_17692_n6613) );
  AND2X2 AND2X2_2592 ( .A(_abc_17692_n6608), .B(_abc_17692_n6613), .Y(_abc_17692_n6614) );
  AND2X2 AND2X2_2593 ( .A(_abc_17692_n6615), .B(_abc_17692_n1863_bF_buf8), .Y(_abc_17692_n6616) );
  AND2X2 AND2X2_2594 ( .A(_abc_17692_n6617), .B(state_6_bF_buf1), .Y(_abc_17692_n6618) );
  AND2X2 AND2X2_2595 ( .A(_abc_17692_n6415), .B(_abc_17692_n6395), .Y(_abc_17692_n6619) );
  AND2X2 AND2X2_2596 ( .A(_abc_17692_n6622), .B(_abc_17692_n1863_bF_buf7), .Y(_abc_17692_n6623) );
  AND2X2 AND2X2_2597 ( .A(_abc_17692_n6623), .B(_abc_17692_n6621), .Y(_abc_17692_n6624) );
  AND2X2 AND2X2_2598 ( .A(_abc_17692_n6625), .B(workunit2_22_), .Y(_abc_17692_n6626) );
  AND2X2 AND2X2_2599 ( .A(_abc_17692_n6627), .B(_abc_17692_n6510), .Y(_abc_17692_n6628) );
  AND2X2 AND2X2_26 ( .A(_abc_17692_n683), .B(x_5_), .Y(_abc_17692_n688) );
  AND2X2 AND2X2_260 ( .A(_abc_17692_n1279), .B(_abc_17692_n1281), .Y(_abc_17692_n1282) );
  AND2X2 AND2X2_2600 ( .A(_abc_17692_n6629), .B(_abc_17692_n6514), .Y(_abc_17692_n6630) );
  AND2X2 AND2X2_2601 ( .A(_abc_17692_n6631), .B(_abc_17692_n1877_bF_buf8), .Y(_abc_17692_n6632) );
  AND2X2 AND2X2_2602 ( .A(_abc_17692_n6354), .B(workunit2_22_), .Y(_abc_17692_n6633) );
  AND2X2 AND2X2_2603 ( .A(_abc_17692_n6442), .B(_abc_17692_n6634), .Y(_abc_17692_n6635) );
  AND2X2 AND2X2_2604 ( .A(_abc_17692_n6638), .B(_abc_17692_n1846_bF_buf8), .Y(_abc_17692_n6639) );
  AND2X2 AND2X2_2605 ( .A(_abc_17692_n6639), .B(_abc_17692_n6637), .Y(_abc_17692_n6640) );
  AND2X2 AND2X2_2606 ( .A(_abc_17692_n6645), .B(_abc_17692_n1830_bF_buf8), .Y(_abc_17692_n6646) );
  AND2X2 AND2X2_2607 ( .A(_abc_17692_n6646), .B(_abc_17692_n6644_1), .Y(_abc_17692_n6647_1) );
  AND2X2 AND2X2_2608 ( .A(_abc_17692_n6650), .B(state_7_bF_buf0), .Y(_abc_17692_n6651) );
  AND2X2 AND2X2_2609 ( .A(_abc_17692_n1885_bF_buf1), .B(workunit2_23_), .Y(_abc_17692_n6652_1) );
  AND2X2 AND2X2_261 ( .A(_abc_17692_n1283), .B(_abc_17692_n1278), .Y(_abc_17692_n1285) );
  AND2X2 AND2X2_2610 ( .A(state_8_bF_buf6), .B(\data_in2[23] ), .Y(_abc_17692_n6653) );
  AND2X2 AND2X2_2611 ( .A(_abc_17692_n6658_1), .B(_abc_17692_n6660_1), .Y(_abc_17692_n6661) );
  AND2X2 AND2X2_2612 ( .A(_abc_17692_n6662), .B(workunit1_24_), .Y(_abc_17692_n6663) );
  AND2X2 AND2X2_2613 ( .A(_abc_17692_n6661), .B(_abc_17692_n5598), .Y(_abc_17692_n6664) );
  AND2X2 AND2X2_2614 ( .A(_abc_17692_n6479), .B(_abc_17692_n6473), .Y(_abc_17692_n6667) );
  AND2X2 AND2X2_2615 ( .A(_abc_17692_n6249), .B(_abc_17692_n6476), .Y(_abc_17692_n6670) );
  AND2X2 AND2X2_2616 ( .A(_abc_17692_n6668), .B(_abc_17692_n6253), .Y(_abc_17692_n6672) );
  AND2X2 AND2X2_2617 ( .A(_abc_17692_n6674), .B(_abc_17692_n6671), .Y(_abc_17692_n6675) );
  AND2X2 AND2X2_2618 ( .A(_abc_17692_n6675), .B(_abc_17692_n6666), .Y(_abc_17692_n6676) );
  AND2X2 AND2X2_2619 ( .A(_abc_17692_n6252), .B(_abc_17692_n6672), .Y(_abc_17692_n6678) );
  AND2X2 AND2X2_262 ( .A(_abc_17692_n1286), .B(state_3_bF_buf0), .Y(_abc_17692_n1287) );
  AND2X2 AND2X2_2620 ( .A(_abc_17692_n6679), .B(_abc_17692_n6665), .Y(_abc_17692_n6680) );
  AND2X2 AND2X2_2621 ( .A(sum_24_), .B(\key_in[120] ), .Y(_abc_17692_n6682) );
  AND2X2 AND2X2_2622 ( .A(_abc_17692_n6683), .B(_abc_17692_n6684), .Y(_abc_17692_n6685) );
  AND2X2 AND2X2_2623 ( .A(_abc_17692_n6586), .B(_abc_17692_n6380), .Y(_abc_17692_n6686) );
  AND2X2 AND2X2_2624 ( .A(_abc_17692_n6688), .B(_abc_17692_n6377), .Y(_abc_17692_n6689) );
  AND2X2 AND2X2_2625 ( .A(_abc_17692_n6383), .B(_abc_17692_n6587), .Y(_abc_17692_n6692) );
  AND2X2 AND2X2_2626 ( .A(_abc_17692_n6691), .B(_abc_17692_n6693), .Y(_abc_17692_n6694) );
  AND2X2 AND2X2_2627 ( .A(_abc_17692_n6694), .B(_abc_17692_n6685), .Y(_abc_17692_n6695) );
  AND2X2 AND2X2_2628 ( .A(_abc_17692_n6697), .B(_abc_17692_n6696), .Y(_abc_17692_n6698) );
  AND2X2 AND2X2_2629 ( .A(_abc_17692_n6701), .B(_abc_17692_n6703), .Y(_abc_17692_n6704) );
  AND2X2 AND2X2_263 ( .A(_abc_17692_n1287), .B(_abc_17692_n1284), .Y(_abc_17692_n1288) );
  AND2X2 AND2X2_2630 ( .A(_abc_17692_n6705), .B(_abc_17692_n6657_1), .Y(_abc_17692_n6706) );
  AND2X2 AND2X2_2631 ( .A(_abc_17692_n6704), .B(workunit2_24_), .Y(_abc_17692_n6707) );
  AND2X2 AND2X2_2632 ( .A(_abc_17692_n6605), .B(_abc_17692_n6398), .Y(_abc_17692_n6710) );
  AND2X2 AND2X2_2633 ( .A(_abc_17692_n6401), .B(_abc_17692_n6710), .Y(_abc_17692_n6711) );
  AND2X2 AND2X2_2634 ( .A(_abc_17692_n6603), .B(workunit2_23_), .Y(_abc_17692_n6712) );
  AND2X2 AND2X2_2635 ( .A(_abc_17692_n6605), .B(_abc_17692_n6607), .Y(_abc_17692_n6713) );
  AND2X2 AND2X2_2636 ( .A(_abc_17692_n6710), .B(_abc_17692_n6402), .Y(_abc_17692_n6717) );
  AND2X2 AND2X2_2637 ( .A(_abc_17692_n6719), .B(_abc_17692_n6716), .Y(_abc_17692_n6720) );
  AND2X2 AND2X2_2638 ( .A(_abc_17692_n6721), .B(_abc_17692_n6709), .Y(_abc_17692_n6722) );
  AND2X2 AND2X2_2639 ( .A(_abc_17692_n6723), .B(_abc_17692_n6724), .Y(_abc_17692_n6725) );
  AND2X2 AND2X2_264 ( .A(_abc_17692_n723), .B(sum_14_), .Y(_abc_17692_n1289) );
  AND2X2 AND2X2_2640 ( .A(sum_24_), .B(\key_in[24] ), .Y(_abc_17692_n6727) );
  AND2X2 AND2X2_2641 ( .A(_abc_17692_n6728), .B(_abc_17692_n6729), .Y(_abc_17692_n6730) );
  AND2X2 AND2X2_2642 ( .A(_abc_17692_n6553), .B(_abc_17692_n6301), .Y(_abc_17692_n6731) );
  AND2X2 AND2X2_2643 ( .A(_abc_17692_n6733), .B(_abc_17692_n6298), .Y(_abc_17692_n6734) );
  AND2X2 AND2X2_2644 ( .A(_abc_17692_n6304), .B(_abc_17692_n6554), .Y(_abc_17692_n6737) );
  AND2X2 AND2X2_2645 ( .A(_abc_17692_n6736), .B(_abc_17692_n6738), .Y(_abc_17692_n6739) );
  AND2X2 AND2X2_2646 ( .A(_abc_17692_n6739), .B(_abc_17692_n6730), .Y(_abc_17692_n6740) );
  AND2X2 AND2X2_2647 ( .A(_abc_17692_n6307), .B(_abc_17692_n6734), .Y(_abc_17692_n6742) );
  AND2X2 AND2X2_2648 ( .A(_abc_17692_n6744), .B(_abc_17692_n6741), .Y(_abc_17692_n6745) );
  AND2X2 AND2X2_2649 ( .A(_abc_17692_n6749), .B(_abc_17692_n6748), .Y(_abc_17692_n6750) );
  AND2X2 AND2X2_265 ( .A(_abc_17692_n1246), .B(sum_13_), .Y(_abc_17692_n1291) );
  AND2X2 AND2X2_2650 ( .A(_abc_17692_n6751), .B(_abc_17692_n6657_1), .Y(_abc_17692_n6752) );
  AND2X2 AND2X2_2651 ( .A(_abc_17692_n6750), .B(workunit2_24_), .Y(_abc_17692_n6753) );
  AND2X2 AND2X2_2652 ( .A(_abc_17692_n6572), .B(_abc_17692_n6320), .Y(_abc_17692_n6756) );
  AND2X2 AND2X2_2653 ( .A(_abc_17692_n6756), .B(_abc_17692_n6324), .Y(_abc_17692_n6757) );
  AND2X2 AND2X2_2654 ( .A(_abc_17692_n6323), .B(_abc_17692_n6756), .Y(_abc_17692_n6761) );
  AND2X2 AND2X2_2655 ( .A(_abc_17692_n6565), .B(workunit2_23_), .Y(_abc_17692_n6762) );
  AND2X2 AND2X2_2656 ( .A(_abc_17692_n6572), .B(_abc_17692_n6573), .Y(_abc_17692_n6763) );
  AND2X2 AND2X2_2657 ( .A(_abc_17692_n6766), .B(_abc_17692_n6760), .Y(_abc_17692_n6767) );
  AND2X2 AND2X2_2658 ( .A(_abc_17692_n6759), .B(_abc_17692_n6767), .Y(_abc_17692_n6768) );
  AND2X2 AND2X2_2659 ( .A(_abc_17692_n6769), .B(_abc_17692_n6755), .Y(_abc_17692_n6771) );
  AND2X2 AND2X2_266 ( .A(_abc_17692_n1264), .B(_abc_17692_n1293), .Y(_abc_17692_n1294) );
  AND2X2 AND2X2_2660 ( .A(_abc_17692_n6772), .B(_abc_17692_n1830_bF_buf7), .Y(_abc_17692_n6773) );
  AND2X2 AND2X2_2661 ( .A(_abc_17692_n6773), .B(_abc_17692_n6770), .Y(_abc_17692_n6774) );
  AND2X2 AND2X2_2662 ( .A(sum_24_), .B(\key_in[88] ), .Y(_abc_17692_n6775) );
  AND2X2 AND2X2_2663 ( .A(_abc_17692_n6776), .B(_abc_17692_n6777), .Y(_abc_17692_n6778) );
  AND2X2 AND2X2_2664 ( .A(_abc_17692_n6488), .B(_abc_17692_n6265), .Y(_abc_17692_n6779) );
  AND2X2 AND2X2_2665 ( .A(_abc_17692_n6781), .B(_abc_17692_n6262), .Y(_abc_17692_n6782) );
  AND2X2 AND2X2_2666 ( .A(_abc_17692_n6259), .B(_abc_17692_n6782), .Y(_abc_17692_n6783) );
  AND2X2 AND2X2_2667 ( .A(_abc_17692_n6268), .B(_abc_17692_n6489), .Y(_abc_17692_n6784) );
  AND2X2 AND2X2_2668 ( .A(_abc_17692_n6788), .B(_abc_17692_n6778), .Y(_abc_17692_n6789) );
  AND2X2 AND2X2_2669 ( .A(_abc_17692_n6787), .B(_abc_17692_n6790), .Y(_abc_17692_n6791) );
  AND2X2 AND2X2_267 ( .A(_abc_17692_n1295), .B(_abc_17692_n1290), .Y(_abc_17692_n1296) );
  AND2X2 AND2X2_2670 ( .A(_abc_17692_n6794), .B(_abc_17692_n6795), .Y(_abc_17692_n6796) );
  AND2X2 AND2X2_2671 ( .A(_abc_17692_n6797), .B(workunit2_24_), .Y(_abc_17692_n6798) );
  AND2X2 AND2X2_2672 ( .A(_abc_17692_n6796), .B(_abc_17692_n6657_1), .Y(_abc_17692_n6799) );
  AND2X2 AND2X2_2673 ( .A(_abc_17692_n6510), .B(_abc_17692_n6281), .Y(_abc_17692_n6801) );
  AND2X2 AND2X2_2674 ( .A(_abc_17692_n6801), .B(_abc_17692_n6285), .Y(_abc_17692_n6802) );
  AND2X2 AND2X2_2675 ( .A(_abc_17692_n5877), .B(_abc_17692_n6802), .Y(_abc_17692_n6803) );
  AND2X2 AND2X2_2676 ( .A(_abc_17692_n6801), .B(_abc_17692_n6284), .Y(_abc_17692_n6806) );
  AND2X2 AND2X2_2677 ( .A(_abc_17692_n6508), .B(workunit2_23_), .Y(_abc_17692_n6808) );
  AND2X2 AND2X2_2678 ( .A(_abc_17692_n6510), .B(_abc_17692_n6278), .Y(_abc_17692_n6809) );
  AND2X2 AND2X2_2679 ( .A(_abc_17692_n6811), .B(_abc_17692_n6807), .Y(_abc_17692_n6812) );
  AND2X2 AND2X2_268 ( .A(_abc_17692_n1298), .B(state_15_bF_buf0), .Y(_abc_17692_n1299) );
  AND2X2 AND2X2_2680 ( .A(_abc_17692_n6805), .B(_abc_17692_n6812), .Y(_abc_17692_n6813) );
  AND2X2 AND2X2_2681 ( .A(_abc_17692_n6815), .B(_abc_17692_n6800), .Y(_abc_17692_n6816) );
  AND2X2 AND2X2_2682 ( .A(_abc_17692_n6818), .B(_abc_17692_n1877_bF_buf7), .Y(_abc_17692_n6819) );
  AND2X2 AND2X2_2683 ( .A(_abc_17692_n6819), .B(_abc_17692_n6817), .Y(_abc_17692_n6820) );
  AND2X2 AND2X2_2684 ( .A(sum_24_), .B(\key_in[56] ), .Y(_abc_17692_n6821) );
  AND2X2 AND2X2_2685 ( .A(_abc_17692_n6822), .B(_abc_17692_n6823), .Y(_abc_17692_n6824) );
  AND2X2 AND2X2_2686 ( .A(_abc_17692_n6522), .B(_abc_17692_n6339), .Y(_abc_17692_n6825) );
  AND2X2 AND2X2_2687 ( .A(_abc_17692_n6827), .B(_abc_17692_n6336), .Y(_abc_17692_n6828) );
  AND2X2 AND2X2_2688 ( .A(_abc_17692_n6342), .B(_abc_17692_n6523_1), .Y(_abc_17692_n6831) );
  AND2X2 AND2X2_2689 ( .A(_abc_17692_n6830), .B(_abc_17692_n6832), .Y(_abc_17692_n6833) );
  AND2X2 AND2X2_269 ( .A(_abc_17692_n1299), .B(_abc_17692_n1297), .Y(_abc_17692_n1300) );
  AND2X2 AND2X2_2690 ( .A(_abc_17692_n6833), .B(_abc_17692_n6824), .Y(_abc_17692_n6834) );
  AND2X2 AND2X2_2691 ( .A(_abc_17692_n6345), .B(_abc_17692_n6828), .Y(_abc_17692_n6836) );
  AND2X2 AND2X2_2692 ( .A(_abc_17692_n6838), .B(_abc_17692_n6835), .Y(_abc_17692_n6839) );
  AND2X2 AND2X2_2693 ( .A(_abc_17692_n6843), .B(_abc_17692_n6842), .Y(_abc_17692_n6844) );
  AND2X2 AND2X2_2694 ( .A(_abc_17692_n6845), .B(_abc_17692_n6657_1), .Y(_abc_17692_n6846) );
  AND2X2 AND2X2_2695 ( .A(_abc_17692_n6844), .B(workunit2_24_), .Y(_abc_17692_n6847) );
  AND2X2 AND2X2_2696 ( .A(_abc_17692_n6534), .B(workunit2_23_), .Y(_abc_17692_n6855) );
  AND2X2 AND2X2_2697 ( .A(_abc_17692_n6857), .B(_abc_17692_n6856), .Y(_abc_17692_n6858) );
  AND2X2 AND2X2_2698 ( .A(_abc_17692_n6854), .B(_abc_17692_n6858), .Y(_abc_17692_n6859) );
  AND2X2 AND2X2_2699 ( .A(_abc_17692_n6853), .B(_abc_17692_n6859), .Y(_abc_17692_n6860) );
  AND2X2 AND2X2_27 ( .A(_abc_17692_n689), .B(_abc_17692_n687), .Y(x_5__FF_INPUT) );
  AND2X2 AND2X2_270 ( .A(_abc_17692_n1303), .B(delta_15_), .Y(_abc_17692_n1304) );
  AND2X2 AND2X2_2700 ( .A(_abc_17692_n6852), .B(_abc_17692_n6860), .Y(_abc_17692_n6861) );
  AND2X2 AND2X2_2701 ( .A(_abc_17692_n6862), .B(_abc_17692_n6849), .Y(_abc_17692_n6863) );
  AND2X2 AND2X2_2702 ( .A(_abc_17692_n6865), .B(_abc_17692_n1846_bF_buf7), .Y(_abc_17692_n6866) );
  AND2X2 AND2X2_2703 ( .A(_abc_17692_n6866), .B(_abc_17692_n6864), .Y(_abc_17692_n6867) );
  AND2X2 AND2X2_2704 ( .A(_abc_17692_n6870), .B(state_6_bF_buf0), .Y(_abc_17692_n6871) );
  AND2X2 AND2X2_2705 ( .A(_abc_17692_n6726), .B(_abc_17692_n6871), .Y(_abc_17692_n6872) );
  AND2X2 AND2X2_2706 ( .A(_abc_17692_n6184), .B(_abc_17692_n5823), .Y(_abc_17692_n6873) );
  AND2X2 AND2X2_2707 ( .A(_abc_17692_n6613), .B(_abc_17692_n6397), .Y(_abc_17692_n6874) );
  AND2X2 AND2X2_2708 ( .A(_abc_17692_n6874), .B(_abc_17692_n6873), .Y(_abc_17692_n6875) );
  AND2X2 AND2X2_2709 ( .A(_abc_17692_n6875), .B(_abc_17692_n5989), .Y(_abc_17692_n6876) );
  AND2X2 AND2X2_271 ( .A(_abc_17692_n1305), .B(_abc_17692_n1306), .Y(_abc_17692_n1307) );
  AND2X2 AND2X2_2710 ( .A(_abc_17692_n6877), .B(_abc_17692_n6183), .Y(_abc_17692_n6878) );
  AND2X2 AND2X2_2711 ( .A(_abc_17692_n6874), .B(_abc_17692_n6878), .Y(_abc_17692_n6879) );
  AND2X2 AND2X2_2712 ( .A(_abc_17692_n6611), .B(_abc_17692_n6395), .Y(_abc_17692_n6880) );
  AND2X2 AND2X2_2713 ( .A(_abc_17692_n5991), .B(_abc_17692_n6875), .Y(_abc_17692_n6885) );
  AND2X2 AND2X2_2714 ( .A(_abc_17692_n6886), .B(_abc_17692_n6708), .Y(_abc_17692_n6888) );
  AND2X2 AND2X2_2715 ( .A(_abc_17692_n6889), .B(_abc_17692_n1863_bF_buf5), .Y(_abc_17692_n6890) );
  AND2X2 AND2X2_2716 ( .A(_abc_17692_n6890), .B(_abc_17692_n6887), .Y(_abc_17692_n6891) );
  AND2X2 AND2X2_2717 ( .A(_abc_17692_n6898), .B(_abc_17692_n6897), .Y(_abc_17692_n6899) );
  AND2X2 AND2X2_2718 ( .A(_abc_17692_n6896), .B(_abc_17692_n6900), .Y(_abc_17692_n6901) );
  AND2X2 AND2X2_2719 ( .A(_abc_17692_n6895), .B(_abc_17692_n6901), .Y(_abc_17692_n6902) );
  AND2X2 AND2X2_272 ( .A(delta_14_), .B(sum_14_), .Y(_abc_17692_n1308_1) );
  AND2X2 AND2X2_2720 ( .A(_abc_17692_n6894), .B(_abc_17692_n6902), .Y(_abc_17692_n6903) );
  AND2X2 AND2X2_2721 ( .A(_abc_17692_n6907), .B(_abc_17692_n1877_bF_buf6), .Y(_abc_17692_n6908) );
  AND2X2 AND2X2_2722 ( .A(_abc_17692_n6908), .B(_abc_17692_n6904), .Y(_abc_17692_n6909) );
  AND2X2 AND2X2_2723 ( .A(_abc_17692_n6540), .B(_abc_17692_n6357), .Y(_abc_17692_n6910) );
  AND2X2 AND2X2_2724 ( .A(_abc_17692_n6910), .B(_abc_17692_n6438), .Y(_abc_17692_n6911) );
  AND2X2 AND2X2_2725 ( .A(_abc_17692_n6026), .B(_abc_17692_n6911), .Y(_abc_17692_n6912) );
  AND2X2 AND2X2_2726 ( .A(_abc_17692_n6910), .B(_abc_17692_n6436), .Y(_abc_17692_n6913) );
  AND2X2 AND2X2_2727 ( .A(_abc_17692_n6915), .B(_abc_17692_n6539), .Y(_abc_17692_n6916) );
  AND2X2 AND2X2_2728 ( .A(_abc_17692_n6029), .B(_abc_17692_n6911), .Y(_abc_17692_n6919) );
  AND2X2 AND2X2_2729 ( .A(_abc_17692_n6920), .B(_abc_17692_n6848), .Y(_abc_17692_n6922) );
  AND2X2 AND2X2_273 ( .A(_abc_17692_n1286), .B(_abc_17692_n1309), .Y(_abc_17692_n1310) );
  AND2X2 AND2X2_2730 ( .A(_abc_17692_n6923), .B(_abc_17692_n1846_bF_buf6), .Y(_abc_17692_n6924) );
  AND2X2 AND2X2_2731 ( .A(_abc_17692_n6924), .B(_abc_17692_n6921), .Y(_abc_17692_n6925) );
  AND2X2 AND2X2_2732 ( .A(_abc_17692_n6571), .B(_abc_17692_n6319_1), .Y(_abc_17692_n6926) );
  AND2X2 AND2X2_2733 ( .A(_abc_17692_n6449), .B(_abc_17692_n6926), .Y(_abc_17692_n6927) );
  AND2X2 AND2X2_2734 ( .A(_abc_17692_n6927), .B(_abc_17692_n6044), .Y(_abc_17692_n6928) );
  AND2X2 AND2X2_2735 ( .A(_abc_17692_n6926), .B(_abc_17692_n6448), .Y(_abc_17692_n6929) );
  AND2X2 AND2X2_2736 ( .A(_abc_17692_n6570), .B(_abc_17692_n6641), .Y(_abc_17692_n6931) );
  AND2X2 AND2X2_2737 ( .A(_abc_17692_n6927), .B(_abc_17692_n6045), .Y(_abc_17692_n6935) );
  AND2X2 AND2X2_2738 ( .A(_abc_17692_n5187), .B(_abc_17692_n6935), .Y(_abc_17692_n6936) );
  AND2X2 AND2X2_2739 ( .A(_abc_17692_n6937), .B(_abc_17692_n6754), .Y(_abc_17692_n6938) );
  AND2X2 AND2X2_274 ( .A(_abc_17692_n1314), .B(state_3_bF_buf4), .Y(_abc_17692_n1315) );
  AND2X2 AND2X2_2740 ( .A(_abc_17692_n6940), .B(_abc_17692_n1830_bF_buf6), .Y(_abc_17692_n6941) );
  AND2X2 AND2X2_2741 ( .A(_abc_17692_n6941), .B(_abc_17692_n6939), .Y(_abc_17692_n6942) );
  AND2X2 AND2X2_2742 ( .A(_abc_17692_n6945), .B(state_7_bF_buf4), .Y(_abc_17692_n6946) );
  AND2X2 AND2X2_2743 ( .A(_abc_17692_n1885_bF_buf0), .B(workunit2_24_), .Y(_abc_17692_n6947) );
  AND2X2 AND2X2_2744 ( .A(state_8_bF_buf5), .B(\data_in2[24] ), .Y(_abc_17692_n6948) );
  AND2X2 AND2X2_2745 ( .A(_abc_17692_n6955), .B(_abc_17692_n6957), .Y(_abc_17692_n6958) );
  AND2X2 AND2X2_2746 ( .A(_abc_17692_n6959), .B(workunit1_25_), .Y(_abc_17692_n6960) );
  AND2X2 AND2X2_2747 ( .A(_abc_17692_n6958), .B(_abc_17692_n5782), .Y(_abc_17692_n6962) );
  AND2X2 AND2X2_2748 ( .A(_abc_17692_n6961), .B(_abc_17692_n6963), .Y(_abc_17692_n6964) );
  AND2X2 AND2X2_2749 ( .A(_abc_17692_n6954), .B(_abc_17692_n6964), .Y(_abc_17692_n6965) );
  AND2X2 AND2X2_275 ( .A(_abc_17692_n1315), .B(_abc_17692_n1311_1), .Y(_abc_17692_n1316) );
  AND2X2 AND2X2_2750 ( .A(_abc_17692_n6966), .B(_abc_17692_n6967), .Y(_abc_17692_n6968) );
  AND2X2 AND2X2_2751 ( .A(sum_25_), .B(\key_in[121] ), .Y(_abc_17692_n6971) );
  AND2X2 AND2X2_2752 ( .A(_abc_17692_n6972), .B(_abc_17692_n6973), .Y(_abc_17692_n6974) );
  AND2X2 AND2X2_2753 ( .A(_abc_17692_n6970), .B(_abc_17692_n6974), .Y(_abc_17692_n6975) );
  AND2X2 AND2X2_2754 ( .A(_abc_17692_n6982), .B(_abc_17692_n6976), .Y(_abc_17692_n6983) );
  AND2X2 AND2X2_2755 ( .A(_abc_17692_n6979), .B(_abc_17692_n6984), .Y(_abc_17692_n6985) );
  AND2X2 AND2X2_2756 ( .A(_abc_17692_n6985), .B(_abc_17692_n6952), .Y(_abc_17692_n6987) );
  AND2X2 AND2X2_2757 ( .A(_abc_17692_n6988), .B(_abc_17692_n6986), .Y(_abc_17692_n6989) );
  AND2X2 AND2X2_2758 ( .A(_abc_17692_n6723), .B(_abc_17692_n6990), .Y(_abc_17692_n6991) );
  AND2X2 AND2X2_2759 ( .A(_abc_17692_n6992), .B(_abc_17692_n6989), .Y(_abc_17692_n6993) );
  AND2X2 AND2X2_276 ( .A(_abc_17692_n723), .B(sum_15_), .Y(_abc_17692_n1317) );
  AND2X2 AND2X2_2760 ( .A(_abc_17692_n6991), .B(_abc_17692_n6994), .Y(_abc_17692_n6995) );
  AND2X2 AND2X2_2761 ( .A(sum_25_), .B(\key_in[89] ), .Y(_abc_17692_n6999) );
  AND2X2 AND2X2_2762 ( .A(_abc_17692_n7000), .B(_abc_17692_n7001), .Y(_abc_17692_n7002) );
  AND2X2 AND2X2_2763 ( .A(_abc_17692_n6998), .B(_abc_17692_n7003), .Y(_abc_17692_n7005) );
  AND2X2 AND2X2_2764 ( .A(_abc_17692_n7006), .B(_abc_17692_n7004), .Y(_abc_17692_n7007) );
  AND2X2 AND2X2_2765 ( .A(_abc_17692_n7011), .B(_abc_17692_n7008), .Y(_abc_17692_n7012) );
  AND2X2 AND2X2_2766 ( .A(_abc_17692_n7012), .B(workunit2_25_), .Y(_abc_17692_n7013) );
  AND2X2 AND2X2_2767 ( .A(_abc_17692_n7014), .B(_abc_17692_n6952), .Y(_abc_17692_n7015) );
  AND2X2 AND2X2_2768 ( .A(_abc_17692_n6796), .B(workunit2_24_), .Y(_abc_17692_n7018) );
  AND2X2 AND2X2_2769 ( .A(_abc_17692_n6817), .B(_abc_17692_n7019), .Y(_abc_17692_n7020) );
  AND2X2 AND2X2_277 ( .A(_abc_17692_n1297), .B(_abc_17692_n1276), .Y(_abc_17692_n1318) );
  AND2X2 AND2X2_2770 ( .A(_abc_17692_n7023), .B(_abc_17692_n1877_bF_buf5), .Y(_abc_17692_n7024) );
  AND2X2 AND2X2_2771 ( .A(_abc_17692_n7024), .B(_abc_17692_n7021), .Y(_abc_17692_n7025) );
  AND2X2 AND2X2_2772 ( .A(sum_25_), .B(\key_in[25] ), .Y(_abc_17692_n7028) );
  AND2X2 AND2X2_2773 ( .A(_abc_17692_n7029), .B(_abc_17692_n7030), .Y(_abc_17692_n7031) );
  AND2X2 AND2X2_2774 ( .A(_abc_17692_n7027), .B(_abc_17692_n7031), .Y(_abc_17692_n7032) );
  AND2X2 AND2X2_2775 ( .A(_abc_17692_n7033), .B(_abc_17692_n7034), .Y(_abc_17692_n7035) );
  AND2X2 AND2X2_2776 ( .A(_abc_17692_n7039), .B(_abc_17692_n7036), .Y(_abc_17692_n7040) );
  AND2X2 AND2X2_2777 ( .A(_abc_17692_n7040), .B(workunit2_25_), .Y(_abc_17692_n7041) );
  AND2X2 AND2X2_2778 ( .A(_abc_17692_n7043), .B(_abc_17692_n6952), .Y(_abc_17692_n7044) );
  AND2X2 AND2X2_2779 ( .A(_abc_17692_n7045), .B(_abc_17692_n7042), .Y(_abc_17692_n7046) );
  AND2X2 AND2X2_278 ( .A(_abc_17692_n1321), .B(state_15_bF_buf4), .Y(_abc_17692_n1322) );
  AND2X2 AND2X2_2780 ( .A(_abc_17692_n6772), .B(_abc_17692_n7048), .Y(_abc_17692_n7049) );
  AND2X2 AND2X2_2781 ( .A(_abc_17692_n7052), .B(_abc_17692_n1830_bF_buf5), .Y(_abc_17692_n7053) );
  AND2X2 AND2X2_2782 ( .A(_abc_17692_n7053), .B(_abc_17692_n7051), .Y(_abc_17692_n7054) );
  AND2X2 AND2X2_2783 ( .A(sum_25_), .B(\key_in[57] ), .Y(_abc_17692_n7057) );
  AND2X2 AND2X2_2784 ( .A(_abc_17692_n7058), .B(_abc_17692_n7059), .Y(_abc_17692_n7060) );
  AND2X2 AND2X2_2785 ( .A(_abc_17692_n7056), .B(_abc_17692_n7060), .Y(_abc_17692_n7061) );
  AND2X2 AND2X2_2786 ( .A(_abc_17692_n7062), .B(_abc_17692_n7063), .Y(_abc_17692_n7064) );
  AND2X2 AND2X2_2787 ( .A(_abc_17692_n6981), .B(_abc_17692_n7065), .Y(_abc_17692_n7066) );
  AND2X2 AND2X2_2788 ( .A(_abc_17692_n6968), .B(_abc_17692_n7064), .Y(_abc_17692_n7067) );
  AND2X2 AND2X2_2789 ( .A(_abc_17692_n7071), .B(_abc_17692_n7070), .Y(_abc_17692_n7072) );
  AND2X2 AND2X2_279 ( .A(_abc_17692_n1322), .B(_abc_17692_n1320_1), .Y(_abc_17692_n1323) );
  AND2X2 AND2X2_2790 ( .A(_abc_17692_n7073), .B(_abc_17692_n7069), .Y(_abc_17692_n7074) );
  AND2X2 AND2X2_2791 ( .A(_abc_17692_n6864), .B(_abc_17692_n7076), .Y(_abc_17692_n7077) );
  AND2X2 AND2X2_2792 ( .A(_abc_17692_n7080), .B(_abc_17692_n1846_bF_buf5), .Y(_abc_17692_n7081) );
  AND2X2 AND2X2_2793 ( .A(_abc_17692_n7081), .B(_abc_17692_n7079), .Y(_abc_17692_n7082) );
  AND2X2 AND2X2_2794 ( .A(_abc_17692_n7085), .B(state_6_bF_buf4), .Y(_abc_17692_n7086) );
  AND2X2 AND2X2_2795 ( .A(_abc_17692_n7086), .B(_abc_17692_n6997), .Y(_abc_17692_n7087) );
  AND2X2 AND2X2_2796 ( .A(_abc_17692_n6705), .B(workunit2_24_), .Y(_abc_17692_n7088) );
  AND2X2 AND2X2_2797 ( .A(_abc_17692_n6889), .B(_abc_17692_n7089), .Y(_abc_17692_n7090) );
  AND2X2 AND2X2_2798 ( .A(_abc_17692_n7093), .B(_abc_17692_n1863_bF_buf3), .Y(_abc_17692_n7094) );
  AND2X2 AND2X2_2799 ( .A(_abc_17692_n7094), .B(_abc_17692_n7092), .Y(_abc_17692_n7095) );
  AND2X2 AND2X2_28 ( .A(_abc_17692_n688), .B(x_6_), .Y(_abc_17692_n692_1) );
  AND2X2 AND2X2_280 ( .A(delta_16_), .B(sum_16_), .Y(_abc_17692_n1326) );
  AND2X2 AND2X2_2800 ( .A(_abc_17692_n6904), .B(_abc_17692_n7096), .Y(_abc_17692_n7097) );
  AND2X2 AND2X2_2801 ( .A(_abc_17692_n7098), .B(_abc_17692_n7016), .Y(_abc_17692_n7099) );
  AND2X2 AND2X2_2802 ( .A(_abc_17692_n7097), .B(_abc_17692_n7017), .Y(_abc_17692_n7100) );
  AND2X2 AND2X2_2803 ( .A(_abc_17692_n7101), .B(_abc_17692_n1877_bF_buf4), .Y(_abc_17692_n7102) );
  AND2X2 AND2X2_2804 ( .A(_abc_17692_n6845), .B(workunit2_24_), .Y(_abc_17692_n7103) );
  AND2X2 AND2X2_2805 ( .A(_abc_17692_n6923), .B(_abc_17692_n7104), .Y(_abc_17692_n7105) );
  AND2X2 AND2X2_2806 ( .A(_abc_17692_n7108), .B(_abc_17692_n1846_bF_buf4), .Y(_abc_17692_n7109) );
  AND2X2 AND2X2_2807 ( .A(_abc_17692_n7109), .B(_abc_17692_n7107), .Y(_abc_17692_n7110) );
  AND2X2 AND2X2_2808 ( .A(_abc_17692_n6751), .B(workunit2_24_), .Y(_abc_17692_n7111) );
  AND2X2 AND2X2_2809 ( .A(_abc_17692_n6939), .B(_abc_17692_n7112), .Y(_abc_17692_n7113) );
  AND2X2 AND2X2_281 ( .A(_abc_17692_n1327), .B(_abc_17692_n1328), .Y(_abc_17692_n1329) );
  AND2X2 AND2X2_2810 ( .A(_abc_17692_n7116), .B(_abc_17692_n1830_bF_buf4), .Y(_abc_17692_n7117) );
  AND2X2 AND2X2_2811 ( .A(_abc_17692_n7117), .B(_abc_17692_n7114), .Y(_abc_17692_n7118) );
  AND2X2 AND2X2_2812 ( .A(_abc_17692_n7121), .B(state_7_bF_buf3), .Y(_abc_17692_n7122) );
  AND2X2 AND2X2_2813 ( .A(_abc_17692_n1885_bF_buf4), .B(workunit2_25_), .Y(_abc_17692_n7123) );
  AND2X2 AND2X2_2814 ( .A(state_8_bF_buf4), .B(\data_in2[25] ), .Y(_abc_17692_n7124) );
  AND2X2 AND2X2_2815 ( .A(_abc_17692_n6666), .B(_abc_17692_n6964), .Y(_abc_17692_n7129) );
  AND2X2 AND2X2_2816 ( .A(_abc_17692_n6675), .B(_abc_17692_n7129), .Y(_abc_17692_n7130) );
  AND2X2 AND2X2_2817 ( .A(_abc_17692_n6963), .B(_abc_17692_n6663), .Y(_abc_17692_n7131) );
  AND2X2 AND2X2_2818 ( .A(_abc_17692_n7134), .B(_abc_17692_n7136), .Y(_abc_17692_n7137) );
  AND2X2 AND2X2_2819 ( .A(_abc_17692_n7138), .B(workunit1_26_), .Y(_abc_17692_n7139) );
  AND2X2 AND2X2_282 ( .A(_abc_17692_n1312), .B(_abc_17692_n1278), .Y(_abc_17692_n1332) );
  AND2X2 AND2X2_2820 ( .A(_abc_17692_n7137), .B(_abc_17692_n6065), .Y(_abc_17692_n7140) );
  AND2X2 AND2X2_2821 ( .A(_abc_17692_n7133), .B(_abc_17692_n7142), .Y(_abc_17692_n7143) );
  AND2X2 AND2X2_2822 ( .A(_abc_17692_n7145), .B(_abc_17692_n7146), .Y(_abc_17692_n7147) );
  AND2X2 AND2X2_2823 ( .A(_abc_17692_n7147), .B(_abc_17692_n7141), .Y(_abc_17692_n7148) );
  AND2X2 AND2X2_2824 ( .A(_abc_17692_n6730), .B(_abc_17692_n7031), .Y(_abc_17692_n7151) );
  AND2X2 AND2X2_2825 ( .A(_abc_17692_n6739), .B(_abc_17692_n7151), .Y(_abc_17692_n7152) );
  AND2X2 AND2X2_2826 ( .A(_abc_17692_n7030), .B(_abc_17692_n6727), .Y(_abc_17692_n7153) );
  AND2X2 AND2X2_2827 ( .A(sum_26_), .B(\key_in[26] ), .Y(_abc_17692_n7156) );
  AND2X2 AND2X2_2828 ( .A(_abc_17692_n7157), .B(_abc_17692_n7158), .Y(_abc_17692_n7159) );
  AND2X2 AND2X2_2829 ( .A(_abc_17692_n7155), .B(_abc_17692_n7159), .Y(_abc_17692_n7160) );
  AND2X2 AND2X2_283 ( .A(_abc_17692_n1312), .B(_abc_17692_n1308_1), .Y(_abc_17692_n1335) );
  AND2X2 AND2X2_2830 ( .A(_abc_17692_n7161), .B(_abc_17692_n7162), .Y(_abc_17692_n7163) );
  AND2X2 AND2X2_2831 ( .A(_abc_17692_n7163), .B(_abc_17692_n7164), .Y(_abc_17692_n7165) );
  AND2X2 AND2X2_2832 ( .A(_abc_17692_n7150), .B(_abc_17692_n7166), .Y(_abc_17692_n7167) );
  AND2X2 AND2X2_2833 ( .A(_abc_17692_n7168), .B(_abc_17692_n7149), .Y(_abc_17692_n7169) );
  AND2X2 AND2X2_2834 ( .A(_abc_17692_n7172), .B(_abc_17692_n7173), .Y(_abc_17692_n7174) );
  AND2X2 AND2X2_2835 ( .A(_abc_17692_n7043), .B(workunit2_25_), .Y(_abc_17692_n7176) );
  AND2X2 AND2X2_2836 ( .A(_abc_17692_n7178), .B(_abc_17692_n7177), .Y(_abc_17692_n7179) );
  AND2X2 AND2X2_2837 ( .A(_abc_17692_n6769), .B(_abc_17692_n7182), .Y(_abc_17692_n7183) );
  AND2X2 AND2X2_2838 ( .A(_abc_17692_n7184), .B(_abc_17692_n7175), .Y(_abc_17692_n7186) );
  AND2X2 AND2X2_2839 ( .A(_abc_17692_n7187), .B(_abc_17692_n1830_bF_buf3), .Y(_abc_17692_n7188) );
  AND2X2 AND2X2_284 ( .A(delta_15_), .B(sum_15_), .Y(_abc_17692_n1336) );
  AND2X2 AND2X2_2840 ( .A(_abc_17692_n7188), .B(_abc_17692_n7185), .Y(_abc_17692_n7189) );
  AND2X2 AND2X2_2841 ( .A(_abc_17692_n6778), .B(_abc_17692_n7002), .Y(_abc_17692_n7190) );
  AND2X2 AND2X2_2842 ( .A(_abc_17692_n7001), .B(_abc_17692_n6775), .Y(_abc_17692_n7193) );
  AND2X2 AND2X2_2843 ( .A(_abc_17692_n7192), .B(_abc_17692_n7195), .Y(_abc_17692_n7196) );
  AND2X2 AND2X2_2844 ( .A(sum_26_), .B(\key_in[90] ), .Y(_abc_17692_n7198) );
  AND2X2 AND2X2_2845 ( .A(_abc_17692_n7199), .B(_abc_17692_n7200), .Y(_abc_17692_n7201) );
  AND2X2 AND2X2_2846 ( .A(_abc_17692_n7197), .B(_abc_17692_n7201), .Y(_abc_17692_n7202) );
  AND2X2 AND2X2_2847 ( .A(_abc_17692_n7196), .B(_abc_17692_n7203), .Y(_abc_17692_n7204) );
  AND2X2 AND2X2_2848 ( .A(_abc_17692_n7207), .B(_abc_17692_n7208), .Y(_abc_17692_n7209) );
  AND2X2 AND2X2_2849 ( .A(_abc_17692_n7209), .B(workunit2_26_), .Y(_abc_17692_n7210) );
  AND2X2 AND2X2_285 ( .A(_abc_17692_n1334), .B(_abc_17692_n1338), .Y(_abc_17692_n1339) );
  AND2X2 AND2X2_2850 ( .A(_abc_17692_n7211), .B(_abc_17692_n7212), .Y(_abc_17692_n7213) );
  AND2X2 AND2X2_2851 ( .A(_abc_17692_n7014), .B(workunit2_25_), .Y(_abc_17692_n7214) );
  AND2X2 AND2X2_2852 ( .A(_abc_17692_n7016), .B(_abc_17692_n7018), .Y(_abc_17692_n7215) );
  AND2X2 AND2X2_2853 ( .A(_abc_17692_n7016), .B(_abc_17692_n6800), .Y(_abc_17692_n7217) );
  AND2X2 AND2X2_2854 ( .A(_abc_17692_n6815), .B(_abc_17692_n7217), .Y(_abc_17692_n7218) );
  AND2X2 AND2X2_2855 ( .A(_abc_17692_n7219), .B(_abc_17692_n7213), .Y(_abc_17692_n7220) );
  AND2X2 AND2X2_2856 ( .A(_abc_17692_n7222), .B(_abc_17692_n1877_bF_buf3), .Y(_abc_17692_n7223) );
  AND2X2 AND2X2_2857 ( .A(_abc_17692_n7223), .B(_abc_17692_n7221), .Y(_abc_17692_n7224) );
  AND2X2 AND2X2_2858 ( .A(_abc_17692_n6824), .B(_abc_17692_n7060), .Y(_abc_17692_n7225) );
  AND2X2 AND2X2_2859 ( .A(_abc_17692_n6833), .B(_abc_17692_n7225), .Y(_abc_17692_n7226) );
  AND2X2 AND2X2_286 ( .A(_abc_17692_n1340), .B(_abc_17692_n1339), .Y(_abc_17692_n1341) );
  AND2X2 AND2X2_2860 ( .A(_abc_17692_n7059), .B(_abc_17692_n6821), .Y(_abc_17692_n7227) );
  AND2X2 AND2X2_2861 ( .A(sum_26_), .B(\key_in[58] ), .Y(_abc_17692_n7230) );
  AND2X2 AND2X2_2862 ( .A(_abc_17692_n7231), .B(_abc_17692_n7232), .Y(_abc_17692_n7233) );
  AND2X2 AND2X2_2863 ( .A(_abc_17692_n7229), .B(_abc_17692_n7233), .Y(_abc_17692_n7234) );
  AND2X2 AND2X2_2864 ( .A(_abc_17692_n7235), .B(_abc_17692_n7236), .Y(_abc_17692_n7237) );
  AND2X2 AND2X2_2865 ( .A(_abc_17692_n7240), .B(_abc_17692_n7238), .Y(_abc_17692_n7241) );
  AND2X2 AND2X2_2866 ( .A(_abc_17692_n7244), .B(_abc_17692_n7242), .Y(_abc_17692_n7245) );
  AND2X2 AND2X2_2867 ( .A(_abc_17692_n7068), .B(workunit2_25_), .Y(_abc_17692_n7247) );
  AND2X2 AND2X2_2868 ( .A(_abc_17692_n7249), .B(_abc_17692_n7248), .Y(_abc_17692_n7250) );
  AND2X2 AND2X2_2869 ( .A(_abc_17692_n7252), .B(_abc_17692_n7250), .Y(_abc_17692_n7253) );
  AND2X2 AND2X2_287 ( .A(_abc_17692_n1342), .B(_abc_17692_n1331_1), .Y(_abc_17692_n1344) );
  AND2X2 AND2X2_2870 ( .A(_abc_17692_n7256), .B(_abc_17692_n1846_bF_buf3), .Y(_abc_17692_n7257) );
  AND2X2 AND2X2_2871 ( .A(_abc_17692_n7257), .B(_abc_17692_n7255), .Y(_abc_17692_n7258) );
  AND2X2 AND2X2_2872 ( .A(_abc_17692_n6685), .B(_abc_17692_n6974), .Y(_abc_17692_n7262) );
  AND2X2 AND2X2_2873 ( .A(_abc_17692_n6694), .B(_abc_17692_n7262), .Y(_abc_17692_n7263) );
  AND2X2 AND2X2_2874 ( .A(_abc_17692_n6973), .B(_abc_17692_n6682), .Y(_abc_17692_n7264) );
  AND2X2 AND2X2_2875 ( .A(sum_26_), .B(\key_in[122] ), .Y(_abc_17692_n7267) );
  AND2X2 AND2X2_2876 ( .A(_abc_17692_n7268), .B(_abc_17692_n7269), .Y(_abc_17692_n7270) );
  AND2X2 AND2X2_2877 ( .A(_abc_17692_n7266), .B(_abc_17692_n7270), .Y(_abc_17692_n7271) );
  AND2X2 AND2X2_2878 ( .A(_abc_17692_n7272), .B(_abc_17692_n7273), .Y(_abc_17692_n7274) );
  AND2X2 AND2X2_2879 ( .A(_abc_17692_n7277), .B(_abc_17692_n7275), .Y(_abc_17692_n7278) );
  AND2X2 AND2X2_288 ( .A(_abc_17692_n1345), .B(state_3_bF_buf3), .Y(_abc_17692_n1346) );
  AND2X2 AND2X2_2880 ( .A(_abc_17692_n7281), .B(_abc_17692_n7279), .Y(_abc_17692_n7282) );
  AND2X2 AND2X2_2881 ( .A(_abc_17692_n6985), .B(workunit2_25_), .Y(_abc_17692_n7283) );
  AND2X2 AND2X2_2882 ( .A(_abc_17692_n6994), .B(_abc_17692_n6707), .Y(_abc_17692_n7284) );
  AND2X2 AND2X2_2883 ( .A(_abc_17692_n6994), .B(_abc_17692_n6709), .Y(_abc_17692_n7287) );
  AND2X2 AND2X2_2884 ( .A(_abc_17692_n7289), .B(_abc_17692_n7286), .Y(_abc_17692_n7290) );
  AND2X2 AND2X2_2885 ( .A(_abc_17692_n7294), .B(_abc_17692_n7291), .Y(_abc_17692_n7295) );
  AND2X2 AND2X2_2886 ( .A(_abc_17692_n7296), .B(state_6_bF_buf3), .Y(_abc_17692_n7297) );
  AND2X2 AND2X2_2887 ( .A(_abc_17692_n7297), .B(_abc_17692_n7261), .Y(_abc_17692_n7298) );
  AND2X2 AND2X2_2888 ( .A(_abc_17692_n6986), .B(_abc_17692_n7089), .Y(_abc_17692_n7299) );
  AND2X2 AND2X2_2889 ( .A(_abc_17692_n6989), .B(_abc_17692_n6708), .Y(_abc_17692_n7302) );
  AND2X2 AND2X2_289 ( .A(_abc_17692_n1346), .B(_abc_17692_n1343_1), .Y(_abc_17692_n1347) );
  AND2X2 AND2X2_2890 ( .A(_abc_17692_n6886), .B(_abc_17692_n7302), .Y(_abc_17692_n7303) );
  AND2X2 AND2X2_2891 ( .A(_abc_17692_n7304), .B(_abc_17692_n7282), .Y(_abc_17692_n7305) );
  AND2X2 AND2X2_2892 ( .A(_abc_17692_n7307), .B(_abc_17692_n1863_bF_buf1), .Y(_abc_17692_n7308) );
  AND2X2 AND2X2_2893 ( .A(_abc_17692_n7308), .B(_abc_17692_n7306), .Y(_abc_17692_n7309) );
  AND2X2 AND2X2_2894 ( .A(_abc_17692_n6906), .B(_abc_17692_n7316), .Y(_abc_17692_n7317) );
  AND2X2 AND2X2_2895 ( .A(_abc_17692_n7318), .B(_abc_17692_n7310), .Y(_abc_17692_n7319) );
  AND2X2 AND2X2_2896 ( .A(_abc_17692_n7321), .B(_abc_17692_n1877_bF_buf2), .Y(_abc_17692_n7322) );
  AND2X2 AND2X2_2897 ( .A(_abc_17692_n7322), .B(_abc_17692_n7320), .Y(_abc_17692_n7323) );
  AND2X2 AND2X2_2898 ( .A(_abc_17692_n7325), .B(_abc_17692_n7073), .Y(_abc_17692_n7326) );
  AND2X2 AND2X2_2899 ( .A(_abc_17692_n7074), .B(_abc_17692_n6848), .Y(_abc_17692_n7327) );
  AND2X2 AND2X2_29 ( .A(_abc_17692_n693_1), .B(_abc_17692_n691), .Y(x_6__FF_INPUT) );
  AND2X2 AND2X2_290 ( .A(_abc_17692_n1290), .B(_abc_17692_n1307), .Y(_abc_17692_n1348) );
  AND2X2 AND2X2_2900 ( .A(_abc_17692_n6920), .B(_abc_17692_n7327), .Y(_abc_17692_n7328) );
  AND2X2 AND2X2_2901 ( .A(_abc_17692_n7329), .B(_abc_17692_n7245), .Y(_abc_17692_n7330) );
  AND2X2 AND2X2_2902 ( .A(_abc_17692_n7332), .B(_abc_17692_n1846_bF_buf2), .Y(_abc_17692_n7333) );
  AND2X2 AND2X2_2903 ( .A(_abc_17692_n7333), .B(_abc_17692_n7331), .Y(_abc_17692_n7334) );
  AND2X2 AND2X2_2904 ( .A(_abc_17692_n7045), .B(_abc_17692_n7335), .Y(_abc_17692_n7336) );
  AND2X2 AND2X2_2905 ( .A(_abc_17692_n7046), .B(_abc_17692_n6754), .Y(_abc_17692_n7337) );
  AND2X2 AND2X2_2906 ( .A(_abc_17692_n6937), .B(_abc_17692_n7337), .Y(_abc_17692_n7338) );
  AND2X2 AND2X2_2907 ( .A(_abc_17692_n7339), .B(_abc_17692_n7174), .Y(_abc_17692_n7340) );
  AND2X2 AND2X2_2908 ( .A(_abc_17692_n7342), .B(_abc_17692_n1830_bF_buf2), .Y(_abc_17692_n7343) );
  AND2X2 AND2X2_2909 ( .A(_abc_17692_n7343), .B(_abc_17692_n7341), .Y(_abc_17692_n7344) );
  AND2X2 AND2X2_291 ( .A(_abc_17692_n1292), .B(_abc_17692_n1348), .Y(_abc_17692_n1349) );
  AND2X2 AND2X2_2910 ( .A(_abc_17692_n7347), .B(state_7_bF_buf2), .Y(_abc_17692_n7348) );
  AND2X2 AND2X2_2911 ( .A(_abc_17692_n1885_bF_buf3), .B(workunit2_26_), .Y(_abc_17692_n7349) );
  AND2X2 AND2X2_2912 ( .A(state_8_bF_buf3), .B(\data_in2[26] ), .Y(_abc_17692_n7350) );
  AND2X2 AND2X2_2913 ( .A(_abc_17692_n7355), .B(_abc_17692_n7354), .Y(_abc_17692_n7356) );
  AND2X2 AND2X2_2914 ( .A(workunit1_23_), .B(workunit1_27_), .Y(_abc_17692_n7357) );
  AND2X2 AND2X2_2915 ( .A(_abc_17692_n5378), .B(_abc_17692_n6242), .Y(_abc_17692_n7358) );
  AND2X2 AND2X2_2916 ( .A(_abc_17692_n7361), .B(_abc_17692_n7363), .Y(_abc_17692_n7364) );
  AND2X2 AND2X2_2917 ( .A(sum_27_), .B(\key_in[123] ), .Y(_abc_17692_n7366) );
  AND2X2 AND2X2_2918 ( .A(_abc_17692_n7367), .B(_abc_17692_n7368), .Y(_abc_17692_n7369) );
  AND2X2 AND2X2_2919 ( .A(_abc_17692_n7365), .B(_abc_17692_n7370), .Y(_abc_17692_n7372) );
  AND2X2 AND2X2_292 ( .A(_abc_17692_n1348), .B(_abc_17692_n1262), .Y(_abc_17692_n1350) );
  AND2X2 AND2X2_2920 ( .A(_abc_17692_n7373), .B(_abc_17692_n7371), .Y(_abc_17692_n7374) );
  AND2X2 AND2X2_2921 ( .A(_abc_17692_n7362), .B(_abc_17692_n7359), .Y(_abc_17692_n7376) );
  AND2X2 AND2X2_2922 ( .A(_abc_17692_n7356), .B(_abc_17692_n7360), .Y(_abc_17692_n7377) );
  AND2X2 AND2X2_2923 ( .A(_abc_17692_n7379), .B(_abc_17692_n7369), .Y(_abc_17692_n7380) );
  AND2X2 AND2X2_2924 ( .A(_abc_17692_n7382), .B(_abc_17692_n7375), .Y(_abc_17692_n7383) );
  AND2X2 AND2X2_2925 ( .A(_abc_17692_n7383), .B(workunit2_27_), .Y(_abc_17692_n7384) );
  AND2X2 AND2X2_2926 ( .A(_abc_17692_n7386), .B(_abc_17692_n7387), .Y(_abc_17692_n7388) );
  AND2X2 AND2X2_2927 ( .A(_abc_17692_n7388), .B(_abc_17692_n7385), .Y(_abc_17692_n7389) );
  AND2X2 AND2X2_2928 ( .A(_abc_17692_n7395), .B(_abc_17692_n7396), .Y(_abc_17692_n7397) );
  AND2X2 AND2X2_2929 ( .A(_abc_17692_n7398), .B(_abc_17692_n1863_bF_buf0), .Y(_abc_17692_n7399) );
  AND2X2 AND2X2_293 ( .A(_abc_17692_n1231), .B(_abc_17692_n1350), .Y(_abc_17692_n1351) );
  AND2X2 AND2X2_2930 ( .A(_abc_17692_n7399), .B(_abc_17692_n7394), .Y(_abc_17692_n7400) );
  AND2X2 AND2X2_2931 ( .A(_abc_17692_n7401), .B(_abc_17692_n7199), .Y(_abc_17692_n7402) );
  AND2X2 AND2X2_2932 ( .A(sum_27_), .B(\key_in[91] ), .Y(_abc_17692_n7403) );
  AND2X2 AND2X2_2933 ( .A(_abc_17692_n7404), .B(_abc_17692_n7405), .Y(_abc_17692_n7406) );
  AND2X2 AND2X2_2934 ( .A(_abc_17692_n7402), .B(_abc_17692_n7406), .Y(_abc_17692_n7407) );
  AND2X2 AND2X2_2935 ( .A(_abc_17692_n7408), .B(_abc_17692_n7409), .Y(_abc_17692_n7410) );
  AND2X2 AND2X2_2936 ( .A(_abc_17692_n7412), .B(_abc_17692_n7413), .Y(_abc_17692_n7414) );
  AND2X2 AND2X2_2937 ( .A(_abc_17692_n7416), .B(_abc_17692_n7411), .Y(_abc_17692_n7417) );
  AND2X2 AND2X2_2938 ( .A(_abc_17692_n7417), .B(workunit2_27_), .Y(_abc_17692_n7418) );
  AND2X2 AND2X2_2939 ( .A(_abc_17692_n7419), .B(_abc_17692_n7420), .Y(_abc_17692_n7421) );
  AND2X2 AND2X2_294 ( .A(_abc_17692_n1352), .B(_abc_17692_n1350), .Y(_abc_17692_n1353) );
  AND2X2 AND2X2_2940 ( .A(_abc_17692_n7421), .B(_abc_17692_n7385), .Y(_abc_17692_n7422) );
  AND2X2 AND2X2_2941 ( .A(_abc_17692_n7425), .B(workunit2_26_), .Y(_abc_17692_n7426) );
  AND2X2 AND2X2_2942 ( .A(_abc_17692_n7320), .B(_abc_17692_n7427), .Y(_abc_17692_n7428) );
  AND2X2 AND2X2_2943 ( .A(_abc_17692_n7431), .B(_abc_17692_n1877_bF_buf1), .Y(_abc_17692_n7432) );
  AND2X2 AND2X2_2944 ( .A(_abc_17692_n7432), .B(_abc_17692_n7430), .Y(_abc_17692_n7433) );
  AND2X2 AND2X2_2945 ( .A(_abc_17692_n7235), .B(_abc_17692_n7231), .Y(_abc_17692_n7434) );
  AND2X2 AND2X2_2946 ( .A(sum_27_), .B(\key_in[59] ), .Y(_abc_17692_n7435) );
  AND2X2 AND2X2_2947 ( .A(_abc_17692_n7436), .B(_abc_17692_n7437), .Y(_abc_17692_n7438) );
  AND2X2 AND2X2_2948 ( .A(_abc_17692_n7434), .B(_abc_17692_n7438), .Y(_abc_17692_n7439) );
  AND2X2 AND2X2_2949 ( .A(_abc_17692_n7440), .B(_abc_17692_n7441), .Y(_abc_17692_n7442) );
  AND2X2 AND2X2_295 ( .A(_abc_17692_n1354), .B(_abc_17692_n1306), .Y(_abc_17692_n1355_1) );
  AND2X2 AND2X2_2950 ( .A(_abc_17692_n7446), .B(_abc_17692_n7445), .Y(_abc_17692_n7447) );
  AND2X2 AND2X2_2951 ( .A(_abc_17692_n7444), .B(_abc_17692_n7448), .Y(_abc_17692_n7449) );
  AND2X2 AND2X2_2952 ( .A(_abc_17692_n7451), .B(_abc_17692_n7452), .Y(_abc_17692_n7453) );
  AND2X2 AND2X2_2953 ( .A(_abc_17692_n7450), .B(_abc_17692_n7454), .Y(_abc_17692_n7455) );
  AND2X2 AND2X2_2954 ( .A(_abc_17692_n7331), .B(_abc_17692_n7242), .Y(_abc_17692_n7456) );
  AND2X2 AND2X2_2955 ( .A(_abc_17692_n7460), .B(_abc_17692_n1846_bF_buf1), .Y(_abc_17692_n7461) );
  AND2X2 AND2X2_2956 ( .A(_abc_17692_n7461), .B(_abc_17692_n7458), .Y(_abc_17692_n7462) );
  AND2X2 AND2X2_2957 ( .A(_abc_17692_n7463), .B(_abc_17692_n7157), .Y(_abc_17692_n7464) );
  AND2X2 AND2X2_2958 ( .A(sum_27_), .B(\key_in[27] ), .Y(_abc_17692_n7465) );
  AND2X2 AND2X2_2959 ( .A(_abc_17692_n7466), .B(_abc_17692_n7467), .Y(_abc_17692_n7468) );
  AND2X2 AND2X2_296 ( .A(_abc_17692_n1359), .B(_abc_17692_n1330), .Y(_abc_17692_n1360) );
  AND2X2 AND2X2_2960 ( .A(_abc_17692_n7464), .B(_abc_17692_n7468), .Y(_abc_17692_n7469) );
  AND2X2 AND2X2_2961 ( .A(_abc_17692_n7470), .B(_abc_17692_n7471), .Y(_abc_17692_n7472) );
  AND2X2 AND2X2_2962 ( .A(_abc_17692_n7476), .B(_abc_17692_n7475), .Y(_abc_17692_n7477) );
  AND2X2 AND2X2_2963 ( .A(_abc_17692_n7474), .B(_abc_17692_n7478), .Y(_abc_17692_n7479) );
  AND2X2 AND2X2_2964 ( .A(_abc_17692_n7481), .B(_abc_17692_n7482), .Y(_abc_17692_n7483) );
  AND2X2 AND2X2_2965 ( .A(_abc_17692_n7480), .B(_abc_17692_n7484), .Y(_abc_17692_n7485) );
  AND2X2 AND2X2_2966 ( .A(_abc_17692_n7341), .B(_abc_17692_n7172), .Y(_abc_17692_n7487) );
  AND2X2 AND2X2_2967 ( .A(_abc_17692_n7490), .B(_abc_17692_n1830_bF_buf1), .Y(_abc_17692_n7491) );
  AND2X2 AND2X2_2968 ( .A(_abc_17692_n7491), .B(_abc_17692_n7488), .Y(_abc_17692_n7492) );
  AND2X2 AND2X2_2969 ( .A(_abc_17692_n7495), .B(state_7_bF_buf1), .Y(_abc_17692_n7496) );
  AND2X2 AND2X2_297 ( .A(_abc_17692_n1362), .B(state_15_bF_buf3), .Y(_abc_17692_n1363) );
  AND2X2 AND2X2_2970 ( .A(_abc_17692_n7291), .B(_abc_17692_n7497), .Y(_abc_17692_n7498) );
  AND2X2 AND2X2_2971 ( .A(_abc_17692_n7499), .B(_abc_17692_n7397), .Y(_abc_17692_n7500) );
  AND2X2 AND2X2_2972 ( .A(_abc_17692_n7498), .B(_abc_17692_n7390), .Y(_abc_17692_n7501) );
  AND2X2 AND2X2_2973 ( .A(_abc_17692_n7507), .B(_abc_17692_n1877_bF_buf0), .Y(_abc_17692_n7508) );
  AND2X2 AND2X2_2974 ( .A(_abc_17692_n7508), .B(_abc_17692_n7506), .Y(_abc_17692_n7509) );
  AND2X2 AND2X2_2975 ( .A(_abc_17692_n7171), .B(workunit2_26_), .Y(_abc_17692_n7510) );
  AND2X2 AND2X2_2976 ( .A(_abc_17692_n7514), .B(_abc_17692_n1830_bF_buf0), .Y(_abc_17692_n7515) );
  AND2X2 AND2X2_2977 ( .A(_abc_17692_n7515), .B(_abc_17692_n7513), .Y(_abc_17692_n7516) );
  AND2X2 AND2X2_2978 ( .A(_abc_17692_n7241), .B(workunit2_26_), .Y(_abc_17692_n7517) );
  AND2X2 AND2X2_2979 ( .A(_abc_17692_n7256), .B(_abc_17692_n7518), .Y(_abc_17692_n7519) );
  AND2X2 AND2X2_298 ( .A(_abc_17692_n1363), .B(_abc_17692_n1361), .Y(_abc_17692_n1364) );
  AND2X2 AND2X2_2980 ( .A(_abc_17692_n7522), .B(_abc_17692_n1846_bF_buf0), .Y(_abc_17692_n7523) );
  AND2X2 AND2X2_2981 ( .A(_abc_17692_n7523), .B(_abc_17692_n7521), .Y(_abc_17692_n7524) );
  AND2X2 AND2X2_2982 ( .A(_abc_17692_n7527), .B(state_6_bF_buf2), .Y(_abc_17692_n7528) );
  AND2X2 AND2X2_2983 ( .A(_abc_17692_n7528), .B(_abc_17692_n7503), .Y(_abc_17692_n7529) );
  AND2X2 AND2X2_2984 ( .A(_abc_17692_n1885_bF_buf2), .B(workunit2_27_), .Y(_abc_17692_n7530) );
  AND2X2 AND2X2_2985 ( .A(state_8_bF_buf2), .B(\data_in2[27] ), .Y(_abc_17692_n7531) );
  AND2X2 AND2X2_2986 ( .A(_abc_17692_n7142), .B(_abc_17692_n7360), .Y(_abc_17692_n7536) );
  AND2X2 AND2X2_2987 ( .A(_abc_17692_n7130), .B(_abc_17692_n7536), .Y(_abc_17692_n7537) );
  AND2X2 AND2X2_2988 ( .A(_abc_17692_n7536), .B(_abc_17692_n7132), .Y(_abc_17692_n7538) );
  AND2X2 AND2X2_2989 ( .A(_abc_17692_n7139), .B(_abc_17692_n7360), .Y(_abc_17692_n7539) );
  AND2X2 AND2X2_299 ( .A(_abc_17692_n722_bF_buf0), .B(sum_16_), .Y(_abc_17692_n1365) );
  AND2X2 AND2X2_2990 ( .A(workunit1_24_), .B(workunit1_28_), .Y(_abc_17692_n7543) );
  AND2X2 AND2X2_2991 ( .A(_abc_17692_n5598), .B(_abc_17692_n6468_1), .Y(_abc_17692_n7544) );
  AND2X2 AND2X2_2992 ( .A(_abc_17692_n7542), .B(_abc_17692_n7546), .Y(_abc_17692_n7547) );
  AND2X2 AND2X2_2993 ( .A(_abc_17692_n7548), .B(_abc_17692_n7549), .Y(_abc_17692_n7550) );
  AND2X2 AND2X2_2994 ( .A(sum_28_), .B(\key_in[124] ), .Y(_abc_17692_n7551) );
  AND2X2 AND2X2_2995 ( .A(_abc_17692_n7552), .B(_abc_17692_n7553), .Y(_abc_17692_n7554) );
  AND2X2 AND2X2_2996 ( .A(_abc_17692_n7268), .B(_abc_17692_n7367), .Y(_abc_17692_n7555) );
  AND2X2 AND2X2_2997 ( .A(_abc_17692_n7557), .B(_abc_17692_n7368), .Y(_abc_17692_n7558) );
  AND2X2 AND2X2_2998 ( .A(_abc_17692_n7558), .B(_abc_17692_n7554), .Y(_abc_17692_n7559) );
  AND2X2 AND2X2_2999 ( .A(_abc_17692_n7561), .B(_abc_17692_n7560), .Y(_abc_17692_n7562) );
  AND2X2 AND2X2_3 ( .A(_abc_17692_n633), .B(_abc_17692_n631), .Y(modereg_FF_INPUT) );
  AND2X2 AND2X2_30 ( .A(_abc_17692_n692_1), .B(x_7_), .Y(_abc_17692_n696) );
  AND2X2 AND2X2_300 ( .A(delta_17_), .B(sum_17_), .Y(_abc_17692_n1369) );
  AND2X2 AND2X2_3000 ( .A(_abc_17692_n7563), .B(_abc_17692_n7550), .Y(_abc_17692_n7564) );
  AND2X2 AND2X2_3001 ( .A(_abc_17692_n7566), .B(_abc_17692_n7565), .Y(_abc_17692_n7567) );
  AND2X2 AND2X2_3002 ( .A(_abc_17692_n7571), .B(_abc_17692_n7569), .Y(_abc_17692_n7572) );
  AND2X2 AND2X2_3003 ( .A(_abc_17692_n7390), .B(_abc_17692_n7292), .Y(_abc_17692_n7573) );
  AND2X2 AND2X2_3004 ( .A(_abc_17692_n7573), .B(_abc_17692_n7287), .Y(_abc_17692_n7574) );
  AND2X2 AND2X2_3005 ( .A(_abc_17692_n7285), .B(_abc_17692_n7573), .Y(_abc_17692_n7577) );
  AND2X2 AND2X2_3006 ( .A(_abc_17692_n7388), .B(workunit2_27_), .Y(_abc_17692_n7579) );
  AND2X2 AND2X2_3007 ( .A(_abc_17692_n7581), .B(_abc_17692_n7580), .Y(_abc_17692_n7582) );
  AND2X2 AND2X2_3008 ( .A(_abc_17692_n7578), .B(_abc_17692_n7582), .Y(_abc_17692_n7583) );
  AND2X2 AND2X2_3009 ( .A(_abc_17692_n7576), .B(_abc_17692_n7583), .Y(_abc_17692_n7584) );
  AND2X2 AND2X2_301 ( .A(_abc_17692_n1371), .B(_abc_17692_n1372), .Y(_abc_17692_n1373) );
  AND2X2 AND2X2_3010 ( .A(_abc_17692_n7586), .B(_abc_17692_n7588), .Y(_abc_17692_n7589) );
  AND2X2 AND2X2_3011 ( .A(sum_28_), .B(\key_in[28] ), .Y(_abc_17692_n7591) );
  AND2X2 AND2X2_3012 ( .A(_abc_17692_n7592), .B(_abc_17692_n7593), .Y(_abc_17692_n7594) );
  AND2X2 AND2X2_3013 ( .A(_abc_17692_n7157), .B(_abc_17692_n7466), .Y(_abc_17692_n7595) );
  AND2X2 AND2X2_3014 ( .A(_abc_17692_n7597), .B(_abc_17692_n7467), .Y(_abc_17692_n7598) );
  AND2X2 AND2X2_3015 ( .A(_abc_17692_n7598), .B(_abc_17692_n7594), .Y(_abc_17692_n7599) );
  AND2X2 AND2X2_3016 ( .A(_abc_17692_n7601), .B(_abc_17692_n7600), .Y(_abc_17692_n7602) );
  AND2X2 AND2X2_3017 ( .A(_abc_17692_n7603), .B(_abc_17692_n7550), .Y(_abc_17692_n7604) );
  AND2X2 AND2X2_3018 ( .A(_abc_17692_n7605), .B(_abc_17692_n7565), .Y(_abc_17692_n7606) );
  AND2X2 AND2X2_3019 ( .A(_abc_17692_n7609), .B(_abc_17692_n7610), .Y(_abc_17692_n7611) );
  AND2X2 AND2X2_302 ( .A(_abc_17692_n1374), .B(_abc_17692_n1370), .Y(_abc_17692_n1375) );
  AND2X2 AND2X2_3020 ( .A(_abc_17692_n7486), .B(_abc_17692_n7175), .Y(_abc_17692_n7613) );
  AND2X2 AND2X2_3021 ( .A(_abc_17692_n7182), .B(_abc_17692_n7613), .Y(_abc_17692_n7614) );
  AND2X2 AND2X2_3022 ( .A(_abc_17692_n7479), .B(workunit2_27_), .Y(_abc_17692_n7619) );
  AND2X2 AND2X2_3023 ( .A(_abc_17692_n7486), .B(_abc_17692_n7510), .Y(_abc_17692_n7620) );
  AND2X2 AND2X2_3024 ( .A(_abc_17692_n7618), .B(_abc_17692_n7622), .Y(_abc_17692_n7623) );
  AND2X2 AND2X2_3025 ( .A(_abc_17692_n7616), .B(_abc_17692_n7623), .Y(_abc_17692_n7624) );
  AND2X2 AND2X2_3026 ( .A(_abc_17692_n7625), .B(_abc_17692_n7612), .Y(_abc_17692_n7627) );
  AND2X2 AND2X2_3027 ( .A(_abc_17692_n7628), .B(_abc_17692_n1830_bF_buf10), .Y(_abc_17692_n7629) );
  AND2X2 AND2X2_3028 ( .A(_abc_17692_n7629), .B(_abc_17692_n7626), .Y(_abc_17692_n7630) );
  AND2X2 AND2X2_3029 ( .A(sum_28_), .B(\key_in[92] ), .Y(_abc_17692_n7631) );
  AND2X2 AND2X2_303 ( .A(_abc_17692_n1345), .B(_abc_17692_n1376), .Y(_abc_17692_n1377) );
  AND2X2 AND2X2_3030 ( .A(_abc_17692_n7632), .B(_abc_17692_n7633), .Y(_abc_17692_n7634) );
  AND2X2 AND2X2_3031 ( .A(_abc_17692_n7199), .B(_abc_17692_n7404), .Y(_abc_17692_n7636) );
  AND2X2 AND2X2_3032 ( .A(_abc_17692_n7401), .B(_abc_17692_n7636), .Y(_abc_17692_n7637) );
  AND2X2 AND2X2_3033 ( .A(_abc_17692_n7639), .B(_abc_17692_n7634), .Y(_abc_17692_n7640) );
  AND2X2 AND2X2_3034 ( .A(_abc_17692_n7638), .B(_abc_17692_n7641), .Y(_abc_17692_n7642) );
  AND2X2 AND2X2_3035 ( .A(_abc_17692_n7645), .B(_abc_17692_n7646), .Y(_abc_17692_n7647) );
  AND2X2 AND2X2_3036 ( .A(_abc_17692_n7647), .B(workunit2_28_), .Y(_abc_17692_n7648) );
  AND2X2 AND2X2_3037 ( .A(_abc_17692_n7649), .B(_abc_17692_n7650), .Y(_abc_17692_n7651) );
  AND2X2 AND2X2_3038 ( .A(_abc_17692_n7655), .B(_abc_17692_n6815), .Y(_abc_17692_n7656) );
  AND2X2 AND2X2_3039 ( .A(_abc_17692_n7421), .B(workunit2_27_), .Y(_abc_17692_n7659) );
  AND2X2 AND2X2_304 ( .A(_abc_17692_n1381), .B(state_3_bF_buf2), .Y(_abc_17692_n1382) );
  AND2X2 AND2X2_3040 ( .A(_abc_17692_n7423), .B(_abc_17692_n7210), .Y(_abc_17692_n7660) );
  AND2X2 AND2X2_3041 ( .A(_abc_17692_n7658), .B(_abc_17692_n7662), .Y(_abc_17692_n7663) );
  AND2X2 AND2X2_3042 ( .A(_abc_17692_n7665), .B(_abc_17692_n7651), .Y(_abc_17692_n7666) );
  AND2X2 AND2X2_3043 ( .A(_abc_17692_n7668), .B(_abc_17692_n1877_bF_buf10), .Y(_abc_17692_n7669) );
  AND2X2 AND2X2_3044 ( .A(_abc_17692_n7669), .B(_abc_17692_n7667), .Y(_abc_17692_n7670) );
  AND2X2 AND2X2_3045 ( .A(sum_28_), .B(\key_in[60] ), .Y(_abc_17692_n7671) );
  AND2X2 AND2X2_3046 ( .A(_abc_17692_n7672), .B(_abc_17692_n7673), .Y(_abc_17692_n7674) );
  AND2X2 AND2X2_3047 ( .A(_abc_17692_n7231), .B(_abc_17692_n7436), .Y(_abc_17692_n7675) );
  AND2X2 AND2X2_3048 ( .A(_abc_17692_n7677), .B(_abc_17692_n7437), .Y(_abc_17692_n7678) );
  AND2X2 AND2X2_3049 ( .A(_abc_17692_n7678), .B(_abc_17692_n7674), .Y(_abc_17692_n7679) );
  AND2X2 AND2X2_305 ( .A(_abc_17692_n1382), .B(_abc_17692_n1379), .Y(_abc_17692_n1383) );
  AND2X2 AND2X2_3050 ( .A(_abc_17692_n7681), .B(_abc_17692_n7680), .Y(_abc_17692_n7682) );
  AND2X2 AND2X2_3051 ( .A(_abc_17692_n7683), .B(_abc_17692_n7550), .Y(_abc_17692_n7684) );
  AND2X2 AND2X2_3052 ( .A(_abc_17692_n7685), .B(_abc_17692_n7565), .Y(_abc_17692_n7686) );
  AND2X2 AND2X2_3053 ( .A(_abc_17692_n7689), .B(_abc_17692_n7690), .Y(_abc_17692_n7691) );
  AND2X2 AND2X2_3054 ( .A(_abc_17692_n7449), .B(workunit2_27_), .Y(_abc_17692_n7697) );
  AND2X2 AND2X2_3055 ( .A(_abc_17692_n7699), .B(_abc_17692_n7698), .Y(_abc_17692_n7700) );
  AND2X2 AND2X2_3056 ( .A(_abc_17692_n7696), .B(_abc_17692_n7700), .Y(_abc_17692_n7701) );
  AND2X2 AND2X2_3057 ( .A(_abc_17692_n7695), .B(_abc_17692_n7701), .Y(_abc_17692_n7702) );
  AND2X2 AND2X2_3058 ( .A(_abc_17692_n7703), .B(_abc_17692_n7692), .Y(_abc_17692_n7704) );
  AND2X2 AND2X2_3059 ( .A(_abc_17692_n7706), .B(_abc_17692_n1846_bF_buf10), .Y(_abc_17692_n7707) );
  AND2X2 AND2X2_306 ( .A(_abc_17692_n1327), .B(sum_16_), .Y(_abc_17692_n1384) );
  AND2X2 AND2X2_3060 ( .A(_abc_17692_n7707), .B(_abc_17692_n7705), .Y(_abc_17692_n7708) );
  AND2X2 AND2X2_3061 ( .A(_abc_17692_n7711), .B(state_6_bF_buf1), .Y(_abc_17692_n7712) );
  AND2X2 AND2X2_3062 ( .A(_abc_17692_n7712), .B(_abc_17692_n7590), .Y(_abc_17692_n7713) );
  AND2X2 AND2X2_3063 ( .A(_abc_17692_n7397), .B(_abc_17692_n7282), .Y(_abc_17692_n7714) );
  AND2X2 AND2X2_3064 ( .A(_abc_17692_n7714), .B(_abc_17692_n7302), .Y(_abc_17692_n7715) );
  AND2X2 AND2X2_3065 ( .A(_abc_17692_n6886), .B(_abc_17692_n7715), .Y(_abc_17692_n7716) );
  AND2X2 AND2X2_3066 ( .A(_abc_17692_n7714), .B(_abc_17692_n7301), .Y(_abc_17692_n7717) );
  AND2X2 AND2X2_3067 ( .A(_abc_17692_n7396), .B(_abc_17692_n7391), .Y(_abc_17692_n7718) );
  AND2X2 AND2X2_3068 ( .A(_abc_17692_n7721), .B(_abc_17692_n7587), .Y(_abc_17692_n7723) );
  AND2X2 AND2X2_3069 ( .A(_abc_17692_n7724), .B(_abc_17692_n1863_bF_buf8), .Y(_abc_17692_n7725) );
  AND2X2 AND2X2_307 ( .A(_abc_17692_n1360), .B(_abc_17692_n1380), .Y(_abc_17692_n1387) );
  AND2X2 AND2X2_3070 ( .A(_abc_17692_n7725), .B(_abc_17692_n7722), .Y(_abc_17692_n7726) );
  AND2X2 AND2X2_3071 ( .A(_abc_17692_n7733), .B(_abc_17692_n7732), .Y(_abc_17692_n7734) );
  AND2X2 AND2X2_3072 ( .A(_abc_17692_n7731), .B(_abc_17692_n7735), .Y(_abc_17692_n7736) );
  AND2X2 AND2X2_3073 ( .A(_abc_17692_n7730), .B(_abc_17692_n7736), .Y(_abc_17692_n7737) );
  AND2X2 AND2X2_3074 ( .A(_abc_17692_n7738), .B(_abc_17692_n7727), .Y(_abc_17692_n7739) );
  AND2X2 AND2X2_3075 ( .A(_abc_17692_n7741), .B(_abc_17692_n1877_bF_buf9), .Y(_abc_17692_n7742) );
  AND2X2 AND2X2_3076 ( .A(_abc_17692_n7742), .B(_abc_17692_n7740), .Y(_abc_17692_n7743) );
  AND2X2 AND2X2_3077 ( .A(_abc_17692_n7455), .B(_abc_17692_n7245), .Y(_abc_17692_n7744) );
  AND2X2 AND2X2_3078 ( .A(_abc_17692_n7744), .B(_abc_17692_n7327), .Y(_abc_17692_n7745) );
  AND2X2 AND2X2_3079 ( .A(_abc_17692_n6920), .B(_abc_17692_n7745), .Y(_abc_17692_n7746) );
  AND2X2 AND2X2_308 ( .A(_abc_17692_n1380), .B(_abc_17692_n1384), .Y(_abc_17692_n1389_1) );
  AND2X2 AND2X2_3080 ( .A(_abc_17692_n7744), .B(_abc_17692_n7326), .Y(_abc_17692_n7747) );
  AND2X2 AND2X2_3081 ( .A(_abc_17692_n7750), .B(_abc_17692_n7454), .Y(_abc_17692_n7751) );
  AND2X2 AND2X2_3082 ( .A(_abc_17692_n7753), .B(_abc_17692_n7691), .Y(_abc_17692_n7755) );
  AND2X2 AND2X2_3083 ( .A(_abc_17692_n7756), .B(_abc_17692_n1846_bF_buf9), .Y(_abc_17692_n7757) );
  AND2X2 AND2X2_3084 ( .A(_abc_17692_n7757), .B(_abc_17692_n7754), .Y(_abc_17692_n7758) );
  AND2X2 AND2X2_3085 ( .A(_abc_17692_n7485), .B(_abc_17692_n7174), .Y(_abc_17692_n7759) );
  AND2X2 AND2X2_3086 ( .A(_abc_17692_n7759), .B(_abc_17692_n7337), .Y(_abc_17692_n7760) );
  AND2X2 AND2X2_3087 ( .A(_abc_17692_n6937), .B(_abc_17692_n7760), .Y(_abc_17692_n7761) );
  AND2X2 AND2X2_3088 ( .A(_abc_17692_n7759), .B(_abc_17692_n7336), .Y(_abc_17692_n7762) );
  AND2X2 AND2X2_3089 ( .A(_abc_17692_n7484), .B(_abc_17692_n7764), .Y(_abc_17692_n7765) );
  AND2X2 AND2X2_309 ( .A(_abc_17692_n1390), .B(state_15_bF_buf2), .Y(_abc_17692_n1391) );
  AND2X2 AND2X2_3090 ( .A(_abc_17692_n7768), .B(_abc_17692_n7611), .Y(_abc_17692_n7769) );
  AND2X2 AND2X2_3091 ( .A(_abc_17692_n7771), .B(_abc_17692_n1830_bF_buf9), .Y(_abc_17692_n7772) );
  AND2X2 AND2X2_3092 ( .A(_abc_17692_n7772), .B(_abc_17692_n7770), .Y(_abc_17692_n7773) );
  AND2X2 AND2X2_3093 ( .A(_abc_17692_n7776), .B(state_7_bF_buf0), .Y(_abc_17692_n7777) );
  AND2X2 AND2X2_3094 ( .A(_abc_17692_n1885_bF_buf1), .B(workunit2_28_), .Y(_abc_17692_n7778) );
  AND2X2 AND2X2_3095 ( .A(state_8_bF_buf1), .B(\data_in2[28] ), .Y(_abc_17692_n7779) );
  AND2X2 AND2X2_3096 ( .A(workunit1_25_), .B(workunit1_29_), .Y(_abc_17692_n7784) );
  AND2X2 AND2X2_3097 ( .A(_abc_17692_n5782), .B(_abc_17692_n6659_1), .Y(_abc_17692_n7786) );
  AND2X2 AND2X2_3098 ( .A(_abc_17692_n7787), .B(_abc_17692_n7785), .Y(_abc_17692_n7788) );
  AND2X2 AND2X2_3099 ( .A(_abc_17692_n7783), .B(_abc_17692_n7788), .Y(_abc_17692_n7790) );
  AND2X2 AND2X2_31 ( .A(_abc_17692_n697), .B(_abc_17692_n695), .Y(x_7__FF_INPUT) );
  AND2X2 AND2X2_310 ( .A(_abc_17692_n1388), .B(_abc_17692_n1391), .Y(_abc_17692_n1392_1) );
  AND2X2 AND2X2_3100 ( .A(_abc_17692_n7791), .B(_abc_17692_n7789), .Y(_abc_17692_n7792) );
  AND2X2 AND2X2_3101 ( .A(_abc_17692_n7793), .B(_abc_17692_n7632), .Y(_abc_17692_n7794) );
  AND2X2 AND2X2_3102 ( .A(sum_29_), .B(\key_in[93] ), .Y(_abc_17692_n7795) );
  AND2X2 AND2X2_3103 ( .A(_abc_17692_n7796), .B(_abc_17692_n7797), .Y(_abc_17692_n7798) );
  AND2X2 AND2X2_3104 ( .A(_abc_17692_n7794), .B(_abc_17692_n7799), .Y(_abc_17692_n7800) );
  AND2X2 AND2X2_3105 ( .A(_abc_17692_n7801), .B(_abc_17692_n7802), .Y(_abc_17692_n7803) );
  AND2X2 AND2X2_3106 ( .A(_abc_17692_n7806), .B(_abc_17692_n7798), .Y(_abc_17692_n7807) );
  AND2X2 AND2X2_3107 ( .A(_abc_17692_n7809), .B(_abc_17692_n7804), .Y(_abc_17692_n7810) );
  AND2X2 AND2X2_3108 ( .A(_abc_17692_n7810), .B(workunit2_29_), .Y(_abc_17692_n7811) );
  AND2X2 AND2X2_3109 ( .A(_abc_17692_n7808), .B(_abc_17692_n7805), .Y(_abc_17692_n7813) );
  AND2X2 AND2X2_311 ( .A(_abc_17692_n1392_1), .B(_abc_17692_n1386), .Y(_abc_17692_n1393) );
  AND2X2 AND2X2_3110 ( .A(_abc_17692_n7803), .B(_abc_17692_n7792), .Y(_abc_17692_n7814) );
  AND2X2 AND2X2_3111 ( .A(_abc_17692_n7815), .B(_abc_17692_n7812), .Y(_abc_17692_n7816) );
  AND2X2 AND2X2_3112 ( .A(_abc_17692_n7667), .B(_abc_17692_n7649), .Y(_abc_17692_n7819) );
  AND2X2 AND2X2_3113 ( .A(_abc_17692_n7822), .B(_abc_17692_n1877_bF_buf8), .Y(_abc_17692_n7823) );
  AND2X2 AND2X2_3114 ( .A(_abc_17692_n7823), .B(_abc_17692_n7820), .Y(_abc_17692_n7824) );
  AND2X2 AND2X2_3115 ( .A(sum_29_), .B(\key_in[29] ), .Y(_abc_17692_n7827) );
  AND2X2 AND2X2_3116 ( .A(_abc_17692_n7828), .B(_abc_17692_n7829), .Y(_abc_17692_n7830) );
  AND2X2 AND2X2_3117 ( .A(_abc_17692_n7826), .B(_abc_17692_n7831), .Y(_abc_17692_n7832) );
  AND2X2 AND2X2_3118 ( .A(_abc_17692_n7825), .B(_abc_17692_n7830), .Y(_abc_17692_n7833) );
  AND2X2 AND2X2_3119 ( .A(_abc_17692_n7834), .B(_abc_17692_n7805), .Y(_abc_17692_n7835) );
  AND2X2 AND2X2_312 ( .A(_abc_17692_n722_bF_buf3), .B(sum_17_), .Y(_abc_17692_n1394) );
  AND2X2 AND2X2_3120 ( .A(_abc_17692_n7837), .B(_abc_17692_n7836), .Y(_abc_17692_n7838) );
  AND2X2 AND2X2_3121 ( .A(_abc_17692_n7838), .B(_abc_17692_n7792), .Y(_abc_17692_n7839) );
  AND2X2 AND2X2_3122 ( .A(_abc_17692_n7843), .B(_abc_17692_n7842), .Y(_abc_17692_n7844) );
  AND2X2 AND2X2_3123 ( .A(_abc_17692_n7841), .B(_abc_17692_n7845), .Y(_abc_17692_n7846) );
  AND2X2 AND2X2_3124 ( .A(_abc_17692_n7608), .B(workunit2_28_), .Y(_abc_17692_n7848) );
  AND2X2 AND2X2_3125 ( .A(_abc_17692_n7628), .B(_abc_17692_n7849), .Y(_abc_17692_n7850) );
  AND2X2 AND2X2_3126 ( .A(_abc_17692_n7853), .B(_abc_17692_n1830_bF_buf8), .Y(_abc_17692_n7854) );
  AND2X2 AND2X2_3127 ( .A(_abc_17692_n7854), .B(_abc_17692_n7852), .Y(_abc_17692_n7855) );
  AND2X2 AND2X2_3128 ( .A(sum_29_), .B(\key_in[61] ), .Y(_abc_17692_n7858) );
  AND2X2 AND2X2_3129 ( .A(_abc_17692_n7859), .B(_abc_17692_n7860), .Y(_abc_17692_n7861) );
  AND2X2 AND2X2_313 ( .A(delta_18_), .B(sum_18_), .Y(_abc_17692_n1398) );
  AND2X2 AND2X2_3130 ( .A(_abc_17692_n7857), .B(_abc_17692_n7862), .Y(_abc_17692_n7863) );
  AND2X2 AND2X2_3131 ( .A(_abc_17692_n7856), .B(_abc_17692_n7861), .Y(_abc_17692_n7864) );
  AND2X2 AND2X2_3132 ( .A(_abc_17692_n7865), .B(_abc_17692_n7805), .Y(_abc_17692_n7866) );
  AND2X2 AND2X2_3133 ( .A(_abc_17692_n7868), .B(_abc_17692_n7867), .Y(_abc_17692_n7869) );
  AND2X2 AND2X2_3134 ( .A(_abc_17692_n7869), .B(_abc_17692_n7792), .Y(_abc_17692_n7870) );
  AND2X2 AND2X2_3135 ( .A(_abc_17692_n7874), .B(_abc_17692_n7873), .Y(_abc_17692_n7875) );
  AND2X2 AND2X2_3136 ( .A(_abc_17692_n7872), .B(_abc_17692_n7876), .Y(_abc_17692_n7877) );
  AND2X2 AND2X2_3137 ( .A(_abc_17692_n7688), .B(workunit2_28_), .Y(_abc_17692_n7878) );
  AND2X2 AND2X2_3138 ( .A(_abc_17692_n7705), .B(_abc_17692_n7879), .Y(_abc_17692_n7880) );
  AND2X2 AND2X2_3139 ( .A(_abc_17692_n7884), .B(_abc_17692_n1846_bF_buf8), .Y(_abc_17692_n7885) );
  AND2X2 AND2X2_314 ( .A(_abc_17692_n1399), .B(_abc_17692_n1400), .Y(_abc_17692_n1401) );
  AND2X2 AND2X2_3140 ( .A(_abc_17692_n7885), .B(_abc_17692_n7881), .Y(_abc_17692_n7886) );
  AND2X2 AND2X2_3141 ( .A(sum_29_), .B(\key_in[125] ), .Y(_abc_17692_n7891) );
  AND2X2 AND2X2_3142 ( .A(_abc_17692_n7892), .B(_abc_17692_n7893), .Y(_abc_17692_n7894) );
  AND2X2 AND2X2_3143 ( .A(_abc_17692_n7890), .B(_abc_17692_n7894), .Y(_abc_17692_n7897) );
  AND2X2 AND2X2_3144 ( .A(_abc_17692_n7898), .B(_abc_17692_n7805), .Y(_abc_17692_n7899) );
  AND2X2 AND2X2_3145 ( .A(_abc_17692_n7900), .B(_abc_17692_n7895), .Y(_abc_17692_n7901) );
  AND2X2 AND2X2_3146 ( .A(_abc_17692_n7901), .B(_abc_17692_n7792), .Y(_abc_17692_n7902) );
  AND2X2 AND2X2_3147 ( .A(_abc_17692_n7906), .B(_abc_17692_n7905), .Y(_abc_17692_n7907) );
  AND2X2 AND2X2_3148 ( .A(_abc_17692_n7904), .B(_abc_17692_n7908), .Y(_abc_17692_n7909) );
  AND2X2 AND2X2_3149 ( .A(_abc_17692_n7588), .B(_abc_17692_n7569), .Y(_abc_17692_n7910) );
  AND2X2 AND2X2_315 ( .A(_abc_17692_n1331_1), .B(_abc_17692_n1375), .Y(_abc_17692_n1404) );
  AND2X2 AND2X2_3150 ( .A(_abc_17692_n7911), .B(_abc_17692_n7909), .Y(_abc_17692_n7912) );
  AND2X2 AND2X2_3151 ( .A(_abc_17692_n7907), .B(workunit2_29_), .Y(_abc_17692_n7913) );
  AND2X2 AND2X2_3152 ( .A(_abc_17692_n7903), .B(_abc_17692_n7812), .Y(_abc_17692_n7914) );
  AND2X2 AND2X2_3153 ( .A(_abc_17692_n7910), .B(_abc_17692_n7915), .Y(_abc_17692_n7916) );
  AND2X2 AND2X2_3154 ( .A(_abc_17692_n7918), .B(state_6_bF_buf0), .Y(_abc_17692_n7919) );
  AND2X2 AND2X2_3155 ( .A(_abc_17692_n7919), .B(_abc_17692_n7889), .Y(_abc_17692_n7920) );
  AND2X2 AND2X2_3156 ( .A(_abc_17692_n7921), .B(workunit2_28_), .Y(_abc_17692_n7922) );
  AND2X2 AND2X2_3157 ( .A(_abc_17692_n7923), .B(_abc_17692_n7817), .Y(_abc_17692_n7924) );
  AND2X2 AND2X2_3158 ( .A(_abc_17692_n7925), .B(_abc_17692_n7818), .Y(_abc_17692_n7926) );
  AND2X2 AND2X2_3159 ( .A(_abc_17692_n7927), .B(_abc_17692_n1877_bF_buf7), .Y(_abc_17692_n7928) );
  AND2X2 AND2X2_316 ( .A(_abc_17692_n1376), .B(_abc_17692_n1370), .Y(_abc_17692_n1407) );
  AND2X2 AND2X2_3160 ( .A(_abc_17692_n7934), .B(_abc_17692_n1863_bF_buf6), .Y(_abc_17692_n7935) );
  AND2X2 AND2X2_3161 ( .A(_abc_17692_n7935), .B(_abc_17692_n7933), .Y(_abc_17692_n7936) );
  AND2X2 AND2X2_3162 ( .A(_abc_17692_n7941), .B(_abc_17692_n1830_bF_buf7), .Y(_abc_17692_n7942) );
  AND2X2 AND2X2_3163 ( .A(_abc_17692_n7942), .B(_abc_17692_n7940), .Y(_abc_17692_n7943) );
  AND2X2 AND2X2_3164 ( .A(_abc_17692_n7948), .B(_abc_17692_n1846_bF_buf7), .Y(_abc_17692_n7949) );
  AND2X2 AND2X2_3165 ( .A(_abc_17692_n7949), .B(_abc_17692_n7947), .Y(_abc_17692_n7950) );
  AND2X2 AND2X2_3166 ( .A(_abc_17692_n7953), .B(state_7_bF_buf4), .Y(_abc_17692_n7954) );
  AND2X2 AND2X2_3167 ( .A(_abc_17692_n1885_bF_buf0), .B(workunit2_29_), .Y(_abc_17692_n7955) );
  AND2X2 AND2X2_3168 ( .A(state_8_bF_buf0), .B(\data_in2[29] ), .Y(_abc_17692_n7956) );
  AND2X2 AND2X2_3169 ( .A(_abc_17692_n7840), .B(workunit2_29_), .Y(_abc_17692_n7962) );
  AND2X2 AND2X2_317 ( .A(_abc_17692_n1406), .B(_abc_17692_n1408), .Y(_abc_17692_n1409) );
  AND2X2 AND2X2_3170 ( .A(_abc_17692_n7847), .B(_abc_17692_n7848), .Y(_abc_17692_n7963) );
  AND2X2 AND2X2_3171 ( .A(_abc_17692_n7961), .B(_abc_17692_n7965), .Y(_abc_17692_n7966) );
  AND2X2 AND2X2_3172 ( .A(workunit1_26_), .B(workunit1_30_), .Y(_abc_17692_n7969) );
  AND2X2 AND2X2_3173 ( .A(_abc_17692_n6065), .B(_abc_17692_n6956), .Y(_abc_17692_n7970) );
  AND2X2 AND2X2_3174 ( .A(_abc_17692_n7783), .B(_abc_17692_n7787), .Y(_abc_17692_n7973) );
  AND2X2 AND2X2_3175 ( .A(_abc_17692_n7974), .B(_abc_17692_n7972), .Y(_abc_17692_n7975) );
  AND2X2 AND2X2_3176 ( .A(_abc_17692_n7976), .B(_abc_17692_n7977), .Y(_abc_17692_n7978) );
  AND2X2 AND2X2_3177 ( .A(sum_30_), .B(\key_in[30] ), .Y(_abc_17692_n7979) );
  AND2X2 AND2X2_3178 ( .A(_abc_17692_n7980), .B(_abc_17692_n7981), .Y(_abc_17692_n7982) );
  AND2X2 AND2X2_3179 ( .A(_abc_17692_n7826), .B(_abc_17692_n7828), .Y(_abc_17692_n7985) );
  AND2X2 AND2X2_318 ( .A(_abc_17692_n1410), .B(_abc_17692_n1403_1), .Y(_abc_17692_n1412) );
  AND2X2 AND2X2_3180 ( .A(_abc_17692_n7986), .B(_abc_17692_n7983), .Y(_abc_17692_n7987) );
  AND2X2 AND2X2_3181 ( .A(_abc_17692_n7988), .B(_abc_17692_n7989), .Y(_abc_17692_n7990) );
  AND2X2 AND2X2_3182 ( .A(_abc_17692_n7990), .B(_abc_17692_n7978), .Y(_abc_17692_n7993) );
  AND2X2 AND2X2_3183 ( .A(_abc_17692_n7996), .B(_abc_17692_n7991), .Y(_abc_17692_n7997) );
  AND2X2 AND2X2_3184 ( .A(_abc_17692_n7995), .B(_abc_17692_n7998), .Y(_abc_17692_n7999) );
  AND2X2 AND2X2_3185 ( .A(_abc_17692_n8002), .B(_abc_17692_n1830_bF_buf6), .Y(_abc_17692_n8003) );
  AND2X2 AND2X2_3186 ( .A(_abc_17692_n8003), .B(_abc_17692_n8001), .Y(_abc_17692_n8004) );
  AND2X2 AND2X2_3187 ( .A(_abc_17692_n7817), .B(_abc_17692_n7651), .Y(_abc_17692_n8005) );
  AND2X2 AND2X2_3188 ( .A(_abc_17692_n7665), .B(_abc_17692_n8005), .Y(_abc_17692_n8006) );
  AND2X2 AND2X2_3189 ( .A(_abc_17692_n7815), .B(workunit2_29_), .Y(_abc_17692_n8007) );
  AND2X2 AND2X2_319 ( .A(_abc_17692_n1413), .B(state_3_bF_buf1), .Y(_abc_17692_n1414) );
  AND2X2 AND2X2_3190 ( .A(_abc_17692_n7817), .B(_abc_17692_n7648), .Y(_abc_17692_n8008) );
  AND2X2 AND2X2_3191 ( .A(sum_30_), .B(\key_in[94] ), .Y(_abc_17692_n8012) );
  AND2X2 AND2X2_3192 ( .A(_abc_17692_n8013), .B(_abc_17692_n8014), .Y(_abc_17692_n8015) );
  AND2X2 AND2X2_3193 ( .A(_abc_17692_n7794), .B(_abc_17692_n7796), .Y(_abc_17692_n8018) );
  AND2X2 AND2X2_3194 ( .A(_abc_17692_n8019), .B(_abc_17692_n8016), .Y(_abc_17692_n8020) );
  AND2X2 AND2X2_3195 ( .A(_abc_17692_n8021), .B(_abc_17692_n8022), .Y(_abc_17692_n8023) );
  AND2X2 AND2X2_3196 ( .A(_abc_17692_n8024), .B(_abc_17692_n8011), .Y(_abc_17692_n8025) );
  AND2X2 AND2X2_3197 ( .A(_abc_17692_n8023), .B(_abc_17692_n7978), .Y(_abc_17692_n8026) );
  AND2X2 AND2X2_3198 ( .A(_abc_17692_n8030), .B(_abc_17692_n8028), .Y(_abc_17692_n8031) );
  AND2X2 AND2X2_3199 ( .A(_abc_17692_n8010), .B(_abc_17692_n8031), .Y(_abc_17692_n8033) );
  AND2X2 AND2X2_32 ( .A(_abc_17692_n701), .B(_abc_17692_n702), .Y(_abc_17692_n703) );
  AND2X2 AND2X2_320 ( .A(_abc_17692_n1414), .B(_abc_17692_n1411), .Y(_abc_17692_n1415) );
  AND2X2 AND2X2_3200 ( .A(_abc_17692_n8034), .B(_abc_17692_n1877_bF_buf6), .Y(_abc_17692_n8035) );
  AND2X2 AND2X2_3201 ( .A(_abc_17692_n8035), .B(_abc_17692_n8032), .Y(_abc_17692_n8036) );
  AND2X2 AND2X2_3202 ( .A(_abc_17692_n7871), .B(workunit2_29_), .Y(_abc_17692_n8039) );
  AND2X2 AND2X2_3203 ( .A(_abc_17692_n8041), .B(_abc_17692_n8040), .Y(_abc_17692_n8042) );
  AND2X2 AND2X2_3204 ( .A(_abc_17692_n8038), .B(_abc_17692_n8042), .Y(_abc_17692_n8043) );
  AND2X2 AND2X2_3205 ( .A(sum_30_), .B(\key_in[62] ), .Y(_abc_17692_n8045) );
  AND2X2 AND2X2_3206 ( .A(_abc_17692_n8046), .B(_abc_17692_n8047), .Y(_abc_17692_n8048) );
  AND2X2 AND2X2_3207 ( .A(_abc_17692_n7857), .B(_abc_17692_n7859), .Y(_abc_17692_n8051) );
  AND2X2 AND2X2_3208 ( .A(_abc_17692_n8052), .B(_abc_17692_n8049), .Y(_abc_17692_n8053) );
  AND2X2 AND2X2_3209 ( .A(_abc_17692_n8054), .B(_abc_17692_n8055), .Y(_abc_17692_n8056) );
  AND2X2 AND2X2_321 ( .A(_abc_17692_n1371), .B(sum_17_), .Y(_abc_17692_n1416) );
  AND2X2 AND2X2_3210 ( .A(_abc_17692_n8059), .B(_abc_17692_n8057), .Y(_abc_17692_n8060) );
  AND2X2 AND2X2_3211 ( .A(_abc_17692_n8062), .B(_abc_17692_n8063), .Y(_abc_17692_n8064) );
  AND2X2 AND2X2_3212 ( .A(_abc_17692_n8061), .B(_abc_17692_n8065), .Y(_abc_17692_n8066) );
  AND2X2 AND2X2_3213 ( .A(_abc_17692_n8069), .B(_abc_17692_n1846_bF_buf6), .Y(_abc_17692_n8070) );
  AND2X2 AND2X2_3214 ( .A(_abc_17692_n8070), .B(_abc_17692_n8068), .Y(_abc_17692_n8071) );
  AND2X2 AND2X2_3215 ( .A(_abc_17692_n7915), .B(_abc_17692_n7572), .Y(_abc_17692_n8075) );
  AND2X2 AND2X2_3216 ( .A(_abc_17692_n7903), .B(workunit2_29_), .Y(_abc_17692_n8078) );
  AND2X2 AND2X2_3217 ( .A(_abc_17692_n8080), .B(_abc_17692_n8079), .Y(_abc_17692_n8081) );
  AND2X2 AND2X2_3218 ( .A(_abc_17692_n8077), .B(_abc_17692_n8081), .Y(_abc_17692_n8082) );
  AND2X2 AND2X2_3219 ( .A(sum_30_), .B(\key_in[126] ), .Y(_abc_17692_n8084) );
  AND2X2 AND2X2_322 ( .A(_abc_17692_n1390), .B(_abc_17692_n1417), .Y(_abc_17692_n1418) );
  AND2X2 AND2X2_3220 ( .A(_abc_17692_n8085), .B(_abc_17692_n8086), .Y(_abc_17692_n8087) );
  AND2X2 AND2X2_3221 ( .A(_abc_17692_n8089), .B(_abc_17692_n7893), .Y(_abc_17692_n8090) );
  AND2X2 AND2X2_3222 ( .A(_abc_17692_n8091), .B(_abc_17692_n8088), .Y(_abc_17692_n8092) );
  AND2X2 AND2X2_3223 ( .A(_abc_17692_n8090), .B(_abc_17692_n8087), .Y(_abc_17692_n8093) );
  AND2X2 AND2X2_3224 ( .A(_abc_17692_n8094), .B(_abc_17692_n8011), .Y(_abc_17692_n8095) );
  AND2X2 AND2X2_3225 ( .A(_abc_17692_n8096), .B(_abc_17692_n7978), .Y(_abc_17692_n8097) );
  AND2X2 AND2X2_3226 ( .A(_abc_17692_n8100), .B(_abc_17692_n8101), .Y(_abc_17692_n8102) );
  AND2X2 AND2X2_3227 ( .A(_abc_17692_n8105), .B(_abc_17692_n8104), .Y(_abc_17692_n8106) );
  AND2X2 AND2X2_3228 ( .A(_abc_17692_n8103), .B(_abc_17692_n8107), .Y(_abc_17692_n8108) );
  AND2X2 AND2X2_3229 ( .A(_abc_17692_n8109), .B(state_6_bF_buf4), .Y(_abc_17692_n8110) );
  AND2X2 AND2X2_323 ( .A(_abc_17692_n1388), .B(_abc_17692_n1418), .Y(_abc_17692_n1419) );
  AND2X2 AND2X2_3230 ( .A(_abc_17692_n8110), .B(_abc_17692_n8074), .Y(_abc_17692_n8111) );
  AND2X2 AND2X2_3231 ( .A(_abc_17692_n7909), .B(_abc_17692_n7587), .Y(_abc_17692_n8112) );
  AND2X2 AND2X2_3232 ( .A(_abc_17692_n7721), .B(_abc_17692_n8112), .Y(_abc_17692_n8113) );
  AND2X2 AND2X2_3233 ( .A(_abc_17692_n7904), .B(_abc_17692_n7929), .Y(_abc_17692_n8114) );
  AND2X2 AND2X2_3234 ( .A(_abc_17692_n8120), .B(_abc_17692_n6881), .Y(_abc_17692_n8121) );
  AND2X2 AND2X2_3235 ( .A(_abc_17692_n8119), .B(_abc_17692_n8121), .Y(_abc_17692_n8122) );
  AND2X2 AND2X2_3236 ( .A(_abc_17692_n8122), .B(_abc_17692_n8129), .Y(_abc_17692_n8130) );
  AND2X2 AND2X2_3237 ( .A(_abc_17692_n8135), .B(_abc_17692_n8136), .Y(_abc_17692_n8137) );
  AND2X2 AND2X2_3238 ( .A(_abc_17692_n8134), .B(_abc_17692_n8137), .Y(_abc_17692_n8138) );
  AND2X2 AND2X2_3239 ( .A(_abc_17692_n8140), .B(_abc_17692_n8115), .Y(_abc_17692_n8141) );
  AND2X2 AND2X2_324 ( .A(_abc_17692_n1420), .B(_abc_17692_n1402), .Y(_abc_17692_n1421_1) );
  AND2X2 AND2X2_3240 ( .A(_abc_17692_n8142), .B(_abc_17692_n1863_bF_buf4), .Y(_abc_17692_n8143) );
  AND2X2 AND2X2_3241 ( .A(_abc_17692_n8143), .B(_abc_17692_n8118), .Y(_abc_17692_n8144) );
  AND2X2 AND2X2_3242 ( .A(_abc_17692_n8149), .B(_abc_17692_n8148), .Y(_abc_17692_n8150) );
  AND2X2 AND2X2_3243 ( .A(_abc_17692_n8147), .B(_abc_17692_n8151), .Y(_abc_17692_n8152) );
  AND2X2 AND2X2_3244 ( .A(_abc_17692_n8155), .B(_abc_17692_n1877_bF_buf5), .Y(_abc_17692_n8156) );
  AND2X2 AND2X2_3245 ( .A(_abc_17692_n8156), .B(_abc_17692_n8154), .Y(_abc_17692_n8157) );
  AND2X2 AND2X2_3246 ( .A(_abc_17692_n7877), .B(_abc_17692_n7691), .Y(_abc_17692_n8158) );
  AND2X2 AND2X2_3247 ( .A(_abc_17692_n7753), .B(_abc_17692_n8158), .Y(_abc_17692_n8159) );
  AND2X2 AND2X2_3248 ( .A(_abc_17692_n7876), .B(_abc_17692_n7944), .Y(_abc_17692_n8161) );
  AND2X2 AND2X2_3249 ( .A(_abc_17692_n8163), .B(_abc_17692_n8066), .Y(_abc_17692_n8164) );
  AND2X2 AND2X2_325 ( .A(_abc_17692_n1423), .B(state_15_bF_buf1), .Y(_abc_17692_n1424) );
  AND2X2 AND2X2_3250 ( .A(_abc_17692_n8166), .B(_abc_17692_n1846_bF_buf5), .Y(_abc_17692_n8167) );
  AND2X2 AND2X2_3251 ( .A(_abc_17692_n8167), .B(_abc_17692_n8165), .Y(_abc_17692_n8168) );
  AND2X2 AND2X2_3252 ( .A(_abc_17692_n7846), .B(_abc_17692_n7611), .Y(_abc_17692_n8169) );
  AND2X2 AND2X2_3253 ( .A(_abc_17692_n7768), .B(_abc_17692_n8169), .Y(_abc_17692_n8170) );
  AND2X2 AND2X2_3254 ( .A(_abc_17692_n7845), .B(_abc_17692_n7937), .Y(_abc_17692_n8172) );
  AND2X2 AND2X2_3255 ( .A(_abc_17692_n8174), .B(_abc_17692_n7999), .Y(_abc_17692_n8175) );
  AND2X2 AND2X2_3256 ( .A(_abc_17692_n8177), .B(_abc_17692_n1830_bF_buf5), .Y(_abc_17692_n8178) );
  AND2X2 AND2X2_3257 ( .A(_abc_17692_n8178), .B(_abc_17692_n8176), .Y(_abc_17692_n8179) );
  AND2X2 AND2X2_3258 ( .A(_abc_17692_n8182), .B(state_7_bF_buf3), .Y(_abc_17692_n8183) );
  AND2X2 AND2X2_3259 ( .A(_abc_17692_n1885_bF_buf4), .B(workunit2_30_), .Y(_abc_17692_n8184) );
  AND2X2 AND2X2_326 ( .A(_abc_17692_n1424), .B(_abc_17692_n1422), .Y(_abc_17692_n1425) );
  AND2X2 AND2X2_3260 ( .A(state_8_bF_buf9), .B(\data_in2[30] ), .Y(_abc_17692_n8185) );
  AND2X2 AND2X2_3261 ( .A(_abc_17692_n8107), .B(_abc_17692_n8100), .Y(_abc_17692_n8189) );
  AND2X2 AND2X2_3262 ( .A(_abc_17692_n8191), .B(_abc_17692_n8085), .Y(_abc_17692_n8192) );
  AND2X2 AND2X2_3263 ( .A(_abc_17692_n8193), .B(_abc_17692_n8195), .Y(_abc_17692_n8196) );
  AND2X2 AND2X2_3264 ( .A(_abc_17692_n8192), .B(_abc_17692_n8197), .Y(_abc_17692_n8198) );
  AND2X2 AND2X2_3265 ( .A(_abc_17692_n8199), .B(_abc_17692_n8200), .Y(_abc_17692_n8201) );
  AND2X2 AND2X2_3266 ( .A(workunit1_27_), .B(workunit1_31_), .Y(_abc_17692_n8205) );
  AND2X2 AND2X2_3267 ( .A(_abc_17692_n6242), .B(_abc_17692_n7135), .Y(_abc_17692_n8206) );
  AND2X2 AND2X2_3268 ( .A(_abc_17692_n8204), .B(_abc_17692_n8207), .Y(_abc_17692_n8208) );
  AND2X2 AND2X2_3269 ( .A(_abc_17692_n8209), .B(_abc_17692_n8210), .Y(_abc_17692_n8211) );
  AND2X2 AND2X2_327 ( .A(_abc_17692_n722_bF_buf2), .B(sum_18_), .Y(_abc_17692_n1426) );
  AND2X2 AND2X2_3270 ( .A(_abc_17692_n8211), .B(_abc_17692_n8202), .Y(_abc_17692_n8212) );
  AND2X2 AND2X2_3271 ( .A(_abc_17692_n8219), .B(_abc_17692_n8216), .Y(_abc_17692_n8220) );
  AND2X2 AND2X2_3272 ( .A(_abc_17692_n8190), .B(_abc_17692_n8221), .Y(_abc_17692_n8222) );
  AND2X2 AND2X2_3273 ( .A(_abc_17692_n8189), .B(_abc_17692_n8220), .Y(_abc_17692_n8223) );
  AND2X2 AND2X2_3274 ( .A(_abc_17692_n8022), .B(_abc_17692_n8013), .Y(_abc_17692_n8229) );
  AND2X2 AND2X2_3275 ( .A(_abc_17692_n8230), .B(_abc_17692_n8232), .Y(_abc_17692_n8233) );
  AND2X2 AND2X2_3276 ( .A(_abc_17692_n8229), .B(_abc_17692_n8234), .Y(_abc_17692_n8235) );
  AND2X2 AND2X2_3277 ( .A(_abc_17692_n8236), .B(_abc_17692_n8237), .Y(_abc_17692_n8238) );
  AND2X2 AND2X2_3278 ( .A(_abc_17692_n8241), .B(_abc_17692_n8239), .Y(_abc_17692_n8242) );
  AND2X2 AND2X2_3279 ( .A(_abc_17692_n8245), .B(_abc_17692_n1877_bF_buf4), .Y(_abc_17692_n8246) );
  AND2X2 AND2X2_328 ( .A(delta_19_), .B(sum_19_), .Y(_abc_17692_n1430) );
  AND2X2 AND2X2_3280 ( .A(_abc_17692_n8246), .B(_abc_17692_n8244), .Y(_abc_17692_n8247) );
  AND2X2 AND2X2_3281 ( .A(_abc_17692_n7994), .B(workunit2_30_), .Y(_abc_17692_n8248) );
  AND2X2 AND2X2_3282 ( .A(_abc_17692_n8002), .B(_abc_17692_n8249), .Y(_abc_17692_n8250) );
  AND2X2 AND2X2_3283 ( .A(_abc_17692_n7989), .B(_abc_17692_n7980), .Y(_abc_17692_n8252) );
  AND2X2 AND2X2_3284 ( .A(_abc_17692_n8253), .B(_abc_17692_n8255), .Y(_abc_17692_n8256) );
  AND2X2 AND2X2_3285 ( .A(_abc_17692_n8252), .B(_abc_17692_n8257), .Y(_abc_17692_n8258) );
  AND2X2 AND2X2_3286 ( .A(_abc_17692_n8259), .B(_abc_17692_n8260), .Y(_abc_17692_n8261) );
  AND2X2 AND2X2_3287 ( .A(_abc_17692_n8262), .B(_abc_17692_n8264), .Y(_abc_17692_n8265) );
  AND2X2 AND2X2_3288 ( .A(_abc_17692_n8268), .B(_abc_17692_n1830_bF_buf4), .Y(_abc_17692_n8269) );
  AND2X2 AND2X2_3289 ( .A(_abc_17692_n8269), .B(_abc_17692_n8267), .Y(_abc_17692_n8270) );
  AND2X2 AND2X2_329 ( .A(_abc_17692_n1432), .B(_abc_17692_n1433), .Y(_abc_17692_n1434) );
  AND2X2 AND2X2_3290 ( .A(_abc_17692_n8060), .B(workunit2_30_), .Y(_abc_17692_n8271) );
  AND2X2 AND2X2_3291 ( .A(_abc_17692_n8069), .B(_abc_17692_n8272), .Y(_abc_17692_n8273) );
  AND2X2 AND2X2_3292 ( .A(_abc_17692_n8055), .B(_abc_17692_n8046), .Y(_abc_17692_n8275) );
  AND2X2 AND2X2_3293 ( .A(_abc_17692_n8276), .B(_abc_17692_n8278), .Y(_abc_17692_n8279) );
  AND2X2 AND2X2_3294 ( .A(_abc_17692_n8275), .B(_abc_17692_n8280), .Y(_abc_17692_n8281) );
  AND2X2 AND2X2_3295 ( .A(_abc_17692_n8282), .B(_abc_17692_n8283), .Y(_abc_17692_n8284) );
  AND2X2 AND2X2_3296 ( .A(_abc_17692_n8285), .B(_abc_17692_n8287), .Y(_abc_17692_n8288) );
  AND2X2 AND2X2_3297 ( .A(_abc_17692_n8291), .B(_abc_17692_n1846_bF_buf4), .Y(_abc_17692_n8292) );
  AND2X2 AND2X2_3298 ( .A(_abc_17692_n8292), .B(_abc_17692_n8290), .Y(_abc_17692_n8293) );
  AND2X2 AND2X2_3299 ( .A(_abc_17692_n8296), .B(state_6_bF_buf3), .Y(_abc_17692_n8297) );
  AND2X2 AND2X2_33 ( .A(_abc_17692_n703), .B(_abc_17692_n700), .Y(_abc_17692_n704) );
  AND2X2 AND2X2_330 ( .A(_abc_17692_n1435), .B(_abc_17692_n1431), .Y(_abc_17692_n1436) );
  AND2X2 AND2X2_3300 ( .A(_abc_17692_n8297), .B(_abc_17692_n8225), .Y(_abc_17692_n8298) );
  AND2X2 AND2X2_3301 ( .A(_abc_17692_n8142), .B(_abc_17692_n8104), .Y(_abc_17692_n8299) );
  AND2X2 AND2X2_3302 ( .A(_abc_17692_n8299), .B(_abc_17692_n8221), .Y(_abc_17692_n8300) );
  AND2X2 AND2X2_3303 ( .A(_abc_17692_n8117), .B(_abc_17692_n8106), .Y(_abc_17692_n8302) );
  AND2X2 AND2X2_3304 ( .A(_abc_17692_n8303), .B(_abc_17692_n8220), .Y(_abc_17692_n8304) );
  AND2X2 AND2X2_3305 ( .A(_abc_17692_n8305), .B(_abc_17692_n1863_bF_buf2), .Y(_abc_17692_n8306) );
  AND2X2 AND2X2_3306 ( .A(_abc_17692_n8029), .B(workunit2_30_), .Y(_abc_17692_n8307) );
  AND2X2 AND2X2_3307 ( .A(_abc_17692_n8155), .B(_abc_17692_n8308), .Y(_abc_17692_n8309) );
  AND2X2 AND2X2_3308 ( .A(_abc_17692_n8312), .B(_abc_17692_n1877_bF_buf3), .Y(_abc_17692_n8313) );
  AND2X2 AND2X2_3309 ( .A(_abc_17692_n8313), .B(_abc_17692_n8311), .Y(_abc_17692_n8314) );
  AND2X2 AND2X2_331 ( .A(_abc_17692_n1441_1), .B(state_3_bF_buf0), .Y(_abc_17692_n1442) );
  AND2X2 AND2X2_3310 ( .A(_abc_17692_n8319), .B(_abc_17692_n1846_bF_buf3), .Y(_abc_17692_n8320) );
  AND2X2 AND2X2_3311 ( .A(_abc_17692_n8320), .B(_abc_17692_n8318), .Y(_abc_17692_n8321) );
  AND2X2 AND2X2_3312 ( .A(_abc_17692_n8326), .B(_abc_17692_n1830_bF_buf3), .Y(_abc_17692_n8327) );
  AND2X2 AND2X2_3313 ( .A(_abc_17692_n8327), .B(_abc_17692_n8325), .Y(_abc_17692_n8328) );
  AND2X2 AND2X2_3314 ( .A(_abc_17692_n8331), .B(state_7_bF_buf2), .Y(_abc_17692_n8332) );
  AND2X2 AND2X2_3315 ( .A(_abc_17692_n1885_bF_buf3), .B(workunit2_31_), .Y(_abc_17692_n8333) );
  AND2X2 AND2X2_3316 ( .A(state_8_bF_buf8), .B(\data_in2[31] ), .Y(_abc_17692_n8334) );
  AND2X2 AND2X2_3317 ( .A(workunit2_0_), .B(workunit2_5_), .Y(_abc_17692_n8339) );
  AND2X2 AND2X2_3318 ( .A(_abc_17692_n1814), .B(_abc_17692_n2633), .Y(_abc_17692_n8340) );
  AND2X2 AND2X2_3319 ( .A(_abc_17692_n1824), .B(_abc_17692_n8341), .Y(_abc_17692_n8342) );
  AND2X2 AND2X2_332 ( .A(_abc_17692_n1442), .B(_abc_17692_n1440), .Y(_abc_17692_n1443) );
  AND2X2 AND2X2_3320 ( .A(_abc_17692_n8343), .B(_abc_17692_n1823), .Y(_abc_17692_n8344) );
  AND2X2 AND2X2_3321 ( .A(_abc_17692_n8346), .B(workunit1_0_), .Y(_abc_17692_n8347) );
  AND2X2 AND2X2_3322 ( .A(_abc_17692_n8349), .B(_abc_17692_n1830_bF_buf2), .Y(_abc_17692_n8350) );
  AND2X2 AND2X2_3323 ( .A(_abc_17692_n8350), .B(_abc_17692_n8348), .Y(_abc_17692_n8351) );
  AND2X2 AND2X2_3324 ( .A(_abc_17692_n1839), .B(_abc_17692_n8341), .Y(_abc_17692_n8352) );
  AND2X2 AND2X2_3325 ( .A(_abc_17692_n8343), .B(_abc_17692_n1838), .Y(_abc_17692_n8353) );
  AND2X2 AND2X2_3326 ( .A(_abc_17692_n8355), .B(workunit1_0_), .Y(_abc_17692_n8357) );
  AND2X2 AND2X2_3327 ( .A(_abc_17692_n8358), .B(_abc_17692_n1846_bF_buf2), .Y(_abc_17692_n8359) );
  AND2X2 AND2X2_3328 ( .A(_abc_17692_n8359), .B(_abc_17692_n8356), .Y(_abc_17692_n8360) );
  AND2X2 AND2X2_3329 ( .A(_abc_17692_n1855_1), .B(_abc_17692_n8341), .Y(_abc_17692_n8362) );
  AND2X2 AND2X2_333 ( .A(_abc_17692_n1399), .B(sum_18_), .Y(_abc_17692_n1444) );
  AND2X2 AND2X2_3330 ( .A(_abc_17692_n8343), .B(_abc_17692_n1854), .Y(_abc_17692_n8363) );
  AND2X2 AND2X2_3331 ( .A(_abc_17692_n8365), .B(workunit1_0_), .Y(_abc_17692_n8366) );
  AND2X2 AND2X2_3332 ( .A(_abc_17692_n8368), .B(_abc_17692_n1863_bF_buf1), .Y(_abc_17692_n8369) );
  AND2X2 AND2X2_3333 ( .A(_abc_17692_n8369), .B(_abc_17692_n8367), .Y(_abc_17692_n8370) );
  AND2X2 AND2X2_3334 ( .A(_abc_17692_n1871), .B(_abc_17692_n8341), .Y(_abc_17692_n8371) );
  AND2X2 AND2X2_3335 ( .A(_abc_17692_n8343), .B(_abc_17692_n1870), .Y(_abc_17692_n8372) );
  AND2X2 AND2X2_3336 ( .A(_abc_17692_n8374), .B(workunit1_0_), .Y(_abc_17692_n8376) );
  AND2X2 AND2X2_3337 ( .A(_abc_17692_n8377), .B(_abc_17692_n1877_bF_buf2), .Y(_abc_17692_n8378) );
  AND2X2 AND2X2_3338 ( .A(_abc_17692_n8378), .B(_abc_17692_n8375), .Y(_abc_17692_n8379) );
  AND2X2 AND2X2_3339 ( .A(_abc_17692_n8381), .B(_abc_17692_n8338), .Y(_abc_17692_n8382) );
  AND2X2 AND2X2_334 ( .A(_abc_17692_n1422), .B(_abc_17692_n1445), .Y(_abc_17692_n1446) );
  AND2X2 AND2X2_3340 ( .A(_abc_17692_n713), .B(_abc_17692_n632), .Y(_abc_17692_n8383) );
  AND2X2 AND2X2_3341 ( .A(_abc_17692_n8383_bF_buf4), .B(workunit1_0_), .Y(_abc_17692_n8384) );
  AND2X2 AND2X2_3342 ( .A(state_8_bF_buf7), .B(\data_in1[0] ), .Y(_abc_17692_n8385) );
  AND2X2 AND2X2_3343 ( .A(_abc_17692_n8346), .B(_abc_17692_n1816), .Y(_abc_17692_n8388) );
  AND2X2 AND2X2_3344 ( .A(workunit2_1_bF_buf0), .B(workunit2_6_), .Y(_abc_17692_n8390) );
  AND2X2 AND2X2_3345 ( .A(_abc_17692_n8391), .B(_abc_17692_n8392), .Y(_abc_17692_n8393) );
  AND2X2 AND2X2_3346 ( .A(_abc_17692_n8393), .B(_abc_17692_n8339), .Y(_abc_17692_n8394) );
  AND2X2 AND2X2_3347 ( .A(_abc_17692_n1919_1), .B(_abc_17692_n2862), .Y(_abc_17692_n8396) );
  AND2X2 AND2X2_3348 ( .A(_abc_17692_n8397), .B(_abc_17692_n8395), .Y(_abc_17692_n8398) );
  AND2X2 AND2X2_3349 ( .A(_abc_17692_n1946), .B(_abc_17692_n8399), .Y(_abc_17692_n8400) );
  AND2X2 AND2X2_335 ( .A(_abc_17692_n1449), .B(state_15_bF_buf0), .Y(_abc_17692_n1450) );
  AND2X2 AND2X2_3350 ( .A(_abc_17692_n8401), .B(_abc_17692_n8402), .Y(_abc_17692_n8403) );
  AND2X2 AND2X2_3351 ( .A(_abc_17692_n1942), .B(_abc_17692_n8403), .Y(_abc_17692_n8404) );
  AND2X2 AND2X2_3352 ( .A(_abc_17692_n8405), .B(workunit1_1_bF_buf1), .Y(_abc_17692_n8406) );
  AND2X2 AND2X2_3353 ( .A(_abc_17692_n8407), .B(_abc_17692_n8408), .Y(_abc_17692_n8409) );
  AND2X2 AND2X2_3354 ( .A(_abc_17692_n8410), .B(_abc_17692_n8389), .Y(_abc_17692_n8411) );
  AND2X2 AND2X2_3355 ( .A(_abc_17692_n8413), .B(_abc_17692_n1830_bF_buf1), .Y(_abc_17692_n8414) );
  AND2X2 AND2X2_3356 ( .A(_abc_17692_n8414), .B(_abc_17692_n8412), .Y(_abc_17692_n8415) );
  AND2X2 AND2X2_3357 ( .A(_abc_17692_n8416), .B(_abc_17692_n8417), .Y(_abc_17692_n8418) );
  AND2X2 AND2X2_3358 ( .A(_abc_17692_n8418), .B(workunit1_1_bF_buf3), .Y(_abc_17692_n8419) );
  AND2X2 AND2X2_3359 ( .A(_abc_17692_n8420), .B(_abc_17692_n8421), .Y(_abc_17692_n8422) );
  AND2X2 AND2X2_336 ( .A(_abc_17692_n1450), .B(_abc_17692_n1448), .Y(_abc_17692_n1451) );
  AND2X2 AND2X2_3360 ( .A(_abc_17692_n8422), .B(_abc_17692_n2637), .Y(_abc_17692_n8423) );
  AND2X2 AND2X2_3361 ( .A(_abc_17692_n8374), .B(_abc_17692_n1816), .Y(_abc_17692_n8425) );
  AND2X2 AND2X2_3362 ( .A(_abc_17692_n8424), .B(_abc_17692_n8426), .Y(_abc_17692_n8428) );
  AND2X2 AND2X2_3363 ( .A(_abc_17692_n8429), .B(_abc_17692_n1877_bF_buf1), .Y(_abc_17692_n8430) );
  AND2X2 AND2X2_3364 ( .A(_abc_17692_n8430), .B(_abc_17692_n8427), .Y(_abc_17692_n8431) );
  AND2X2 AND2X2_3365 ( .A(_abc_17692_n8355), .B(_abc_17692_n1816), .Y(_abc_17692_n8432) );
  AND2X2 AND2X2_3366 ( .A(_abc_17692_n1978), .B(_abc_17692_n8399), .Y(_abc_17692_n8434) );
  AND2X2 AND2X2_3367 ( .A(_abc_17692_n1974_1), .B(_abc_17692_n8403), .Y(_abc_17692_n8435) );
  AND2X2 AND2X2_3368 ( .A(_abc_17692_n8436), .B(workunit1_1_bF_buf2), .Y(_abc_17692_n8437) );
  AND2X2 AND2X2_3369 ( .A(_abc_17692_n8438), .B(_abc_17692_n8439), .Y(_abc_17692_n8440) );
  AND2X2 AND2X2_337 ( .A(_abc_17692_n722_bF_buf1), .B(sum_19_), .Y(_abc_17692_n1452) );
  AND2X2 AND2X2_3370 ( .A(_abc_17692_n8443), .B(_abc_17692_n1846_bF_buf1), .Y(_abc_17692_n8444) );
  AND2X2 AND2X2_3371 ( .A(_abc_17692_n8444), .B(_abc_17692_n8442), .Y(_abc_17692_n8445) );
  AND2X2 AND2X2_3372 ( .A(_abc_17692_n8365), .B(_abc_17692_n1816), .Y(_abc_17692_n8448) );
  AND2X2 AND2X2_3373 ( .A(_abc_17692_n2007), .B(_abc_17692_n8403), .Y(_abc_17692_n8451) );
  AND2X2 AND2X2_3374 ( .A(_abc_17692_n8452), .B(_abc_17692_n8450), .Y(_abc_17692_n8453) );
  AND2X2 AND2X2_3375 ( .A(_abc_17692_n2002), .B(_abc_17692_n8399), .Y(_abc_17692_n8455) );
  AND2X2 AND2X2_3376 ( .A(_abc_17692_n8454), .B(_abc_17692_n8457), .Y(_abc_17692_n8458) );
  AND2X2 AND2X2_3377 ( .A(_abc_17692_n8459), .B(_abc_17692_n8449), .Y(_abc_17692_n8460) );
  AND2X2 AND2X2_3378 ( .A(_abc_17692_n8462), .B(_abc_17692_n1863_bF_buf0), .Y(_abc_17692_n8463) );
  AND2X2 AND2X2_3379 ( .A(_abc_17692_n8463), .B(_abc_17692_n8461), .Y(_abc_17692_n8464) );
  AND2X2 AND2X2_338 ( .A(_abc_17692_n1456), .B(delta_20_), .Y(_abc_17692_n1457) );
  AND2X2 AND2X2_3380 ( .A(_abc_17692_n8465), .B(state_10_bF_buf3), .Y(_abc_17692_n8466) );
  AND2X2 AND2X2_3381 ( .A(_abc_17692_n8469), .B(_abc_17692_n1877_bF_buf0), .Y(_abc_17692_n8470) );
  AND2X2 AND2X2_3382 ( .A(_abc_17692_n8470), .B(_abc_17692_n8468), .Y(_abc_17692_n8471) );
  AND2X2 AND2X2_3383 ( .A(_abc_17692_n8409), .B(_abc_17692_n8347), .Y(_abc_17692_n8472) );
  AND2X2 AND2X2_3384 ( .A(_abc_17692_n8474), .B(_abc_17692_n1830_bF_buf0), .Y(_abc_17692_n8475) );
  AND2X2 AND2X2_3385 ( .A(_abc_17692_n8475), .B(_abc_17692_n8473), .Y(_abc_17692_n8476) );
  AND2X2 AND2X2_3386 ( .A(_abc_17692_n8458), .B(_abc_17692_n8366), .Y(_abc_17692_n8478) );
  AND2X2 AND2X2_3387 ( .A(_abc_17692_n8480), .B(_abc_17692_n1863_bF_buf10), .Y(_abc_17692_n8481) );
  AND2X2 AND2X2_3388 ( .A(_abc_17692_n8481), .B(_abc_17692_n8479), .Y(_abc_17692_n8482) );
  AND2X2 AND2X2_3389 ( .A(_abc_17692_n8440), .B(_abc_17692_n8357), .Y(_abc_17692_n8483) );
  AND2X2 AND2X2_339 ( .A(_abc_17692_n1403_1), .B(_abc_17692_n1436), .Y(_abc_17692_n1461) );
  AND2X2 AND2X2_3390 ( .A(_abc_17692_n8485), .B(_abc_17692_n1846_bF_buf0), .Y(_abc_17692_n8486) );
  AND2X2 AND2X2_3391 ( .A(_abc_17692_n8486), .B(_abc_17692_n8484), .Y(_abc_17692_n8487) );
  AND2X2 AND2X2_3392 ( .A(_abc_17692_n8489), .B(state_14_bF_buf3), .Y(_abc_17692_n8490) );
  AND2X2 AND2X2_3393 ( .A(_abc_17692_n8383_bF_buf3), .B(workunit1_1_bF_buf3), .Y(_abc_17692_n8491) );
  AND2X2 AND2X2_3394 ( .A(state_8_bF_buf6), .B(\data_in1[1] ), .Y(_abc_17692_n8492) );
  AND2X2 AND2X2_3395 ( .A(_abc_17692_n8401), .B(_abc_17692_n8391), .Y(_abc_17692_n8496) );
  AND2X2 AND2X2_3396 ( .A(workunit2_2_), .B(workunit2_7_), .Y(_abc_17692_n8497) );
  AND2X2 AND2X2_3397 ( .A(_abc_17692_n2091), .B(_abc_17692_n3060), .Y(_abc_17692_n8498) );
  AND2X2 AND2X2_3398 ( .A(_abc_17692_n8500), .B(_abc_17692_n8503), .Y(_abc_17692_n8504) );
  AND2X2 AND2X2_3399 ( .A(_abc_17692_n8501), .B(_abc_17692_n8502), .Y(_abc_17692_n8506) );
  AND2X2 AND2X2_34 ( .A(_abc_17692_n705), .B(_abc_17692_n706), .Y(while_flag_FF_INPUT) );
  AND2X2 AND2X2_340 ( .A(_abc_17692_n1435), .B(_abc_17692_n1398), .Y(_abc_17692_n1464) );
  AND2X2 AND2X2_3400 ( .A(_abc_17692_n8496), .B(_abc_17692_n8499), .Y(_abc_17692_n8507) );
  AND2X2 AND2X2_3401 ( .A(_abc_17692_n8505), .B(_abc_17692_n8509), .Y(_abc_17692_n8510) );
  AND2X2 AND2X2_3402 ( .A(_abc_17692_n8512), .B(_abc_17692_n8513), .Y(_abc_17692_n8514) );
  AND2X2 AND2X2_3403 ( .A(_abc_17692_n8511), .B(_abc_17692_n8515), .Y(_abc_17692_n8516) );
  AND2X2 AND2X2_3404 ( .A(_abc_17692_n8422), .B(workunit1_1_bF_buf2), .Y(_abc_17692_n8517) );
  AND2X2 AND2X2_3405 ( .A(_abc_17692_n8518), .B(_abc_17692_n8516), .Y(_abc_17692_n8519) );
  AND2X2 AND2X2_3406 ( .A(_abc_17692_n8521), .B(_abc_17692_n1877_bF_buf10), .Y(_abc_17692_n8522) );
  AND2X2 AND2X2_3407 ( .A(_abc_17692_n8522), .B(_abc_17692_n8520), .Y(_abc_17692_n8523) );
  AND2X2 AND2X2_3408 ( .A(_abc_17692_n2117), .B(_abc_17692_n8508), .Y(_abc_17692_n8524) );
  AND2X2 AND2X2_3409 ( .A(_abc_17692_n2113), .B(_abc_17692_n8504), .Y(_abc_17692_n8526) );
  AND2X2 AND2X2_341 ( .A(_abc_17692_n1463), .B(_abc_17692_n1466), .Y(_abc_17692_n1467) );
  AND2X2 AND2X2_3410 ( .A(_abc_17692_n8525), .B(_abc_17692_n8527), .Y(_abc_17692_n8528) );
  AND2X2 AND2X2_3411 ( .A(_abc_17692_n8529), .B(_abc_17692_n8531), .Y(_abc_17692_n8532) );
  AND2X2 AND2X2_3412 ( .A(_abc_17692_n8534), .B(_abc_17692_n8535), .Y(_abc_17692_n8536) );
  AND2X2 AND2X2_3413 ( .A(_abc_17692_n8536), .B(workunit1_1_bF_buf1), .Y(_abc_17692_n8537) );
  AND2X2 AND2X2_3414 ( .A(_abc_17692_n8443), .B(_abc_17692_n8538), .Y(_abc_17692_n8539) );
  AND2X2 AND2X2_3415 ( .A(_abc_17692_n8542), .B(_abc_17692_n1846_bF_buf10), .Y(_abc_17692_n8543) );
  AND2X2 AND2X2_3416 ( .A(_abc_17692_n8543), .B(_abc_17692_n8541), .Y(_abc_17692_n8544) );
  AND2X2 AND2X2_3417 ( .A(_abc_17692_n2141), .B(_abc_17692_n8508), .Y(_abc_17692_n8545) );
  AND2X2 AND2X2_3418 ( .A(_abc_17692_n2146), .B(_abc_17692_n8504), .Y(_abc_17692_n8546) );
  AND2X2 AND2X2_3419 ( .A(_abc_17692_n8547), .B(workunit1_2_), .Y(_abc_17692_n8548) );
  AND2X2 AND2X2_342 ( .A(_abc_17692_n1468), .B(_abc_17692_n1467), .Y(_abc_17692_n1469) );
  AND2X2 AND2X2_3420 ( .A(_abc_17692_n8549), .B(_abc_17692_n8550), .Y(_abc_17692_n8551) );
  AND2X2 AND2X2_3421 ( .A(_abc_17692_n8553), .B(workunit1_1_bF_buf0), .Y(_abc_17692_n8554) );
  AND2X2 AND2X2_3422 ( .A(_abc_17692_n8552), .B(_abc_17692_n8555), .Y(_abc_17692_n8556) );
  AND2X2 AND2X2_3423 ( .A(_abc_17692_n8558), .B(_abc_17692_n1830_bF_buf10), .Y(_abc_17692_n8559) );
  AND2X2 AND2X2_3424 ( .A(_abc_17692_n8559), .B(_abc_17692_n8557), .Y(_abc_17692_n8560) );
  AND2X2 AND2X2_3425 ( .A(_abc_17692_n8563), .B(_abc_17692_n8564), .Y(_abc_17692_n8565) );
  AND2X2 AND2X2_3426 ( .A(_abc_17692_n8567), .B(_abc_17692_n8568), .Y(_abc_17692_n8569) );
  AND2X2 AND2X2_3427 ( .A(_abc_17692_n8566), .B(_abc_17692_n8570), .Y(_abc_17692_n8571) );
  AND2X2 AND2X2_3428 ( .A(_abc_17692_n8453), .B(workunit1_1_bF_buf3), .Y(_abc_17692_n8573) );
  AND2X2 AND2X2_3429 ( .A(_abc_17692_n8574), .B(_abc_17692_n8572), .Y(_abc_17692_n8575) );
  AND2X2 AND2X2_343 ( .A(_abc_17692_n1470), .B(_abc_17692_n1460), .Y(_abc_17692_n1472) );
  AND2X2 AND2X2_3430 ( .A(_abc_17692_n8577), .B(_abc_17692_n1863_bF_buf9), .Y(_abc_17692_n8578) );
  AND2X2 AND2X2_3431 ( .A(_abc_17692_n8578), .B(_abc_17692_n8576), .Y(_abc_17692_n8579) );
  AND2X2 AND2X2_3432 ( .A(_abc_17692_n8580), .B(state_10_bF_buf2), .Y(_abc_17692_n8581) );
  AND2X2 AND2X2_3433 ( .A(_abc_17692_n8469), .B(_abc_17692_n8583), .Y(_abc_17692_n8584) );
  AND2X2 AND2X2_3434 ( .A(_abc_17692_n8587), .B(_abc_17692_n1877_bF_buf9), .Y(_abc_17692_n8588) );
  AND2X2 AND2X2_3435 ( .A(_abc_17692_n8588), .B(_abc_17692_n8586), .Y(_abc_17692_n8589) );
  AND2X2 AND2X2_3436 ( .A(_abc_17692_n8551), .B(_abc_17692_n8590), .Y(_abc_17692_n8591) );
  AND2X2 AND2X2_3437 ( .A(_abc_17692_n8593), .B(_abc_17692_n1830_bF_buf9), .Y(_abc_17692_n8594) );
  AND2X2 AND2X2_3438 ( .A(_abc_17692_n8594), .B(_abc_17692_n8592), .Y(_abc_17692_n8595) );
  AND2X2 AND2X2_3439 ( .A(_abc_17692_n8598), .B(_abc_17692_n8571), .Y(_abc_17692_n8599) );
  AND2X2 AND2X2_344 ( .A(_abc_17692_n1473), .B(state_3_bF_buf4), .Y(_abc_17692_n1474) );
  AND2X2 AND2X2_3440 ( .A(_abc_17692_n8601), .B(_abc_17692_n1863_bF_buf8), .Y(_abc_17692_n8602) );
  AND2X2 AND2X2_3441 ( .A(_abc_17692_n8602), .B(_abc_17692_n8600), .Y(_abc_17692_n8603) );
  AND2X2 AND2X2_3442 ( .A(_abc_17692_n8604), .B(_abc_17692_n8532), .Y(_abc_17692_n8605) );
  AND2X2 AND2X2_3443 ( .A(_abc_17692_n8607), .B(_abc_17692_n1846_bF_buf9), .Y(_abc_17692_n8608) );
  AND2X2 AND2X2_3444 ( .A(_abc_17692_n8608), .B(_abc_17692_n8606), .Y(_abc_17692_n8609) );
  AND2X2 AND2X2_3445 ( .A(_abc_17692_n8611), .B(state_14_bF_buf2), .Y(_abc_17692_n8612) );
  AND2X2 AND2X2_3446 ( .A(_abc_17692_n8383_bF_buf2), .B(workunit1_2_), .Y(_abc_17692_n8613) );
  AND2X2 AND2X2_3447 ( .A(state_8_bF_buf5), .B(\data_in1[2] ), .Y(_abc_17692_n8614) );
  AND2X2 AND2X2_3448 ( .A(workunit2_3_), .B(workunit2_8_bF_buf1), .Y(_abc_17692_n8618) );
  AND2X2 AND2X2_3449 ( .A(_abc_17692_n2246), .B(_abc_17692_n3198), .Y(_abc_17692_n8619) );
  AND2X2 AND2X2_345 ( .A(_abc_17692_n1474), .B(_abc_17692_n1471), .Y(_abc_17692_n1475) );
  AND2X2 AND2X2_3450 ( .A(_abc_17692_n8500), .B(_abc_17692_n8621), .Y(_abc_17692_n8622) );
  AND2X2 AND2X2_3451 ( .A(_abc_17692_n8622), .B(_abc_17692_n8620), .Y(_abc_17692_n8623) );
  AND2X2 AND2X2_3452 ( .A(_abc_17692_n8625), .B(_abc_17692_n8624), .Y(_abc_17692_n8626) );
  AND2X2 AND2X2_3453 ( .A(_abc_17692_n8630), .B(_abc_17692_n8629), .Y(_abc_17692_n8631) );
  AND2X2 AND2X2_3454 ( .A(_abc_17692_n8632), .B(_abc_17692_n8628), .Y(_abc_17692_n8633) );
  AND2X2 AND2X2_3455 ( .A(_abc_17692_n8635), .B(_abc_17692_n8636), .Y(_abc_17692_n8637) );
  AND2X2 AND2X2_3456 ( .A(_abc_17692_n8634), .B(_abc_17692_n8638), .Y(_abc_17692_n8639) );
  AND2X2 AND2X2_3457 ( .A(_abc_17692_n8639), .B(_abc_17692_n8641), .Y(_abc_17692_n8642) );
  AND2X2 AND2X2_3458 ( .A(_abc_17692_n8644), .B(_abc_17692_n1877_bF_buf8), .Y(_abc_17692_n8645) );
  AND2X2 AND2X2_3459 ( .A(_abc_17692_n8645), .B(_abc_17692_n8643), .Y(_abc_17692_n8646) );
  AND2X2 AND2X2_346 ( .A(_abc_17692_n723), .B(sum_20_), .Y(_abc_17692_n1476) );
  AND2X2 AND2X2_3460 ( .A(_abc_17692_n8647), .B(_abc_17692_n8648), .Y(_abc_17692_n8649) );
  AND2X2 AND2X2_3461 ( .A(_abc_17692_n8652), .B(_abc_17692_n8651), .Y(_abc_17692_n8653) );
  AND2X2 AND2X2_3462 ( .A(_abc_17692_n8650), .B(_abc_17692_n8654), .Y(_abc_17692_n8655) );
  AND2X2 AND2X2_3463 ( .A(_abc_17692_n8528), .B(workunit1_2_), .Y(_abc_17692_n8657) );
  AND2X2 AND2X2_3464 ( .A(_abc_17692_n8542), .B(_abc_17692_n8658), .Y(_abc_17692_n8659) );
  AND2X2 AND2X2_3465 ( .A(_abc_17692_n8662), .B(_abc_17692_n1846_bF_buf8), .Y(_abc_17692_n8663) );
  AND2X2 AND2X2_3466 ( .A(_abc_17692_n8663), .B(_abc_17692_n8661), .Y(_abc_17692_n8664) );
  AND2X2 AND2X2_3467 ( .A(_abc_17692_n8665), .B(_abc_17692_n8666), .Y(_abc_17692_n8667) );
  AND2X2 AND2X2_3468 ( .A(_abc_17692_n8669), .B(_abc_17692_n8670), .Y(_abc_17692_n8671) );
  AND2X2 AND2X2_3469 ( .A(_abc_17692_n8674), .B(_abc_17692_n8671), .Y(_abc_17692_n8675) );
  AND2X2 AND2X2_347 ( .A(_abc_17692_n1437), .B(_abc_17692_n1402), .Y(_abc_17692_n1478) );
  AND2X2 AND2X2_3470 ( .A(_abc_17692_n8677), .B(_abc_17692_n1830_bF_buf8), .Y(_abc_17692_n8678) );
  AND2X2 AND2X2_3471 ( .A(_abc_17692_n8678), .B(_abc_17692_n8676), .Y(_abc_17692_n8679) );
  AND2X2 AND2X2_3472 ( .A(_abc_17692_n8682), .B(_abc_17692_n8683), .Y(_abc_17692_n8684) );
  AND2X2 AND2X2_3473 ( .A(_abc_17692_n8687), .B(_abc_17692_n8686), .Y(_abc_17692_n8688) );
  AND2X2 AND2X2_3474 ( .A(_abc_17692_n8685), .B(_abc_17692_n8689), .Y(_abc_17692_n8690) );
  AND2X2 AND2X2_3475 ( .A(_abc_17692_n8576), .B(_abc_17692_n8692), .Y(_abc_17692_n8693) );
  AND2X2 AND2X2_3476 ( .A(_abc_17692_n8694), .B(_abc_17692_n8691), .Y(_abc_17692_n8696) );
  AND2X2 AND2X2_3477 ( .A(_abc_17692_n8697), .B(_abc_17692_n1863_bF_buf7), .Y(_abc_17692_n8698) );
  AND2X2 AND2X2_3478 ( .A(_abc_17692_n8698), .B(_abc_17692_n8695), .Y(_abc_17692_n8699) );
  AND2X2 AND2X2_3479 ( .A(_abc_17692_n8700), .B(state_10_bF_buf1), .Y(_abc_17692_n8701) );
  AND2X2 AND2X2_348 ( .A(_abc_17692_n1387), .B(_abc_17692_n1478), .Y(_abc_17692_n1479) );
  AND2X2 AND2X2_3480 ( .A(_abc_17692_n8587), .B(_abc_17692_n8703), .Y(_abc_17692_n8704) );
  AND2X2 AND2X2_3481 ( .A(_abc_17692_n8707), .B(_abc_17692_n1877_bF_buf7), .Y(_abc_17692_n8708) );
  AND2X2 AND2X2_3482 ( .A(_abc_17692_n8708), .B(_abc_17692_n8706), .Y(_abc_17692_n8709) );
  AND2X2 AND2X2_3483 ( .A(_abc_17692_n8711), .B(_abc_17692_n8710), .Y(_abc_17692_n8712) );
  AND2X2 AND2X2_3484 ( .A(_abc_17692_n8712), .B(_abc_17692_n8713), .Y(_abc_17692_n8714) );
  AND2X2 AND2X2_3485 ( .A(_abc_17692_n8716), .B(_abc_17692_n1830_bF_buf7), .Y(_abc_17692_n8717) );
  AND2X2 AND2X2_3486 ( .A(_abc_17692_n8717), .B(_abc_17692_n8715), .Y(_abc_17692_n8718) );
  AND2X2 AND2X2_3487 ( .A(_abc_17692_n8721), .B(_abc_17692_n8690), .Y(_abc_17692_n8722) );
  AND2X2 AND2X2_3488 ( .A(_abc_17692_n8724), .B(_abc_17692_n1863_bF_buf6), .Y(_abc_17692_n8725) );
  AND2X2 AND2X2_3489 ( .A(_abc_17692_n8725), .B(_abc_17692_n8723), .Y(_abc_17692_n8726) );
  AND2X2 AND2X2_349 ( .A(_abc_17692_n1480), .B(_abc_17692_n1478), .Y(_abc_17692_n1481) );
  AND2X2 AND2X2_3490 ( .A(_abc_17692_n8728), .B(_abc_17692_n8655), .Y(_abc_17692_n8729) );
  AND2X2 AND2X2_3491 ( .A(_abc_17692_n8731), .B(_abc_17692_n1846_bF_buf7), .Y(_abc_17692_n8732) );
  AND2X2 AND2X2_3492 ( .A(_abc_17692_n8732), .B(_abc_17692_n8730), .Y(_abc_17692_n8733) );
  AND2X2 AND2X2_3493 ( .A(_abc_17692_n8735), .B(state_14_bF_buf1), .Y(_abc_17692_n8736) );
  AND2X2 AND2X2_3494 ( .A(_abc_17692_n8383_bF_buf1), .B(workunit1_3_), .Y(_abc_17692_n8737) );
  AND2X2 AND2X2_3495 ( .A(state_8_bF_buf4), .B(\data_in1[3] ), .Y(_abc_17692_n8738) );
  AND2X2 AND2X2_3496 ( .A(_abc_17692_n8742), .B(_abc_17692_n8743), .Y(_abc_17692_n8744) );
  AND2X2 AND2X2_3497 ( .A(_abc_17692_n3471), .B(workunit2_0_), .Y(_abc_17692_n8746) );
  AND2X2 AND2X2_3498 ( .A(_abc_17692_n1814), .B(workunit2_9_), .Y(_abc_17692_n8747) );
  AND2X2 AND2X2_3499 ( .A(_abc_17692_n8749), .B(_abc_17692_n8745), .Y(_abc_17692_n8750) );
  AND2X2 AND2X2_35 ( .A(_abc_17692_n627), .B(_abc_17692_n712), .Y(_abc_17692_n713) );
  AND2X2 AND2X2_350 ( .A(_abc_17692_n1437), .B(_abc_17692_n1444), .Y(_abc_17692_n1482) );
  AND2X2 AND2X2_3500 ( .A(_abc_17692_n8501), .B(_abc_17692_n8752), .Y(_abc_17692_n8753) );
  AND2X2 AND2X2_3501 ( .A(_abc_17692_n8624), .B(_abc_17692_n8497), .Y(_abc_17692_n8754) );
  AND2X2 AND2X2_3502 ( .A(_abc_17692_n8756), .B(_abc_17692_n8750), .Y(_abc_17692_n8757) );
  AND2X2 AND2X2_3503 ( .A(_abc_17692_n8748), .B(workunit2_4_), .Y(_abc_17692_n8758) );
  AND2X2 AND2X2_3504 ( .A(_abc_17692_n8744), .B(_abc_17692_n2482), .Y(_abc_17692_n8759) );
  AND2X2 AND2X2_3505 ( .A(_abc_17692_n8762), .B(_abc_17692_n8761), .Y(_abc_17692_n8763) );
  AND2X2 AND2X2_3506 ( .A(_abc_17692_n8763), .B(_abc_17692_n8760), .Y(_abc_17692_n8764) );
  AND2X2 AND2X2_3507 ( .A(_abc_17692_n2478), .B(_abc_17692_n8765), .Y(_abc_17692_n8766) );
  AND2X2 AND2X2_3508 ( .A(_abc_17692_n8767), .B(_abc_17692_n2476), .Y(_abc_17692_n8768) );
  AND2X2 AND2X2_3509 ( .A(_abc_17692_n8769), .B(workunit1_4_), .Y(_abc_17692_n8770) );
  AND2X2 AND2X2_351 ( .A(_abc_17692_n1432), .B(sum_19_), .Y(_abc_17692_n1483) );
  AND2X2 AND2X2_3510 ( .A(_abc_17692_n8771), .B(_abc_17692_n2433), .Y(_abc_17692_n8772) );
  AND2X2 AND2X2_3511 ( .A(_abc_17692_n8775), .B(_abc_17692_n8773), .Y(_abc_17692_n8776) );
  AND2X2 AND2X2_3512 ( .A(_abc_17692_n8778), .B(_abc_17692_n1830_bF_buf6), .Y(_abc_17692_n8779) );
  AND2X2 AND2X2_3513 ( .A(_abc_17692_n8779), .B(_abc_17692_n8777), .Y(_abc_17692_n8780) );
  AND2X2 AND2X2_3514 ( .A(_abc_17692_n2510), .B(_abc_17692_n8765), .Y(_abc_17692_n8781) );
  AND2X2 AND2X2_3515 ( .A(_abc_17692_n8767), .B(_abc_17692_n2508), .Y(_abc_17692_n8782) );
  AND2X2 AND2X2_3516 ( .A(_abc_17692_n8785), .B(_abc_17692_n8786), .Y(_abc_17692_n8787) );
  AND2X2 AND2X2_3517 ( .A(_abc_17692_n8789), .B(_abc_17692_n8787), .Y(_abc_17692_n8791) );
  AND2X2 AND2X2_3518 ( .A(_abc_17692_n8792), .B(_abc_17692_n1877_bF_buf6), .Y(_abc_17692_n8793) );
  AND2X2 AND2X2_3519 ( .A(_abc_17692_n8793), .B(_abc_17692_n8790), .Y(_abc_17692_n8794) );
  AND2X2 AND2X2_352 ( .A(_abc_17692_n1486), .B(_abc_17692_n1477), .Y(_abc_17692_n1487) );
  AND2X2 AND2X2_3520 ( .A(_abc_17692_n2543), .B(_abc_17692_n8765), .Y(_abc_17692_n8795) );
  AND2X2 AND2X2_3521 ( .A(_abc_17692_n8767), .B(_abc_17692_n2541), .Y(_abc_17692_n8796) );
  AND2X2 AND2X2_3522 ( .A(_abc_17692_n8797), .B(workunit1_4_), .Y(_abc_17692_n8798) );
  AND2X2 AND2X2_3523 ( .A(_abc_17692_n8799), .B(_abc_17692_n2433), .Y(_abc_17692_n8800) );
  AND2X2 AND2X2_3524 ( .A(_abc_17692_n8649), .B(workunit1_3_), .Y(_abc_17692_n8802) );
  AND2X2 AND2X2_3525 ( .A(_abc_17692_n8662), .B(_abc_17692_n8803), .Y(_abc_17692_n8804) );
  AND2X2 AND2X2_3526 ( .A(_abc_17692_n8805), .B(_abc_17692_n8801), .Y(_abc_17692_n8806) );
  AND2X2 AND2X2_3527 ( .A(_abc_17692_n8808), .B(_abc_17692_n1846_bF_buf6), .Y(_abc_17692_n8809) );
  AND2X2 AND2X2_3528 ( .A(_abc_17692_n8809), .B(_abc_17692_n8807), .Y(_abc_17692_n8810) );
  AND2X2 AND2X2_3529 ( .A(_abc_17692_n8813), .B(_abc_17692_n8814), .Y(_abc_17692_n8815) );
  AND2X2 AND2X2_353 ( .A(_abc_17692_n1489), .B(state_15_bF_buf4), .Y(_abc_17692_n1490) );
  AND2X2 AND2X2_3530 ( .A(_abc_17692_n8817), .B(_abc_17692_n8818), .Y(_abc_17692_n8819) );
  AND2X2 AND2X2_3531 ( .A(_abc_17692_n8820), .B(_abc_17692_n8816), .Y(_abc_17692_n8821) );
  AND2X2 AND2X2_3532 ( .A(_abc_17692_n8825), .B(_abc_17692_n8822), .Y(_abc_17692_n8826) );
  AND2X2 AND2X2_3533 ( .A(_abc_17692_n8828), .B(_abc_17692_n1863_bF_buf5), .Y(_abc_17692_n8829) );
  AND2X2 AND2X2_3534 ( .A(_abc_17692_n8829), .B(_abc_17692_n8827), .Y(_abc_17692_n8830) );
  AND2X2 AND2X2_3535 ( .A(_abc_17692_n8831), .B(state_10_bF_buf0), .Y(_abc_17692_n8832) );
  AND2X2 AND2X2_3536 ( .A(_abc_17692_n8707), .B(_abc_17692_n8834), .Y(_abc_17692_n8835) );
  AND2X2 AND2X2_3537 ( .A(_abc_17692_n8838), .B(_abc_17692_n1877_bF_buf5), .Y(_abc_17692_n8839) );
  AND2X2 AND2X2_3538 ( .A(_abc_17692_n8839), .B(_abc_17692_n8837), .Y(_abc_17692_n8840) );
  AND2X2 AND2X2_3539 ( .A(_abc_17692_n8843), .B(_abc_17692_n8841), .Y(_abc_17692_n8844) );
  AND2X2 AND2X2_354 ( .A(_abc_17692_n1490), .B(_abc_17692_n1488), .Y(_abc_17692_n1491) );
  AND2X2 AND2X2_3540 ( .A(_abc_17692_n8846), .B(_abc_17692_n1830_bF_buf5), .Y(_abc_17692_n8847) );
  AND2X2 AND2X2_3541 ( .A(_abc_17692_n8847), .B(_abc_17692_n8845), .Y(_abc_17692_n8848) );
  AND2X2 AND2X2_3542 ( .A(_abc_17692_n8851), .B(_abc_17692_n8821), .Y(_abc_17692_n8852) );
  AND2X2 AND2X2_3543 ( .A(_abc_17692_n8854), .B(_abc_17692_n1863_bF_buf4), .Y(_abc_17692_n8855) );
  AND2X2 AND2X2_3544 ( .A(_abc_17692_n8855), .B(_abc_17692_n8853), .Y(_abc_17692_n8856) );
  AND2X2 AND2X2_3545 ( .A(_abc_17692_n8859), .B(_abc_17692_n8857), .Y(_abc_17692_n8860) );
  AND2X2 AND2X2_3546 ( .A(_abc_17692_n8862), .B(_abc_17692_n1846_bF_buf5), .Y(_abc_17692_n8863) );
  AND2X2 AND2X2_3547 ( .A(_abc_17692_n8863), .B(_abc_17692_n8861), .Y(_abc_17692_n8864) );
  AND2X2 AND2X2_3548 ( .A(_abc_17692_n8866), .B(state_14_bF_buf0), .Y(_abc_17692_n8867) );
  AND2X2 AND2X2_3549 ( .A(_abc_17692_n8383_bF_buf0), .B(workunit1_4_), .Y(_abc_17692_n8868) );
  AND2X2 AND2X2_355 ( .A(delta_21_), .B(sum_21_), .Y(_abc_17692_n1494) );
  AND2X2 AND2X2_3550 ( .A(state_8_bF_buf3), .B(\data_in1[4] ), .Y(_abc_17692_n8869) );
  AND2X2 AND2X2_3551 ( .A(_abc_17692_n8873), .B(_abc_17692_n8745), .Y(_abc_17692_n8874) );
  AND2X2 AND2X2_3552 ( .A(workunit2_1_bF_buf2), .B(workunit2_10_bF_buf3), .Y(_abc_17692_n8875) );
  AND2X2 AND2X2_3553 ( .A(_abc_17692_n1919_1), .B(_abc_17692_n3751), .Y(_abc_17692_n8876) );
  AND2X2 AND2X2_3554 ( .A(_abc_17692_n8879), .B(_abc_17692_n8880), .Y(_abc_17692_n8881) );
  AND2X2 AND2X2_3555 ( .A(_abc_17692_n8878), .B(_abc_17692_n8882), .Y(_abc_17692_n8883) );
  AND2X2 AND2X2_3556 ( .A(_abc_17692_n8874), .B(_abc_17692_n8883), .Y(_abc_17692_n8884) );
  AND2X2 AND2X2_3557 ( .A(_abc_17692_n8881), .B(workunit2_5_), .Y(_abc_17692_n8886) );
  AND2X2 AND2X2_3558 ( .A(_abc_17692_n8877), .B(_abc_17692_n2633), .Y(_abc_17692_n8887) );
  AND2X2 AND2X2_3559 ( .A(_abc_17692_n8885), .B(_abc_17692_n8888), .Y(_abc_17692_n8889) );
  AND2X2 AND2X2_356 ( .A(_abc_17692_n1496), .B(_abc_17692_n1497), .Y(_abc_17692_n1498) );
  AND2X2 AND2X2_3560 ( .A(_abc_17692_n2664), .B(_abc_17692_n8890), .Y(_abc_17692_n8891) );
  AND2X2 AND2X2_3561 ( .A(_abc_17692_n8893), .B(_abc_17692_n8892), .Y(_abc_17692_n8894) );
  AND2X2 AND2X2_3562 ( .A(_abc_17692_n2663), .B(_abc_17692_n8894), .Y(_abc_17692_n8895) );
  AND2X2 AND2X2_3563 ( .A(_abc_17692_n8898), .B(_abc_17692_n8899), .Y(_abc_17692_n8900) );
  AND2X2 AND2X2_3564 ( .A(_abc_17692_n8902), .B(_abc_17692_n8900), .Y(_abc_17692_n8903) );
  AND2X2 AND2X2_3565 ( .A(_abc_17692_n8905), .B(_abc_17692_n1877_bF_buf4), .Y(_abc_17692_n8906) );
  AND2X2 AND2X2_3566 ( .A(_abc_17692_n8906), .B(_abc_17692_n8904), .Y(_abc_17692_n8907) );
  AND2X2 AND2X2_3567 ( .A(_abc_17692_n8909), .B(_abc_17692_n8908), .Y(_abc_17692_n8910) );
  AND2X2 AND2X2_3568 ( .A(_abc_17692_n8911), .B(workunit1_5_), .Y(_abc_17692_n8912) );
  AND2X2 AND2X2_3569 ( .A(_abc_17692_n8913), .B(_abc_17692_n8914), .Y(_abc_17692_n8915) );
  AND2X2 AND2X2_357 ( .A(_abc_17692_n1499), .B(_abc_17692_n1495), .Y(_abc_17692_n1500) );
  AND2X2 AND2X2_3570 ( .A(_abc_17692_n8771), .B(workunit1_4_), .Y(_abc_17692_n8916) );
  AND2X2 AND2X2_3571 ( .A(_abc_17692_n8917), .B(_abc_17692_n8915), .Y(_abc_17692_n8918) );
  AND2X2 AND2X2_3572 ( .A(_abc_17692_n8920), .B(_abc_17692_n1830_bF_buf4), .Y(_abc_17692_n8921) );
  AND2X2 AND2X2_3573 ( .A(_abc_17692_n8921), .B(_abc_17692_n8919), .Y(_abc_17692_n8922) );
  AND2X2 AND2X2_3574 ( .A(_abc_17692_n8890), .B(_abc_17692_n2720), .Y(_abc_17692_n8923) );
  AND2X2 AND2X2_3575 ( .A(_abc_17692_n8894), .B(_abc_17692_n2724), .Y(_abc_17692_n8924) );
  AND2X2 AND2X2_3576 ( .A(_abc_17692_n8927), .B(_abc_17692_n8928), .Y(_abc_17692_n8929) );
  AND2X2 AND2X2_3577 ( .A(_abc_17692_n8926), .B(_abc_17692_n8930), .Y(_abc_17692_n8931) );
  AND2X2 AND2X2_3578 ( .A(_abc_17692_n8799), .B(workunit1_4_), .Y(_abc_17692_n8933) );
  AND2X2 AND2X2_3579 ( .A(_abc_17692_n8934), .B(_abc_17692_n8932), .Y(_abc_17692_n8936) );
  AND2X2 AND2X2_358 ( .A(delta_20_), .B(sum_20_), .Y(_abc_17692_n1501) );
  AND2X2 AND2X2_3580 ( .A(_abc_17692_n8937), .B(_abc_17692_n1846_bF_buf4), .Y(_abc_17692_n8938) );
  AND2X2 AND2X2_3581 ( .A(_abc_17692_n8938), .B(_abc_17692_n8935), .Y(_abc_17692_n8939) );
  AND2X2 AND2X2_3582 ( .A(_abc_17692_n8942), .B(_abc_17692_n8943), .Y(_abc_17692_n8944) );
  AND2X2 AND2X2_3583 ( .A(_abc_17692_n8946), .B(_abc_17692_n8947), .Y(_abc_17692_n8948) );
  AND2X2 AND2X2_3584 ( .A(_abc_17692_n8945), .B(_abc_17692_n8949), .Y(_abc_17692_n8950) );
  AND2X2 AND2X2_3585 ( .A(_abc_17692_n8954), .B(_abc_17692_n8951), .Y(_abc_17692_n8955) );
  AND2X2 AND2X2_3586 ( .A(_abc_17692_n8957), .B(_abc_17692_n1863_bF_buf3), .Y(_abc_17692_n8958) );
  AND2X2 AND2X2_3587 ( .A(_abc_17692_n8958), .B(_abc_17692_n8956), .Y(_abc_17692_n8959) );
  AND2X2 AND2X2_3588 ( .A(_abc_17692_n8960), .B(state_10_bF_buf4), .Y(_abc_17692_n8961) );
  AND2X2 AND2X2_3589 ( .A(_abc_17692_n8783), .B(workunit1_4_), .Y(_abc_17692_n8963) );
  AND2X2 AND2X2_359 ( .A(_abc_17692_n1473), .B(_abc_17692_n1502), .Y(_abc_17692_n1503) );
  AND2X2 AND2X2_3590 ( .A(_abc_17692_n8838), .B(_abc_17692_n8964), .Y(_abc_17692_n8965) );
  AND2X2 AND2X2_3591 ( .A(_abc_17692_n8968), .B(_abc_17692_n1877_bF_buf3), .Y(_abc_17692_n8969) );
  AND2X2 AND2X2_3592 ( .A(_abc_17692_n8969), .B(_abc_17692_n8967), .Y(_abc_17692_n8970) );
  AND2X2 AND2X2_3593 ( .A(_abc_17692_n8972), .B(_abc_17692_n8971), .Y(_abc_17692_n8973) );
  AND2X2 AND2X2_3594 ( .A(_abc_17692_n8975), .B(_abc_17692_n1830_bF_buf3), .Y(_abc_17692_n8976) );
  AND2X2 AND2X2_3595 ( .A(_abc_17692_n8976), .B(_abc_17692_n8974), .Y(_abc_17692_n8977) );
  AND2X2 AND2X2_3596 ( .A(_abc_17692_n8980), .B(_abc_17692_n8950), .Y(_abc_17692_n8981) );
  AND2X2 AND2X2_3597 ( .A(_abc_17692_n8983), .B(_abc_17692_n1863_bF_buf2), .Y(_abc_17692_n8984) );
  AND2X2 AND2X2_3598 ( .A(_abc_17692_n8984), .B(_abc_17692_n8982), .Y(_abc_17692_n8985) );
  AND2X2 AND2X2_3599 ( .A(_abc_17692_n8986), .B(_abc_17692_n8931), .Y(_abc_17692_n8987) );
  AND2X2 AND2X2_36 ( .A(_abc_17692_n715_1), .B(_abc_17692_n713), .Y(_abc_17692_n716) );
  AND2X2 AND2X2_360 ( .A(_abc_17692_n1507), .B(state_3_bF_buf3), .Y(_abc_17692_n1508) );
  AND2X2 AND2X2_3600 ( .A(_abc_17692_n8989), .B(_abc_17692_n1846_bF_buf3), .Y(_abc_17692_n8990) );
  AND2X2 AND2X2_3601 ( .A(_abc_17692_n8990), .B(_abc_17692_n8988), .Y(_abc_17692_n8991) );
  AND2X2 AND2X2_3602 ( .A(_abc_17692_n8993), .B(state_14_bF_buf4), .Y(_abc_17692_n8994) );
  AND2X2 AND2X2_3603 ( .A(_abc_17692_n8383_bF_buf4), .B(workunit1_5_), .Y(_abc_17692_n8995) );
  AND2X2 AND2X2_3604 ( .A(state_8_bF_buf2), .B(\data_in1[5] ), .Y(_abc_17692_n8996) );
  AND2X2 AND2X2_3605 ( .A(_abc_17692_n9002), .B(_abc_17692_n8878), .Y(_abc_17692_n9003) );
  AND2X2 AND2X2_3606 ( .A(_abc_17692_n9001), .B(_abc_17692_n9003), .Y(_abc_17692_n9004) );
  AND2X2 AND2X2_3607 ( .A(workunit2_2_), .B(workunit2_11_), .Y(_abc_17692_n9005) );
  AND2X2 AND2X2_3608 ( .A(_abc_17692_n9006), .B(_abc_17692_n9007), .Y(_abc_17692_n9008) );
  AND2X2 AND2X2_3609 ( .A(_abc_17692_n9008), .B(workunit2_6_), .Y(_abc_17692_n9009) );
  AND2X2 AND2X2_361 ( .A(_abc_17692_n1508), .B(_abc_17692_n1505), .Y(_abc_17692_n1509) );
  AND2X2 AND2X2_3610 ( .A(_abc_17692_n2091), .B(_abc_17692_n3905), .Y(_abc_17692_n9010) );
  AND2X2 AND2X2_3611 ( .A(_abc_17692_n9011), .B(_abc_17692_n2862), .Y(_abc_17692_n9012) );
  AND2X2 AND2X2_3612 ( .A(_abc_17692_n9004), .B(_abc_17692_n9013), .Y(_abc_17692_n9014) );
  AND2X2 AND2X2_3613 ( .A(_abc_17692_n8750), .B(_abc_17692_n8883), .Y(_abc_17692_n9015) );
  AND2X2 AND2X2_3614 ( .A(_abc_17692_n8756), .B(_abc_17692_n9015), .Y(_abc_17692_n9016) );
  AND2X2 AND2X2_3615 ( .A(_abc_17692_n9017), .B(_abc_17692_n8882), .Y(_abc_17692_n9018) );
  AND2X2 AND2X2_3616 ( .A(_abc_17692_n9020), .B(_abc_17692_n9021), .Y(_abc_17692_n9022) );
  AND2X2 AND2X2_3617 ( .A(_abc_17692_n9019), .B(_abc_17692_n9022), .Y(_abc_17692_n9023) );
  AND2X2 AND2X2_3618 ( .A(_abc_17692_n2890), .B(_abc_17692_n9024), .Y(_abc_17692_n9025) );
  AND2X2 AND2X2_3619 ( .A(_abc_17692_n9026), .B(_abc_17692_n2888), .Y(_abc_17692_n9027) );
  AND2X2 AND2X2_362 ( .A(_abc_17692_n1477), .B(_abc_17692_n1506), .Y(_abc_17692_n1512) );
  AND2X2 AND2X2_3620 ( .A(_abc_17692_n9028), .B(workunit1_6_), .Y(_abc_17692_n9029) );
  AND2X2 AND2X2_3621 ( .A(_abc_17692_n9030), .B(_abc_17692_n2821), .Y(_abc_17692_n9031) );
  AND2X2 AND2X2_3622 ( .A(_abc_17692_n9033), .B(_abc_17692_n9032), .Y(_abc_17692_n9034) );
  AND2X2 AND2X2_3623 ( .A(_abc_17692_n9036), .B(_abc_17692_n1830_bF_buf2), .Y(_abc_17692_n9037) );
  AND2X2 AND2X2_3624 ( .A(_abc_17692_n9037), .B(_abc_17692_n9035), .Y(_abc_17692_n9038) );
  AND2X2 AND2X2_3625 ( .A(_abc_17692_n2856), .B(_abc_17692_n9024), .Y(_abc_17692_n9039) );
  AND2X2 AND2X2_3626 ( .A(_abc_17692_n2857), .B(_abc_17692_n9026), .Y(_abc_17692_n9040) );
  AND2X2 AND2X2_3627 ( .A(_abc_17692_n9041), .B(workunit1_6_), .Y(_abc_17692_n9042) );
  AND2X2 AND2X2_3628 ( .A(_abc_17692_n9043), .B(_abc_17692_n2821), .Y(_abc_17692_n9044) );
  AND2X2 AND2X2_3629 ( .A(_abc_17692_n9047), .B(_abc_17692_n9045), .Y(_abc_17692_n9049) );
  AND2X2 AND2X2_363 ( .A(_abc_17692_n1486), .B(_abc_17692_n1512), .Y(_abc_17692_n1513) );
  AND2X2 AND2X2_3630 ( .A(_abc_17692_n9050), .B(_abc_17692_n1877_bF_buf2), .Y(_abc_17692_n9051) );
  AND2X2 AND2X2_3631 ( .A(_abc_17692_n9051), .B(_abc_17692_n9048), .Y(_abc_17692_n9052) );
  AND2X2 AND2X2_3632 ( .A(_abc_17692_n2925), .B(_abc_17692_n9024), .Y(_abc_17692_n9053) );
  AND2X2 AND2X2_3633 ( .A(_abc_17692_n9026), .B(_abc_17692_n2923), .Y(_abc_17692_n9054) );
  AND2X2 AND2X2_3634 ( .A(_abc_17692_n9056), .B(workunit1_6_), .Y(_abc_17692_n9057) );
  AND2X2 AND2X2_3635 ( .A(_abc_17692_n9055), .B(_abc_17692_n2821), .Y(_abc_17692_n9058) );
  AND2X2 AND2X2_3636 ( .A(_abc_17692_n8925), .B(workunit1_5_), .Y(_abc_17692_n9063) );
  AND2X2 AND2X2_3637 ( .A(_abc_17692_n9066), .B(_abc_17692_n9064), .Y(_abc_17692_n9067) );
  AND2X2 AND2X2_3638 ( .A(_abc_17692_n9062), .B(_abc_17692_n9067), .Y(_abc_17692_n9068) );
  AND2X2 AND2X2_3639 ( .A(_abc_17692_n9069), .B(_abc_17692_n9060), .Y(_abc_17692_n9071) );
  AND2X2 AND2X2_364 ( .A(_abc_17692_n1506), .B(_abc_17692_n1459_1), .Y(_abc_17692_n1515) );
  AND2X2 AND2X2_3640 ( .A(_abc_17692_n9072), .B(_abc_17692_n1846_bF_buf2), .Y(_abc_17692_n9073) );
  AND2X2 AND2X2_3641 ( .A(_abc_17692_n9073), .B(_abc_17692_n9070), .Y(_abc_17692_n9074) );
  AND2X2 AND2X2_3642 ( .A(_abc_17692_n2962), .B(_abc_17692_n9024), .Y(_abc_17692_n9077) );
  AND2X2 AND2X2_3643 ( .A(_abc_17692_n2963), .B(_abc_17692_n9026), .Y(_abc_17692_n9078) );
  AND2X2 AND2X2_3644 ( .A(_abc_17692_n9082), .B(_abc_17692_n9080), .Y(_abc_17692_n9083) );
  AND2X2 AND2X2_3645 ( .A(_abc_17692_n9086), .B(_abc_17692_n9083), .Y(_abc_17692_n9088) );
  AND2X2 AND2X2_3646 ( .A(_abc_17692_n9089), .B(_abc_17692_n1863_bF_buf1), .Y(_abc_17692_n9090) );
  AND2X2 AND2X2_3647 ( .A(_abc_17692_n9090), .B(_abc_17692_n9087), .Y(_abc_17692_n9091) );
  AND2X2 AND2X2_3648 ( .A(_abc_17692_n9092), .B(state_10_bF_buf3), .Y(_abc_17692_n9093) );
  AND2X2 AND2X2_3649 ( .A(_abc_17692_n9097), .B(_abc_17692_n9094), .Y(_abc_17692_n9098) );
  AND2X2 AND2X2_365 ( .A(_abc_17692_n1516), .B(state_15_bF_buf3), .Y(_abc_17692_n1517_1) );
  AND2X2 AND2X2_3650 ( .A(_abc_17692_n9100), .B(_abc_17692_n1830_bF_buf1), .Y(_abc_17692_n9101) );
  AND2X2 AND2X2_3651 ( .A(_abc_17692_n9101), .B(_abc_17692_n9099), .Y(_abc_17692_n9102) );
  AND2X2 AND2X2_3652 ( .A(_abc_17692_n9104), .B(_abc_17692_n9059), .Y(_abc_17692_n9106) );
  AND2X2 AND2X2_3653 ( .A(_abc_17692_n9107), .B(_abc_17692_n1846_bF_buf1), .Y(_abc_17692_n9108) );
  AND2X2 AND2X2_3654 ( .A(_abc_17692_n9108), .B(_abc_17692_n9105), .Y(_abc_17692_n9109) );
  AND2X2 AND2X2_3655 ( .A(_abc_17692_n9113), .B(_abc_17692_n9111), .Y(_abc_17692_n9114) );
  AND2X2 AND2X2_3656 ( .A(_abc_17692_n9116), .B(_abc_17692_n1863_bF_buf0), .Y(_abc_17692_n9117) );
  AND2X2 AND2X2_3657 ( .A(_abc_17692_n9117), .B(_abc_17692_n9115), .Y(_abc_17692_n9118) );
  AND2X2 AND2X2_3658 ( .A(_abc_17692_n8897), .B(workunit1_5_), .Y(_abc_17692_n9119) );
  AND2X2 AND2X2_3659 ( .A(_abc_17692_n8968), .B(_abc_17692_n9120), .Y(_abc_17692_n9121) );
  AND2X2 AND2X2_366 ( .A(_abc_17692_n1514), .B(_abc_17692_n1517_1), .Y(_abc_17692_n1518) );
  AND2X2 AND2X2_3660 ( .A(_abc_17692_n9125), .B(_abc_17692_n1877_bF_buf1), .Y(_abc_17692_n9126) );
  AND2X2 AND2X2_3661 ( .A(_abc_17692_n9126), .B(_abc_17692_n9122), .Y(_abc_17692_n9127) );
  AND2X2 AND2X2_3662 ( .A(_abc_17692_n9129), .B(state_14_bF_buf3), .Y(_abc_17692_n9130) );
  AND2X2 AND2X2_3663 ( .A(_abc_17692_n8383_bF_buf3), .B(workunit1_6_), .Y(_abc_17692_n9131) );
  AND2X2 AND2X2_3664 ( .A(state_8_bF_buf1), .B(\data_in1[6] ), .Y(_abc_17692_n9132) );
  AND2X2 AND2X2_3665 ( .A(_abc_17692_n9136), .B(_abc_17692_n9020), .Y(_abc_17692_n9137) );
  AND2X2 AND2X2_3666 ( .A(workunit2_3_), .B(workunit2_12_bF_buf1), .Y(_abc_17692_n9138) );
  AND2X2 AND2X2_3667 ( .A(_abc_17692_n9139), .B(_abc_17692_n9140), .Y(_abc_17692_n9141) );
  AND2X2 AND2X2_3668 ( .A(_abc_17692_n9141), .B(workunit2_7_), .Y(_abc_17692_n9142) );
  AND2X2 AND2X2_3669 ( .A(_abc_17692_n9143), .B(_abc_17692_n9144), .Y(_abc_17692_n9145) );
  AND2X2 AND2X2_367 ( .A(_abc_17692_n1518), .B(_abc_17692_n1511), .Y(_abc_17692_n1519) );
  AND2X2 AND2X2_3670 ( .A(_abc_17692_n9145), .B(_abc_17692_n3060), .Y(_abc_17692_n9146) );
  AND2X2 AND2X2_3671 ( .A(_abc_17692_n9137), .B(_abc_17692_n9147), .Y(_abc_17692_n9148) );
  AND2X2 AND2X2_3672 ( .A(_abc_17692_n9150), .B(_abc_17692_n9151), .Y(_abc_17692_n9152) );
  AND2X2 AND2X2_3673 ( .A(_abc_17692_n9149), .B(_abc_17692_n9152), .Y(_abc_17692_n9153) );
  AND2X2 AND2X2_3674 ( .A(_abc_17692_n9157), .B(_abc_17692_n9156), .Y(_abc_17692_n9158) );
  AND2X2 AND2X2_3675 ( .A(_abc_17692_n9155), .B(_abc_17692_n9159), .Y(_abc_17692_n9160) );
  AND2X2 AND2X2_3676 ( .A(_abc_17692_n9162), .B(_abc_17692_n9163), .Y(_abc_17692_n9164) );
  AND2X2 AND2X2_3677 ( .A(_abc_17692_n9161), .B(_abc_17692_n9165), .Y(_abc_17692_n9166) );
  AND2X2 AND2X2_3678 ( .A(_abc_17692_n9072), .B(_abc_17692_n9168), .Y(_abc_17692_n9169) );
  AND2X2 AND2X2_3679 ( .A(_abc_17692_n9172), .B(_abc_17692_n1846_bF_buf0), .Y(_abc_17692_n9173) );
  AND2X2 AND2X2_368 ( .A(_abc_17692_n722_bF_buf0), .B(sum_21_), .Y(_abc_17692_n1520_1) );
  AND2X2 AND2X2_3680 ( .A(_abc_17692_n9173), .B(_abc_17692_n9171), .Y(_abc_17692_n9174) );
  AND2X2 AND2X2_3681 ( .A(_abc_17692_n3081), .B(_abc_17692_n9154), .Y(_abc_17692_n9175) );
  AND2X2 AND2X2_3682 ( .A(_abc_17692_n3082), .B(_abc_17692_n9158), .Y(_abc_17692_n9176) );
  AND2X2 AND2X2_3683 ( .A(_abc_17692_n9178), .B(workunit1_7_), .Y(_abc_17692_n9179) );
  AND2X2 AND2X2_3684 ( .A(_abc_17692_n9177), .B(_abc_17692_n2063), .Y(_abc_17692_n9180) );
  AND2X2 AND2X2_3685 ( .A(_abc_17692_n9043), .B(workunit1_6_), .Y(_abc_17692_n9182) );
  AND2X2 AND2X2_3686 ( .A(_abc_17692_n9183), .B(_abc_17692_n9181), .Y(_abc_17692_n9184) );
  AND2X2 AND2X2_3687 ( .A(_abc_17692_n9186), .B(_abc_17692_n1877_bF_buf0), .Y(_abc_17692_n9187) );
  AND2X2 AND2X2_3688 ( .A(_abc_17692_n9187), .B(_abc_17692_n9185), .Y(_abc_17692_n9188) );
  AND2X2 AND2X2_3689 ( .A(_abc_17692_n9030), .B(workunit1_6_), .Y(_abc_17692_n9189) );
  AND2X2 AND2X2_369 ( .A(delta_22_), .B(sum_22_), .Y(_abc_17692_n1524) );
  AND2X2 AND2X2_3690 ( .A(_abc_17692_n3056), .B(_abc_17692_n9154), .Y(_abc_17692_n9190) );
  AND2X2 AND2X2_3691 ( .A(_abc_17692_n3051), .B(_abc_17692_n9158), .Y(_abc_17692_n9191) );
  AND2X2 AND2X2_3692 ( .A(_abc_17692_n9193), .B(workunit1_7_), .Y(_abc_17692_n9194) );
  AND2X2 AND2X2_3693 ( .A(_abc_17692_n9192), .B(_abc_17692_n2063), .Y(_abc_17692_n9195) );
  AND2X2 AND2X2_3694 ( .A(_abc_17692_n9034), .B(_abc_17692_n9196), .Y(_abc_17692_n9199) );
  AND2X2 AND2X2_3695 ( .A(_abc_17692_n9196), .B(_abc_17692_n9189), .Y(_abc_17692_n9201) );
  AND2X2 AND2X2_3696 ( .A(_abc_17692_n9202), .B(_abc_17692_n1830_bF_buf0), .Y(_abc_17692_n9203) );
  AND2X2 AND2X2_3697 ( .A(_abc_17692_n9200), .B(_abc_17692_n9203), .Y(_abc_17692_n9204) );
  AND2X2 AND2X2_3698 ( .A(_abc_17692_n9204), .B(_abc_17692_n9198), .Y(_abc_17692_n9205) );
  AND2X2 AND2X2_3699 ( .A(_abc_17692_n3141_1), .B(_abc_17692_n9154), .Y(_abc_17692_n9208) );
  AND2X2 AND2X2_37 ( .A(_abc_17692_n711), .B(_abc_17692_n716), .Y(_abc_17692_n717) );
  AND2X2 AND2X2_370 ( .A(_abc_17692_n1525), .B(_abc_17692_n1526_1), .Y(_abc_17692_n1527) );
  AND2X2 AND2X2_3700 ( .A(_abc_17692_n3142), .B(_abc_17692_n9158), .Y(_abc_17692_n9209) );
  AND2X2 AND2X2_3701 ( .A(_abc_17692_n9211), .B(_abc_17692_n2063), .Y(_abc_17692_n9212) );
  AND2X2 AND2X2_3702 ( .A(_abc_17692_n9210), .B(workunit1_7_), .Y(_abc_17692_n9213) );
  AND2X2 AND2X2_3703 ( .A(_abc_17692_n9217), .B(_abc_17692_n9215), .Y(_abc_17692_n9219) );
  AND2X2 AND2X2_3704 ( .A(_abc_17692_n9220), .B(_abc_17692_n1863_bF_buf10), .Y(_abc_17692_n9221) );
  AND2X2 AND2X2_3705 ( .A(_abc_17692_n9221), .B(_abc_17692_n9218), .Y(_abc_17692_n9222) );
  AND2X2 AND2X2_3706 ( .A(_abc_17692_n9223), .B(state_10_bF_buf2), .Y(_abc_17692_n9224) );
  AND2X2 AND2X2_3707 ( .A(_abc_17692_n9099), .B(_abc_17692_n9225), .Y(_abc_17692_n9226) );
  AND2X2 AND2X2_3708 ( .A(_abc_17692_n9228), .B(_abc_17692_n9229), .Y(_abc_17692_n9230) );
  AND2X2 AND2X2_3709 ( .A(_abc_17692_n9232), .B(_abc_17692_n1830_bF_buf10), .Y(_abc_17692_n9233) );
  AND2X2 AND2X2_371 ( .A(_abc_17692_n1495), .B(_abc_17692_n1502), .Y(_abc_17692_n1530) );
  AND2X2 AND2X2_3710 ( .A(_abc_17692_n9233), .B(_abc_17692_n9227), .Y(_abc_17692_n9234) );
  AND2X2 AND2X2_3711 ( .A(_abc_17692_n9055), .B(workunit1_6_), .Y(_abc_17692_n9235) );
  AND2X2 AND2X2_3712 ( .A(_abc_17692_n9107), .B(_abc_17692_n9236), .Y(_abc_17692_n9237) );
  AND2X2 AND2X2_3713 ( .A(_abc_17692_n9240), .B(_abc_17692_n1846_bF_buf10), .Y(_abc_17692_n9241) );
  AND2X2 AND2X2_3714 ( .A(_abc_17692_n9241), .B(_abc_17692_n9239), .Y(_abc_17692_n9242) );
  AND2X2 AND2X2_3715 ( .A(_abc_17692_n9246), .B(_abc_17692_n9214), .Y(_abc_17692_n9248) );
  AND2X2 AND2X2_3716 ( .A(_abc_17692_n9249), .B(_abc_17692_n1863_bF_buf9), .Y(_abc_17692_n9250) );
  AND2X2 AND2X2_3717 ( .A(_abc_17692_n9250), .B(_abc_17692_n9247), .Y(_abc_17692_n9251) );
  AND2X2 AND2X2_3718 ( .A(_abc_17692_n9258), .B(_abc_17692_n1877_bF_buf10), .Y(_abc_17692_n9259) );
  AND2X2 AND2X2_3719 ( .A(_abc_17692_n9256), .B(_abc_17692_n9259), .Y(_abc_17692_n9260) );
  AND2X2 AND2X2_372 ( .A(_abc_17692_n1460), .B(_abc_17692_n1500), .Y(_abc_17692_n1533) );
  AND2X2 AND2X2_3720 ( .A(_abc_17692_n9260), .B(_abc_17692_n9255), .Y(_abc_17692_n9261) );
  AND2X2 AND2X2_3721 ( .A(_abc_17692_n9263), .B(state_14_bF_buf2), .Y(_abc_17692_n9264) );
  AND2X2 AND2X2_3722 ( .A(_abc_17692_n8383_bF_buf2), .B(workunit1_7_), .Y(_abc_17692_n9265) );
  AND2X2 AND2X2_3723 ( .A(state_8_bF_buf0), .B(\data_in1[7] ), .Y(_abc_17692_n9266) );
  AND2X2 AND2X2_3724 ( .A(_abc_17692_n9022), .B(_abc_17692_n9152), .Y(_abc_17692_n9270) );
  AND2X2 AND2X2_3725 ( .A(_abc_17692_n9015), .B(_abc_17692_n9270), .Y(_abc_17692_n9271) );
  AND2X2 AND2X2_3726 ( .A(_abc_17692_n9271), .B(_abc_17692_n8756), .Y(_abc_17692_n9272) );
  AND2X2 AND2X2_3727 ( .A(_abc_17692_n9018), .B(_abc_17692_n9270), .Y(_abc_17692_n9273) );
  AND2X2 AND2X2_3728 ( .A(_abc_17692_n9020), .B(_abc_17692_n9150), .Y(_abc_17692_n9274) );
  AND2X2 AND2X2_3729 ( .A(_abc_17692_n4351), .B(workunit2_4_), .Y(_abc_17692_n9279) );
  AND2X2 AND2X2_373 ( .A(_abc_17692_n1470), .B(_abc_17692_n1533), .Y(_abc_17692_n1534) );
  AND2X2 AND2X2_3730 ( .A(_abc_17692_n2482), .B(workunit2_13_), .Y(_abc_17692_n9280) );
  AND2X2 AND2X2_3731 ( .A(_abc_17692_n9281), .B(workunit2_8_bF_buf0), .Y(_abc_17692_n9282) );
  AND2X2 AND2X2_3732 ( .A(_abc_17692_n9283), .B(_abc_17692_n9284), .Y(_abc_17692_n9285) );
  AND2X2 AND2X2_3733 ( .A(_abc_17692_n9285), .B(_abc_17692_n3198), .Y(_abc_17692_n9286) );
  AND2X2 AND2X2_3734 ( .A(_abc_17692_n9278), .B(_abc_17692_n9288), .Y(_abc_17692_n9289) );
  AND2X2 AND2X2_3735 ( .A(_abc_17692_n9293), .B(_abc_17692_n9275), .Y(_abc_17692_n9294) );
  AND2X2 AND2X2_3736 ( .A(_abc_17692_n9292), .B(_abc_17692_n9294), .Y(_abc_17692_n9295) );
  AND2X2 AND2X2_3737 ( .A(_abc_17692_n9295), .B(_abc_17692_n9287), .Y(_abc_17692_n9296) );
  AND2X2 AND2X2_3738 ( .A(_abc_17692_n9300), .B(_abc_17692_n9299), .Y(_abc_17692_n9301) );
  AND2X2 AND2X2_3739 ( .A(_abc_17692_n9301), .B(workunit1_8_bF_buf2), .Y(_abc_17692_n9302) );
  AND2X2 AND2X2_374 ( .A(_abc_17692_n1535), .B(_abc_17692_n1529), .Y(_abc_17692_n1537) );
  AND2X2 AND2X2_3740 ( .A(_abc_17692_n9303), .B(_abc_17692_n9304), .Y(_abc_17692_n9305) );
  AND2X2 AND2X2_3741 ( .A(_abc_17692_n9309), .B(_abc_17692_n9310), .Y(_abc_17692_n9311) );
  AND2X2 AND2X2_3742 ( .A(_abc_17692_n9314), .B(_abc_17692_n9313), .Y(_abc_17692_n9315) );
  AND2X2 AND2X2_3743 ( .A(_abc_17692_n9316), .B(_abc_17692_n2250), .Y(_abc_17692_n9317) );
  AND2X2 AND2X2_3744 ( .A(_abc_17692_n9315), .B(workunit1_8_bF_buf0), .Y(_abc_17692_n9318) );
  AND2X2 AND2X2_3745 ( .A(_abc_17692_n9177), .B(workunit1_7_), .Y(_abc_17692_n9321) );
  AND2X2 AND2X2_3746 ( .A(_abc_17692_n9322), .B(_abc_17692_n9320), .Y(_abc_17692_n9324) );
  AND2X2 AND2X2_3747 ( .A(_abc_17692_n9325), .B(_abc_17692_n1877_bF_buf9), .Y(_abc_17692_n9326) );
  AND2X2 AND2X2_3748 ( .A(_abc_17692_n9326), .B(_abc_17692_n9323), .Y(_abc_17692_n9327) );
  AND2X2 AND2X2_3749 ( .A(_abc_17692_n9328), .B(_abc_17692_n9329), .Y(_abc_17692_n9330) );
  AND2X2 AND2X2_375 ( .A(_abc_17692_n1538_1), .B(state_3_bF_buf2), .Y(_abc_17692_n1539) );
  AND2X2 AND2X2_3750 ( .A(_abc_17692_n9330), .B(workunit1_8_bF_buf3), .Y(_abc_17692_n9331) );
  AND2X2 AND2X2_3751 ( .A(_abc_17692_n9332), .B(_abc_17692_n9333), .Y(_abc_17692_n9334) );
  AND2X2 AND2X2_3752 ( .A(_abc_17692_n9192), .B(workunit1_7_), .Y(_abc_17692_n9335) );
  AND2X2 AND2X2_3753 ( .A(_abc_17692_n9337), .B(_abc_17692_n9334), .Y(_abc_17692_n9339) );
  AND2X2 AND2X2_3754 ( .A(_abc_17692_n9340), .B(_abc_17692_n1830_bF_buf9), .Y(_abc_17692_n9341) );
  AND2X2 AND2X2_3755 ( .A(_abc_17692_n9341), .B(_abc_17692_n9338), .Y(_abc_17692_n9342) );
  AND2X2 AND2X2_3756 ( .A(_abc_17692_n9343), .B(_abc_17692_n9344), .Y(_abc_17692_n9345) );
  AND2X2 AND2X2_3757 ( .A(_abc_17692_n9345), .B(workunit1_8_bF_buf1), .Y(_abc_17692_n9346) );
  AND2X2 AND2X2_3758 ( .A(_abc_17692_n9347), .B(_abc_17692_n9348), .Y(_abc_17692_n9349) );
  AND2X2 AND2X2_3759 ( .A(_abc_17692_n9160), .B(workunit1_7_), .Y(_abc_17692_n9351) );
  AND2X2 AND2X2_376 ( .A(_abc_17692_n1539), .B(_abc_17692_n1536), .Y(_abc_17692_n1540) );
  AND2X2 AND2X2_3760 ( .A(_abc_17692_n9350), .B(_abc_17692_n9352), .Y(_abc_17692_n9353) );
  AND2X2 AND2X2_3761 ( .A(_abc_17692_n9355), .B(_abc_17692_n9353), .Y(_abc_17692_n9356) );
  AND2X2 AND2X2_3762 ( .A(_abc_17692_n9357), .B(_abc_17692_n9349), .Y(_abc_17692_n9359) );
  AND2X2 AND2X2_3763 ( .A(_abc_17692_n9360), .B(_abc_17692_n1846_bF_buf9), .Y(_abc_17692_n9361) );
  AND2X2 AND2X2_3764 ( .A(_abc_17692_n9361), .B(_abc_17692_n9358), .Y(_abc_17692_n9362) );
  AND2X2 AND2X2_3765 ( .A(_abc_17692_n9365), .B(state_10_bF_buf1), .Y(_abc_17692_n9366) );
  AND2X2 AND2X2_3766 ( .A(_abc_17692_n9366), .B(_abc_17692_n9312), .Y(_abc_17692_n9367) );
  AND2X2 AND2X2_3767 ( .A(_abc_17692_n9211), .B(workunit1_7_), .Y(_abc_17692_n9368) );
  AND2X2 AND2X2_3768 ( .A(_abc_17692_n9369), .B(_abc_17692_n9306), .Y(_abc_17692_n9371) );
  AND2X2 AND2X2_3769 ( .A(_abc_17692_n9372), .B(_abc_17692_n1863_bF_buf7), .Y(_abc_17692_n9373) );
  AND2X2 AND2X2_377 ( .A(_abc_17692_n1496), .B(sum_21_), .Y(_abc_17692_n1541) );
  AND2X2 AND2X2_3770 ( .A(_abc_17692_n9373), .B(_abc_17692_n9370), .Y(_abc_17692_n9374) );
  AND2X2 AND2X2_3771 ( .A(_abc_17692_n9258), .B(_abc_17692_n9375), .Y(_abc_17692_n9376) );
  AND2X2 AND2X2_3772 ( .A(_abc_17692_n9256), .B(_abc_17692_n9376), .Y(_abc_17692_n9377) );
  AND2X2 AND2X2_3773 ( .A(_abc_17692_n9378), .B(_abc_17692_n9319), .Y(_abc_17692_n9379) );
  AND2X2 AND2X2_3774 ( .A(_abc_17692_n9381), .B(_abc_17692_n1877_bF_buf8), .Y(_abc_17692_n9382) );
  AND2X2 AND2X2_3775 ( .A(_abc_17692_n9382), .B(_abc_17692_n9380), .Y(_abc_17692_n9383) );
  AND2X2 AND2X2_3776 ( .A(_abc_17692_n9166), .B(_abc_17692_n9235), .Y(_abc_17692_n9386) );
  AND2X2 AND2X2_3777 ( .A(_abc_17692_n9166), .B(_abc_17692_n9059), .Y(_abc_17692_n9388) );
  AND2X2 AND2X2_3778 ( .A(_abc_17692_n9104), .B(_abc_17692_n9388), .Y(_abc_17692_n9389) );
  AND2X2 AND2X2_3779 ( .A(_abc_17692_n9390), .B(_abc_17692_n9384), .Y(_abc_17692_n9392) );
  AND2X2 AND2X2_378 ( .A(_abc_17692_n1514), .B(_abc_17692_n1543), .Y(_abc_17692_n1544) );
  AND2X2 AND2X2_3780 ( .A(_abc_17692_n9393), .B(_abc_17692_n1846_bF_buf8), .Y(_abc_17692_n9394) );
  AND2X2 AND2X2_3781 ( .A(_abc_17692_n9394), .B(_abc_17692_n9391), .Y(_abc_17692_n9395) );
  AND2X2 AND2X2_3782 ( .A(_abc_17692_n9230), .B(_abc_17692_n9029), .Y(_abc_17692_n9397) );
  AND2X2 AND2X2_3783 ( .A(_abc_17692_n9400), .B(_abc_17692_n9097), .Y(_abc_17692_n9401) );
  AND2X2 AND2X2_3784 ( .A(_abc_17692_n9402), .B(_abc_17692_n9396), .Y(_abc_17692_n9403) );
  AND2X2 AND2X2_3785 ( .A(_abc_17692_n9405), .B(_abc_17692_n1830_bF_buf8), .Y(_abc_17692_n9406) );
  AND2X2 AND2X2_3786 ( .A(_abc_17692_n9406), .B(_abc_17692_n9404), .Y(_abc_17692_n9407) );
  AND2X2 AND2X2_3787 ( .A(_abc_17692_n9410), .B(state_14_bF_buf1), .Y(_abc_17692_n9411) );
  AND2X2 AND2X2_3788 ( .A(_abc_17692_n8383_bF_buf1), .B(workunit1_8_bF_buf3), .Y(_abc_17692_n9412) );
  AND2X2 AND2X2_3789 ( .A(state_8_bF_buf9), .B(\data_in1[8] ), .Y(_abc_17692_n9413) );
  AND2X2 AND2X2_379 ( .A(_abc_17692_n1545), .B(_abc_17692_n1528), .Y(_abc_17692_n1546) );
  AND2X2 AND2X2_3790 ( .A(_abc_17692_n9325), .B(_abc_17692_n9417), .Y(_abc_17692_n9418) );
  AND2X2 AND2X2_3791 ( .A(workunit2_5_), .B(workunit2_14_bF_buf1), .Y(_abc_17692_n9421) );
  AND2X2 AND2X2_3792 ( .A(_abc_17692_n9422), .B(_abc_17692_n9423), .Y(_abc_17692_n9424) );
  AND2X2 AND2X2_3793 ( .A(_abc_17692_n9424), .B(workunit2_9_), .Y(_abc_17692_n9425) );
  AND2X2 AND2X2_3794 ( .A(_abc_17692_n9427), .B(_abc_17692_n3471), .Y(_abc_17692_n9428) );
  AND2X2 AND2X2_3795 ( .A(_abc_17692_n9420), .B(_abc_17692_n9430), .Y(_abc_17692_n9431) );
  AND2X2 AND2X2_3796 ( .A(_abc_17692_n9419), .B(_abc_17692_n9429), .Y(_abc_17692_n9432) );
  AND2X2 AND2X2_3797 ( .A(_abc_17692_n9435), .B(_abc_17692_n9436), .Y(_abc_17692_n9437) );
  AND2X2 AND2X2_3798 ( .A(_abc_17692_n9437), .B(workunit1_9_), .Y(_abc_17692_n9438) );
  AND2X2 AND2X2_3799 ( .A(_abc_17692_n9439), .B(_abc_17692_n2435), .Y(_abc_17692_n9440) );
  AND2X2 AND2X2_38 ( .A(_abc_17692_n722_bF_buf3), .B(_abc_17692_n632), .Y(_abc_17692_n723) );
  AND2X2 AND2X2_380 ( .A(_abc_17692_n1548), .B(state_15_bF_buf2), .Y(_abc_17692_n1549) );
  AND2X2 AND2X2_3800 ( .A(_abc_17692_n9418), .B(_abc_17692_n9441), .Y(_abc_17692_n9442) );
  AND2X2 AND2X2_3801 ( .A(_abc_17692_n9443), .B(_abc_17692_n9444), .Y(_abc_17692_n9445) );
  AND2X2 AND2X2_3802 ( .A(_abc_17692_n9446), .B(_abc_17692_n1877_bF_buf7), .Y(_abc_17692_n9447) );
  AND2X2 AND2X2_3803 ( .A(_abc_17692_n9360), .B(_abc_17692_n9347), .Y(_abc_17692_n9448) );
  AND2X2 AND2X2_3804 ( .A(_abc_17692_n9450), .B(_abc_17692_n9451), .Y(_abc_17692_n9452) );
  AND2X2 AND2X2_3805 ( .A(_abc_17692_n9454), .B(_abc_17692_n9455), .Y(_abc_17692_n9456) );
  AND2X2 AND2X2_3806 ( .A(_abc_17692_n9453), .B(_abc_17692_n9457), .Y(_abc_17692_n9458) );
  AND2X2 AND2X2_3807 ( .A(_abc_17692_n9461), .B(_abc_17692_n1846_bF_buf7), .Y(_abc_17692_n9462) );
  AND2X2 AND2X2_3808 ( .A(_abc_17692_n9462), .B(_abc_17692_n9460), .Y(_abc_17692_n9463) );
  AND2X2 AND2X2_3809 ( .A(_abc_17692_n9340), .B(_abc_17692_n9332), .Y(_abc_17692_n9464) );
  AND2X2 AND2X2_381 ( .A(_abc_17692_n1549), .B(_abc_17692_n1547), .Y(_abc_17692_n1550_1) );
  AND2X2 AND2X2_3810 ( .A(_abc_17692_n9466), .B(_abc_17692_n9467), .Y(_abc_17692_n9468) );
  AND2X2 AND2X2_3811 ( .A(_abc_17692_n9468), .B(workunit1_9_), .Y(_abc_17692_n9469) );
  AND2X2 AND2X2_3812 ( .A(_abc_17692_n9470), .B(_abc_17692_n9471), .Y(_abc_17692_n9472) );
  AND2X2 AND2X2_3813 ( .A(_abc_17692_n9475), .B(_abc_17692_n1830_bF_buf7), .Y(_abc_17692_n9476) );
  AND2X2 AND2X2_3814 ( .A(_abc_17692_n9476), .B(_abc_17692_n9474), .Y(_abc_17692_n9477) );
  AND2X2 AND2X2_3815 ( .A(_abc_17692_n9309), .B(_abc_17692_n9303), .Y(_abc_17692_n9480) );
  AND2X2 AND2X2_3816 ( .A(_abc_17692_n9482), .B(_abc_17692_n9481), .Y(_abc_17692_n9483) );
  AND2X2 AND2X2_3817 ( .A(_abc_17692_n9483), .B(workunit1_9_), .Y(_abc_17692_n9484) );
  AND2X2 AND2X2_3818 ( .A(_abc_17692_n9486), .B(_abc_17692_n2435), .Y(_abc_17692_n9487) );
  AND2X2 AND2X2_3819 ( .A(_abc_17692_n9488), .B(_abc_17692_n9485), .Y(_abc_17692_n9489) );
  AND2X2 AND2X2_382 ( .A(_abc_17692_n722_bF_buf3), .B(sum_22_), .Y(_abc_17692_n1551) );
  AND2X2 AND2X2_3820 ( .A(_abc_17692_n9480), .B(_abc_17692_n9490), .Y(_abc_17692_n9491) );
  AND2X2 AND2X2_3821 ( .A(_abc_17692_n9492), .B(_abc_17692_n9489), .Y(_abc_17692_n9493) );
  AND2X2 AND2X2_3822 ( .A(_abc_17692_n9494), .B(_abc_17692_n1863_bF_buf6), .Y(_abc_17692_n9495) );
  AND2X2 AND2X2_3823 ( .A(_abc_17692_n9496), .B(state_10_bF_buf0), .Y(_abc_17692_n9497) );
  AND2X2 AND2X2_3824 ( .A(_abc_17692_n9498), .B(workunit1_8_bF_buf2), .Y(_abc_17692_n9499) );
  AND2X2 AND2X2_3825 ( .A(_abc_17692_n9372), .B(_abc_17692_n9500), .Y(_abc_17692_n9501) );
  AND2X2 AND2X2_3826 ( .A(_abc_17692_n9502), .B(_abc_17692_n9490), .Y(_abc_17692_n9503) );
  AND2X2 AND2X2_3827 ( .A(_abc_17692_n9501), .B(_abc_17692_n9489), .Y(_abc_17692_n9504) );
  AND2X2 AND2X2_3828 ( .A(_abc_17692_n9505), .B(_abc_17692_n1863_bF_buf5), .Y(_abc_17692_n9506) );
  AND2X2 AND2X2_3829 ( .A(_abc_17692_n9316), .B(workunit1_8_bF_buf1), .Y(_abc_17692_n9507) );
  AND2X2 AND2X2_383 ( .A(delta_23_), .B(sum_23_), .Y(_abc_17692_n1555) );
  AND2X2 AND2X2_3830 ( .A(_abc_17692_n9380), .B(_abc_17692_n9508), .Y(_abc_17692_n9509) );
  AND2X2 AND2X2_3831 ( .A(_abc_17692_n9512), .B(_abc_17692_n1877_bF_buf6), .Y(_abc_17692_n9513) );
  AND2X2 AND2X2_3832 ( .A(_abc_17692_n9513), .B(_abc_17692_n9511), .Y(_abc_17692_n9514) );
  AND2X2 AND2X2_3833 ( .A(_abc_17692_n9515), .B(workunit1_8_bF_buf0), .Y(_abc_17692_n9516) );
  AND2X2 AND2X2_3834 ( .A(_abc_17692_n9404), .B(_abc_17692_n9517), .Y(_abc_17692_n9518) );
  AND2X2 AND2X2_3835 ( .A(_abc_17692_n9521), .B(_abc_17692_n1830_bF_buf6), .Y(_abc_17692_n9522) );
  AND2X2 AND2X2_3836 ( .A(_abc_17692_n9522), .B(_abc_17692_n9519), .Y(_abc_17692_n9523) );
  AND2X2 AND2X2_3837 ( .A(_abc_17692_n9524), .B(workunit1_8_bF_buf3), .Y(_abc_17692_n9525) );
  AND2X2 AND2X2_3838 ( .A(_abc_17692_n9393), .B(_abc_17692_n9526), .Y(_abc_17692_n9527) );
  AND2X2 AND2X2_3839 ( .A(_abc_17692_n9530), .B(_abc_17692_n1846_bF_buf6), .Y(_abc_17692_n9531) );
  AND2X2 AND2X2_384 ( .A(_abc_17692_n1557), .B(_abc_17692_n1558), .Y(_abc_17692_n1559) );
  AND2X2 AND2X2_3840 ( .A(_abc_17692_n9531), .B(_abc_17692_n9529), .Y(_abc_17692_n9532) );
  AND2X2 AND2X2_3841 ( .A(_abc_17692_n9535), .B(state_14_bF_buf0), .Y(_abc_17692_n9536) );
  AND2X2 AND2X2_3842 ( .A(_abc_17692_n8383_bF_buf0), .B(workunit1_9_), .Y(_abc_17692_n9537) );
  AND2X2 AND2X2_3843 ( .A(state_8_bF_buf8), .B(\data_in1[9] ), .Y(_abc_17692_n9538) );
  AND2X2 AND2X2_3844 ( .A(_abc_17692_n9546), .B(_abc_17692_n9544), .Y(_abc_17692_n9547) );
  AND2X2 AND2X2_3845 ( .A(_abc_17692_n9543), .B(_abc_17692_n9547), .Y(_abc_17692_n9548) );
  AND2X2 AND2X2_3846 ( .A(_abc_17692_n4765), .B(workunit2_6_), .Y(_abc_17692_n9549) );
  AND2X2 AND2X2_3847 ( .A(_abc_17692_n2862), .B(workunit2_15_), .Y(_abc_17692_n9550) );
  AND2X2 AND2X2_3848 ( .A(_abc_17692_n9551), .B(workunit2_10_bF_buf1), .Y(_abc_17692_n9552) );
  AND2X2 AND2X2_3849 ( .A(_abc_17692_n9553), .B(_abc_17692_n9554), .Y(_abc_17692_n9555) );
  AND2X2 AND2X2_385 ( .A(_abc_17692_n1560), .B(_abc_17692_n1556), .Y(_abc_17692_n1561) );
  AND2X2 AND2X2_3850 ( .A(_abc_17692_n9555), .B(_abc_17692_n3751), .Y(_abc_17692_n9556) );
  AND2X2 AND2X2_3851 ( .A(_abc_17692_n9548), .B(_abc_17692_n9557), .Y(_abc_17692_n9558) );
  AND2X2 AND2X2_3852 ( .A(_abc_17692_n9278), .B(_abc_17692_n9559), .Y(_abc_17692_n9560) );
  AND2X2 AND2X2_3853 ( .A(_abc_17692_n9562), .B(_abc_17692_n9561), .Y(_abc_17692_n9563) );
  AND2X2 AND2X2_3854 ( .A(_abc_17692_n9566), .B(_abc_17692_n9565), .Y(_abc_17692_n9567) );
  AND2X2 AND2X2_3855 ( .A(_abc_17692_n9564), .B(_abc_17692_n9567), .Y(_abc_17692_n9568) );
  AND2X2 AND2X2_3856 ( .A(_abc_17692_n3768), .B(_abc_17692_n9569), .Y(_abc_17692_n9570) );
  AND2X2 AND2X2_3857 ( .A(_abc_17692_n3767), .B(_abc_17692_n9571), .Y(_abc_17692_n9572) );
  AND2X2 AND2X2_3858 ( .A(_abc_17692_n9575), .B(_abc_17692_n9576), .Y(_abc_17692_n9577) );
  AND2X2 AND2X2_3859 ( .A(_abc_17692_n9486), .B(workunit1_9_), .Y(_abc_17692_n9579) );
  AND2X2 AND2X2_386 ( .A(_abc_17692_n1566), .B(state_3_bF_buf1), .Y(_abc_17692_n1567) );
  AND2X2 AND2X2_3860 ( .A(_abc_17692_n9490), .B(_abc_17692_n9302), .Y(_abc_17692_n9580) );
  AND2X2 AND2X2_3861 ( .A(_abc_17692_n9490), .B(_abc_17692_n9305), .Y(_abc_17692_n9583) );
  AND2X2 AND2X2_3862 ( .A(_abc_17692_n9307), .B(_abc_17692_n9583), .Y(_abc_17692_n9584) );
  AND2X2 AND2X2_3863 ( .A(_abc_17692_n9585), .B(_abc_17692_n9582), .Y(_abc_17692_n9586) );
  AND2X2 AND2X2_3864 ( .A(_abc_17692_n9587), .B(_abc_17692_n9578), .Y(_abc_17692_n9588) );
  AND2X2 AND2X2_3865 ( .A(_abc_17692_n9589), .B(_abc_17692_n9590), .Y(_abc_17692_n9591) );
  AND2X2 AND2X2_3866 ( .A(_abc_17692_n9594), .B(_abc_17692_n9593), .Y(_abc_17692_n9595) );
  AND2X2 AND2X2_3867 ( .A(_abc_17692_n9595), .B(workunit1_10_), .Y(_abc_17692_n9596) );
  AND2X2 AND2X2_3868 ( .A(_abc_17692_n9597), .B(_abc_17692_n2638), .Y(_abc_17692_n9598) );
  AND2X2 AND2X2_3869 ( .A(_abc_17692_n9441), .B(_abc_17692_n9320), .Y(_abc_17692_n9601) );
  AND2X2 AND2X2_387 ( .A(_abc_17692_n1567), .B(_abc_17692_n1565), .Y(_abc_17692_n1568) );
  AND2X2 AND2X2_3870 ( .A(_abc_17692_n9322), .B(_abc_17692_n9601), .Y(_abc_17692_n9602) );
  AND2X2 AND2X2_3871 ( .A(_abc_17692_n9439), .B(workunit1_9_), .Y(_abc_17692_n9603) );
  AND2X2 AND2X2_3872 ( .A(_abc_17692_n9441), .B(_abc_17692_n9318), .Y(_abc_17692_n9604) );
  AND2X2 AND2X2_3873 ( .A(_abc_17692_n9606), .B(_abc_17692_n9600), .Y(_abc_17692_n9607) );
  AND2X2 AND2X2_3874 ( .A(_abc_17692_n9609), .B(_abc_17692_n1877_bF_buf5), .Y(_abc_17692_n9610) );
  AND2X2 AND2X2_3875 ( .A(_abc_17692_n9610), .B(_abc_17692_n9608), .Y(_abc_17692_n9611) );
  AND2X2 AND2X2_3876 ( .A(_abc_17692_n3727), .B(_abc_17692_n9569), .Y(_abc_17692_n9612) );
  AND2X2 AND2X2_3877 ( .A(_abc_17692_n9571), .B(_abc_17692_n3726), .Y(_abc_17692_n9613) );
  AND2X2 AND2X2_3878 ( .A(_abc_17692_n9616), .B(_abc_17692_n9617), .Y(_abc_17692_n9618) );
  AND2X2 AND2X2_3879 ( .A(_abc_17692_n9473), .B(_abc_17692_n9334), .Y(_abc_17692_n9621) );
  AND2X2 AND2X2_388 ( .A(_abc_17692_n1525), .B(sum_22_), .Y(_abc_17692_n1569) );
  AND2X2 AND2X2_3880 ( .A(_abc_17692_n9624), .B(workunit1_9_), .Y(_abc_17692_n9625) );
  AND2X2 AND2X2_3881 ( .A(_abc_17692_n9473), .B(_abc_17692_n9331), .Y(_abc_17692_n9626) );
  AND2X2 AND2X2_3882 ( .A(_abc_17692_n9623), .B(_abc_17692_n9628), .Y(_abc_17692_n9629) );
  AND2X2 AND2X2_3883 ( .A(_abc_17692_n9630), .B(_abc_17692_n9619), .Y(_abc_17692_n9631) );
  AND2X2 AND2X2_3884 ( .A(_abc_17692_n9633), .B(_abc_17692_n1830_bF_buf5), .Y(_abc_17692_n9634) );
  AND2X2 AND2X2_3885 ( .A(_abc_17692_n9634), .B(_abc_17692_n9632), .Y(_abc_17692_n9635) );
  AND2X2 AND2X2_3886 ( .A(_abc_17692_n3692), .B(_abc_17692_n9569), .Y(_abc_17692_n9636) );
  AND2X2 AND2X2_3887 ( .A(_abc_17692_n9571), .B(_abc_17692_n3690), .Y(_abc_17692_n9637) );
  AND2X2 AND2X2_3888 ( .A(_abc_17692_n9640), .B(_abc_17692_n9641), .Y(_abc_17692_n9642) );
  AND2X2 AND2X2_3889 ( .A(_abc_17692_n9452), .B(workunit1_9_), .Y(_abc_17692_n9646) );
  AND2X2 AND2X2_389 ( .A(_abc_17692_n1547), .B(_abc_17692_n1570), .Y(_abc_17692_n1571) );
  AND2X2 AND2X2_3890 ( .A(_abc_17692_n9648), .B(_abc_17692_n9647), .Y(_abc_17692_n9649) );
  AND2X2 AND2X2_3891 ( .A(_abc_17692_n9645), .B(_abc_17692_n9649), .Y(_abc_17692_n9650) );
  AND2X2 AND2X2_3892 ( .A(_abc_17692_n9651), .B(_abc_17692_n9643), .Y(_abc_17692_n9652) );
  AND2X2 AND2X2_3893 ( .A(_abc_17692_n9654), .B(_abc_17692_n1846_bF_buf5), .Y(_abc_17692_n9655) );
  AND2X2 AND2X2_3894 ( .A(_abc_17692_n9655), .B(_abc_17692_n9653), .Y(_abc_17692_n9656) );
  AND2X2 AND2X2_3895 ( .A(_abc_17692_n9659), .B(state_10_bF_buf4), .Y(_abc_17692_n9660) );
  AND2X2 AND2X2_3896 ( .A(_abc_17692_n9660), .B(_abc_17692_n9592), .Y(_abc_17692_n9661) );
  AND2X2 AND2X2_3897 ( .A(_abc_17692_n9489), .B(_abc_17692_n9306), .Y(_abc_17692_n9662) );
  AND2X2 AND2X2_3898 ( .A(_abc_17692_n9369), .B(_abc_17692_n9662), .Y(_abc_17692_n9663) );
  AND2X2 AND2X2_3899 ( .A(_abc_17692_n9488), .B(_abc_17692_n9664), .Y(_abc_17692_n9665) );
  AND2X2 AND2X2_39 ( .A(_abc_17692_n720), .B(_abc_17692_n723), .Y(_abc_17692_n724) );
  AND2X2 AND2X2_390 ( .A(_abc_17692_n1574), .B(state_15_bF_buf1), .Y(_abc_17692_n1575) );
  AND2X2 AND2X2_3900 ( .A(_abc_17692_n9666), .B(_abc_17692_n9577), .Y(_abc_17692_n9668) );
  AND2X2 AND2X2_3901 ( .A(_abc_17692_n9669), .B(_abc_17692_n1863_bF_buf3), .Y(_abc_17692_n9670) );
  AND2X2 AND2X2_3902 ( .A(_abc_17692_n9670), .B(_abc_17692_n9667), .Y(_abc_17692_n9671) );
  AND2X2 AND2X2_3903 ( .A(_abc_17692_n9444), .B(_abc_17692_n9319), .Y(_abc_17692_n9672) );
  AND2X2 AND2X2_3904 ( .A(_abc_17692_n9676), .B(_abc_17692_n9675), .Y(_abc_17692_n9677) );
  AND2X2 AND2X2_3905 ( .A(_abc_17692_n9674), .B(_abc_17692_n9677), .Y(_abc_17692_n9678) );
  AND2X2 AND2X2_3906 ( .A(_abc_17692_n9679), .B(_abc_17692_n9599), .Y(_abc_17692_n9680) );
  AND2X2 AND2X2_3907 ( .A(_abc_17692_n9682), .B(_abc_17692_n1877_bF_buf4), .Y(_abc_17692_n9683) );
  AND2X2 AND2X2_3908 ( .A(_abc_17692_n9683), .B(_abc_17692_n9681), .Y(_abc_17692_n9684) );
  AND2X2 AND2X2_3909 ( .A(_abc_17692_n9458), .B(_abc_17692_n9384), .Y(_abc_17692_n9685) );
  AND2X2 AND2X2_391 ( .A(_abc_17692_n1575), .B(_abc_17692_n1572), .Y(_abc_17692_n1576) );
  AND2X2 AND2X2_3910 ( .A(_abc_17692_n9390), .B(_abc_17692_n9685), .Y(_abc_17692_n9686) );
  AND2X2 AND2X2_3911 ( .A(_abc_17692_n9688), .B(_abc_17692_n9457), .Y(_abc_17692_n9689) );
  AND2X2 AND2X2_3912 ( .A(_abc_17692_n9690), .B(_abc_17692_n9642), .Y(_abc_17692_n9692) );
  AND2X2 AND2X2_3913 ( .A(_abc_17692_n9693), .B(_abc_17692_n1846_bF_buf4), .Y(_abc_17692_n9694) );
  AND2X2 AND2X2_3914 ( .A(_abc_17692_n9694), .B(_abc_17692_n9691), .Y(_abc_17692_n9695) );
  AND2X2 AND2X2_3915 ( .A(_abc_17692_n9472), .B(_abc_17692_n9396), .Y(_abc_17692_n9696) );
  AND2X2 AND2X2_3916 ( .A(_abc_17692_n9402), .B(_abc_17692_n9696), .Y(_abc_17692_n9697) );
  AND2X2 AND2X2_3917 ( .A(_abc_17692_n9698), .B(_abc_17692_n9471), .Y(_abc_17692_n9699) );
  AND2X2 AND2X2_3918 ( .A(_abc_17692_n9700), .B(_abc_17692_n9618), .Y(_abc_17692_n9701) );
  AND2X2 AND2X2_3919 ( .A(_abc_17692_n9703), .B(_abc_17692_n1830_bF_buf4), .Y(_abc_17692_n9704) );
  AND2X2 AND2X2_392 ( .A(_abc_17692_n722_bF_buf2), .B(sum_23_), .Y(_abc_17692_n1577) );
  AND2X2 AND2X2_3920 ( .A(_abc_17692_n9704), .B(_abc_17692_n9702), .Y(_abc_17692_n9705) );
  AND2X2 AND2X2_3921 ( .A(_abc_17692_n9708), .B(state_14_bF_buf4), .Y(_abc_17692_n9709) );
  AND2X2 AND2X2_3922 ( .A(_abc_17692_n8383_bF_buf4), .B(workunit1_10_), .Y(_abc_17692_n9710) );
  AND2X2 AND2X2_3923 ( .A(state_8_bF_buf7), .B(\data_in1[10] ), .Y(_abc_17692_n9711) );
  AND2X2 AND2X2_3924 ( .A(_abc_17692_n9716), .B(_abc_17692_n9718), .Y(_abc_17692_n9719) );
  AND2X2 AND2X2_3925 ( .A(_abc_17692_n9717), .B(workunit2_7_), .Y(_abc_17692_n9721) );
  AND2X2 AND2X2_3926 ( .A(_abc_17692_n3060), .B(workunit2_16_bF_buf3), .Y(_abc_17692_n9722) );
  AND2X2 AND2X2_3927 ( .A(_abc_17692_n9724), .B(_abc_17692_n9720), .Y(_abc_17692_n9725) );
  AND2X2 AND2X2_3928 ( .A(_abc_17692_n9727), .B(_abc_17692_n9565), .Y(_abc_17692_n9728) );
  AND2X2 AND2X2_3929 ( .A(_abc_17692_n9723), .B(workunit2_11_), .Y(_abc_17692_n9729) );
  AND2X2 AND2X2_393 ( .A(_abc_17692_n1581), .B(delta_24_), .Y(_abc_17692_n1582) );
  AND2X2 AND2X2_3930 ( .A(_abc_17692_n9719), .B(_abc_17692_n3905), .Y(_abc_17692_n9730) );
  AND2X2 AND2X2_3931 ( .A(_abc_17692_n9732), .B(_abc_17692_n9726), .Y(_abc_17692_n9733) );
  AND2X2 AND2X2_3932 ( .A(_abc_17692_n9728), .B(_abc_17692_n9731), .Y(_abc_17692_n9735) );
  AND2X2 AND2X2_3933 ( .A(_abc_17692_n9715), .B(_abc_17692_n9725), .Y(_abc_17692_n9736) );
  AND2X2 AND2X2_3934 ( .A(_abc_17692_n9738), .B(_abc_17692_n9734), .Y(_abc_17692_n9739) );
  AND2X2 AND2X2_3935 ( .A(_abc_17692_n9739), .B(_abc_17692_n2823), .Y(_abc_17692_n9740) );
  AND2X2 AND2X2_3936 ( .A(_abc_17692_n3896), .B(_abc_17692_n9737), .Y(_abc_17692_n9742) );
  AND2X2 AND2X2_3937 ( .A(_abc_17692_n3901), .B(_abc_17692_n9733), .Y(_abc_17692_n9743) );
  AND2X2 AND2X2_3938 ( .A(_abc_17692_n9744), .B(workunit1_11_bF_buf0), .Y(_abc_17692_n9745) );
  AND2X2 AND2X2_3939 ( .A(_abc_17692_n9741), .B(_abc_17692_n9746), .Y(_abc_17692_n9747) );
  AND2X2 AND2X2_394 ( .A(_abc_17692_n1529), .B(_abc_17692_n1561), .Y(_abc_17692_n1586) );
  AND2X2 AND2X2_3940 ( .A(_abc_17692_n9608), .B(_abc_17692_n9749), .Y(_abc_17692_n9750) );
  AND2X2 AND2X2_3941 ( .A(_abc_17692_n9753), .B(_abc_17692_n1877_bF_buf3), .Y(_abc_17692_n9754) );
  AND2X2 AND2X2_3942 ( .A(_abc_17692_n9754), .B(_abc_17692_n9751), .Y(_abc_17692_n9755) );
  AND2X2 AND2X2_3943 ( .A(_abc_17692_n9756), .B(_abc_17692_n9757), .Y(_abc_17692_n9758) );
  AND2X2 AND2X2_3944 ( .A(_abc_17692_n9760), .B(_abc_17692_n9761), .Y(_abc_17692_n9762) );
  AND2X2 AND2X2_3945 ( .A(_abc_17692_n9759), .B(_abc_17692_n9763), .Y(_abc_17692_n9764) );
  AND2X2 AND2X2_3946 ( .A(_abc_17692_n9639), .B(workunit1_10_), .Y(_abc_17692_n9766) );
  AND2X2 AND2X2_3947 ( .A(_abc_17692_n9653), .B(_abc_17692_n9767), .Y(_abc_17692_n9768) );
  AND2X2 AND2X2_3948 ( .A(_abc_17692_n9771), .B(_abc_17692_n1846_bF_buf3), .Y(_abc_17692_n9772) );
  AND2X2 AND2X2_3949 ( .A(_abc_17692_n9772), .B(_abc_17692_n9770), .Y(_abc_17692_n9773) );
  AND2X2 AND2X2_395 ( .A(_abc_17692_n1533), .B(_abc_17692_n1586), .Y(_abc_17692_n1587) );
  AND2X2 AND2X2_3950 ( .A(_abc_17692_n9775), .B(_abc_17692_n9774), .Y(_abc_17692_n9776) );
  AND2X2 AND2X2_3951 ( .A(_abc_17692_n9776), .B(workunit1_11_bF_buf2), .Y(_abc_17692_n9777) );
  AND2X2 AND2X2_3952 ( .A(_abc_17692_n3961), .B(_abc_17692_n9737), .Y(_abc_17692_n9778) );
  AND2X2 AND2X2_3953 ( .A(_abc_17692_n3959), .B(_abc_17692_n9733), .Y(_abc_17692_n9779) );
  AND2X2 AND2X2_3954 ( .A(_abc_17692_n9780), .B(_abc_17692_n2823), .Y(_abc_17692_n9781) );
  AND2X2 AND2X2_3955 ( .A(_abc_17692_n9615), .B(workunit1_10_), .Y(_abc_17692_n9783) );
  AND2X2 AND2X2_3956 ( .A(_abc_17692_n9632), .B(_abc_17692_n9784), .Y(_abc_17692_n9785) );
  AND2X2 AND2X2_3957 ( .A(_abc_17692_n9788), .B(_abc_17692_n9789), .Y(_abc_17692_n9790) );
  AND2X2 AND2X2_3958 ( .A(_abc_17692_n9791), .B(_abc_17692_n1830_bF_buf3), .Y(_abc_17692_n9792) );
  AND2X2 AND2X2_3959 ( .A(_abc_17692_n9792), .B(_abc_17692_n9787), .Y(_abc_17692_n9793) );
  AND2X2 AND2X2_396 ( .A(_abc_17692_n1532), .B(_abc_17692_n1586), .Y(_abc_17692_n1590) );
  AND2X2 AND2X2_3960 ( .A(_abc_17692_n9796), .B(_abc_17692_n9797), .Y(_abc_17692_n9798) );
  AND2X2 AND2X2_3961 ( .A(_abc_17692_n9800), .B(_abc_17692_n9801), .Y(_abc_17692_n9802) );
  AND2X2 AND2X2_3962 ( .A(_abc_17692_n9799), .B(_abc_17692_n9803), .Y(_abc_17692_n9804) );
  AND2X2 AND2X2_3963 ( .A(_abc_17692_n9574), .B(workunit1_10_), .Y(_abc_17692_n9806) );
  AND2X2 AND2X2_3964 ( .A(_abc_17692_n9589), .B(_abc_17692_n9807), .Y(_abc_17692_n9808) );
  AND2X2 AND2X2_3965 ( .A(_abc_17692_n9808), .B(_abc_17692_n9805), .Y(_abc_17692_n9809) );
  AND2X2 AND2X2_3966 ( .A(_abc_17692_n9810), .B(_abc_17692_n9804), .Y(_abc_17692_n9811) );
  AND2X2 AND2X2_3967 ( .A(_abc_17692_n9812), .B(_abc_17692_n1863_bF_buf2), .Y(_abc_17692_n9813) );
  AND2X2 AND2X2_3968 ( .A(_abc_17692_n9814), .B(state_10_bF_buf3), .Y(_abc_17692_n9815) );
  AND2X2 AND2X2_3969 ( .A(_abc_17692_n9669), .B(_abc_17692_n9575), .Y(_abc_17692_n9816) );
  AND2X2 AND2X2_397 ( .A(_abc_17692_n1560), .B(_abc_17692_n1524), .Y(_abc_17692_n1591) );
  AND2X2 AND2X2_3970 ( .A(_abc_17692_n9817), .B(_abc_17692_n9805), .Y(_abc_17692_n9818) );
  AND2X2 AND2X2_3971 ( .A(_abc_17692_n9816), .B(_abc_17692_n9804), .Y(_abc_17692_n9819) );
  AND2X2 AND2X2_3972 ( .A(_abc_17692_n9820), .B(_abc_17692_n1863_bF_buf1), .Y(_abc_17692_n9821) );
  AND2X2 AND2X2_3973 ( .A(_abc_17692_n9597), .B(workunit1_10_), .Y(_abc_17692_n9822) );
  AND2X2 AND2X2_3974 ( .A(_abc_17692_n9681), .B(_abc_17692_n9823), .Y(_abc_17692_n9824) );
  AND2X2 AND2X2_3975 ( .A(_abc_17692_n9827), .B(_abc_17692_n1877_bF_buf2), .Y(_abc_17692_n9828) );
  AND2X2 AND2X2_3976 ( .A(_abc_17692_n9828), .B(_abc_17692_n9826), .Y(_abc_17692_n9829) );
  AND2X2 AND2X2_3977 ( .A(_abc_17692_n9693), .B(_abc_17692_n9640), .Y(_abc_17692_n9830) );
  AND2X2 AND2X2_3978 ( .A(_abc_17692_n9833), .B(_abc_17692_n1846_bF_buf2), .Y(_abc_17692_n9834) );
  AND2X2 AND2X2_3979 ( .A(_abc_17692_n9834), .B(_abc_17692_n9832), .Y(_abc_17692_n9835) );
  AND2X2 AND2X2_398 ( .A(_abc_17692_n1589), .B(_abc_17692_n1594), .Y(_abc_17692_n1595_1) );
  AND2X2 AND2X2_3980 ( .A(_abc_17692_n9702), .B(_abc_17692_n9616), .Y(_abc_17692_n9836) );
  AND2X2 AND2X2_3981 ( .A(_abc_17692_n9839), .B(_abc_17692_n1830_bF_buf2), .Y(_abc_17692_n9840) );
  AND2X2 AND2X2_3982 ( .A(_abc_17692_n9840), .B(_abc_17692_n9838), .Y(_abc_17692_n9841) );
  AND2X2 AND2X2_3983 ( .A(_abc_17692_n9844), .B(state_14_bF_buf3), .Y(_abc_17692_n9845) );
  AND2X2 AND2X2_3984 ( .A(_abc_17692_n8383_bF_buf3), .B(workunit1_11_bF_buf3), .Y(_abc_17692_n9846) );
  AND2X2 AND2X2_3985 ( .A(state_8_bF_buf6), .B(\data_in1[11] ), .Y(_abc_17692_n9847) );
  AND2X2 AND2X2_3986 ( .A(_abc_17692_n9567), .B(_abc_17692_n9725), .Y(_abc_17692_n9851) );
  AND2X2 AND2X2_3987 ( .A(_abc_17692_n9851), .B(_abc_17692_n9563), .Y(_abc_17692_n9852) );
  AND2X2 AND2X2_3988 ( .A(_abc_17692_n9565), .B(_abc_17692_n9720), .Y(_abc_17692_n9853) );
  AND2X2 AND2X2_3989 ( .A(_abc_17692_n9278), .B(_abc_17692_n9859), .Y(_abc_17692_n9860) );
  AND2X2 AND2X2_399 ( .A(_abc_17692_n1596), .B(_abc_17692_n1595_1), .Y(_abc_17692_n1597) );
  AND2X2 AND2X2_3990 ( .A(_abc_17692_n5260), .B(workunit2_8_bF_buf3), .Y(_abc_17692_n9862) );
  AND2X2 AND2X2_3991 ( .A(_abc_17692_n3198), .B(workunit2_17_), .Y(_abc_17692_n9863) );
  AND2X2 AND2X2_3992 ( .A(_abc_17692_n9864), .B(workunit2_12_bF_buf2), .Y(_abc_17692_n9865) );
  AND2X2 AND2X2_3993 ( .A(_abc_17692_n9866), .B(_abc_17692_n9867), .Y(_abc_17692_n9868) );
  AND2X2 AND2X2_3994 ( .A(_abc_17692_n9861), .B(_abc_17692_n9868), .Y(_abc_17692_n9869) );
  AND2X2 AND2X2_3995 ( .A(_abc_17692_n9870), .B(_abc_17692_n9854), .Y(_abc_17692_n9871) );
  AND2X2 AND2X2_3996 ( .A(_abc_17692_n9872), .B(_abc_17692_n9871), .Y(_abc_17692_n9873) );
  AND2X2 AND2X2_3997 ( .A(_abc_17692_n9873), .B(_abc_17692_n9875), .Y(_abc_17692_n9876) );
  AND2X2 AND2X2_3998 ( .A(_abc_17692_n9880), .B(_abc_17692_n9879), .Y(_abc_17692_n9881) );
  AND2X2 AND2X2_3999 ( .A(_abc_17692_n9882), .B(_abc_17692_n3026), .Y(_abc_17692_n9883) );
  AND2X2 AND2X2_4 ( .A(_abc_17692_n632), .B(delta_1_), .Y(delta_1__FF_INPUT) );
  AND2X2 AND2X2_40 ( .A(_abc_17692_n717), .B(_abc_17692_n724), .Y(_abc_17692_n725) );
  AND2X2 AND2X2_400 ( .A(_abc_17692_n1598_1), .B(_abc_17692_n1585), .Y(_abc_17692_n1600) );
  AND2X2 AND2X2_4000 ( .A(_abc_17692_n9881), .B(workunit1_12_bF_buf0), .Y(_abc_17692_n9884) );
  AND2X2 AND2X2_4001 ( .A(_abc_17692_n9747), .B(_abc_17692_n9600), .Y(_abc_17692_n9886) );
  AND2X2 AND2X2_4002 ( .A(_abc_17692_n9886), .B(_abc_17692_n9601), .Y(_abc_17692_n9887) );
  AND2X2 AND2X2_4003 ( .A(_abc_17692_n9322), .B(_abc_17692_n9887), .Y(_abc_17692_n9888) );
  AND2X2 AND2X2_4004 ( .A(_abc_17692_n9746), .B(_abc_17692_n9749), .Y(_abc_17692_n9889) );
  AND2X2 AND2X2_4005 ( .A(_abc_17692_n9886), .B(_abc_17692_n9605), .Y(_abc_17692_n9892) );
  AND2X2 AND2X2_4006 ( .A(_abc_17692_n9895), .B(_abc_17692_n9885), .Y(_abc_17692_n9896) );
  AND2X2 AND2X2_4007 ( .A(_abc_17692_n9894), .B(_abc_17692_n9898), .Y(_abc_17692_n9899) );
  AND2X2 AND2X2_4008 ( .A(_abc_17692_n9902), .B(_abc_17692_n9903), .Y(_abc_17692_n9904) );
  AND2X2 AND2X2_4009 ( .A(_abc_17692_n9904), .B(workunit1_12_bF_buf3), .Y(_abc_17692_n9905) );
  AND2X2 AND2X2_401 ( .A(_abc_17692_n1601), .B(state_3_bF_buf0), .Y(_abc_17692_n1602) );
  AND2X2 AND2X2_4010 ( .A(_abc_17692_n9906), .B(_abc_17692_n9907), .Y(_abc_17692_n9908) );
  AND2X2 AND2X2_4011 ( .A(_abc_17692_n9758), .B(workunit1_11_bF_buf2), .Y(_abc_17692_n9912) );
  AND2X2 AND2X2_4012 ( .A(_abc_17692_n9914), .B(_abc_17692_n9913), .Y(_abc_17692_n9915) );
  AND2X2 AND2X2_4013 ( .A(_abc_17692_n9911), .B(_abc_17692_n9915), .Y(_abc_17692_n9916) );
  AND2X2 AND2X2_4014 ( .A(_abc_17692_n9910), .B(_abc_17692_n9916), .Y(_abc_17692_n9917) );
  AND2X2 AND2X2_4015 ( .A(_abc_17692_n9918), .B(_abc_17692_n9908), .Y(_abc_17692_n9919) );
  AND2X2 AND2X2_4016 ( .A(_abc_17692_n9917), .B(_abc_17692_n9921), .Y(_abc_17692_n9922) );
  AND2X2 AND2X2_4017 ( .A(_abc_17692_n9926), .B(_abc_17692_n9925), .Y(_abc_17692_n9927) );
  AND2X2 AND2X2_4018 ( .A(_abc_17692_n9927), .B(workunit1_12_bF_buf1), .Y(_abc_17692_n9928) );
  AND2X2 AND2X2_4019 ( .A(_abc_17692_n9929), .B(_abc_17692_n9930), .Y(_abc_17692_n9931) );
  AND2X2 AND2X2_402 ( .A(_abc_17692_n1602), .B(_abc_17692_n1599), .Y(_abc_17692_n1603) );
  AND2X2 AND2X2_4020 ( .A(_abc_17692_n9782), .B(_abc_17692_n9619), .Y(_abc_17692_n9933) );
  AND2X2 AND2X2_4021 ( .A(_abc_17692_n9933), .B(_abc_17692_n9621), .Y(_abc_17692_n9934) );
  AND2X2 AND2X2_4022 ( .A(_abc_17692_n9337), .B(_abc_17692_n9934), .Y(_abc_17692_n9935) );
  AND2X2 AND2X2_4023 ( .A(_abc_17692_n9627), .B(_abc_17692_n9933), .Y(_abc_17692_n9936) );
  AND2X2 AND2X2_4024 ( .A(_abc_17692_n9782), .B(_abc_17692_n9783), .Y(_abc_17692_n9937) );
  AND2X2 AND2X2_4025 ( .A(_abc_17692_n9780), .B(workunit1_11_bF_buf1), .Y(_abc_17692_n9938) );
  AND2X2 AND2X2_4026 ( .A(_abc_17692_n9942), .B(_abc_17692_n9932), .Y(_abc_17692_n9943) );
  AND2X2 AND2X2_4027 ( .A(_abc_17692_n9941), .B(_abc_17692_n9931), .Y(_abc_17692_n9945) );
  AND2X2 AND2X2_4028 ( .A(_abc_17692_n9947), .B(_abc_17692_n9924), .Y(_abc_17692_n9948) );
  AND2X2 AND2X2_4029 ( .A(_abc_17692_n9948), .B(_abc_17692_n9901), .Y(_abc_17692_n9949) );
  AND2X2 AND2X2_403 ( .A(_abc_17692_n723), .B(sum_24_), .Y(_abc_17692_n1604) );
  AND2X2 AND2X2_4030 ( .A(_abc_17692_n9951), .B(_abc_17692_n9950), .Y(_abc_17692_n9952) );
  AND2X2 AND2X2_4031 ( .A(_abc_17692_n9952), .B(workunit1_12_bF_buf3), .Y(_abc_17692_n9953) );
  AND2X2 AND2X2_4032 ( .A(_abc_17692_n9954), .B(_abc_17692_n9955), .Y(_abc_17692_n9956) );
  AND2X2 AND2X2_4033 ( .A(_abc_17692_n9805), .B(_abc_17692_n9578), .Y(_abc_17692_n9958) );
  AND2X2 AND2X2_4034 ( .A(_abc_17692_n9584), .B(_abc_17692_n9958), .Y(_abc_17692_n9959) );
  AND2X2 AND2X2_4035 ( .A(_abc_17692_n9581), .B(_abc_17692_n9958), .Y(_abc_17692_n9960) );
  AND2X2 AND2X2_4036 ( .A(_abc_17692_n9805), .B(_abc_17692_n9806), .Y(_abc_17692_n9961) );
  AND2X2 AND2X2_4037 ( .A(_abc_17692_n9798), .B(workunit1_11_bF_buf0), .Y(_abc_17692_n9962) );
  AND2X2 AND2X2_4038 ( .A(_abc_17692_n9966), .B(_abc_17692_n9957), .Y(_abc_17692_n9967) );
  AND2X2 AND2X2_4039 ( .A(_abc_17692_n9965), .B(_abc_17692_n9956), .Y(_abc_17692_n9968) );
  AND2X2 AND2X2_404 ( .A(_abc_17692_n1562_1), .B(_abc_17692_n1528), .Y(_abc_17692_n1606) );
  AND2X2 AND2X2_4040 ( .A(_abc_17692_n9970), .B(_abc_17692_n9949), .Y(_abc_17692_n9971) );
  AND2X2 AND2X2_4041 ( .A(_abc_17692_n9804), .B(_abc_17692_n9577), .Y(_abc_17692_n9973) );
  AND2X2 AND2X2_4042 ( .A(_abc_17692_n9973), .B(_abc_17692_n9662), .Y(_abc_17692_n9974) );
  AND2X2 AND2X2_4043 ( .A(_abc_17692_n9369), .B(_abc_17692_n9974), .Y(_abc_17692_n9975) );
  AND2X2 AND2X2_4044 ( .A(_abc_17692_n9803), .B(_abc_17692_n9977), .Y(_abc_17692_n9978) );
  AND2X2 AND2X2_4045 ( .A(_abc_17692_n9973), .B(_abc_17692_n9665), .Y(_abc_17692_n9980) );
  AND2X2 AND2X2_4046 ( .A(_abc_17692_n9982), .B(_abc_17692_n9957), .Y(_abc_17692_n9983) );
  AND2X2 AND2X2_4047 ( .A(_abc_17692_n9984), .B(_abc_17692_n9956), .Y(_abc_17692_n9985) );
  AND2X2 AND2X2_4048 ( .A(_abc_17692_n9989), .B(_abc_17692_n9672), .Y(_abc_17692_n9990) );
  AND2X2 AND2X2_4049 ( .A(_abc_17692_n9990), .B(_abc_17692_n9378), .Y(_abc_17692_n9991) );
  AND2X2 AND2X2_405 ( .A(_abc_17692_n1542), .B(_abc_17692_n1606), .Y(_abc_17692_n1607) );
  AND2X2 AND2X2_4050 ( .A(_abc_17692_n9739), .B(workunit1_11_bF_buf3), .Y(_abc_17692_n9994) );
  AND2X2 AND2X2_4051 ( .A(_abc_17692_n9996), .B(_abc_17692_n9995), .Y(_abc_17692_n9997) );
  AND2X2 AND2X2_4052 ( .A(_abc_17692_n9993), .B(_abc_17692_n9997), .Y(_abc_17692_n9998) );
  AND2X2 AND2X2_4053 ( .A(_abc_17692_n9992), .B(_abc_17692_n9998), .Y(_abc_17692_n9999) );
  AND2X2 AND2X2_4054 ( .A(_abc_17692_n9999), .B(_abc_17692_n9898), .Y(_abc_17692_n10000) );
  AND2X2 AND2X2_4055 ( .A(_abc_17692_n10002), .B(_abc_17692_n9885), .Y(_abc_17692_n10003) );
  AND2X2 AND2X2_4056 ( .A(_abc_17692_n9764), .B(_abc_17692_n9642), .Y(_abc_17692_n10008) );
  AND2X2 AND2X2_4057 ( .A(_abc_17692_n10014), .B(_abc_17692_n9763), .Y(_abc_17692_n10015) );
  AND2X2 AND2X2_4058 ( .A(_abc_17692_n10018), .B(_abc_17692_n10016), .Y(_abc_17692_n10019) );
  AND2X2 AND2X2_4059 ( .A(_abc_17692_n10011), .B(_abc_17692_n10019), .Y(_abc_17692_n10020) );
  AND2X2 AND2X2_406 ( .A(_abc_17692_n1562_1), .B(_abc_17692_n1569), .Y(_abc_17692_n1608) );
  AND2X2 AND2X2_4060 ( .A(_abc_17692_n10020), .B(_abc_17692_n9908), .Y(_abc_17692_n10021) );
  AND2X2 AND2X2_4061 ( .A(_abc_17692_n10023), .B(_abc_17692_n10024), .Y(_abc_17692_n10025) );
  AND2X2 AND2X2_4062 ( .A(_abc_17692_n10025), .B(_abc_17692_n9921), .Y(_abc_17692_n10026) );
  AND2X2 AND2X2_4063 ( .A(_abc_17692_n9790), .B(_abc_17692_n9618), .Y(_abc_17692_n10029) );
  AND2X2 AND2X2_4064 ( .A(_abc_17692_n10029), .B(_abc_17692_n9696), .Y(_abc_17692_n10030) );
  AND2X2 AND2X2_4065 ( .A(_abc_17692_n10030), .B(_abc_17692_n9402), .Y(_abc_17692_n10031) );
  AND2X2 AND2X2_4066 ( .A(_abc_17692_n10032), .B(_abc_17692_n9788), .Y(_abc_17692_n10033) );
  AND2X2 AND2X2_4067 ( .A(_abc_17692_n10029), .B(_abc_17692_n9699), .Y(_abc_17692_n10035) );
  AND2X2 AND2X2_4068 ( .A(_abc_17692_n10037), .B(_abc_17692_n9932), .Y(_abc_17692_n10038) );
  AND2X2 AND2X2_4069 ( .A(_abc_17692_n10039), .B(_abc_17692_n9228), .Y(_abc_17692_n10040) );
  AND2X2 AND2X2_407 ( .A(_abc_17692_n1557), .B(sum_23_), .Y(_abc_17692_n1609) );
  AND2X2 AND2X2_4070 ( .A(_abc_17692_n8974), .B(_abc_17692_n9095), .Y(_abc_17692_n10041) );
  AND2X2 AND2X2_4071 ( .A(_abc_17692_n10042), .B(_abc_17692_n10040), .Y(_abc_17692_n10043) );
  AND2X2 AND2X2_4072 ( .A(_abc_17692_n10049), .B(_abc_17692_n10033), .Y(_abc_17692_n10050) );
  AND2X2 AND2X2_4073 ( .A(_abc_17692_n10047), .B(_abc_17692_n10050), .Y(_abc_17692_n10051) );
  AND2X2 AND2X2_4074 ( .A(_abc_17692_n10051), .B(_abc_17692_n9931), .Y(_abc_17692_n10052) );
  AND2X2 AND2X2_4075 ( .A(_abc_17692_n10028), .B(_abc_17692_n10054), .Y(_abc_17692_n10055) );
  AND2X2 AND2X2_4076 ( .A(_abc_17692_n10055), .B(_abc_17692_n10005), .Y(_abc_17692_n10056) );
  AND2X2 AND2X2_4077 ( .A(_abc_17692_n10056), .B(_abc_17692_n9987), .Y(_abc_17692_n10057) );
  AND2X2 AND2X2_4078 ( .A(state_8_bF_buf5), .B(\data_in1[12] ), .Y(_abc_17692_n10061) );
  AND2X2 AND2X2_4079 ( .A(_abc_17692_n10060), .B(_abc_17692_n10062), .Y(_abc_17692_n10063) );
  AND2X2 AND2X2_408 ( .A(_abc_17692_n1512), .B(_abc_17692_n1606), .Y(_abc_17692_n1612) );
  AND2X2 AND2X2_4080 ( .A(_abc_17692_n10058), .B(_abc_17692_n10063), .Y(_abc_17692_n10064) );
  AND2X2 AND2X2_4081 ( .A(_abc_17692_n9972), .B(_abc_17692_n10064), .Y(_abc_17692_n10065) );
  AND2X2 AND2X2_4082 ( .A(_abc_17692_n5430), .B(workunit2_9_), .Y(_abc_17692_n10068) );
  AND2X2 AND2X2_4083 ( .A(_abc_17692_n3471), .B(workunit2_18_), .Y(_abc_17692_n10069) );
  AND2X2 AND2X2_4084 ( .A(_abc_17692_n10070), .B(workunit2_13_), .Y(_abc_17692_n10071) );
  AND2X2 AND2X2_4085 ( .A(_abc_17692_n10067), .B(_abc_17692_n10074), .Y(_abc_17692_n10075) );
  AND2X2 AND2X2_4086 ( .A(_abc_17692_n10076), .B(_abc_17692_n10077), .Y(_abc_17692_n10078) );
  AND2X2 AND2X2_4087 ( .A(_abc_17692_n10081), .B(_abc_17692_n10079), .Y(_abc_17692_n10082) );
  AND2X2 AND2X2_4088 ( .A(_abc_17692_n10082), .B(workunit1_13_bF_buf0), .Y(_abc_17692_n10083) );
  AND2X2 AND2X2_4089 ( .A(_abc_17692_n10084), .B(_abc_17692_n3208), .Y(_abc_17692_n10085) );
  AND2X2 AND2X2_409 ( .A(_abc_17692_n1486), .B(_abc_17692_n1612), .Y(_abc_17692_n1613_1) );
  AND2X2 AND2X2_4090 ( .A(_abc_17692_n10088), .B(_abc_17692_n10087), .Y(_abc_17692_n10089) );
  AND2X2 AND2X2_4091 ( .A(_abc_17692_n10090), .B(_abc_17692_n10086), .Y(_abc_17692_n10091) );
  AND2X2 AND2X2_4092 ( .A(_abc_17692_n10094), .B(_abc_17692_n10095), .Y(_abc_17692_n10096) );
  AND2X2 AND2X2_4093 ( .A(_abc_17692_n10096), .B(workunit1_13_bF_buf3), .Y(_abc_17692_n10097) );
  AND2X2 AND2X2_4094 ( .A(_abc_17692_n10098), .B(_abc_17692_n3208), .Y(_abc_17692_n10099) );
  AND2X2 AND2X2_4095 ( .A(_abc_17692_n10105), .B(_abc_17692_n1877_bF_buf0), .Y(_abc_17692_n10106) );
  AND2X2 AND2X2_4096 ( .A(_abc_17692_n10106), .B(_abc_17692_n10104), .Y(_abc_17692_n10107) );
  AND2X2 AND2X2_4097 ( .A(_abc_17692_n10109), .B(_abc_17692_n10108), .Y(_abc_17692_n10110) );
  AND2X2 AND2X2_4098 ( .A(_abc_17692_n10110), .B(workunit1_13_bF_buf2), .Y(_abc_17692_n10111) );
  AND2X2 AND2X2_4099 ( .A(_abc_17692_n10112), .B(_abc_17692_n10113), .Y(_abc_17692_n10114) );
  AND2X2 AND2X2_41 ( .A(_abc_17692_n728), .B(_abc_17692_n726), .Y(data_out2_0__FF_INPUT) );
  AND2X2 AND2X2_410 ( .A(_abc_17692_n1614), .B(_abc_17692_n1605), .Y(_abc_17692_n1615) );
  AND2X2 AND2X2_4100 ( .A(_abc_17692_n10119), .B(_abc_17692_n1830_bF_buf0), .Y(_abc_17692_n10120) );
  AND2X2 AND2X2_4101 ( .A(_abc_17692_n10120), .B(_abc_17692_n10117), .Y(_abc_17692_n10121) );
  AND2X2 AND2X2_4102 ( .A(_abc_17692_n10122), .B(_abc_17692_n10123), .Y(_abc_17692_n10124) );
  AND2X2 AND2X2_4103 ( .A(_abc_17692_n10127), .B(_abc_17692_n10126), .Y(_abc_17692_n10128) );
  AND2X2 AND2X2_4104 ( .A(_abc_17692_n10129), .B(_abc_17692_n10125), .Y(_abc_17692_n10130) );
  AND2X2 AND2X2_4105 ( .A(_abc_17692_n10132), .B(_abc_17692_n9906), .Y(_abc_17692_n10133) );
  AND2X2 AND2X2_4106 ( .A(_abc_17692_n10136), .B(_abc_17692_n1846_bF_buf0), .Y(_abc_17692_n10137) );
  AND2X2 AND2X2_4107 ( .A(_abc_17692_n10137), .B(_abc_17692_n10135), .Y(_abc_17692_n10138) );
  AND2X2 AND2X2_4108 ( .A(_abc_17692_n10141), .B(state_10_bF_buf2), .Y(_abc_17692_n10142) );
  AND2X2 AND2X2_4109 ( .A(_abc_17692_n10142), .B(_abc_17692_n10093), .Y(_abc_17692_n10143) );
  AND2X2 AND2X2_411 ( .A(_abc_17692_n1617), .B(state_15_bF_buf0), .Y(_abc_17692_n1618) );
  AND2X2 AND2X2_4110 ( .A(_abc_17692_n10144), .B(workunit1_12_bF_buf1), .Y(_abc_17692_n10145) );
  AND2X2 AND2X2_4111 ( .A(_abc_17692_n10146), .B(_abc_17692_n10086), .Y(_abc_17692_n10147) );
  AND2X2 AND2X2_4112 ( .A(_abc_17692_n10148), .B(_abc_17692_n10087), .Y(_abc_17692_n10149) );
  AND2X2 AND2X2_4113 ( .A(_abc_17692_n10150), .B(_abc_17692_n1863_bF_buf10), .Y(_abc_17692_n10151) );
  AND2X2 AND2X2_4114 ( .A(_abc_17692_n9882), .B(workunit1_12_bF_buf0), .Y(_abc_17692_n10152) );
  AND2X2 AND2X2_4115 ( .A(_abc_17692_n10156), .B(_abc_17692_n1877_bF_buf10), .Y(_abc_17692_n10157) );
  AND2X2 AND2X2_4116 ( .A(_abc_17692_n10157), .B(_abc_17692_n10154), .Y(_abc_17692_n10158) );
  AND2X2 AND2X2_4117 ( .A(_abc_17692_n10159), .B(workunit1_12_bF_buf3), .Y(_abc_17692_n10160) );
  AND2X2 AND2X2_4118 ( .A(_abc_17692_n10164), .B(_abc_17692_n1830_bF_buf10), .Y(_abc_17692_n10165) );
  AND2X2 AND2X2_4119 ( .A(_abc_17692_n10165), .B(_abc_17692_n10163), .Y(_abc_17692_n10166) );
  AND2X2 AND2X2_412 ( .A(_abc_17692_n1618), .B(_abc_17692_n1616), .Y(_abc_17692_n1619) );
  AND2X2 AND2X2_4120 ( .A(_abc_17692_n10167), .B(workunit1_12_bF_buf2), .Y(_abc_17692_n10168) );
  AND2X2 AND2X2_4121 ( .A(_abc_17692_n10169), .B(_abc_17692_n10131), .Y(_abc_17692_n10170) );
  AND2X2 AND2X2_4122 ( .A(_abc_17692_n10171), .B(_abc_17692_n10130), .Y(_abc_17692_n10172) );
  AND2X2 AND2X2_4123 ( .A(_abc_17692_n10173), .B(_abc_17692_n1846_bF_buf10), .Y(_abc_17692_n10174) );
  AND2X2 AND2X2_4124 ( .A(_abc_17692_n10177), .B(state_14_bF_buf2), .Y(_abc_17692_n10178) );
  AND2X2 AND2X2_4125 ( .A(_abc_17692_n8383_bF_buf1), .B(workunit1_13_bF_buf3), .Y(_abc_17692_n10179) );
  AND2X2 AND2X2_4126 ( .A(state_8_bF_buf4), .B(\data_in1[13] ), .Y(_abc_17692_n10180) );
  AND2X2 AND2X2_4127 ( .A(_abc_17692_n10184), .B(_abc_17692_n10072), .Y(_abc_17692_n10185) );
  AND2X2 AND2X2_4128 ( .A(_abc_17692_n9868), .B(_abc_17692_n10185), .Y(_abc_17692_n10186) );
  AND2X2 AND2X2_4129 ( .A(_abc_17692_n10189), .B(_abc_17692_n10072), .Y(_abc_17692_n10190) );
  AND2X2 AND2X2_413 ( .A(delta_25_), .B(sum_25_), .Y(_abc_17692_n1622) );
  AND2X2 AND2X2_4130 ( .A(_abc_17692_n10188), .B(_abc_17692_n10191), .Y(_abc_17692_n10192) );
  AND2X2 AND2X2_4131 ( .A(_abc_17692_n5626), .B(workunit2_10_bF_buf3), .Y(_abc_17692_n10193) );
  AND2X2 AND2X2_4132 ( .A(_abc_17692_n3751), .B(workunit2_19_), .Y(_abc_17692_n10194) );
  AND2X2 AND2X2_4133 ( .A(_abc_17692_n10195), .B(workunit2_14_bF_buf3), .Y(_abc_17692_n10196) );
  AND2X2 AND2X2_4134 ( .A(_abc_17692_n10192), .B(_abc_17692_n10199), .Y(_abc_17692_n10200) );
  AND2X2 AND2X2_4135 ( .A(_abc_17692_n9861), .B(_abc_17692_n10186), .Y(_abc_17692_n10201) );
  AND2X2 AND2X2_4136 ( .A(_abc_17692_n10203), .B(_abc_17692_n10197), .Y(_abc_17692_n10204) );
  AND2X2 AND2X2_4137 ( .A(_abc_17692_n10202), .B(_abc_17692_n10204), .Y(_abc_17692_n10205) );
  AND2X2 AND2X2_4138 ( .A(_abc_17692_n4528), .B(_abc_17692_n10206), .Y(_abc_17692_n10207) );
  AND2X2 AND2X2_4139 ( .A(_abc_17692_n4527), .B(_abc_17692_n10208), .Y(_abc_17692_n10209) );
  AND2X2 AND2X2_414 ( .A(_abc_17692_n1624), .B(_abc_17692_n1625), .Y(_abc_17692_n1626) );
  AND2X2 AND2X2_4140 ( .A(_abc_17692_n10212), .B(_abc_17692_n10213), .Y(_abc_17692_n10214) );
  AND2X2 AND2X2_4141 ( .A(_abc_17692_n10215), .B(_abc_17692_n10216), .Y(_abc_17692_n10217) );
  AND2X2 AND2X2_4142 ( .A(_abc_17692_n10087), .B(_abc_17692_n9957), .Y(_abc_17692_n10218) );
  AND2X2 AND2X2_4143 ( .A(_abc_17692_n9982), .B(_abc_17692_n10218), .Y(_abc_17692_n10219) );
  AND2X2 AND2X2_4144 ( .A(_abc_17692_n10220), .B(_abc_17692_n10214), .Y(_abc_17692_n10222) );
  AND2X2 AND2X2_4145 ( .A(_abc_17692_n10223), .B(_abc_17692_n1863_bF_buf9), .Y(_abc_17692_n10224) );
  AND2X2 AND2X2_4146 ( .A(_abc_17692_n10224), .B(_abc_17692_n10221), .Y(_abc_17692_n10225) );
  AND2X2 AND2X2_4147 ( .A(_abc_17692_n10227), .B(_abc_17692_n10226), .Y(_abc_17692_n10228) );
  AND2X2 AND2X2_4148 ( .A(_abc_17692_n10228), .B(workunit1_14_bF_buf3), .Y(_abc_17692_n10229) );
  AND2X2 AND2X2_4149 ( .A(_abc_17692_n10230), .B(_abc_17692_n10231), .Y(_abc_17692_n10232) );
  AND2X2 AND2X2_415 ( .A(_abc_17692_n1627), .B(_abc_17692_n1623), .Y(_abc_17692_n1628) );
  AND2X2 AND2X2_4150 ( .A(_abc_17692_n10234), .B(_abc_17692_n10235), .Y(_abc_17692_n10236) );
  AND2X2 AND2X2_4151 ( .A(_abc_17692_n10101), .B(_abc_17692_n9885), .Y(_abc_17692_n10237) );
  AND2X2 AND2X2_4152 ( .A(_abc_17692_n10002), .B(_abc_17692_n10237), .Y(_abc_17692_n10238) );
  AND2X2 AND2X2_4153 ( .A(_abc_17692_n10239), .B(_abc_17692_n10233), .Y(_abc_17692_n10240) );
  AND2X2 AND2X2_4154 ( .A(_abc_17692_n10242), .B(_abc_17692_n1877_bF_buf9), .Y(_abc_17692_n10243) );
  AND2X2 AND2X2_4155 ( .A(_abc_17692_n10243), .B(_abc_17692_n10241), .Y(_abc_17692_n10244) );
  AND2X2 AND2X2_4156 ( .A(_abc_17692_n4642), .B(_abc_17692_n10206), .Y(_abc_17692_n10245) );
  AND2X2 AND2X2_4157 ( .A(_abc_17692_n10208), .B(_abc_17692_n4640), .Y(_abc_17692_n10246) );
  AND2X2 AND2X2_4158 ( .A(_abc_17692_n10249), .B(_abc_17692_n10250), .Y(_abc_17692_n10251) );
  AND2X2 AND2X2_4159 ( .A(_abc_17692_n10253), .B(_abc_17692_n10129), .Y(_abc_17692_n10254) );
  AND2X2 AND2X2_416 ( .A(delta_24_), .B(sum_24_), .Y(_abc_17692_n1630) );
  AND2X2 AND2X2_4160 ( .A(_abc_17692_n10130), .B(_abc_17692_n9921), .Y(_abc_17692_n10255) );
  AND2X2 AND2X2_4161 ( .A(_abc_17692_n10025), .B(_abc_17692_n10255), .Y(_abc_17692_n10256) );
  AND2X2 AND2X2_4162 ( .A(_abc_17692_n10257), .B(_abc_17692_n10251), .Y(_abc_17692_n10258) );
  AND2X2 AND2X2_4163 ( .A(_abc_17692_n10260), .B(_abc_17692_n1846_bF_buf9), .Y(_abc_17692_n10261) );
  AND2X2 AND2X2_4164 ( .A(_abc_17692_n10261), .B(_abc_17692_n10259), .Y(_abc_17692_n10262) );
  AND2X2 AND2X2_4165 ( .A(_abc_17692_n4601), .B(_abc_17692_n10206), .Y(_abc_17692_n10263) );
  AND2X2 AND2X2_4166 ( .A(_abc_17692_n10208), .B(_abc_17692_n4600), .Y(_abc_17692_n10264) );
  AND2X2 AND2X2_4167 ( .A(_abc_17692_n10267), .B(_abc_17692_n10268), .Y(_abc_17692_n10269) );
  AND2X2 AND2X2_4168 ( .A(_abc_17692_n10270), .B(_abc_17692_n10113), .Y(_abc_17692_n10271) );
  AND2X2 AND2X2_4169 ( .A(_abc_17692_n10114), .B(_abc_17692_n9932), .Y(_abc_17692_n10272) );
  AND2X2 AND2X2_417 ( .A(_abc_17692_n1634), .B(state_3_bF_buf4), .Y(_abc_17692_n1635) );
  AND2X2 AND2X2_4170 ( .A(_abc_17692_n10037), .B(_abc_17692_n10272), .Y(_abc_17692_n10273) );
  AND2X2 AND2X2_4171 ( .A(_abc_17692_n10274), .B(_abc_17692_n10269), .Y(_abc_17692_n10275) );
  AND2X2 AND2X2_4172 ( .A(_abc_17692_n10277), .B(_abc_17692_n1830_bF_buf9), .Y(_abc_17692_n10278) );
  AND2X2 AND2X2_4173 ( .A(_abc_17692_n10278), .B(_abc_17692_n10276), .Y(_abc_17692_n10279) );
  AND2X2 AND2X2_4174 ( .A(_abc_17692_n10282), .B(state_14_bF_buf1), .Y(_abc_17692_n10283) );
  AND2X2 AND2X2_4175 ( .A(_abc_17692_n10098), .B(workunit1_13_bF_buf2), .Y(_abc_17692_n10284) );
  AND2X2 AND2X2_4176 ( .A(_abc_17692_n10100), .B(_abc_17692_n9884), .Y(_abc_17692_n10285) );
  AND2X2 AND2X2_4177 ( .A(_abc_17692_n10100), .B(_abc_17692_n9898), .Y(_abc_17692_n10287) );
  AND2X2 AND2X2_4178 ( .A(_abc_17692_n9894), .B(_abc_17692_n10287), .Y(_abc_17692_n10288) );
  AND2X2 AND2X2_4179 ( .A(_abc_17692_n10289), .B(_abc_17692_n10232), .Y(_abc_17692_n10290) );
  AND2X2 AND2X2_418 ( .A(_abc_17692_n1635), .B(_abc_17692_n1633), .Y(_abc_17692_n1636_1) );
  AND2X2 AND2X2_4180 ( .A(_abc_17692_n10292), .B(_abc_17692_n1877_bF_buf8), .Y(_abc_17692_n10293) );
  AND2X2 AND2X2_4181 ( .A(_abc_17692_n10293), .B(_abc_17692_n10291), .Y(_abc_17692_n10294) );
  AND2X2 AND2X2_4182 ( .A(_abc_17692_n10124), .B(workunit1_13_bF_buf1), .Y(_abc_17692_n10296) );
  AND2X2 AND2X2_4183 ( .A(_abc_17692_n10298), .B(_abc_17692_n10297), .Y(_abc_17692_n10299) );
  AND2X2 AND2X2_4184 ( .A(_abc_17692_n9918), .B(_abc_17692_n10302), .Y(_abc_17692_n10303) );
  AND2X2 AND2X2_4185 ( .A(_abc_17692_n10304), .B(_abc_17692_n10295), .Y(_abc_17692_n10305) );
  AND2X2 AND2X2_4186 ( .A(_abc_17692_n10307), .B(_abc_17692_n1846_bF_buf8), .Y(_abc_17692_n10308) );
  AND2X2 AND2X2_4187 ( .A(_abc_17692_n10308), .B(_abc_17692_n10306), .Y(_abc_17692_n10309) );
  AND2X2 AND2X2_4188 ( .A(_abc_17692_n10311), .B(workunit1_13_bF_buf0), .Y(_abc_17692_n10312) );
  AND2X2 AND2X2_4189 ( .A(_abc_17692_n10115), .B(_abc_17692_n9928), .Y(_abc_17692_n10313) );
  AND2X2 AND2X2_419 ( .A(_abc_17692_n1605), .B(_abc_17692_n1629), .Y(_abc_17692_n1639) );
  AND2X2 AND2X2_4190 ( .A(_abc_17692_n10115), .B(_abc_17692_n9931), .Y(_abc_17692_n10315) );
  AND2X2 AND2X2_4191 ( .A(_abc_17692_n9941), .B(_abc_17692_n10315), .Y(_abc_17692_n10316) );
  AND2X2 AND2X2_4192 ( .A(_abc_17692_n10317), .B(_abc_17692_n10310), .Y(_abc_17692_n10318) );
  AND2X2 AND2X2_4193 ( .A(_abc_17692_n10320), .B(_abc_17692_n1830_bF_buf8), .Y(_abc_17692_n10321) );
  AND2X2 AND2X2_4194 ( .A(_abc_17692_n10321), .B(_abc_17692_n10319), .Y(_abc_17692_n10322) );
  AND2X2 AND2X2_4195 ( .A(_abc_17692_n10084), .B(workunit1_13_bF_buf3), .Y(_abc_17692_n10326) );
  AND2X2 AND2X2_4196 ( .A(_abc_17692_n10086), .B(_abc_17692_n9953), .Y(_abc_17692_n10327) );
  AND2X2 AND2X2_4197 ( .A(_abc_17692_n10086), .B(_abc_17692_n9956), .Y(_abc_17692_n10329) );
  AND2X2 AND2X2_4198 ( .A(_abc_17692_n9965), .B(_abc_17692_n10329), .Y(_abc_17692_n10330) );
  AND2X2 AND2X2_4199 ( .A(_abc_17692_n10331), .B(_abc_17692_n10325), .Y(_abc_17692_n10332) );
  AND2X2 AND2X2_42 ( .A(_abc_17692_n731_1), .B(_abc_17692_n730_1), .Y(data_out2_1__FF_INPUT) );
  AND2X2 AND2X2_420 ( .A(_abc_17692_n1614), .B(_abc_17692_n1639), .Y(_abc_17692_n1640) );
  AND2X2 AND2X2_4200 ( .A(_abc_17692_n10334), .B(_abc_17692_n1863_bF_buf8), .Y(_abc_17692_n10335) );
  AND2X2 AND2X2_4201 ( .A(_abc_17692_n10335), .B(_abc_17692_n10333), .Y(_abc_17692_n10336) );
  AND2X2 AND2X2_4202 ( .A(_abc_17692_n10337), .B(state_10_bF_buf1), .Y(_abc_17692_n10338) );
  AND2X2 AND2X2_4203 ( .A(_abc_17692_n8383_bF_buf0), .B(workunit1_14_bF_buf3), .Y(_abc_17692_n10339) );
  AND2X2 AND2X2_4204 ( .A(state_8_bF_buf3), .B(\data_in1[14] ), .Y(_abc_17692_n10340) );
  AND2X2 AND2X2_4205 ( .A(_abc_17692_n5769), .B(workunit2_11_), .Y(_abc_17692_n10345) );
  AND2X2 AND2X2_4206 ( .A(_abc_17692_n3905), .B(workunit2_20_), .Y(_abc_17692_n10346) );
  AND2X2 AND2X2_4207 ( .A(_abc_17692_n10347), .B(workunit2_15_), .Y(_abc_17692_n10348) );
  AND2X2 AND2X2_4208 ( .A(_abc_17692_n10349), .B(_abc_17692_n10350), .Y(_abc_17692_n10351) );
  AND2X2 AND2X2_4209 ( .A(_abc_17692_n10353), .B(_abc_17692_n10203), .Y(_abc_17692_n10354) );
  AND2X2 AND2X2_421 ( .A(_abc_17692_n1629), .B(_abc_17692_n1584), .Y(_abc_17692_n1642) );
  AND2X2 AND2X2_4210 ( .A(_abc_17692_n10357), .B(_abc_17692_n10352), .Y(_abc_17692_n10358) );
  AND2X2 AND2X2_4211 ( .A(_abc_17692_n10354), .B(_abc_17692_n10356), .Y(_abc_17692_n10360) );
  AND2X2 AND2X2_4212 ( .A(_abc_17692_n10344), .B(_abc_17692_n10351), .Y(_abc_17692_n10361) );
  AND2X2 AND2X2_4213 ( .A(_abc_17692_n10363), .B(_abc_17692_n10359), .Y(_abc_17692_n10364) );
  AND2X2 AND2X2_4214 ( .A(_abc_17692_n10366), .B(_abc_17692_n10367), .Y(_abc_17692_n10368) );
  AND2X2 AND2X2_4215 ( .A(_abc_17692_n10370), .B(workunit1_14_bF_buf2), .Y(_abc_17692_n10371) );
  AND2X2 AND2X2_4216 ( .A(_abc_17692_n10241), .B(_abc_17692_n10372), .Y(_abc_17692_n10373) );
  AND2X2 AND2X2_4217 ( .A(_abc_17692_n10373), .B(_abc_17692_n10369), .Y(_abc_17692_n10374) );
  AND2X2 AND2X2_4218 ( .A(_abc_17692_n10375), .B(_abc_17692_n10368), .Y(_abc_17692_n10376) );
  AND2X2 AND2X2_4219 ( .A(_abc_17692_n10377), .B(_abc_17692_n1877_bF_buf7), .Y(_abc_17692_n10378) );
  AND2X2 AND2X2_422 ( .A(_abc_17692_n1643), .B(state_15_bF_buf4), .Y(_abc_17692_n1644) );
  AND2X2 AND2X2_4220 ( .A(_abc_17692_n10379), .B(_abc_17692_n10380), .Y(_abc_17692_n10381) );
  AND2X2 AND2X2_4221 ( .A(_abc_17692_n10383), .B(_abc_17692_n10384), .Y(_abc_17692_n10385) );
  AND2X2 AND2X2_4222 ( .A(_abc_17692_n10382), .B(_abc_17692_n10386), .Y(_abc_17692_n10387) );
  AND2X2 AND2X2_4223 ( .A(_abc_17692_n10223), .B(_abc_17692_n10212), .Y(_abc_17692_n10388) );
  AND2X2 AND2X2_4224 ( .A(_abc_17692_n10392), .B(_abc_17692_n1863_bF_buf7), .Y(_abc_17692_n10393) );
  AND2X2 AND2X2_4225 ( .A(_abc_17692_n10393), .B(_abc_17692_n10390), .Y(_abc_17692_n10394) );
  AND2X2 AND2X2_4226 ( .A(_abc_17692_n10395), .B(_abc_17692_n10396), .Y(_abc_17692_n10397) );
  AND2X2 AND2X2_4227 ( .A(_abc_17692_n10399), .B(_abc_17692_n10400), .Y(_abc_17692_n10401) );
  AND2X2 AND2X2_4228 ( .A(_abc_17692_n10398), .B(_abc_17692_n10402), .Y(_abc_17692_n10403) );
  AND2X2 AND2X2_4229 ( .A(_abc_17692_n10259), .B(_abc_17692_n10249), .Y(_abc_17692_n10404) );
  AND2X2 AND2X2_423 ( .A(_abc_17692_n1641), .B(_abc_17692_n1644), .Y(_abc_17692_n1645) );
  AND2X2 AND2X2_4230 ( .A(_abc_17692_n10408), .B(_abc_17692_n1846_bF_buf7), .Y(_abc_17692_n10409) );
  AND2X2 AND2X2_4231 ( .A(_abc_17692_n10409), .B(_abc_17692_n10406), .Y(_abc_17692_n10410) );
  AND2X2 AND2X2_4232 ( .A(_abc_17692_n10412), .B(_abc_17692_n10411), .Y(_abc_17692_n10413) );
  AND2X2 AND2X2_4233 ( .A(_abc_17692_n10413), .B(workunit1_15_), .Y(_abc_17692_n10414) );
  AND2X2 AND2X2_4234 ( .A(_abc_17692_n4789_1), .B(_abc_17692_n10362), .Y(_abc_17692_n10415) );
  AND2X2 AND2X2_4235 ( .A(_abc_17692_n4787), .B(_abc_17692_n10358), .Y(_abc_17692_n10416) );
  AND2X2 AND2X2_4236 ( .A(_abc_17692_n10417), .B(_abc_17692_n3614), .Y(_abc_17692_n10418) );
  AND2X2 AND2X2_4237 ( .A(_abc_17692_n10276), .B(_abc_17692_n10267), .Y(_abc_17692_n10420) );
  AND2X2 AND2X2_4238 ( .A(_abc_17692_n10422), .B(_abc_17692_n10423), .Y(_abc_17692_n10424) );
  AND2X2 AND2X2_4239 ( .A(_abc_17692_n10426), .B(_abc_17692_n1830_bF_buf7), .Y(_abc_17692_n10427) );
  AND2X2 AND2X2_424 ( .A(_abc_17692_n1645), .B(_abc_17692_n1638), .Y(_abc_17692_n1646) );
  AND2X2 AND2X2_4240 ( .A(_abc_17692_n10427), .B(_abc_17692_n10421), .Y(_abc_17692_n10428) );
  AND2X2 AND2X2_4241 ( .A(_abc_17692_n10431), .B(state_14_bF_buf0), .Y(_abc_17692_n10432) );
  AND2X2 AND2X2_4242 ( .A(_abc_17692_n10291), .B(_abc_17692_n10230), .Y(_abc_17692_n10433) );
  AND2X2 AND2X2_4243 ( .A(_abc_17692_n10436), .B(_abc_17692_n1877_bF_buf6), .Y(_abc_17692_n10437) );
  AND2X2 AND2X2_4244 ( .A(_abc_17692_n10437), .B(_abc_17692_n10434), .Y(_abc_17692_n10438) );
  AND2X2 AND2X2_4245 ( .A(_abc_17692_n10266), .B(workunit1_14_bF_buf1), .Y(_abc_17692_n10439) );
  AND2X2 AND2X2_4246 ( .A(_abc_17692_n10319), .B(_abc_17692_n10440), .Y(_abc_17692_n10441) );
  AND2X2 AND2X2_4247 ( .A(_abc_17692_n10444), .B(_abc_17692_n1830_bF_buf6), .Y(_abc_17692_n10445) );
  AND2X2 AND2X2_4248 ( .A(_abc_17692_n10445), .B(_abc_17692_n10443), .Y(_abc_17692_n10446) );
  AND2X2 AND2X2_4249 ( .A(_abc_17692_n10248), .B(workunit1_14_bF_buf0), .Y(_abc_17692_n10447) );
  AND2X2 AND2X2_425 ( .A(_abc_17692_n722_bF_buf1), .B(sum_25_), .Y(_abc_17692_n1647) );
  AND2X2 AND2X2_4250 ( .A(_abc_17692_n10306), .B(_abc_17692_n10448), .Y(_abc_17692_n10449) );
  AND2X2 AND2X2_4251 ( .A(_abc_17692_n10452), .B(_abc_17692_n1846_bF_buf6), .Y(_abc_17692_n10453) );
  AND2X2 AND2X2_4252 ( .A(_abc_17692_n10453), .B(_abc_17692_n10451), .Y(_abc_17692_n10454) );
  AND2X2 AND2X2_4253 ( .A(_abc_17692_n10211), .B(workunit1_14_bF_buf3), .Y(_abc_17692_n10457) );
  AND2X2 AND2X2_4254 ( .A(_abc_17692_n10333), .B(_abc_17692_n10458), .Y(_abc_17692_n10459) );
  AND2X2 AND2X2_4255 ( .A(_abc_17692_n10462), .B(_abc_17692_n1863_bF_buf6), .Y(_abc_17692_n10463) );
  AND2X2 AND2X2_4256 ( .A(_abc_17692_n10463), .B(_abc_17692_n10461), .Y(_abc_17692_n10464) );
  AND2X2 AND2X2_4257 ( .A(_abc_17692_n10465), .B(state_10_bF_buf0), .Y(_abc_17692_n10466) );
  AND2X2 AND2X2_4258 ( .A(_abc_17692_n8383_bF_buf4), .B(workunit1_15_), .Y(_abc_17692_n10467) );
  AND2X2 AND2X2_4259 ( .A(state_8_bF_buf2), .B(\data_in1[15] ), .Y(_abc_17692_n10468) );
  AND2X2 AND2X2_426 ( .A(delta_26_), .B(sum_26_), .Y(_abc_17692_n1651) );
  AND2X2 AND2X2_4260 ( .A(_abc_17692_n10204), .B(_abc_17692_n10351), .Y(_abc_17692_n10472) );
  AND2X2 AND2X2_4261 ( .A(_abc_17692_n10186), .B(_abc_17692_n10472), .Y(_abc_17692_n10473) );
  AND2X2 AND2X2_4262 ( .A(_abc_17692_n10472), .B(_abc_17692_n10190), .Y(_abc_17692_n10478) );
  AND2X2 AND2X2_4263 ( .A(_abc_17692_n10350), .B(_abc_17692_n10196), .Y(_abc_17692_n10479) );
  AND2X2 AND2X2_4264 ( .A(_abc_17692_n10477), .B(_abc_17692_n10482), .Y(_abc_17692_n10483) );
  AND2X2 AND2X2_4265 ( .A(_abc_17692_n10476), .B(_abc_17692_n10483), .Y(_abc_17692_n10484) );
  AND2X2 AND2X2_4266 ( .A(_abc_17692_n10485), .B(_abc_17692_n10486), .Y(_abc_17692_n10487) );
  AND2X2 AND2X2_4267 ( .A(_abc_17692_n10488), .B(workunit2_16_bF_buf2), .Y(_abc_17692_n10489) );
  AND2X2 AND2X2_4268 ( .A(_abc_17692_n10487), .B(_abc_17692_n9717), .Y(_abc_17692_n10490) );
  AND2X2 AND2X2_4269 ( .A(_abc_17692_n10484), .B(_abc_17692_n10491), .Y(_abc_17692_n10492) );
  AND2X2 AND2X2_427 ( .A(_abc_17692_n1652), .B(_abc_17692_n1653), .Y(_abc_17692_n1654) );
  AND2X2 AND2X2_4270 ( .A(_abc_17692_n9859), .B(_abc_17692_n10473), .Y(_abc_17692_n10493) );
  AND2X2 AND2X2_4271 ( .A(_abc_17692_n9278), .B(_abc_17692_n10493), .Y(_abc_17692_n10494) );
  AND2X2 AND2X2_4272 ( .A(_abc_17692_n9856), .B(_abc_17692_n10473), .Y(_abc_17692_n10495) );
  AND2X2 AND2X2_4273 ( .A(_abc_17692_n10497), .B(_abc_17692_n10498), .Y(_abc_17692_n10499) );
  AND2X2 AND2X2_4274 ( .A(_abc_17692_n10503), .B(_abc_17692_n10502), .Y(_abc_17692_n10504) );
  AND2X2 AND2X2_4275 ( .A(_abc_17692_n10504), .B(workunit1_16_bF_buf1), .Y(_abc_17692_n10505) );
  AND2X2 AND2X2_4276 ( .A(_abc_17692_n10506), .B(_abc_17692_n10507), .Y(_abc_17692_n10508) );
  AND2X2 AND2X2_4277 ( .A(_abc_17692_n10368), .B(_abc_17692_n10232), .Y(_abc_17692_n10509) );
  AND2X2 AND2X2_4278 ( .A(_abc_17692_n10509), .B(_abc_17692_n10286), .Y(_abc_17692_n10510) );
  AND2X2 AND2X2_4279 ( .A(_abc_17692_n10366), .B(_abc_17692_n10229), .Y(_abc_17692_n10512) );
  AND2X2 AND2X2_428 ( .A(_abc_17692_n1585), .B(_abc_17692_n1628), .Y(_abc_17692_n1657) );
  AND2X2 AND2X2_4280 ( .A(_abc_17692_n10509), .B(_abc_17692_n10287), .Y(_abc_17692_n10515) );
  AND2X2 AND2X2_4281 ( .A(_abc_17692_n9894), .B(_abc_17692_n10515), .Y(_abc_17692_n10516) );
  AND2X2 AND2X2_4282 ( .A(_abc_17692_n10517), .B(_abc_17692_n10508), .Y(_abc_17692_n10518) );
  AND2X2 AND2X2_4283 ( .A(_abc_17692_n10520), .B(_abc_17692_n1877_bF_buf5), .Y(_abc_17692_n10521) );
  AND2X2 AND2X2_4284 ( .A(_abc_17692_n10521), .B(_abc_17692_n10519), .Y(_abc_17692_n10522) );
  AND2X2 AND2X2_4285 ( .A(_abc_17692_n10523), .B(_abc_17692_n10524), .Y(_abc_17692_n10525) );
  AND2X2 AND2X2_4286 ( .A(_abc_17692_n10525), .B(workunit1_16_bF_buf3), .Y(_abc_17692_n10526) );
  AND2X2 AND2X2_4287 ( .A(_abc_17692_n10527), .B(_abc_17692_n10528), .Y(_abc_17692_n10529) );
  AND2X2 AND2X2_4288 ( .A(_abc_17692_n10397), .B(workunit1_15_), .Y(_abc_17692_n10532) );
  AND2X2 AND2X2_4289 ( .A(_abc_17692_n10534), .B(_abc_17692_n10533), .Y(_abc_17692_n10535) );
  AND2X2 AND2X2_429 ( .A(_abc_17692_n1627), .B(_abc_17692_n1630), .Y(_abc_17692_n1660_1) );
  AND2X2 AND2X2_4290 ( .A(_abc_17692_n10531), .B(_abc_17692_n10535), .Y(_abc_17692_n10536) );
  AND2X2 AND2X2_4291 ( .A(_abc_17692_n10538), .B(_abc_17692_n10536), .Y(_abc_17692_n10539) );
  AND2X2 AND2X2_4292 ( .A(_abc_17692_n10540), .B(_abc_17692_n10529), .Y(_abc_17692_n10542) );
  AND2X2 AND2X2_4293 ( .A(_abc_17692_n10543), .B(_abc_17692_n1846_bF_buf5), .Y(_abc_17692_n10544) );
  AND2X2 AND2X2_4294 ( .A(_abc_17692_n10544), .B(_abc_17692_n10541), .Y(_abc_17692_n10545) );
  AND2X2 AND2X2_4295 ( .A(_abc_17692_n10546), .B(_abc_17692_n10547), .Y(_abc_17692_n10548) );
  AND2X2 AND2X2_4296 ( .A(_abc_17692_n10548), .B(workunit1_16_bF_buf1), .Y(_abc_17692_n10549) );
  AND2X2 AND2X2_4297 ( .A(_abc_17692_n10550), .B(_abc_17692_n10551), .Y(_abc_17692_n10552) );
  AND2X2 AND2X2_4298 ( .A(_abc_17692_n10419), .B(_abc_17692_n10310), .Y(_abc_17692_n10553) );
  AND2X2 AND2X2_4299 ( .A(_abc_17692_n10314), .B(_abc_17692_n10553), .Y(_abc_17692_n10554) );
  AND2X2 AND2X2_43 ( .A(_abc_17692_n734), .B(_abc_17692_n733), .Y(data_out2_2__FF_INPUT) );
  AND2X2 AND2X2_430 ( .A(_abc_17692_n1659), .B(_abc_17692_n1662), .Y(_abc_17692_n1663) );
  AND2X2 AND2X2_4300 ( .A(_abc_17692_n10419), .B(_abc_17692_n10439), .Y(_abc_17692_n10555) );
  AND2X2 AND2X2_4301 ( .A(_abc_17692_n10417), .B(workunit1_15_), .Y(_abc_17692_n10556) );
  AND2X2 AND2X2_4302 ( .A(_abc_17692_n10553), .B(_abc_17692_n10315), .Y(_abc_17692_n10559) );
  AND2X2 AND2X2_4303 ( .A(_abc_17692_n9941), .B(_abc_17692_n10559), .Y(_abc_17692_n10560) );
  AND2X2 AND2X2_4304 ( .A(_abc_17692_n10561), .B(_abc_17692_n10552), .Y(_abc_17692_n10563) );
  AND2X2 AND2X2_4305 ( .A(_abc_17692_n10564), .B(_abc_17692_n1830_bF_buf5), .Y(_abc_17692_n10565) );
  AND2X2 AND2X2_4306 ( .A(_abc_17692_n10565), .B(_abc_17692_n10562), .Y(_abc_17692_n10566) );
  AND2X2 AND2X2_4307 ( .A(_abc_17692_n10570), .B(_abc_17692_n10569), .Y(_abc_17692_n10571) );
  AND2X2 AND2X2_4308 ( .A(_abc_17692_n10571), .B(workunit1_16_bF_buf3), .Y(_abc_17692_n10572) );
  AND2X2 AND2X2_4309 ( .A(_abc_17692_n10573), .B(_abc_17692_n10574), .Y(_abc_17692_n10575) );
  AND2X2 AND2X2_431 ( .A(_abc_17692_n1664), .B(_abc_17692_n1656), .Y(_abc_17692_n1666) );
  AND2X2 AND2X2_4310 ( .A(_abc_17692_n10391), .B(_abc_17692_n10325), .Y(_abc_17692_n10576) );
  AND2X2 AND2X2_4311 ( .A(_abc_17692_n10576), .B(_abc_17692_n10328), .Y(_abc_17692_n10577) );
  AND2X2 AND2X2_4312 ( .A(_abc_17692_n10391), .B(_abc_17692_n10457), .Y(_abc_17692_n10578) );
  AND2X2 AND2X2_4313 ( .A(_abc_17692_n10381), .B(workunit1_15_), .Y(_abc_17692_n10579) );
  AND2X2 AND2X2_4314 ( .A(_abc_17692_n10576), .B(_abc_17692_n10329), .Y(_abc_17692_n10582) );
  AND2X2 AND2X2_4315 ( .A(_abc_17692_n9965), .B(_abc_17692_n10582), .Y(_abc_17692_n10583) );
  AND2X2 AND2X2_4316 ( .A(_abc_17692_n10584), .B(_abc_17692_n10575), .Y(_abc_17692_n10586) );
  AND2X2 AND2X2_4317 ( .A(_abc_17692_n10587), .B(_abc_17692_n1863_bF_buf5), .Y(_abc_17692_n10588) );
  AND2X2 AND2X2_4318 ( .A(_abc_17692_n10588), .B(_abc_17692_n10585), .Y(_abc_17692_n10589) );
  AND2X2 AND2X2_4319 ( .A(_abc_17692_n10590), .B(state_10_bF_buf4), .Y(_abc_17692_n10591) );
  AND2X2 AND2X2_432 ( .A(_abc_17692_n1667), .B(state_3_bF_buf3), .Y(_abc_17692_n1668) );
  AND2X2 AND2X2_4320 ( .A(_abc_17692_n10387), .B(_abc_17692_n10214), .Y(_abc_17692_n10593) );
  AND2X2 AND2X2_4321 ( .A(_abc_17692_n10593), .B(_abc_17692_n10217), .Y(_abc_17692_n10594) );
  AND2X2 AND2X2_4322 ( .A(_abc_17692_n10597), .B(_abc_17692_n10386), .Y(_abc_17692_n10598) );
  AND2X2 AND2X2_4323 ( .A(_abc_17692_n10593), .B(_abc_17692_n10218), .Y(_abc_17692_n10600) );
  AND2X2 AND2X2_4324 ( .A(_abc_17692_n9982), .B(_abc_17692_n10600), .Y(_abc_17692_n10601) );
  AND2X2 AND2X2_4325 ( .A(_abc_17692_n10602), .B(_abc_17692_n10592), .Y(_abc_17692_n10604) );
  AND2X2 AND2X2_4326 ( .A(_abc_17692_n10605), .B(_abc_17692_n1863_bF_buf4), .Y(_abc_17692_n10606) );
  AND2X2 AND2X2_4327 ( .A(_abc_17692_n10606), .B(_abc_17692_n10603), .Y(_abc_17692_n10607) );
  AND2X2 AND2X2_4328 ( .A(_abc_17692_n10364), .B(workunit1_15_), .Y(_abc_17692_n10612) );
  AND2X2 AND2X2_4329 ( .A(_abc_17692_n10614), .B(_abc_17692_n10613), .Y(_abc_17692_n10615) );
  AND2X2 AND2X2_433 ( .A(_abc_17692_n1668), .B(_abc_17692_n1665), .Y(_abc_17692_n1669) );
  AND2X2 AND2X2_4330 ( .A(_abc_17692_n10611), .B(_abc_17692_n10615), .Y(_abc_17692_n10616) );
  AND2X2 AND2X2_4331 ( .A(_abc_17692_n10620), .B(_abc_17692_n10002), .Y(_abc_17692_n10621) );
  AND2X2 AND2X2_4332 ( .A(_abc_17692_n10622), .B(_abc_17692_n10608), .Y(_abc_17692_n10623) );
  AND2X2 AND2X2_4333 ( .A(_abc_17692_n10625), .B(_abc_17692_n1877_bF_buf4), .Y(_abc_17692_n10626) );
  AND2X2 AND2X2_4334 ( .A(_abc_17692_n10626), .B(_abc_17692_n10624), .Y(_abc_17692_n10627) );
  AND2X2 AND2X2_4335 ( .A(_abc_17692_n10424), .B(_abc_17692_n10269), .Y(_abc_17692_n10629) );
  AND2X2 AND2X2_4336 ( .A(_abc_17692_n10629), .B(_abc_17692_n10271), .Y(_abc_17692_n10630) );
  AND2X2 AND2X2_4337 ( .A(_abc_17692_n10631), .B(_abc_17692_n10422), .Y(_abc_17692_n10632) );
  AND2X2 AND2X2_4338 ( .A(_abc_17692_n10629), .B(_abc_17692_n10272), .Y(_abc_17692_n10635) );
  AND2X2 AND2X2_4339 ( .A(_abc_17692_n10037), .B(_abc_17692_n10635), .Y(_abc_17692_n10636) );
  AND2X2 AND2X2_434 ( .A(_abc_17692_n1624), .B(sum_25_), .Y(_abc_17692_n1670) );
  AND2X2 AND2X2_4340 ( .A(_abc_17692_n10637), .B(_abc_17692_n10628), .Y(_abc_17692_n10638) );
  AND2X2 AND2X2_4341 ( .A(_abc_17692_n10640), .B(_abc_17692_n1830_bF_buf4), .Y(_abc_17692_n10641) );
  AND2X2 AND2X2_4342 ( .A(_abc_17692_n10641), .B(_abc_17692_n10639), .Y(_abc_17692_n10642) );
  AND2X2 AND2X2_4343 ( .A(_abc_17692_n10403), .B(_abc_17692_n10251), .Y(_abc_17692_n10644) );
  AND2X2 AND2X2_4344 ( .A(_abc_17692_n10644), .B(_abc_17692_n10254), .Y(_abc_17692_n10645) );
  AND2X2 AND2X2_4345 ( .A(_abc_17692_n10402), .B(_abc_17692_n10646), .Y(_abc_17692_n10647) );
  AND2X2 AND2X2_4346 ( .A(_abc_17692_n10648), .B(_abc_17692_n10398), .Y(_abc_17692_n10649) );
  AND2X2 AND2X2_4347 ( .A(_abc_17692_n10644), .B(_abc_17692_n10255), .Y(_abc_17692_n10652) );
  AND2X2 AND2X2_4348 ( .A(_abc_17692_n10025), .B(_abc_17692_n10652), .Y(_abc_17692_n10653) );
  AND2X2 AND2X2_4349 ( .A(_abc_17692_n10654), .B(_abc_17692_n10643), .Y(_abc_17692_n10656) );
  AND2X2 AND2X2_435 ( .A(_abc_17692_n1672), .B(_abc_17692_n1655), .Y(_abc_17692_n1673) );
  AND2X2 AND2X2_4350 ( .A(_abc_17692_n10657), .B(_abc_17692_n1846_bF_buf4), .Y(_abc_17692_n10658) );
  AND2X2 AND2X2_4351 ( .A(_abc_17692_n10658), .B(_abc_17692_n10655), .Y(_abc_17692_n10659) );
  AND2X2 AND2X2_4352 ( .A(_abc_17692_n10662), .B(state_14_bF_buf4), .Y(_abc_17692_n10663) );
  AND2X2 AND2X2_4353 ( .A(_abc_17692_n8383_bF_buf3), .B(workunit1_16_bF_buf1), .Y(_abc_17692_n10664) );
  AND2X2 AND2X2_4354 ( .A(state_8_bF_buf1), .B(\data_in1[16] ), .Y(_abc_17692_n10665) );
  AND2X2 AND2X2_4355 ( .A(_abc_17692_n10670), .B(_abc_17692_n10671), .Y(_abc_17692_n10672) );
  AND2X2 AND2X2_4356 ( .A(_abc_17692_n10673), .B(workunit2_17_), .Y(_abc_17692_n10674) );
  AND2X2 AND2X2_4357 ( .A(_abc_17692_n10672), .B(_abc_17692_n5260), .Y(_abc_17692_n10676) );
  AND2X2 AND2X2_4358 ( .A(_abc_17692_n10675), .B(_abc_17692_n10677), .Y(_abc_17692_n10678) );
  AND2X2 AND2X2_4359 ( .A(_abc_17692_n10669), .B(_abc_17692_n10679), .Y(_abc_17692_n10681) );
  AND2X2 AND2X2_436 ( .A(_abc_17692_n1675), .B(state_15_bF_buf3), .Y(_abc_17692_n1676) );
  AND2X2 AND2X2_4360 ( .A(_abc_17692_n10682), .B(_abc_17692_n10680), .Y(_abc_17692_n10683) );
  AND2X2 AND2X2_4361 ( .A(_abc_17692_n10686), .B(_abc_17692_n10684), .Y(_abc_17692_n10687) );
  AND2X2 AND2X2_4362 ( .A(_abc_17692_n10687), .B(workunit1_17_), .Y(_abc_17692_n10688) );
  AND2X2 AND2X2_4363 ( .A(_abc_17692_n10690), .B(_abc_17692_n4059), .Y(_abc_17692_n10691) );
  AND2X2 AND2X2_4364 ( .A(_abc_17692_n10692), .B(_abc_17692_n10689), .Y(_abc_17692_n10693) );
  AND2X2 AND2X2_4365 ( .A(_abc_17692_n10587), .B(_abc_17692_n10573), .Y(_abc_17692_n10694) );
  AND2X2 AND2X2_4366 ( .A(_abc_17692_n10695), .B(_abc_17692_n10693), .Y(_abc_17692_n10696) );
  AND2X2 AND2X2_4367 ( .A(_abc_17692_n10694), .B(_abc_17692_n10697), .Y(_abc_17692_n10698) );
  AND2X2 AND2X2_4368 ( .A(_abc_17692_n10702), .B(_abc_17692_n10701), .Y(_abc_17692_n10703) );
  AND2X2 AND2X2_4369 ( .A(_abc_17692_n10703), .B(workunit1_17_), .Y(_abc_17692_n10704) );
  AND2X2 AND2X2_437 ( .A(_abc_17692_n1676), .B(_abc_17692_n1674), .Y(_abc_17692_n1677) );
  AND2X2 AND2X2_4370 ( .A(_abc_17692_n10706), .B(_abc_17692_n4059), .Y(_abc_17692_n10707) );
  AND2X2 AND2X2_4371 ( .A(_abc_17692_n10708), .B(_abc_17692_n10705), .Y(_abc_17692_n10709) );
  AND2X2 AND2X2_4372 ( .A(_abc_17692_n10519), .B(_abc_17692_n10506), .Y(_abc_17692_n10710) );
  AND2X2 AND2X2_4373 ( .A(_abc_17692_n10714), .B(_abc_17692_n1877_bF_buf3), .Y(_abc_17692_n10715) );
  AND2X2 AND2X2_4374 ( .A(_abc_17692_n10715), .B(_abc_17692_n10711), .Y(_abc_17692_n10716) );
  AND2X2 AND2X2_4375 ( .A(_abc_17692_n10717), .B(_abc_17692_n10718), .Y(_abc_17692_n10719) );
  AND2X2 AND2X2_4376 ( .A(_abc_17692_n10720), .B(workunit1_17_), .Y(_abc_17692_n10721) );
  AND2X2 AND2X2_4377 ( .A(_abc_17692_n10719), .B(_abc_17692_n4059), .Y(_abc_17692_n10722) );
  AND2X2 AND2X2_4378 ( .A(_abc_17692_n10564), .B(_abc_17692_n10550), .Y(_abc_17692_n10724) );
  AND2X2 AND2X2_4379 ( .A(_abc_17692_n10728), .B(_abc_17692_n1830_bF_buf3), .Y(_abc_17692_n10729) );
  AND2X2 AND2X2_438 ( .A(_abc_17692_n722_bF_buf0), .B(sum_26_), .Y(_abc_17692_n1678) );
  AND2X2 AND2X2_4380 ( .A(_abc_17692_n10729), .B(_abc_17692_n10726), .Y(_abc_17692_n10730) );
  AND2X2 AND2X2_4381 ( .A(_abc_17692_n5287), .B(_abc_17692_n10685), .Y(_abc_17692_n10731) );
  AND2X2 AND2X2_4382 ( .A(_abc_17692_n5286), .B(_abc_17692_n10683), .Y(_abc_17692_n10732) );
  AND2X2 AND2X2_4383 ( .A(_abc_17692_n10736), .B(_abc_17692_n10734), .Y(_abc_17692_n10737) );
  AND2X2 AND2X2_4384 ( .A(_abc_17692_n10543), .B(_abc_17692_n10527), .Y(_abc_17692_n10738) );
  AND2X2 AND2X2_4385 ( .A(_abc_17692_n10742), .B(_abc_17692_n1846_bF_buf3), .Y(_abc_17692_n10743) );
  AND2X2 AND2X2_4386 ( .A(_abc_17692_n10743), .B(_abc_17692_n10739), .Y(_abc_17692_n10744) );
  AND2X2 AND2X2_4387 ( .A(_abc_17692_n10747), .B(state_10_bF_buf3), .Y(_abc_17692_n10748) );
  AND2X2 AND2X2_4388 ( .A(_abc_17692_n10748), .B(_abc_17692_n10700), .Y(_abc_17692_n10749) );
  AND2X2 AND2X2_4389 ( .A(_abc_17692_n10750), .B(workunit1_16_bF_buf0), .Y(_abc_17692_n10751) );
  AND2X2 AND2X2_439 ( .A(_abc_17692_n1682), .B(delta_27_), .Y(_abc_17692_n1683) );
  AND2X2 AND2X2_4390 ( .A(_abc_17692_n10605), .B(_abc_17692_n10752), .Y(_abc_17692_n10753) );
  AND2X2 AND2X2_4391 ( .A(_abc_17692_n10754), .B(_abc_17692_n10697), .Y(_abc_17692_n10755) );
  AND2X2 AND2X2_4392 ( .A(_abc_17692_n10753), .B(_abc_17692_n10693), .Y(_abc_17692_n10756) );
  AND2X2 AND2X2_4393 ( .A(_abc_17692_n10757), .B(_abc_17692_n1863_bF_buf2), .Y(_abc_17692_n10758) );
  AND2X2 AND2X2_4394 ( .A(_abc_17692_n10759), .B(workunit1_16_bF_buf3), .Y(_abc_17692_n10760) );
  AND2X2 AND2X2_4395 ( .A(_abc_17692_n10624), .B(_abc_17692_n10761), .Y(_abc_17692_n10762) );
  AND2X2 AND2X2_4396 ( .A(_abc_17692_n10765), .B(_abc_17692_n10763), .Y(_abc_17692_n10766) );
  AND2X2 AND2X2_4397 ( .A(_abc_17692_n10766), .B(_abc_17692_n1877_bF_buf2), .Y(_abc_17692_n10767) );
  AND2X2 AND2X2_4398 ( .A(_abc_17692_n10768), .B(workunit1_16_bF_buf2), .Y(_abc_17692_n10769) );
  AND2X2 AND2X2_4399 ( .A(_abc_17692_n10657), .B(_abc_17692_n10770), .Y(_abc_17692_n10771) );
  AND2X2 AND2X2_44 ( .A(_abc_17692_n737), .B(_abc_17692_n736), .Y(data_out2_3__FF_INPUT) );
  AND2X2 AND2X2_440 ( .A(_abc_17692_n1686), .B(_abc_17692_n1656), .Y(_abc_17692_n1689) );
  AND2X2 AND2X2_4400 ( .A(_abc_17692_n10774), .B(_abc_17692_n1846_bF_buf2), .Y(_abc_17692_n10775) );
  AND2X2 AND2X2_4401 ( .A(_abc_17692_n10775), .B(_abc_17692_n10773), .Y(_abc_17692_n10776) );
  AND2X2 AND2X2_4402 ( .A(_abc_17692_n10777), .B(workunit1_16_bF_buf1), .Y(_abc_17692_n10778) );
  AND2X2 AND2X2_4403 ( .A(_abc_17692_n10639), .B(_abc_17692_n10779), .Y(_abc_17692_n10780) );
  AND2X2 AND2X2_4404 ( .A(_abc_17692_n10783), .B(_abc_17692_n1830_bF_buf2), .Y(_abc_17692_n10784) );
  AND2X2 AND2X2_4405 ( .A(_abc_17692_n10784), .B(_abc_17692_n10781), .Y(_abc_17692_n10785) );
  AND2X2 AND2X2_4406 ( .A(_abc_17692_n10788), .B(state_14_bF_buf3), .Y(_abc_17692_n10789) );
  AND2X2 AND2X2_4407 ( .A(_abc_17692_n8383_bF_buf2), .B(workunit1_17_), .Y(_abc_17692_n10790) );
  AND2X2 AND2X2_4408 ( .A(state_8_bF_buf0), .B(\data_in1[17] ), .Y(_abc_17692_n10791) );
  AND2X2 AND2X2_4409 ( .A(_abc_17692_n10677), .B(_abc_17692_n10489), .Y(_abc_17692_n10795) );
  AND2X2 AND2X2_441 ( .A(_abc_17692_n1686), .B(_abc_17692_n1651), .Y(_abc_17692_n1692) );
  AND2X2 AND2X2_4410 ( .A(_abc_17692_n10498), .B(_abc_17692_n10678), .Y(_abc_17692_n10797) );
  AND2X2 AND2X2_4411 ( .A(_abc_17692_n10497), .B(_abc_17692_n10797), .Y(_abc_17692_n10798) );
  AND2X2 AND2X2_4412 ( .A(_abc_17692_n10800), .B(_abc_17692_n10801), .Y(_abc_17692_n10802) );
  AND2X2 AND2X2_4413 ( .A(_abc_17692_n10803), .B(workunit2_18_), .Y(_abc_17692_n10804) );
  AND2X2 AND2X2_4414 ( .A(_abc_17692_n10802), .B(_abc_17692_n5430), .Y(_abc_17692_n10805) );
  AND2X2 AND2X2_4415 ( .A(_abc_17692_n10799), .B(_abc_17692_n10807), .Y(_abc_17692_n10808) );
  AND2X2 AND2X2_4416 ( .A(_abc_17692_n10809), .B(_abc_17692_n10806), .Y(_abc_17692_n10810) );
  AND2X2 AND2X2_4417 ( .A(_abc_17692_n10814), .B(_abc_17692_n10813), .Y(_abc_17692_n10815) );
  AND2X2 AND2X2_4418 ( .A(_abc_17692_n10816), .B(_abc_17692_n4322), .Y(_abc_17692_n10817) );
  AND2X2 AND2X2_4419 ( .A(_abc_17692_n10815), .B(workunit1_18_), .Y(_abc_17692_n10818) );
  AND2X2 AND2X2_442 ( .A(_abc_17692_n1693), .B(state_3_bF_buf2), .Y(_abc_17692_n1694) );
  AND2X2 AND2X2_4420 ( .A(_abc_17692_n10692), .B(_abc_17692_n10820), .Y(_abc_17692_n10821) );
  AND2X2 AND2X2_4421 ( .A(_abc_17692_n10693), .B(_abc_17692_n10592), .Y(_abc_17692_n10822) );
  AND2X2 AND2X2_4422 ( .A(_abc_17692_n10602), .B(_abc_17692_n10822), .Y(_abc_17692_n10823) );
  AND2X2 AND2X2_4423 ( .A(_abc_17692_n10824), .B(_abc_17692_n10819), .Y(_abc_17692_n10826) );
  AND2X2 AND2X2_4424 ( .A(_abc_17692_n10827), .B(_abc_17692_n1863_bF_buf1), .Y(_abc_17692_n10828) );
  AND2X2 AND2X2_4425 ( .A(_abc_17692_n10828), .B(_abc_17692_n10825), .Y(_abc_17692_n10829) );
  AND2X2 AND2X2_4426 ( .A(_abc_17692_n10831), .B(_abc_17692_n10830), .Y(_abc_17692_n10832) );
  AND2X2 AND2X2_4427 ( .A(_abc_17692_n10832), .B(workunit1_18_), .Y(_abc_17692_n10833) );
  AND2X2 AND2X2_4428 ( .A(_abc_17692_n10834), .B(_abc_17692_n10835), .Y(_abc_17692_n10836) );
  AND2X2 AND2X2_4429 ( .A(_abc_17692_n10708), .B(_abc_17692_n10838), .Y(_abc_17692_n10839) );
  AND2X2 AND2X2_443 ( .A(_abc_17692_n1691), .B(_abc_17692_n1694), .Y(_abc_17692_n1695) );
  AND2X2 AND2X2_4430 ( .A(_abc_17692_n10709), .B(_abc_17692_n10608), .Y(_abc_17692_n10840) );
  AND2X2 AND2X2_4431 ( .A(_abc_17692_n10622), .B(_abc_17692_n10840), .Y(_abc_17692_n10841) );
  AND2X2 AND2X2_4432 ( .A(_abc_17692_n10842), .B(_abc_17692_n10837), .Y(_abc_17692_n10843) );
  AND2X2 AND2X2_4433 ( .A(_abc_17692_n10845), .B(_abc_17692_n1877_bF_buf1), .Y(_abc_17692_n10846) );
  AND2X2 AND2X2_4434 ( .A(_abc_17692_n10846), .B(_abc_17692_n10844), .Y(_abc_17692_n10847) );
  AND2X2 AND2X2_4435 ( .A(_abc_17692_n10848), .B(_abc_17692_n10849), .Y(_abc_17692_n10850) );
  AND2X2 AND2X2_4436 ( .A(_abc_17692_n10853), .B(_abc_17692_n10851), .Y(_abc_17692_n10854) );
  AND2X2 AND2X2_4437 ( .A(_abc_17692_n10856), .B(_abc_17692_n10855), .Y(_abc_17692_n10857) );
  AND2X2 AND2X2_4438 ( .A(_abc_17692_n10727), .B(_abc_17692_n10628), .Y(_abc_17692_n10858) );
  AND2X2 AND2X2_4439 ( .A(_abc_17692_n10637), .B(_abc_17692_n10858), .Y(_abc_17692_n10859) );
  AND2X2 AND2X2_444 ( .A(_abc_17692_n1688), .B(_abc_17692_n1695), .Y(_abc_17692_n1696) );
  AND2X2 AND2X2_4440 ( .A(_abc_17692_n10860), .B(_abc_17692_n10854), .Y(_abc_17692_n10861) );
  AND2X2 AND2X2_4441 ( .A(_abc_17692_n10863), .B(_abc_17692_n1830_bF_buf1), .Y(_abc_17692_n10864) );
  AND2X2 AND2X2_4442 ( .A(_abc_17692_n10864), .B(_abc_17692_n10862), .Y(_abc_17692_n10865) );
  AND2X2 AND2X2_4443 ( .A(_abc_17692_n10866), .B(_abc_17692_n10867), .Y(_abc_17692_n10868) );
  AND2X2 AND2X2_4444 ( .A(_abc_17692_n10868), .B(workunit1_18_), .Y(_abc_17692_n10870) );
  AND2X2 AND2X2_4445 ( .A(_abc_17692_n10871), .B(_abc_17692_n10869), .Y(_abc_17692_n10872) );
  AND2X2 AND2X2_4446 ( .A(_abc_17692_n10734), .B(_abc_17692_n10770), .Y(_abc_17692_n10875) );
  AND2X2 AND2X2_4447 ( .A(_abc_17692_n10879), .B(_abc_17692_n10877), .Y(_abc_17692_n10880) );
  AND2X2 AND2X2_4448 ( .A(_abc_17692_n10737), .B(_abc_17692_n10643), .Y(_abc_17692_n10881) );
  AND2X2 AND2X2_4449 ( .A(_abc_17692_n10883), .B(_abc_17692_n10876), .Y(_abc_17692_n10884) );
  AND2X2 AND2X2_445 ( .A(_abc_17692_n723), .B(sum_27_), .Y(_abc_17692_n1697) );
  AND2X2 AND2X2_4450 ( .A(_abc_17692_n10885), .B(_abc_17692_n10873), .Y(_abc_17692_n10886) );
  AND2X2 AND2X2_4451 ( .A(_abc_17692_n10888), .B(_abc_17692_n1846_bF_buf1), .Y(_abc_17692_n10889) );
  AND2X2 AND2X2_4452 ( .A(_abc_17692_n10889), .B(_abc_17692_n10887), .Y(_abc_17692_n10890) );
  AND2X2 AND2X2_4453 ( .A(_abc_17692_n10893), .B(state_14_bF_buf2), .Y(_abc_17692_n10894) );
  AND2X2 AND2X2_4454 ( .A(_abc_17692_n10690), .B(workunit1_17_), .Y(_abc_17692_n10896) );
  AND2X2 AND2X2_4455 ( .A(_abc_17692_n10898), .B(_abc_17692_n10897), .Y(_abc_17692_n10899) );
  AND2X2 AND2X2_4456 ( .A(_abc_17692_n10697), .B(_abc_17692_n10575), .Y(_abc_17692_n10901) );
  AND2X2 AND2X2_4457 ( .A(_abc_17692_n10584), .B(_abc_17692_n10901), .Y(_abc_17692_n10902) );
  AND2X2 AND2X2_4458 ( .A(_abc_17692_n10903), .B(_abc_17692_n10895), .Y(_abc_17692_n10905) );
  AND2X2 AND2X2_4459 ( .A(_abc_17692_n10906), .B(_abc_17692_n10904), .Y(_abc_17692_n10907) );
  AND2X2 AND2X2_446 ( .A(_abc_17692_n1652), .B(sum_26_), .Y(_abc_17692_n1699) );
  AND2X2 AND2X2_4460 ( .A(_abc_17692_n10706), .B(workunit1_17_), .Y(_abc_17692_n10909) );
  AND2X2 AND2X2_4461 ( .A(_abc_17692_n10712), .B(_abc_17692_n10505), .Y(_abc_17692_n10910) );
  AND2X2 AND2X2_4462 ( .A(_abc_17692_n10712), .B(_abc_17692_n10508), .Y(_abc_17692_n10912) );
  AND2X2 AND2X2_4463 ( .A(_abc_17692_n10517), .B(_abc_17692_n10912), .Y(_abc_17692_n10913) );
  AND2X2 AND2X2_4464 ( .A(_abc_17692_n10914), .B(_abc_17692_n10836), .Y(_abc_17692_n10916) );
  AND2X2 AND2X2_4465 ( .A(_abc_17692_n10917), .B(_abc_17692_n1877_bF_buf0), .Y(_abc_17692_n10918) );
  AND2X2 AND2X2_4466 ( .A(_abc_17692_n10918), .B(_abc_17692_n10915), .Y(_abc_17692_n10919) );
  AND2X2 AND2X2_4467 ( .A(_abc_17692_n10719), .B(workunit1_17_), .Y(_abc_17692_n10921) );
  AND2X2 AND2X2_4468 ( .A(_abc_17692_n10723), .B(_abc_17692_n10549), .Y(_abc_17692_n10922) );
  AND2X2 AND2X2_4469 ( .A(_abc_17692_n10723), .B(_abc_17692_n10552), .Y(_abc_17692_n10924) );
  AND2X2 AND2X2_447 ( .A(_abc_17692_n1698), .B(_abc_17692_n1655), .Y(_abc_17692_n1702) );
  AND2X2 AND2X2_4470 ( .A(_abc_17692_n10561), .B(_abc_17692_n10924), .Y(_abc_17692_n10925) );
  AND2X2 AND2X2_4471 ( .A(_abc_17692_n10926), .B(_abc_17692_n10920), .Y(_abc_17692_n10927) );
  AND2X2 AND2X2_4472 ( .A(_abc_17692_n10929), .B(_abc_17692_n1830_bF_buf0), .Y(_abc_17692_n10930) );
  AND2X2 AND2X2_4473 ( .A(_abc_17692_n10930), .B(_abc_17692_n10928), .Y(_abc_17692_n10931) );
  AND2X2 AND2X2_4474 ( .A(_abc_17692_n10733), .B(workunit1_17_), .Y(_abc_17692_n10932) );
  AND2X2 AND2X2_4475 ( .A(_abc_17692_n10934), .B(_abc_17692_n10933), .Y(_abc_17692_n10935) );
  AND2X2 AND2X2_4476 ( .A(_abc_17692_n10740), .B(_abc_17692_n10529), .Y(_abc_17692_n10937) );
  AND2X2 AND2X2_4477 ( .A(_abc_17692_n10540), .B(_abc_17692_n10937), .Y(_abc_17692_n10938) );
  AND2X2 AND2X2_4478 ( .A(_abc_17692_n10939), .B(_abc_17692_n10872), .Y(_abc_17692_n10941) );
  AND2X2 AND2X2_4479 ( .A(_abc_17692_n10942), .B(_abc_17692_n1846_bF_buf0), .Y(_abc_17692_n10943) );
  AND2X2 AND2X2_448 ( .A(_abc_17692_n1672), .B(_abc_17692_n1702), .Y(_abc_17692_n1703) );
  AND2X2 AND2X2_4480 ( .A(_abc_17692_n10943), .B(_abc_17692_n10940), .Y(_abc_17692_n10944) );
  AND2X2 AND2X2_4481 ( .A(_abc_17692_n10947), .B(state_10_bF_buf2), .Y(_abc_17692_n10948) );
  AND2X2 AND2X2_4482 ( .A(_abc_17692_n10948), .B(_abc_17692_n10908), .Y(_abc_17692_n10949) );
  AND2X2 AND2X2_4483 ( .A(_abc_17692_n8383_bF_buf1), .B(workunit1_18_), .Y(_abc_17692_n10950) );
  AND2X2 AND2X2_4484 ( .A(state_8_bF_buf9), .B(\data_in1[18] ), .Y(_abc_17692_n10951) );
  AND2X2 AND2X2_4485 ( .A(_abc_17692_n10957), .B(_abc_17692_n10958), .Y(_abc_17692_n10959) );
  AND2X2 AND2X2_4486 ( .A(_abc_17692_n10960), .B(workunit2_19_), .Y(_abc_17692_n10961) );
  AND2X2 AND2X2_4487 ( .A(_abc_17692_n10959), .B(_abc_17692_n5626), .Y(_abc_17692_n10963) );
  AND2X2 AND2X2_4488 ( .A(_abc_17692_n10962), .B(_abc_17692_n10964), .Y(_abc_17692_n10965) );
  AND2X2 AND2X2_4489 ( .A(_abc_17692_n10956), .B(_abc_17692_n10966), .Y(_abc_17692_n10967) );
  AND2X2 AND2X2_449 ( .A(_abc_17692_n1698), .B(_abc_17692_n1699), .Y(_abc_17692_n1705) );
  AND2X2 AND2X2_4490 ( .A(_abc_17692_n10955), .B(_abc_17692_n10965), .Y(_abc_17692_n10969) );
  AND2X2 AND2X2_4491 ( .A(_abc_17692_n10968), .B(_abc_17692_n10970), .Y(_abc_17692_n10971) );
  AND2X2 AND2X2_4492 ( .A(_abc_17692_n10972), .B(_abc_17692_n10974), .Y(_abc_17692_n10975) );
  AND2X2 AND2X2_4493 ( .A(_abc_17692_n10975), .B(_abc_17692_n4494), .Y(_abc_17692_n10976) );
  AND2X2 AND2X2_4494 ( .A(_abc_17692_n10978), .B(_abc_17692_n10977), .Y(_abc_17692_n10979) );
  AND2X2 AND2X2_4495 ( .A(_abc_17692_n10979), .B(workunit1_19_), .Y(_abc_17692_n10980) );
  AND2X2 AND2X2_4496 ( .A(_abc_17692_n10850), .B(workunit1_18_), .Y(_abc_17692_n10982) );
  AND2X2 AND2X2_4497 ( .A(_abc_17692_n10928), .B(_abc_17692_n10983), .Y(_abc_17692_n10984) );
  AND2X2 AND2X2_4498 ( .A(_abc_17692_n10988), .B(_abc_17692_n1830_bF_buf10), .Y(_abc_17692_n10989) );
  AND2X2 AND2X2_4499 ( .A(_abc_17692_n10989), .B(_abc_17692_n10985), .Y(_abc_17692_n10990) );
  AND2X2 AND2X2_45 ( .A(_abc_17692_n740), .B(_abc_17692_n739), .Y(data_out2_4__FF_INPUT) );
  AND2X2 AND2X2_450 ( .A(_abc_17692_n1706), .B(state_15_bF_buf2), .Y(_abc_17692_n1707) );
  AND2X2 AND2X2_4500 ( .A(_abc_17692_n10991), .B(_abc_17692_n10992), .Y(_abc_17692_n10993) );
  AND2X2 AND2X2_4501 ( .A(_abc_17692_n10995), .B(_abc_17692_n10996), .Y(_abc_17692_n10997) );
  AND2X2 AND2X2_4502 ( .A(_abc_17692_n10917), .B(_abc_17692_n10834), .Y(_abc_17692_n10998) );
  AND2X2 AND2X2_4503 ( .A(_abc_17692_n11002), .B(_abc_17692_n1877_bF_buf10), .Y(_abc_17692_n11003) );
  AND2X2 AND2X2_4504 ( .A(_abc_17692_n11003), .B(_abc_17692_n11000), .Y(_abc_17692_n11004) );
  AND2X2 AND2X2_4505 ( .A(_abc_17692_n11006), .B(_abc_17692_n11005), .Y(_abc_17692_n11007) );
  AND2X2 AND2X2_4506 ( .A(_abc_17692_n11009), .B(_abc_17692_n11010), .Y(_abc_17692_n11011) );
  AND2X2 AND2X2_4507 ( .A(_abc_17692_n11012), .B(_abc_17692_n11008), .Y(_abc_17692_n11013) );
  AND2X2 AND2X2_4508 ( .A(_abc_17692_n10942), .B(_abc_17692_n10871), .Y(_abc_17692_n11014) );
  AND2X2 AND2X2_4509 ( .A(_abc_17692_n11011), .B(_abc_17692_n4494), .Y(_abc_17692_n11017) );
  AND2X2 AND2X2_451 ( .A(_abc_17692_n1704), .B(_abc_17692_n1707), .Y(_abc_17692_n1708) );
  AND2X2 AND2X2_4510 ( .A(_abc_17692_n11007), .B(workunit1_19_), .Y(_abc_17692_n11018) );
  AND2X2 AND2X2_4511 ( .A(_abc_17692_n11020), .B(_abc_17692_n1846_bF_buf10), .Y(_abc_17692_n11021) );
  AND2X2 AND2X2_4512 ( .A(_abc_17692_n11021), .B(_abc_17692_n11016), .Y(_abc_17692_n11022) );
  AND2X2 AND2X2_4513 ( .A(_abc_17692_n11025), .B(_abc_17692_n11026), .Y(_abc_17692_n11027) );
  AND2X2 AND2X2_4514 ( .A(_abc_17692_n11027), .B(_abc_17692_n4494), .Y(_abc_17692_n11028) );
  AND2X2 AND2X2_4515 ( .A(_abc_17692_n11029), .B(_abc_17692_n11030), .Y(_abc_17692_n11031) );
  AND2X2 AND2X2_4516 ( .A(_abc_17692_n11031), .B(workunit1_19_), .Y(_abc_17692_n11032) );
  AND2X2 AND2X2_4517 ( .A(_abc_17692_n10906), .B(_abc_17692_n11034), .Y(_abc_17692_n11035) );
  AND2X2 AND2X2_4518 ( .A(_abc_17692_n11036), .B(_abc_17692_n11033), .Y(_abc_17692_n11037) );
  AND2X2 AND2X2_4519 ( .A(_abc_17692_n11038), .B(_abc_17692_n11039), .Y(_abc_17692_n11040) );
  AND2X2 AND2X2_452 ( .A(_abc_17692_n1708), .B(_abc_17692_n1701), .Y(_abc_17692_n1709) );
  AND2X2 AND2X2_4520 ( .A(_abc_17692_n11035), .B(_abc_17692_n11040), .Y(_abc_17692_n11041) );
  AND2X2 AND2X2_4521 ( .A(_abc_17692_n11042), .B(_abc_17692_n1863_bF_buf10), .Y(_abc_17692_n11043) );
  AND2X2 AND2X2_4522 ( .A(_abc_17692_n11044), .B(state_10_bF_buf1), .Y(_abc_17692_n11045) );
  AND2X2 AND2X2_4523 ( .A(_abc_17692_n10816), .B(workunit1_18_), .Y(_abc_17692_n11046) );
  AND2X2 AND2X2_4524 ( .A(_abc_17692_n11050), .B(_abc_17692_n1863_bF_buf9), .Y(_abc_17692_n11051) );
  AND2X2 AND2X2_4525 ( .A(_abc_17692_n11051), .B(_abc_17692_n11049), .Y(_abc_17692_n11052) );
  AND2X2 AND2X2_4526 ( .A(_abc_17692_n11053), .B(workunit1_18_), .Y(_abc_17692_n11054) );
  AND2X2 AND2X2_4527 ( .A(_abc_17692_n10844), .B(_abc_17692_n11055), .Y(_abc_17692_n11056) );
  AND2X2 AND2X2_4528 ( .A(_abc_17692_n11059), .B(_abc_17692_n1877_bF_buf9), .Y(_abc_17692_n11060) );
  AND2X2 AND2X2_4529 ( .A(_abc_17692_n11060), .B(_abc_17692_n11057), .Y(_abc_17692_n11061) );
  AND2X2 AND2X2_453 ( .A(_abc_17692_n1712), .B(delta_28_), .Y(_abc_17692_n1713) );
  AND2X2 AND2X2_4530 ( .A(_abc_17692_n11067), .B(_abc_17692_n1846_bF_buf9), .Y(_abc_17692_n11068) );
  AND2X2 AND2X2_4531 ( .A(_abc_17692_n11068), .B(_abc_17692_n11066), .Y(_abc_17692_n11069) );
  AND2X2 AND2X2_4532 ( .A(_abc_17692_n10862), .B(_abc_17692_n10851), .Y(_abc_17692_n11070) );
  AND2X2 AND2X2_4533 ( .A(_abc_17692_n11073), .B(_abc_17692_n1830_bF_buf9), .Y(_abc_17692_n11074) );
  AND2X2 AND2X2_4534 ( .A(_abc_17692_n11074), .B(_abc_17692_n11072), .Y(_abc_17692_n11075) );
  AND2X2 AND2X2_4535 ( .A(_abc_17692_n11078), .B(state_14_bF_buf1), .Y(_abc_17692_n11079) );
  AND2X2 AND2X2_4536 ( .A(_abc_17692_n8383_bF_buf0), .B(workunit1_19_), .Y(_abc_17692_n11080) );
  AND2X2 AND2X2_4537 ( .A(state_8_bF_buf8), .B(\data_in1[19] ), .Y(_abc_17692_n11081) );
  AND2X2 AND2X2_4538 ( .A(_abc_17692_n10807), .B(_abc_17692_n10965), .Y(_abc_17692_n11085) );
  AND2X2 AND2X2_4539 ( .A(_abc_17692_n10797), .B(_abc_17692_n11085), .Y(_abc_17692_n11086) );
  AND2X2 AND2X2_454 ( .A(delta_27_), .B(sum_27_), .Y(_abc_17692_n1717) );
  AND2X2 AND2X2_4540 ( .A(_abc_17692_n11085), .B(_abc_17692_n10796), .Y(_abc_17692_n11089) );
  AND2X2 AND2X2_4541 ( .A(_abc_17692_n11091), .B(_abc_17692_n10962), .Y(_abc_17692_n11092) );
  AND2X2 AND2X2_4542 ( .A(_abc_17692_n11090), .B(_abc_17692_n11093), .Y(_abc_17692_n11094) );
  AND2X2 AND2X2_4543 ( .A(_abc_17692_n11088), .B(_abc_17692_n11094), .Y(_abc_17692_n11095) );
  AND2X2 AND2X2_4544 ( .A(_abc_17692_n11096), .B(_abc_17692_n11097), .Y(_abc_17692_n11098) );
  AND2X2 AND2X2_4545 ( .A(_abc_17692_n11099), .B(workunit2_20_), .Y(_abc_17692_n11100) );
  AND2X2 AND2X2_4546 ( .A(_abc_17692_n11098), .B(_abc_17692_n5769), .Y(_abc_17692_n11101) );
  AND2X2 AND2X2_4547 ( .A(_abc_17692_n11095), .B(_abc_17692_n11102), .Y(_abc_17692_n11103) );
  AND2X2 AND2X2_4548 ( .A(_abc_17692_n10497), .B(_abc_17692_n11086), .Y(_abc_17692_n11104) );
  AND2X2 AND2X2_4549 ( .A(_abc_17692_n11106), .B(_abc_17692_n11107), .Y(_abc_17692_n11108) );
  AND2X2 AND2X2_455 ( .A(_abc_17692_n1691), .B(_abc_17692_n1719), .Y(_abc_17692_n1720) );
  AND2X2 AND2X2_4550 ( .A(_abc_17692_n11112), .B(_abc_17692_n11111), .Y(_abc_17692_n11113) );
  AND2X2 AND2X2_4551 ( .A(_abc_17692_n11114), .B(_abc_17692_n4730), .Y(_abc_17692_n11115) );
  AND2X2 AND2X2_4552 ( .A(_abc_17692_n11113), .B(workunit1_20_), .Y(_abc_17692_n11116) );
  AND2X2 AND2X2_4553 ( .A(_abc_17692_n11040), .B(_abc_17692_n10895), .Y(_abc_17692_n11119) );
  AND2X2 AND2X2_4554 ( .A(_abc_17692_n11119), .B(_abc_17692_n10901), .Y(_abc_17692_n11120) );
  AND2X2 AND2X2_4555 ( .A(_abc_17692_n10584), .B(_abc_17692_n11120), .Y(_abc_17692_n11121) );
  AND2X2 AND2X2_4556 ( .A(_abc_17692_n11038), .B(_abc_17692_n10818), .Y(_abc_17692_n11124) );
  AND2X2 AND2X2_4557 ( .A(_abc_17692_n11123), .B(_abc_17692_n11126), .Y(_abc_17692_n11127) );
  AND2X2 AND2X2_4558 ( .A(_abc_17692_n11129), .B(_abc_17692_n11118), .Y(_abc_17692_n11130) );
  AND2X2 AND2X2_4559 ( .A(_abc_17692_n11131), .B(_abc_17692_n11132), .Y(_abc_17692_n11133) );
  AND2X2 AND2X2_456 ( .A(_abc_17692_n1724), .B(state_3_bF_buf1), .Y(_abc_17692_n1725) );
  AND2X2 AND2X2_4560 ( .A(_abc_17692_n11136), .B(_abc_17692_n11135), .Y(_abc_17692_n11137) );
  AND2X2 AND2X2_4561 ( .A(_abc_17692_n11137), .B(workunit1_20_), .Y(_abc_17692_n11138) );
  AND2X2 AND2X2_4562 ( .A(_abc_17692_n11139), .B(_abc_17692_n11140), .Y(_abc_17692_n11141) );
  AND2X2 AND2X2_4563 ( .A(_abc_17692_n10997), .B(_abc_17692_n10836), .Y(_abc_17692_n11142) );
  AND2X2 AND2X2_4564 ( .A(_abc_17692_n11142), .B(_abc_17692_n10911), .Y(_abc_17692_n11143) );
  AND2X2 AND2X2_4565 ( .A(_abc_17692_n11145), .B(_abc_17692_n10996), .Y(_abc_17692_n11146) );
  AND2X2 AND2X2_4566 ( .A(_abc_17692_n11142), .B(_abc_17692_n10912), .Y(_abc_17692_n11149) );
  AND2X2 AND2X2_4567 ( .A(_abc_17692_n10517), .B(_abc_17692_n11149), .Y(_abc_17692_n11150) );
  AND2X2 AND2X2_4568 ( .A(_abc_17692_n11151), .B(_abc_17692_n11141), .Y(_abc_17692_n11153) );
  AND2X2 AND2X2_4569 ( .A(_abc_17692_n11154), .B(_abc_17692_n1877_bF_buf8), .Y(_abc_17692_n11155) );
  AND2X2 AND2X2_457 ( .A(_abc_17692_n1725), .B(_abc_17692_n1722), .Y(_abc_17692_n1726) );
  AND2X2 AND2X2_4570 ( .A(_abc_17692_n11155), .B(_abc_17692_n11152), .Y(_abc_17692_n11156) );
  AND2X2 AND2X2_4571 ( .A(_abc_17692_n11157), .B(_abc_17692_n11158), .Y(_abc_17692_n11159) );
  AND2X2 AND2X2_4572 ( .A(_abc_17692_n11160), .B(_abc_17692_n4730), .Y(_abc_17692_n11161) );
  AND2X2 AND2X2_4573 ( .A(_abc_17692_n11159), .B(workunit1_20_), .Y(_abc_17692_n11162) );
  AND2X2 AND2X2_4574 ( .A(_abc_17692_n10986), .B(_abc_17692_n10920), .Y(_abc_17692_n11165) );
  AND2X2 AND2X2_4575 ( .A(_abc_17692_n11165), .B(_abc_17692_n10923), .Y(_abc_17692_n11166) );
  AND2X2 AND2X2_4576 ( .A(_abc_17692_n10986), .B(_abc_17692_n10982), .Y(_abc_17692_n11167) );
  AND2X2 AND2X2_4577 ( .A(_abc_17692_n11165), .B(_abc_17692_n10924), .Y(_abc_17692_n11170) );
  AND2X2 AND2X2_4578 ( .A(_abc_17692_n10561), .B(_abc_17692_n11170), .Y(_abc_17692_n11171) );
  AND2X2 AND2X2_4579 ( .A(_abc_17692_n11172), .B(_abc_17692_n11164), .Y(_abc_17692_n11173) );
  AND2X2 AND2X2_458 ( .A(_abc_17692_n723), .B(sum_28_), .Y(_abc_17692_n1727) );
  AND2X2 AND2X2_4580 ( .A(_abc_17692_n11175), .B(_abc_17692_n1830_bF_buf8), .Y(_abc_17692_n11176) );
  AND2X2 AND2X2_4581 ( .A(_abc_17692_n11176), .B(_abc_17692_n11174), .Y(_abc_17692_n11177) );
  AND2X2 AND2X2_4582 ( .A(_abc_17692_n11178), .B(_abc_17692_n11179), .Y(_abc_17692_n11180) );
  AND2X2 AND2X2_4583 ( .A(_abc_17692_n11181), .B(_abc_17692_n4730), .Y(_abc_17692_n11182) );
  AND2X2 AND2X2_4584 ( .A(_abc_17692_n11180), .B(workunit1_20_), .Y(_abc_17692_n11183) );
  AND2X2 AND2X2_4585 ( .A(_abc_17692_n11188), .B(_abc_17692_n11008), .Y(_abc_17692_n11189) );
  AND2X2 AND2X2_4586 ( .A(_abc_17692_n11187), .B(_abc_17692_n11190), .Y(_abc_17692_n11191) );
  AND2X2 AND2X2_4587 ( .A(_abc_17692_n11192), .B(_abc_17692_n10937), .Y(_abc_17692_n11193) );
  AND2X2 AND2X2_4588 ( .A(_abc_17692_n11195), .B(_abc_17692_n11191), .Y(_abc_17692_n11196) );
  AND2X2 AND2X2_4589 ( .A(_abc_17692_n11197), .B(_abc_17692_n11185), .Y(_abc_17692_n11198) );
  AND2X2 AND2X2_459 ( .A(_abc_17692_n1706), .B(_abc_17692_n1684), .Y(_abc_17692_n1728) );
  AND2X2 AND2X2_4590 ( .A(_abc_17692_n11200), .B(_abc_17692_n1846_bF_buf8), .Y(_abc_17692_n11201) );
  AND2X2 AND2X2_4591 ( .A(_abc_17692_n11201), .B(_abc_17692_n11199), .Y(_abc_17692_n11202) );
  AND2X2 AND2X2_4592 ( .A(_abc_17692_n11205), .B(state_10_bF_buf0), .Y(_abc_17692_n11206) );
  AND2X2 AND2X2_4593 ( .A(_abc_17692_n11134), .B(_abc_17692_n11206), .Y(_abc_17692_n11207) );
  AND2X2 AND2X2_4594 ( .A(_abc_17692_n11033), .B(_abc_17692_n10819), .Y(_abc_17692_n11208) );
  AND2X2 AND2X2_4595 ( .A(_abc_17692_n11208), .B(_abc_17692_n10821), .Y(_abc_17692_n11209) );
  AND2X2 AND2X2_4596 ( .A(_abc_17692_n11033), .B(_abc_17692_n11046), .Y(_abc_17692_n11210) );
  AND2X2 AND2X2_4597 ( .A(_abc_17692_n11027), .B(workunit1_19_), .Y(_abc_17692_n11211) );
  AND2X2 AND2X2_4598 ( .A(_abc_17692_n11208), .B(_abc_17692_n10822), .Y(_abc_17692_n11214) );
  AND2X2 AND2X2_4599 ( .A(_abc_17692_n10602), .B(_abc_17692_n11214), .Y(_abc_17692_n11215) );
  AND2X2 AND2X2_46 ( .A(_abc_17692_n743), .B(_abc_17692_n742), .Y(data_out2_5__FF_INPUT) );
  AND2X2 AND2X2_460 ( .A(_abc_17692_n1730), .B(_abc_17692_n1723), .Y(_abc_17692_n1731) );
  AND2X2 AND2X2_4600 ( .A(_abc_17692_n11216), .B(_abc_17692_n11117), .Y(_abc_17692_n11218) );
  AND2X2 AND2X2_4601 ( .A(_abc_17692_n11219), .B(_abc_17692_n1863_bF_buf7), .Y(_abc_17692_n11220) );
  AND2X2 AND2X2_4602 ( .A(_abc_17692_n11220), .B(_abc_17692_n11217), .Y(_abc_17692_n11221) );
  AND2X2 AND2X2_4603 ( .A(_abc_17692_n10993), .B(workunit1_19_), .Y(_abc_17692_n11226) );
  AND2X2 AND2X2_4604 ( .A(_abc_17692_n11228), .B(_abc_17692_n11227), .Y(_abc_17692_n11229) );
  AND2X2 AND2X2_4605 ( .A(_abc_17692_n11225), .B(_abc_17692_n11229), .Y(_abc_17692_n11230) );
  AND2X2 AND2X2_4606 ( .A(_abc_17692_n11232), .B(_abc_17692_n10840), .Y(_abc_17692_n11233) );
  AND2X2 AND2X2_4607 ( .A(_abc_17692_n10622), .B(_abc_17692_n11233), .Y(_abc_17692_n11234) );
  AND2X2 AND2X2_4608 ( .A(_abc_17692_n11235), .B(_abc_17692_n11222), .Y(_abc_17692_n11236) );
  AND2X2 AND2X2_4609 ( .A(_abc_17692_n11238), .B(_abc_17692_n1877_bF_buf7), .Y(_abc_17692_n11239) );
  AND2X2 AND2X2_461 ( .A(_abc_17692_n1733), .B(state_15_bF_buf1), .Y(_abc_17692_n1734) );
  AND2X2 AND2X2_4610 ( .A(_abc_17692_n11239), .B(_abc_17692_n11237), .Y(_abc_17692_n11240) );
  AND2X2 AND2X2_4611 ( .A(_abc_17692_n11011), .B(workunit1_19_), .Y(_abc_17692_n11243) );
  AND2X2 AND2X2_4612 ( .A(_abc_17692_n11245), .B(_abc_17692_n11244), .Y(_abc_17692_n11246) );
  AND2X2 AND2X2_4613 ( .A(_abc_17692_n11242), .B(_abc_17692_n11246), .Y(_abc_17692_n11247) );
  AND2X2 AND2X2_4614 ( .A(_abc_17692_n10654), .B(_abc_17692_n11250), .Y(_abc_17692_n11251) );
  AND2X2 AND2X2_4615 ( .A(_abc_17692_n11252), .B(_abc_17692_n11184), .Y(_abc_17692_n11254) );
  AND2X2 AND2X2_4616 ( .A(_abc_17692_n11255), .B(_abc_17692_n1846_bF_buf7), .Y(_abc_17692_n11256) );
  AND2X2 AND2X2_4617 ( .A(_abc_17692_n11256), .B(_abc_17692_n11253), .Y(_abc_17692_n11257) );
  AND2X2 AND2X2_4618 ( .A(_abc_17692_n10981), .B(_abc_17692_n10854), .Y(_abc_17692_n11258) );
  AND2X2 AND2X2_4619 ( .A(_abc_17692_n11258), .B(_abc_17692_n10857), .Y(_abc_17692_n11259) );
  AND2X2 AND2X2_462 ( .A(_abc_17692_n1734), .B(_abc_17692_n1732), .Y(_abc_17692_n1735) );
  AND2X2 AND2X2_4620 ( .A(_abc_17692_n10975), .B(workunit1_19_), .Y(_abc_17692_n11260) );
  AND2X2 AND2X2_4621 ( .A(_abc_17692_n10981), .B(_abc_17692_n11261), .Y(_abc_17692_n11262) );
  AND2X2 AND2X2_4622 ( .A(_abc_17692_n11268), .B(_abc_17692_n10632), .Y(_abc_17692_n11269) );
  AND2X2 AND2X2_4623 ( .A(_abc_17692_n11272), .B(_abc_17692_n11269), .Y(_abc_17692_n11273) );
  AND2X2 AND2X2_4624 ( .A(_abc_17692_n11258), .B(_abc_17692_n10858), .Y(_abc_17692_n11274) );
  AND2X2 AND2X2_4625 ( .A(_abc_17692_n11276), .B(_abc_17692_n11265), .Y(_abc_17692_n11277) );
  AND2X2 AND2X2_4626 ( .A(_abc_17692_n11278), .B(_abc_17692_n11163), .Y(_abc_17692_n11279) );
  AND2X2 AND2X2_4627 ( .A(_abc_17692_n11281), .B(_abc_17692_n1830_bF_buf7), .Y(_abc_17692_n11282) );
  AND2X2 AND2X2_4628 ( .A(_abc_17692_n11282), .B(_abc_17692_n11280), .Y(_abc_17692_n11283) );
  AND2X2 AND2X2_4629 ( .A(_abc_17692_n11286), .B(state_14_bF_buf0), .Y(_abc_17692_n11287) );
  AND2X2 AND2X2_463 ( .A(_abc_17692_n1738), .B(delta_29_), .Y(_abc_17692_n1739) );
  AND2X2 AND2X2_4630 ( .A(_abc_17692_n8383_bF_buf4), .B(workunit1_20_), .Y(_abc_17692_n11288) );
  AND2X2 AND2X2_4631 ( .A(state_8_bF_buf7), .B(\data_in1[20] ), .Y(_abc_17692_n11289) );
  AND2X2 AND2X2_4632 ( .A(_abc_17692_n11294), .B(_abc_17692_n11295), .Y(_abc_17692_n11296) );
  AND2X2 AND2X2_4633 ( .A(_abc_17692_n11297), .B(workunit2_21_), .Y(_abc_17692_n11298) );
  AND2X2 AND2X2_4634 ( .A(_abc_17692_n11296), .B(_abc_17692_n6095), .Y(_abc_17692_n11300) );
  AND2X2 AND2X2_4635 ( .A(_abc_17692_n11299), .B(_abc_17692_n11301), .Y(_abc_17692_n11302) );
  AND2X2 AND2X2_4636 ( .A(_abc_17692_n11293), .B(_abc_17692_n11303), .Y(_abc_17692_n11304) );
  AND2X2 AND2X2_4637 ( .A(_abc_17692_n11305), .B(_abc_17692_n11306), .Y(_abc_17692_n11307) );
  AND2X2 AND2X2_4638 ( .A(_abc_17692_n11308), .B(_abc_17692_n11310), .Y(_abc_17692_n11311) );
  AND2X2 AND2X2_4639 ( .A(_abc_17692_n11311), .B(workunit1_21_), .Y(_abc_17692_n11312) );
  AND2X2 AND2X2_464 ( .A(_abc_17692_n1741), .B(sum_29_), .Y(_abc_17692_n1742) );
  AND2X2 AND2X2_4640 ( .A(_abc_17692_n11313), .B(_abc_17692_n4926), .Y(_abc_17692_n11314) );
  AND2X2 AND2X2_4641 ( .A(_abc_17692_n11154), .B(_abc_17692_n11139), .Y(_abc_17692_n11316) );
  AND2X2 AND2X2_4642 ( .A(_abc_17692_n11320), .B(_abc_17692_n1877_bF_buf6), .Y(_abc_17692_n11321) );
  AND2X2 AND2X2_4643 ( .A(_abc_17692_n11321), .B(_abc_17692_n11318), .Y(_abc_17692_n11322) );
  AND2X2 AND2X2_4644 ( .A(_abc_17692_n11324), .B(_abc_17692_n11323), .Y(_abc_17692_n11325) );
  AND2X2 AND2X2_4645 ( .A(_abc_17692_n11325), .B(workunit1_21_), .Y(_abc_17692_n11326) );
  AND2X2 AND2X2_4646 ( .A(_abc_17692_n11327), .B(_abc_17692_n4926), .Y(_abc_17692_n11328) );
  AND2X2 AND2X2_4647 ( .A(_abc_17692_n11329), .B(_abc_17692_n11162), .Y(_abc_17692_n11332) );
  AND2X2 AND2X2_4648 ( .A(_abc_17692_n11331), .B(_abc_17692_n11333), .Y(_abc_17692_n11334) );
  AND2X2 AND2X2_4649 ( .A(_abc_17692_n11336), .B(_abc_17692_n1830_bF_buf6), .Y(_abc_17692_n11337) );
  AND2X2 AND2X2_465 ( .A(_abc_17692_n1740), .B(_abc_17692_n1743), .Y(_abc_17692_n1744) );
  AND2X2 AND2X2_4650 ( .A(_abc_17692_n11334), .B(_abc_17692_n11337), .Y(_abc_17692_n11338) );
  AND2X2 AND2X2_4651 ( .A(_abc_17692_n11339), .B(_abc_17692_n11340), .Y(_abc_17692_n11341) );
  AND2X2 AND2X2_4652 ( .A(_abc_17692_n11344), .B(_abc_17692_n11343), .Y(_abc_17692_n11345) );
  AND2X2 AND2X2_4653 ( .A(_abc_17692_n11342), .B(_abc_17692_n11346), .Y(_abc_17692_n11347) );
  AND2X2 AND2X2_4654 ( .A(_abc_17692_n11199), .B(_abc_17692_n11349), .Y(_abc_17692_n11350) );
  AND2X2 AND2X2_4655 ( .A(_abc_17692_n11353), .B(_abc_17692_n1846_bF_buf6), .Y(_abc_17692_n11354) );
  AND2X2 AND2X2_4656 ( .A(_abc_17692_n11354), .B(_abc_17692_n11352), .Y(_abc_17692_n11355) );
  AND2X2 AND2X2_4657 ( .A(_abc_17692_n6176), .B(_abc_17692_n11309), .Y(_abc_17692_n11358) );
  AND2X2 AND2X2_4658 ( .A(_abc_17692_n6174), .B(_abc_17692_n11307), .Y(_abc_17692_n11359) );
  AND2X2 AND2X2_4659 ( .A(_abc_17692_n11361), .B(workunit1_21_), .Y(_abc_17692_n11362) );
  AND2X2 AND2X2_466 ( .A(delta_28_), .B(sum_28_), .Y(_abc_17692_n1746) );
  AND2X2 AND2X2_4660 ( .A(_abc_17692_n11360), .B(_abc_17692_n4926), .Y(_abc_17692_n11363) );
  AND2X2 AND2X2_4661 ( .A(_abc_17692_n11131), .B(_abc_17692_n11365), .Y(_abc_17692_n11366) );
  AND2X2 AND2X2_4662 ( .A(_abc_17692_n11366), .B(_abc_17692_n11364), .Y(_abc_17692_n11367) );
  AND2X2 AND2X2_4663 ( .A(_abc_17692_n11369), .B(_abc_17692_n11368), .Y(_abc_17692_n11370) );
  AND2X2 AND2X2_4664 ( .A(_abc_17692_n11371), .B(_abc_17692_n1863_bF_buf6), .Y(_abc_17692_n11372) );
  AND2X2 AND2X2_4665 ( .A(_abc_17692_n11373), .B(state_10_bF_buf4), .Y(_abc_17692_n11374) );
  AND2X2 AND2X2_4666 ( .A(_abc_17692_n11114), .B(workunit1_20_), .Y(_abc_17692_n11375) );
  AND2X2 AND2X2_4667 ( .A(_abc_17692_n11376), .B(_abc_17692_n11364), .Y(_abc_17692_n11377) );
  AND2X2 AND2X2_4668 ( .A(_abc_17692_n11378), .B(_abc_17692_n11368), .Y(_abc_17692_n11379) );
  AND2X2 AND2X2_4669 ( .A(_abc_17692_n11380), .B(_abc_17692_n1863_bF_buf5), .Y(_abc_17692_n11381) );
  AND2X2 AND2X2_467 ( .A(_abc_17692_n1724), .B(_abc_17692_n1747), .Y(_abc_17692_n1748) );
  AND2X2 AND2X2_4670 ( .A(_abc_17692_n11382), .B(workunit1_20_), .Y(_abc_17692_n11383) );
  AND2X2 AND2X2_4671 ( .A(_abc_17692_n11237), .B(_abc_17692_n11384), .Y(_abc_17692_n11385) );
  AND2X2 AND2X2_4672 ( .A(_abc_17692_n11388), .B(_abc_17692_n1877_bF_buf5), .Y(_abc_17692_n11389) );
  AND2X2 AND2X2_4673 ( .A(_abc_17692_n11389), .B(_abc_17692_n11387), .Y(_abc_17692_n11390) );
  AND2X2 AND2X2_4674 ( .A(_abc_17692_n11181), .B(workunit1_20_), .Y(_abc_17692_n11391) );
  AND2X2 AND2X2_4675 ( .A(_abc_17692_n11255), .B(_abc_17692_n11392), .Y(_abc_17692_n11393) );
  AND2X2 AND2X2_4676 ( .A(_abc_17692_n11396), .B(_abc_17692_n1846_bF_buf5), .Y(_abc_17692_n11397) );
  AND2X2 AND2X2_4677 ( .A(_abc_17692_n11397), .B(_abc_17692_n11395), .Y(_abc_17692_n11398) );
  AND2X2 AND2X2_4678 ( .A(_abc_17692_n11160), .B(workunit1_20_), .Y(_abc_17692_n11399) );
  AND2X2 AND2X2_4679 ( .A(_abc_17692_n11280), .B(_abc_17692_n11400), .Y(_abc_17692_n11401) );
  AND2X2 AND2X2_468 ( .A(_abc_17692_n1750), .B(_abc_17692_n1751), .Y(_abc_17692_n1752) );
  AND2X2 AND2X2_4680 ( .A(_abc_17692_n11404), .B(_abc_17692_n1830_bF_buf5), .Y(_abc_17692_n11405) );
  AND2X2 AND2X2_4681 ( .A(_abc_17692_n11405), .B(_abc_17692_n11402), .Y(_abc_17692_n11406) );
  AND2X2 AND2X2_4682 ( .A(_abc_17692_n11409), .B(state_14_bF_buf4), .Y(_abc_17692_n11410) );
  AND2X2 AND2X2_4683 ( .A(_abc_17692_n8383_bF_buf3), .B(workunit1_21_), .Y(_abc_17692_n11411) );
  AND2X2 AND2X2_4684 ( .A(state_8_bF_buf6), .B(\data_in1[21] ), .Y(_abc_17692_n11412) );
  AND2X2 AND2X2_4685 ( .A(_abc_17692_n11107), .B(_abc_17692_n11302), .Y(_abc_17692_n11416) );
  AND2X2 AND2X2_4686 ( .A(_abc_17692_n11301), .B(_abc_17692_n11100), .Y(_abc_17692_n11419) );
  AND2X2 AND2X2_4687 ( .A(_abc_17692_n11418), .B(_abc_17692_n11421), .Y(_abc_17692_n11422) );
  AND2X2 AND2X2_4688 ( .A(_abc_17692_n11423), .B(_abc_17692_n11424), .Y(_abc_17692_n11425) );
  AND2X2 AND2X2_4689 ( .A(_abc_17692_n11426), .B(workunit2_22_), .Y(_abc_17692_n11427) );
  AND2X2 AND2X2_469 ( .A(_abc_17692_n1752), .B(state_3_bF_buf0), .Y(_abc_17692_n1753) );
  AND2X2 AND2X2_4690 ( .A(_abc_17692_n11425), .B(_abc_17692_n6293), .Y(_abc_17692_n11428) );
  AND2X2 AND2X2_4691 ( .A(_abc_17692_n11422), .B(_abc_17692_n11429), .Y(_abc_17692_n11430) );
  AND2X2 AND2X2_4692 ( .A(_abc_17692_n11106), .B(_abc_17692_n11416), .Y(_abc_17692_n11431) );
  AND2X2 AND2X2_4693 ( .A(_abc_17692_n11432), .B(_abc_17692_n11433), .Y(_abc_17692_n11434) );
  AND2X2 AND2X2_4694 ( .A(_abc_17692_n11438), .B(_abc_17692_n11437), .Y(_abc_17692_n11439) );
  AND2X2 AND2X2_4695 ( .A(_abc_17692_n11439), .B(workunit1_22_), .Y(_abc_17692_n11440) );
  AND2X2 AND2X2_4696 ( .A(_abc_17692_n11441), .B(_abc_17692_n11442), .Y(_abc_17692_n11443) );
  AND2X2 AND2X2_4697 ( .A(_abc_17692_n11313), .B(workunit1_21_), .Y(_abc_17692_n11444) );
  AND2X2 AND2X2_4698 ( .A(_abc_17692_n11315), .B(_abc_17692_n11138), .Y(_abc_17692_n11445) );
  AND2X2 AND2X2_4699 ( .A(_abc_17692_n11315), .B(_abc_17692_n11141), .Y(_abc_17692_n11447) );
  AND2X2 AND2X2_47 ( .A(_abc_17692_n746), .B(_abc_17692_n745), .Y(data_out2_6__FF_INPUT) );
  AND2X2 AND2X2_470 ( .A(_abc_17692_n723), .B(sum_29_), .Y(_abc_17692_n1754) );
  AND2X2 AND2X2_4700 ( .A(_abc_17692_n11151), .B(_abc_17692_n11447), .Y(_abc_17692_n11448) );
  AND2X2 AND2X2_4701 ( .A(_abc_17692_n11449), .B(_abc_17692_n11443), .Y(_abc_17692_n11450) );
  AND2X2 AND2X2_4702 ( .A(_abc_17692_n11452), .B(_abc_17692_n1877_bF_buf4), .Y(_abc_17692_n11453) );
  AND2X2 AND2X2_4703 ( .A(_abc_17692_n11453), .B(_abc_17692_n11451), .Y(_abc_17692_n11454) );
  AND2X2 AND2X2_4704 ( .A(_abc_17692_n11455), .B(_abc_17692_n11456), .Y(_abc_17692_n11457) );
  AND2X2 AND2X2_4705 ( .A(_abc_17692_n11458), .B(workunit1_22_), .Y(_abc_17692_n11459) );
  AND2X2 AND2X2_4706 ( .A(_abc_17692_n11457), .B(_abc_17692_n5205), .Y(_abc_17692_n11460) );
  AND2X2 AND2X2_4707 ( .A(_abc_17692_n11341), .B(workunit1_21_), .Y(_abc_17692_n11462) );
  AND2X2 AND2X2_4708 ( .A(_abc_17692_n11464), .B(_abc_17692_n11463), .Y(_abc_17692_n11465) );
  AND2X2 AND2X2_4709 ( .A(_abc_17692_n11197), .B(_abc_17692_n11468), .Y(_abc_17692_n11469) );
  AND2X2 AND2X2_471 ( .A(_abc_17692_n1758_1), .B(_abc_17692_n1756), .Y(_abc_17692_n1759) );
  AND2X2 AND2X2_4710 ( .A(_abc_17692_n11470), .B(_abc_17692_n11461), .Y(_abc_17692_n11471) );
  AND2X2 AND2X2_4711 ( .A(_abc_17692_n11473), .B(_abc_17692_n1846_bF_buf4), .Y(_abc_17692_n11474) );
  AND2X2 AND2X2_4712 ( .A(_abc_17692_n11474), .B(_abc_17692_n11472), .Y(_abc_17692_n11475) );
  AND2X2 AND2X2_4713 ( .A(_abc_17692_n6313), .B(_abc_17692_n11435), .Y(_abc_17692_n11476) );
  AND2X2 AND2X2_4714 ( .A(_abc_17692_n11436), .B(_abc_17692_n6311), .Y(_abc_17692_n11477) );
  AND2X2 AND2X2_4715 ( .A(_abc_17692_n11480), .B(_abc_17692_n11481), .Y(_abc_17692_n11482) );
  AND2X2 AND2X2_4716 ( .A(_abc_17692_n11327), .B(workunit1_21_), .Y(_abc_17692_n11484) );
  AND2X2 AND2X2_4717 ( .A(_abc_17692_n11331), .B(_abc_17692_n11486), .Y(_abc_17692_n11487) );
  AND2X2 AND2X2_4718 ( .A(_abc_17692_n11490), .B(_abc_17692_n1830_bF_buf4), .Y(_abc_17692_n11491) );
  AND2X2 AND2X2_4719 ( .A(_abc_17692_n11491), .B(_abc_17692_n11489), .Y(_abc_17692_n11492) );
  AND2X2 AND2X2_472 ( .A(_abc_17692_n1759), .B(state_15_bF_buf0), .Y(_abc_17692_n1760) );
  AND2X2 AND2X2_4720 ( .A(_abc_17692_n6391), .B(_abc_17692_n11435), .Y(_abc_17692_n11495) );
  AND2X2 AND2X2_4721 ( .A(_abc_17692_n6389), .B(_abc_17692_n11436), .Y(_abc_17692_n11496) );
  AND2X2 AND2X2_4722 ( .A(_abc_17692_n11499), .B(_abc_17692_n11500), .Y(_abc_17692_n11501) );
  AND2X2 AND2X2_4723 ( .A(_abc_17692_n11360), .B(workunit1_21_), .Y(_abc_17692_n11503) );
  AND2X2 AND2X2_4724 ( .A(_abc_17692_n11364), .B(_abc_17692_n11116), .Y(_abc_17692_n11504) );
  AND2X2 AND2X2_4725 ( .A(_abc_17692_n11364), .B(_abc_17692_n11118), .Y(_abc_17692_n11506) );
  AND2X2 AND2X2_4726 ( .A(_abc_17692_n11129), .B(_abc_17692_n11506), .Y(_abc_17692_n11507) );
  AND2X2 AND2X2_4727 ( .A(_abc_17692_n11508), .B(_abc_17692_n11502), .Y(_abc_17692_n11509) );
  AND2X2 AND2X2_4728 ( .A(_abc_17692_n11511), .B(_abc_17692_n1863_bF_buf4), .Y(_abc_17692_n11512) );
  AND2X2 AND2X2_4729 ( .A(_abc_17692_n11512), .B(_abc_17692_n11510), .Y(_abc_17692_n11513) );
  AND2X2 AND2X2_473 ( .A(delta_30_), .B(sum_30_), .Y(_abc_17692_n1763) );
  AND2X2 AND2X2_4730 ( .A(_abc_17692_n11514), .B(state_10_bF_buf3), .Y(_abc_17692_n11515) );
  AND2X2 AND2X2_4731 ( .A(_abc_17692_n11517), .B(_abc_17692_n11516), .Y(_abc_17692_n11518) );
  AND2X2 AND2X2_4732 ( .A(_abc_17692_n11216), .B(_abc_17692_n11520), .Y(_abc_17692_n11521) );
  AND2X2 AND2X2_4733 ( .A(_abc_17692_n11522), .B(_abc_17692_n11501), .Y(_abc_17692_n11523) );
  AND2X2 AND2X2_4734 ( .A(_abc_17692_n11525), .B(_abc_17692_n1863_bF_buf3), .Y(_abc_17692_n11526) );
  AND2X2 AND2X2_4735 ( .A(_abc_17692_n11526), .B(_abc_17692_n11524), .Y(_abc_17692_n11527) );
  AND2X2 AND2X2_4736 ( .A(_abc_17692_n11235), .B(_abc_17692_n11530), .Y(_abc_17692_n11531) );
  AND2X2 AND2X2_4737 ( .A(_abc_17692_n11532), .B(_abc_17692_n11384), .Y(_abc_17692_n11533) );
  AND2X2 AND2X2_4738 ( .A(_abc_17692_n11536), .B(_abc_17692_n11528), .Y(_abc_17692_n11537) );
  AND2X2 AND2X2_4739 ( .A(_abc_17692_n11539), .B(_abc_17692_n1877_bF_buf3), .Y(_abc_17692_n11540) );
  AND2X2 AND2X2_474 ( .A(_abc_17692_n1764), .B(_abc_17692_n1765), .Y(_abc_17692_n1766) );
  AND2X2 AND2X2_4740 ( .A(_abc_17692_n11540), .B(_abc_17692_n11538), .Y(_abc_17692_n11541) );
  AND2X2 AND2X2_4741 ( .A(_abc_17692_n11252), .B(_abc_17692_n11544), .Y(_abc_17692_n11545) );
  AND2X2 AND2X2_4742 ( .A(_abc_17692_n11342), .B(_abc_17692_n11392), .Y(_abc_17692_n11547) );
  AND2X2 AND2X2_4743 ( .A(_abc_17692_n11550), .B(_abc_17692_n11542), .Y(_abc_17692_n11552) );
  AND2X2 AND2X2_4744 ( .A(_abc_17692_n11553), .B(_abc_17692_n1846_bF_buf3), .Y(_abc_17692_n11554) );
  AND2X2 AND2X2_4745 ( .A(_abc_17692_n11554), .B(_abc_17692_n11551), .Y(_abc_17692_n11555) );
  AND2X2 AND2X2_4746 ( .A(_abc_17692_n11556), .B(_abc_17692_n11557), .Y(_abc_17692_n11558) );
  AND2X2 AND2X2_4747 ( .A(_abc_17692_n11330), .B(_abc_17692_n11163), .Y(_abc_17692_n11559) );
  AND2X2 AND2X2_4748 ( .A(_abc_17692_n11278), .B(_abc_17692_n11559), .Y(_abc_17692_n11560) );
  AND2X2 AND2X2_4749 ( .A(_abc_17692_n11561), .B(_abc_17692_n11482), .Y(_abc_17692_n11562) );
  AND2X2 AND2X2_475 ( .A(delta_29_), .B(sum_29_), .Y(_abc_17692_n1769) );
  AND2X2 AND2X2_4750 ( .A(_abc_17692_n11564), .B(_abc_17692_n1830_bF_buf3), .Y(_abc_17692_n11565) );
  AND2X2 AND2X2_4751 ( .A(_abc_17692_n11565), .B(_abc_17692_n11563), .Y(_abc_17692_n11566) );
  AND2X2 AND2X2_4752 ( .A(_abc_17692_n11569), .B(state_14_bF_buf3), .Y(_abc_17692_n11570) );
  AND2X2 AND2X2_4753 ( .A(_abc_17692_n8383_bF_buf2), .B(workunit1_22_), .Y(_abc_17692_n11571) );
  AND2X2 AND2X2_4754 ( .A(state_8_bF_buf5), .B(\data_in1[22] ), .Y(_abc_17692_n11572) );
  AND2X2 AND2X2_4755 ( .A(_abc_17692_n11577), .B(_abc_17692_n11576), .Y(_abc_17692_n11578) );
  AND2X2 AND2X2_4756 ( .A(_abc_17692_n11579), .B(_abc_17692_n11580), .Y(_abc_17692_n11581) );
  AND2X2 AND2X2_4757 ( .A(_abc_17692_n11582), .B(workunit2_23_), .Y(_abc_17692_n11583) );
  AND2X2 AND2X2_4758 ( .A(_abc_17692_n11581), .B(_abc_17692_n6505), .Y(_abc_17692_n11585) );
  AND2X2 AND2X2_4759 ( .A(_abc_17692_n11584), .B(_abc_17692_n11586), .Y(_abc_17692_n11587) );
  AND2X2 AND2X2_476 ( .A(_abc_17692_n1741), .B(_abc_17692_n1738), .Y(_abc_17692_n1771) );
  AND2X2 AND2X2_4760 ( .A(_abc_17692_n11578), .B(_abc_17692_n11588), .Y(_abc_17692_n11589) );
  AND2X2 AND2X2_4761 ( .A(_abc_17692_n11590), .B(_abc_17692_n11587), .Y(_abc_17692_n11591) );
  AND2X2 AND2X2_4762 ( .A(_abc_17692_n11595), .B(_abc_17692_n11594), .Y(_abc_17692_n11596) );
  AND2X2 AND2X2_4763 ( .A(_abc_17692_n11593), .B(_abc_17692_n11597), .Y(_abc_17692_n11598) );
  AND2X2 AND2X2_4764 ( .A(_abc_17692_n11600), .B(_abc_17692_n11601), .Y(_abc_17692_n11602) );
  AND2X2 AND2X2_4765 ( .A(_abc_17692_n11599), .B(_abc_17692_n11603), .Y(_abc_17692_n11604) );
  AND2X2 AND2X2_4766 ( .A(_abc_17692_n11451), .B(_abc_17692_n11441), .Y(_abc_17692_n11605) );
  AND2X2 AND2X2_4767 ( .A(_abc_17692_n11609), .B(_abc_17692_n1877_bF_buf2), .Y(_abc_17692_n11610) );
  AND2X2 AND2X2_4768 ( .A(_abc_17692_n11610), .B(_abc_17692_n11607), .Y(_abc_17692_n11611) );
  AND2X2 AND2X2_4769 ( .A(_abc_17692_n11612), .B(_abc_17692_n11613), .Y(_abc_17692_n11614) );
  AND2X2 AND2X2_477 ( .A(_abc_17692_n1772), .B(_abc_17692_n1770), .Y(_abc_17692_n1773) );
  AND2X2 AND2X2_4770 ( .A(_abc_17692_n11614), .B(_abc_17692_n5378), .Y(_abc_17692_n11615) );
  AND2X2 AND2X2_4771 ( .A(_abc_17692_n11616), .B(_abc_17692_n11617), .Y(_abc_17692_n11618) );
  AND2X2 AND2X2_4772 ( .A(_abc_17692_n11618), .B(workunit1_23_), .Y(_abc_17692_n11619) );
  AND2X2 AND2X2_4773 ( .A(_abc_17692_n11479), .B(workunit1_22_), .Y(_abc_17692_n11622) );
  AND2X2 AND2X2_4774 ( .A(_abc_17692_n11490), .B(_abc_17692_n11623), .Y(_abc_17692_n11624) );
  AND2X2 AND2X2_4775 ( .A(_abc_17692_n11627), .B(_abc_17692_n1830_bF_buf2), .Y(_abc_17692_n11628) );
  AND2X2 AND2X2_4776 ( .A(_abc_17692_n11628), .B(_abc_17692_n11626), .Y(_abc_17692_n11629) );
  AND2X2 AND2X2_4777 ( .A(_abc_17692_n11630), .B(_abc_17692_n11631), .Y(_abc_17692_n11632) );
  AND2X2 AND2X2_4778 ( .A(_abc_17692_n11634), .B(_abc_17692_n11635), .Y(_abc_17692_n11636) );
  AND2X2 AND2X2_4779 ( .A(_abc_17692_n11633), .B(_abc_17692_n11637), .Y(_abc_17692_n11638) );
  AND2X2 AND2X2_478 ( .A(_abc_17692_n1776), .B(state_3_bF_buf4), .Y(_abc_17692_n1777) );
  AND2X2 AND2X2_4780 ( .A(_abc_17692_n11472), .B(_abc_17692_n11639), .Y(_abc_17692_n11640) );
  AND2X2 AND2X2_4781 ( .A(_abc_17692_n11636), .B(_abc_17692_n5378), .Y(_abc_17692_n11643) );
  AND2X2 AND2X2_4782 ( .A(_abc_17692_n11632), .B(workunit1_23_), .Y(_abc_17692_n11644) );
  AND2X2 AND2X2_4783 ( .A(_abc_17692_n11646), .B(_abc_17692_n1846_bF_buf2), .Y(_abc_17692_n11647) );
  AND2X2 AND2X2_4784 ( .A(_abc_17692_n11647), .B(_abc_17692_n11642), .Y(_abc_17692_n11648) );
  AND2X2 AND2X2_4785 ( .A(_abc_17692_n11651), .B(_abc_17692_n11652), .Y(_abc_17692_n11653) );
  AND2X2 AND2X2_4786 ( .A(_abc_17692_n11653), .B(_abc_17692_n5378), .Y(_abc_17692_n11654) );
  AND2X2 AND2X2_4787 ( .A(_abc_17692_n11655), .B(_abc_17692_n11656), .Y(_abc_17692_n11657) );
  AND2X2 AND2X2_4788 ( .A(_abc_17692_n11657), .B(workunit1_23_), .Y(_abc_17692_n11658) );
  AND2X2 AND2X2_4789 ( .A(_abc_17692_n11510), .B(_abc_17692_n11660), .Y(_abc_17692_n11661) );
  AND2X2 AND2X2_479 ( .A(_abc_17692_n1777), .B(_abc_17692_n1775_1), .Y(_abc_17692_n1778) );
  AND2X2 AND2X2_4790 ( .A(_abc_17692_n11662), .B(_abc_17692_n11659), .Y(_abc_17692_n11663) );
  AND2X2 AND2X2_4791 ( .A(_abc_17692_n11664), .B(_abc_17692_n11665), .Y(_abc_17692_n11666) );
  AND2X2 AND2X2_4792 ( .A(_abc_17692_n11661), .B(_abc_17692_n11666), .Y(_abc_17692_n11667) );
  AND2X2 AND2X2_4793 ( .A(_abc_17692_n11668), .B(_abc_17692_n1863_bF_buf2), .Y(_abc_17692_n11669) );
  AND2X2 AND2X2_4794 ( .A(_abc_17692_n11670), .B(state_10_bF_buf2), .Y(_abc_17692_n11671) );
  AND2X2 AND2X2_4795 ( .A(_abc_17692_n11676), .B(_abc_17692_n1863_bF_buf1), .Y(_abc_17692_n11677) );
  AND2X2 AND2X2_4796 ( .A(_abc_17692_n11677), .B(_abc_17692_n11675), .Y(_abc_17692_n11678) );
  AND2X2 AND2X2_4797 ( .A(_abc_17692_n11679), .B(workunit1_22_), .Y(_abc_17692_n11680) );
  AND2X2 AND2X2_4798 ( .A(_abc_17692_n11538), .B(_abc_17692_n11681), .Y(_abc_17692_n11682) );
  AND2X2 AND2X2_4799 ( .A(_abc_17692_n11685), .B(_abc_17692_n1877_bF_buf1), .Y(_abc_17692_n11686) );
  AND2X2 AND2X2_48 ( .A(_abc_17692_n749), .B(_abc_17692_n748), .Y(data_out2_7__FF_INPUT) );
  AND2X2 AND2X2_480 ( .A(_abc_17692_n1755_1), .B(_abc_17692_n1740), .Y(_abc_17692_n1779) );
  AND2X2 AND2X2_4800 ( .A(_abc_17692_n11686), .B(_abc_17692_n11684), .Y(_abc_17692_n11687) );
  AND2X2 AND2X2_4801 ( .A(_abc_17692_n11691), .B(_abc_17692_n1846_bF_buf1), .Y(_abc_17692_n11692) );
  AND2X2 AND2X2_4802 ( .A(_abc_17692_n11692), .B(_abc_17692_n11690), .Y(_abc_17692_n11693) );
  AND2X2 AND2X2_4803 ( .A(_abc_17692_n11698), .B(_abc_17692_n1830_bF_buf1), .Y(_abc_17692_n11699) );
  AND2X2 AND2X2_4804 ( .A(_abc_17692_n11699), .B(_abc_17692_n11697), .Y(_abc_17692_n11700) );
  AND2X2 AND2X2_4805 ( .A(_abc_17692_n11703), .B(state_14_bF_buf2), .Y(_abc_17692_n11704) );
  AND2X2 AND2X2_4806 ( .A(_abc_17692_n8383_bF_buf1), .B(workunit1_23_), .Y(_abc_17692_n11705) );
  AND2X2 AND2X2_4807 ( .A(state_8_bF_buf4), .B(\data_in1[23] ), .Y(_abc_17692_n11706) );
  AND2X2 AND2X2_4808 ( .A(_abc_17692_n11710), .B(_abc_17692_n11711), .Y(_abc_17692_n11712) );
  AND2X2 AND2X2_4809 ( .A(_abc_17692_n11713), .B(workunit2_24_), .Y(_abc_17692_n11714) );
  AND2X2 AND2X2_481 ( .A(_abc_17692_n1780), .B(_abc_17692_n1767), .Y(_abc_17692_n1782) );
  AND2X2 AND2X2_4810 ( .A(_abc_17692_n11712), .B(_abc_17692_n6657_1), .Y(_abc_17692_n11715) );
  AND2X2 AND2X2_4811 ( .A(_abc_17692_n11576), .B(_abc_17692_n11584), .Y(_abc_17692_n11718) );
  AND2X2 AND2X2_4812 ( .A(_abc_17692_n11433), .B(_abc_17692_n11587), .Y(_abc_17692_n11720) );
  AND2X2 AND2X2_4813 ( .A(_abc_17692_n11722), .B(_abc_17692_n11719), .Y(_abc_17692_n11723) );
  AND2X2 AND2X2_4814 ( .A(_abc_17692_n11725), .B(_abc_17692_n11723), .Y(_abc_17692_n11726) );
  AND2X2 AND2X2_4815 ( .A(_abc_17692_n11728), .B(_abc_17692_n11726), .Y(_abc_17692_n11729) );
  AND2X2 AND2X2_4816 ( .A(_abc_17692_n11730), .B(_abc_17692_n11717), .Y(_abc_17692_n11731) );
  AND2X2 AND2X2_4817 ( .A(_abc_17692_n11729), .B(_abc_17692_n11716), .Y(_abc_17692_n11732) );
  AND2X2 AND2X2_4818 ( .A(_abc_17692_n11735), .B(_abc_17692_n11736), .Y(_abc_17692_n11737) );
  AND2X2 AND2X2_4819 ( .A(_abc_17692_n11737), .B(workunit1_24_), .Y(_abc_17692_n11738) );
  AND2X2 AND2X2_482 ( .A(_abc_17692_n1783), .B(state_15_bF_buf4), .Y(_abc_17692_n1784) );
  AND2X2 AND2X2_4820 ( .A(_abc_17692_n11739), .B(_abc_17692_n5598), .Y(_abc_17692_n11740) );
  AND2X2 AND2X2_4821 ( .A(_abc_17692_n11666), .B(_abc_17692_n11502), .Y(_abc_17692_n11742) );
  AND2X2 AND2X2_4822 ( .A(_abc_17692_n11505), .B(_abc_17692_n11742), .Y(_abc_17692_n11743) );
  AND2X2 AND2X2_4823 ( .A(_abc_17692_n11745), .B(_abc_17692_n11665), .Y(_abc_17692_n11746) );
  AND2X2 AND2X2_4824 ( .A(_abc_17692_n11744), .B(_abc_17692_n11746), .Y(_abc_17692_n11747) );
  AND2X2 AND2X2_4825 ( .A(_abc_17692_n11742), .B(_abc_17692_n11506), .Y(_abc_17692_n11748) );
  AND2X2 AND2X2_4826 ( .A(_abc_17692_n11750), .B(_abc_17692_n11747), .Y(_abc_17692_n11751) );
  AND2X2 AND2X2_4827 ( .A(_abc_17692_n11748), .B(_abc_17692_n11120), .Y(_abc_17692_n11752) );
  AND2X2 AND2X2_4828 ( .A(_abc_17692_n10584), .B(_abc_17692_n11752), .Y(_abc_17692_n11753) );
  AND2X2 AND2X2_4829 ( .A(_abc_17692_n11754), .B(_abc_17692_n11751), .Y(_abc_17692_n11755) );
  AND2X2 AND2X2_483 ( .A(_abc_17692_n1784), .B(_abc_17692_n1781), .Y(_abc_17692_n1785) );
  AND2X2 AND2X2_4830 ( .A(_abc_17692_n11756), .B(_abc_17692_n11741), .Y(_abc_17692_n11757) );
  AND2X2 AND2X2_4831 ( .A(_abc_17692_n11758), .B(_abc_17692_n11759), .Y(_abc_17692_n11760) );
  AND2X2 AND2X2_4832 ( .A(_abc_17692_n11762), .B(_abc_17692_n11763), .Y(_abc_17692_n11764) );
  AND2X2 AND2X2_4833 ( .A(_abc_17692_n11764), .B(workunit1_24_), .Y(_abc_17692_n11765) );
  AND2X2 AND2X2_4834 ( .A(_abc_17692_n11766), .B(_abc_17692_n11767), .Y(_abc_17692_n11768) );
  AND2X2 AND2X2_4835 ( .A(_abc_17692_n11604), .B(_abc_17692_n11443), .Y(_abc_17692_n11770) );
  AND2X2 AND2X2_4836 ( .A(_abc_17692_n11770), .B(_abc_17692_n11447), .Y(_abc_17692_n11771) );
  AND2X2 AND2X2_4837 ( .A(_abc_17692_n11150), .B(_abc_17692_n11771), .Y(_abc_17692_n11772) );
  AND2X2 AND2X2_4838 ( .A(_abc_17692_n11770), .B(_abc_17692_n11446), .Y(_abc_17692_n11773) );
  AND2X2 AND2X2_4839 ( .A(_abc_17692_n11599), .B(_abc_17692_n11440), .Y(_abc_17692_n11775) );
  AND2X2 AND2X2_484 ( .A(_abc_17692_n722_bF_buf3), .B(sum_30_), .Y(_abc_17692_n1786) );
  AND2X2 AND2X2_4840 ( .A(_abc_17692_n11148), .B(_abc_17692_n11771), .Y(_abc_17692_n11778) );
  AND2X2 AND2X2_4841 ( .A(_abc_17692_n11780), .B(_abc_17692_n11769), .Y(_abc_17692_n11782) );
  AND2X2 AND2X2_4842 ( .A(_abc_17692_n11783), .B(_abc_17692_n1877_bF_buf0), .Y(_abc_17692_n11784) );
  AND2X2 AND2X2_4843 ( .A(_abc_17692_n11784), .B(_abc_17692_n11781), .Y(_abc_17692_n11785) );
  AND2X2 AND2X2_4844 ( .A(_abc_17692_n11786), .B(_abc_17692_n11787), .Y(_abc_17692_n11788) );
  AND2X2 AND2X2_4845 ( .A(_abc_17692_n11788), .B(workunit1_24_), .Y(_abc_17692_n11789) );
  AND2X2 AND2X2_4846 ( .A(_abc_17692_n11790), .B(_abc_17692_n5598), .Y(_abc_17692_n11791) );
  AND2X2 AND2X2_4847 ( .A(_abc_17692_n11621), .B(_abc_17692_n11483), .Y(_abc_17692_n11793) );
  AND2X2 AND2X2_4848 ( .A(_abc_17692_n11793), .B(_abc_17692_n11485), .Y(_abc_17692_n11794) );
  AND2X2 AND2X2_4849 ( .A(_abc_17692_n11621), .B(_abc_17692_n11622), .Y(_abc_17692_n11795) );
  AND2X2 AND2X2_485 ( .A(_abc_17692_n1791), .B(_abc_17692_n1793), .Y(_abc_17692_n1794) );
  AND2X2 AND2X2_4850 ( .A(_abc_17692_n11329), .B(_abc_17692_n11164), .Y(_abc_17692_n11798) );
  AND2X2 AND2X2_4851 ( .A(_abc_17692_n11793), .B(_abc_17692_n11798), .Y(_abc_17692_n11799) );
  AND2X2 AND2X2_4852 ( .A(_abc_17692_n11169), .B(_abc_17692_n11799), .Y(_abc_17692_n11800) );
  AND2X2 AND2X2_4853 ( .A(_abc_17692_n11799), .B(_abc_17692_n11170), .Y(_abc_17692_n11802) );
  AND2X2 AND2X2_4854 ( .A(_abc_17692_n10561), .B(_abc_17692_n11802), .Y(_abc_17692_n11803) );
  AND2X2 AND2X2_4855 ( .A(_abc_17692_n11804), .B(_abc_17692_n11792), .Y(_abc_17692_n11805) );
  AND2X2 AND2X2_4856 ( .A(_abc_17692_n11807), .B(_abc_17692_n1830_bF_buf0), .Y(_abc_17692_n11808) );
  AND2X2 AND2X2_4857 ( .A(_abc_17692_n11808), .B(_abc_17692_n11806), .Y(_abc_17692_n11809) );
  AND2X2 AND2X2_4858 ( .A(_abc_17692_n11810), .B(_abc_17692_n11811), .Y(_abc_17692_n11812) );
  AND2X2 AND2X2_4859 ( .A(_abc_17692_n11812), .B(workunit1_24_), .Y(_abc_17692_n11813) );
  AND2X2 AND2X2_486 ( .A(_abc_17692_n1776), .B(_abc_17692_n1796), .Y(_abc_17692_n1797) );
  AND2X2 AND2X2_4860 ( .A(_abc_17692_n11814), .B(_abc_17692_n5598), .Y(_abc_17692_n11815) );
  AND2X2 AND2X2_4861 ( .A(_abc_17692_n11822), .B(_abc_17692_n11637), .Y(_abc_17692_n11823) );
  AND2X2 AND2X2_4862 ( .A(_abc_17692_n11821), .B(_abc_17692_n11823), .Y(_abc_17692_n11824) );
  AND2X2 AND2X2_4863 ( .A(_abc_17692_n11820), .B(_abc_17692_n11824), .Y(_abc_17692_n11825) );
  AND2X2 AND2X2_4864 ( .A(_abc_17692_n11819), .B(_abc_17692_n11825), .Y(_abc_17692_n11826) );
  AND2X2 AND2X2_4865 ( .A(_abc_17692_n11827), .B(_abc_17692_n11816), .Y(_abc_17692_n11828) );
  AND2X2 AND2X2_4866 ( .A(_abc_17692_n11830), .B(_abc_17692_n1846_bF_buf0), .Y(_abc_17692_n11831) );
  AND2X2 AND2X2_4867 ( .A(_abc_17692_n11831), .B(_abc_17692_n11829), .Y(_abc_17692_n11832) );
  AND2X2 AND2X2_4868 ( .A(_abc_17692_n11835), .B(state_10_bF_buf1), .Y(_abc_17692_n11836) );
  AND2X2 AND2X2_4869 ( .A(_abc_17692_n11836), .B(_abc_17692_n11761), .Y(_abc_17692_n11837) );
  AND2X2 AND2X2_487 ( .A(_abc_17692_n1800), .B(state_3_bF_buf3), .Y(_abc_17692_n1801) );
  AND2X2 AND2X2_4870 ( .A(_abc_17692_n11659), .B(_abc_17692_n11501), .Y(_abc_17692_n11839) );
  AND2X2 AND2X2_4871 ( .A(_abc_17692_n11839), .B(_abc_17692_n11520), .Y(_abc_17692_n11840) );
  AND2X2 AND2X2_4872 ( .A(_abc_17692_n11840), .B(_abc_17692_n11213), .Y(_abc_17692_n11841) );
  AND2X2 AND2X2_4873 ( .A(_abc_17692_n11839), .B(_abc_17692_n11518), .Y(_abc_17692_n11842) );
  AND2X2 AND2X2_4874 ( .A(_abc_17692_n11653), .B(workunit1_23_), .Y(_abc_17692_n11843) );
  AND2X2 AND2X2_4875 ( .A(_abc_17692_n11659), .B(_abc_17692_n11672), .Y(_abc_17692_n11844) );
  AND2X2 AND2X2_4876 ( .A(_abc_17692_n11215), .B(_abc_17692_n11840), .Y(_abc_17692_n11848) );
  AND2X2 AND2X2_4877 ( .A(_abc_17692_n11849), .B(_abc_17692_n11838), .Y(_abc_17692_n11851) );
  AND2X2 AND2X2_4878 ( .A(_abc_17692_n11852), .B(_abc_17692_n1863_bF_buf10), .Y(_abc_17692_n11853) );
  AND2X2 AND2X2_4879 ( .A(_abc_17692_n11853), .B(_abc_17692_n11850), .Y(_abc_17692_n11854) );
  AND2X2 AND2X2_488 ( .A(_abc_17692_n1801), .B(_abc_17692_n1799), .Y(_abc_17692_n1802) );
  AND2X2 AND2X2_4880 ( .A(_abc_17692_n11602), .B(workunit1_23_), .Y(_abc_17692_n11859) );
  AND2X2 AND2X2_4881 ( .A(_abc_17692_n11861), .B(_abc_17692_n11860), .Y(_abc_17692_n11862) );
  AND2X2 AND2X2_4882 ( .A(_abc_17692_n11858), .B(_abc_17692_n11862), .Y(_abc_17692_n11863) );
  AND2X2 AND2X2_4883 ( .A(_abc_17692_n11857), .B(_abc_17692_n11863), .Y(_abc_17692_n11864) );
  AND2X2 AND2X2_4884 ( .A(_abc_17692_n11865), .B(_abc_17692_n10616), .Y(_abc_17692_n11866) );
  AND2X2 AND2X2_4885 ( .A(_abc_17692_n11869), .B(_abc_17692_n11864), .Y(_abc_17692_n11870) );
  AND2X2 AND2X2_4886 ( .A(_abc_17692_n11871), .B(_abc_17692_n11768), .Y(_abc_17692_n11872) );
  AND2X2 AND2X2_4887 ( .A(_abc_17692_n11874), .B(_abc_17692_n1877_bF_buf10), .Y(_abc_17692_n11875) );
  AND2X2 AND2X2_4888 ( .A(_abc_17692_n11875), .B(_abc_17692_n11873), .Y(_abc_17692_n11876) );
  AND2X2 AND2X2_4889 ( .A(_abc_17692_n11636), .B(workunit1_23_), .Y(_abc_17692_n11882) );
  AND2X2 AND2X2_489 ( .A(_abc_17692_n1764), .B(sum_30_), .Y(_abc_17692_n1803) );
  AND2X2 AND2X2_4890 ( .A(_abc_17692_n11885), .B(_abc_17692_n11883), .Y(_abc_17692_n11886) );
  AND2X2 AND2X2_4891 ( .A(_abc_17692_n11881), .B(_abc_17692_n11886), .Y(_abc_17692_n11887) );
  AND2X2 AND2X2_4892 ( .A(_abc_17692_n11880), .B(_abc_17692_n11887), .Y(_abc_17692_n11888) );
  AND2X2 AND2X2_4893 ( .A(_abc_17692_n11890), .B(_abc_17692_n11888), .Y(_abc_17692_n11891) );
  AND2X2 AND2X2_4894 ( .A(_abc_17692_n11894), .B(_abc_17692_n1846_bF_buf10), .Y(_abc_17692_n11895) );
  AND2X2 AND2X2_4895 ( .A(_abc_17692_n11895), .B(_abc_17692_n11893), .Y(_abc_17692_n11896) );
  AND2X2 AND2X2_4896 ( .A(_abc_17692_n11620), .B(_abc_17692_n11482), .Y(_abc_17692_n11897) );
  AND2X2 AND2X2_4897 ( .A(_abc_17692_n11897), .B(_abc_17692_n11559), .Y(_abc_17692_n11898) );
  AND2X2 AND2X2_4898 ( .A(_abc_17692_n11898), .B(_abc_17692_n11274), .Y(_abc_17692_n11899) );
  AND2X2 AND2X2_4899 ( .A(_abc_17692_n10637), .B(_abc_17692_n11899), .Y(_abc_17692_n11900) );
  AND2X2 AND2X2_49 ( .A(_abc_17692_n752), .B(_abc_17692_n751_1), .Y(data_out2_8__FF_INPUT) );
  AND2X2 AND2X2_490 ( .A(_abc_17692_n1807), .B(state_15_bF_buf3), .Y(_abc_17692_n1808) );
  AND2X2 AND2X2_4900 ( .A(_abc_17692_n11264), .B(_abc_17692_n11898), .Y(_abc_17692_n11901) );
  AND2X2 AND2X2_4901 ( .A(_abc_17692_n11897), .B(_abc_17692_n11558), .Y(_abc_17692_n11902) );
  AND2X2 AND2X2_4902 ( .A(_abc_17692_n11614), .B(workunit1_23_), .Y(_abc_17692_n11903) );
  AND2X2 AND2X2_4903 ( .A(_abc_17692_n11620), .B(_abc_17692_n11694), .Y(_abc_17692_n11904) );
  AND2X2 AND2X2_4904 ( .A(_abc_17692_n11912), .B(_abc_17692_n1830_bF_buf10), .Y(_abc_17692_n11913) );
  AND2X2 AND2X2_4905 ( .A(_abc_17692_n11913), .B(_abc_17692_n11910), .Y(_abc_17692_n11914) );
  AND2X2 AND2X2_4906 ( .A(_abc_17692_n11917), .B(state_14_bF_buf1), .Y(_abc_17692_n11918) );
  AND2X2 AND2X2_4907 ( .A(_abc_17692_n8383_bF_buf0), .B(workunit1_24_), .Y(_abc_17692_n11919) );
  AND2X2 AND2X2_4908 ( .A(state_8_bF_buf3), .B(\data_in1[24] ), .Y(_abc_17692_n11920) );
  AND2X2 AND2X2_4909 ( .A(_abc_17692_n11926), .B(_abc_17692_n11927), .Y(_abc_17692_n11928) );
  AND2X2 AND2X2_491 ( .A(_abc_17692_n1808), .B(_abc_17692_n1806), .Y(_abc_17692_n1809) );
  AND2X2 AND2X2_4910 ( .A(_abc_17692_n11929), .B(workunit2_25_), .Y(_abc_17692_n11930) );
  AND2X2 AND2X2_4911 ( .A(_abc_17692_n11928), .B(_abc_17692_n6952), .Y(_abc_17692_n11932) );
  AND2X2 AND2X2_4912 ( .A(_abc_17692_n11931), .B(_abc_17692_n11933), .Y(_abc_17692_n11934) );
  AND2X2 AND2X2_4913 ( .A(_abc_17692_n11925), .B(_abc_17692_n11935), .Y(_abc_17692_n11936) );
  AND2X2 AND2X2_4914 ( .A(_abc_17692_n11924), .B(_abc_17692_n11934), .Y(_abc_17692_n11937) );
  AND2X2 AND2X2_4915 ( .A(_abc_17692_n11939), .B(_abc_17692_n11941), .Y(_abc_17692_n11942) );
  AND2X2 AND2X2_4916 ( .A(_abc_17692_n11944), .B(_abc_17692_n11945), .Y(_abc_17692_n11946) );
  AND2X2 AND2X2_4917 ( .A(_abc_17692_n11943), .B(_abc_17692_n11947), .Y(_abc_17692_n11948) );
  AND2X2 AND2X2_4918 ( .A(_abc_17692_n11950), .B(workunit1_24_), .Y(_abc_17692_n11951) );
  AND2X2 AND2X2_4919 ( .A(_abc_17692_n11783), .B(_abc_17692_n11952), .Y(_abc_17692_n11953) );
  AND2X2 AND2X2_492 ( .A(_abc_17692_n722_bF_buf2), .B(sum_31_), .Y(_abc_17692_n1810) );
  AND2X2 AND2X2_4920 ( .A(_abc_17692_n11956), .B(_abc_17692_n1877_bF_buf9), .Y(_abc_17692_n11957) );
  AND2X2 AND2X2_4921 ( .A(_abc_17692_n11957), .B(_abc_17692_n11954), .Y(_abc_17692_n11958) );
  AND2X2 AND2X2_4922 ( .A(_abc_17692_n11959), .B(_abc_17692_n11960), .Y(_abc_17692_n11961) );
  AND2X2 AND2X2_4923 ( .A(_abc_17692_n11963), .B(_abc_17692_n11964), .Y(_abc_17692_n11965) );
  AND2X2 AND2X2_4924 ( .A(_abc_17692_n11962), .B(_abc_17692_n11966), .Y(_abc_17692_n11967) );
  AND2X2 AND2X2_4925 ( .A(_abc_17692_n11814), .B(workunit1_24_), .Y(_abc_17692_n11968) );
  AND2X2 AND2X2_4926 ( .A(_abc_17692_n11829), .B(_abc_17692_n11969), .Y(_abc_17692_n11970) );
  AND2X2 AND2X2_4927 ( .A(_abc_17692_n11974), .B(_abc_17692_n1846_bF_buf9), .Y(_abc_17692_n11975) );
  AND2X2 AND2X2_4928 ( .A(_abc_17692_n11975), .B(_abc_17692_n11972), .Y(_abc_17692_n11976) );
  AND2X2 AND2X2_4929 ( .A(_abc_17692_n11977), .B(_abc_17692_n11978), .Y(_abc_17692_n11979) );
  AND2X2 AND2X2_493 ( .A(workunit1_0_), .B(workunit1_5_), .Y(_abc_17692_n1815_1) );
  AND2X2 AND2X2_4930 ( .A(_abc_17692_n11979), .B(_abc_17692_n5782), .Y(_abc_17692_n11980) );
  AND2X2 AND2X2_4931 ( .A(_abc_17692_n11981), .B(_abc_17692_n11982), .Y(_abc_17692_n11983) );
  AND2X2 AND2X2_4932 ( .A(_abc_17692_n11983), .B(workunit1_25_), .Y(_abc_17692_n11984) );
  AND2X2 AND2X2_4933 ( .A(_abc_17692_n11790), .B(workunit1_24_), .Y(_abc_17692_n11986) );
  AND2X2 AND2X2_4934 ( .A(_abc_17692_n11806), .B(_abc_17692_n11987), .Y(_abc_17692_n11988) );
  AND2X2 AND2X2_4935 ( .A(_abc_17692_n11992), .B(_abc_17692_n1830_bF_buf9), .Y(_abc_17692_n11993) );
  AND2X2 AND2X2_4936 ( .A(_abc_17692_n11993), .B(_abc_17692_n11989), .Y(_abc_17692_n11994) );
  AND2X2 AND2X2_4937 ( .A(_abc_17692_n11997), .B(_abc_17692_n11998), .Y(_abc_17692_n11999) );
  AND2X2 AND2X2_4938 ( .A(_abc_17692_n11999), .B(_abc_17692_n5782), .Y(_abc_17692_n12000) );
  AND2X2 AND2X2_4939 ( .A(_abc_17692_n12002), .B(_abc_17692_n12003), .Y(_abc_17692_n12004) );
  AND2X2 AND2X2_494 ( .A(_abc_17692_n1816), .B(_abc_17692_n1817), .Y(_abc_17692_n1818) );
  AND2X2 AND2X2_4940 ( .A(_abc_17692_n12004), .B(workunit1_25_), .Y(_abc_17692_n12005) );
  AND2X2 AND2X2_4941 ( .A(_abc_17692_n12001), .B(_abc_17692_n12006), .Y(_abc_17692_n12007) );
  AND2X2 AND2X2_4942 ( .A(_abc_17692_n11739), .B(workunit1_24_), .Y(_abc_17692_n12008) );
  AND2X2 AND2X2_4943 ( .A(_abc_17692_n11758), .B(_abc_17692_n12009), .Y(_abc_17692_n12010) );
  AND2X2 AND2X2_4944 ( .A(_abc_17692_n12010), .B(_abc_17692_n12007), .Y(_abc_17692_n12011) );
  AND2X2 AND2X2_4945 ( .A(_abc_17692_n12013), .B(_abc_17692_n12012), .Y(_abc_17692_n12014) );
  AND2X2 AND2X2_4946 ( .A(_abc_17692_n12015), .B(_abc_17692_n1863_bF_buf9), .Y(_abc_17692_n12016) );
  AND2X2 AND2X2_4947 ( .A(_abc_17692_n12017), .B(state_10_bF_buf0), .Y(_abc_17692_n12018) );
  AND2X2 AND2X2_4948 ( .A(_abc_17692_n11852), .B(_abc_17692_n12019), .Y(_abc_17692_n12020) );
  AND2X2 AND2X2_4949 ( .A(_abc_17692_n12022), .B(_abc_17692_n12023), .Y(_abc_17692_n12024) );
  AND2X2 AND2X2_495 ( .A(sum_0_), .B(\key_in[0] ), .Y(_abc_17692_n1820) );
  AND2X2 AND2X2_4950 ( .A(_abc_17692_n12024), .B(_abc_17692_n1863_bF_buf8), .Y(_abc_17692_n12025) );
  AND2X2 AND2X2_4951 ( .A(_abc_17692_n11873), .B(_abc_17692_n11766), .Y(_abc_17692_n12026) );
  AND2X2 AND2X2_4952 ( .A(_abc_17692_n12029), .B(_abc_17692_n1877_bF_buf8), .Y(_abc_17692_n12030) );
  AND2X2 AND2X2_4953 ( .A(_abc_17692_n12030), .B(_abc_17692_n12028), .Y(_abc_17692_n12031) );
  AND2X2 AND2X2_4954 ( .A(_abc_17692_n11894), .B(_abc_17692_n12032), .Y(_abc_17692_n12033) );
  AND2X2 AND2X2_4955 ( .A(_abc_17692_n12036), .B(_abc_17692_n1846_bF_buf8), .Y(_abc_17692_n12037) );
  AND2X2 AND2X2_4956 ( .A(_abc_17692_n12037), .B(_abc_17692_n12035), .Y(_abc_17692_n12038) );
  AND2X2 AND2X2_4957 ( .A(_abc_17692_n11910), .B(_abc_17692_n12039), .Y(_abc_17692_n12040) );
  AND2X2 AND2X2_4958 ( .A(_abc_17692_n12040), .B(_abc_17692_n11985), .Y(_abc_17692_n12041) );
  AND2X2 AND2X2_4959 ( .A(_abc_17692_n12042), .B(_abc_17692_n11990), .Y(_abc_17692_n12043) );
  AND2X2 AND2X2_496 ( .A(_abc_17692_n1821), .B(_abc_17692_n1822), .Y(_abc_17692_n1823) );
  AND2X2 AND2X2_4960 ( .A(_abc_17692_n12044), .B(_abc_17692_n1830_bF_buf8), .Y(_abc_17692_n12045) );
  AND2X2 AND2X2_4961 ( .A(_abc_17692_n12048), .B(state_14_bF_buf0), .Y(_abc_17692_n12049) );
  AND2X2 AND2X2_4962 ( .A(_abc_17692_n8383_bF_buf4), .B(workunit1_25_), .Y(_abc_17692_n12050) );
  AND2X2 AND2X2_4963 ( .A(state_8_bF_buf2), .B(\data_in1[25] ), .Y(_abc_17692_n12051) );
  AND2X2 AND2X2_4964 ( .A(_abc_17692_n11948), .B(_abc_17692_n11769), .Y(_abc_17692_n12055) );
  AND2X2 AND2X2_4965 ( .A(_abc_17692_n11780), .B(_abc_17692_n12055), .Y(_abc_17692_n12056) );
  AND2X2 AND2X2_4966 ( .A(_abc_17692_n12057), .B(_abc_17692_n11947), .Y(_abc_17692_n12058) );
  AND2X2 AND2X2_4967 ( .A(_abc_17692_n11717), .B(_abc_17692_n11934), .Y(_abc_17692_n12061) );
  AND2X2 AND2X2_4968 ( .A(_abc_17692_n11730), .B(_abc_17692_n12061), .Y(_abc_17692_n12062) );
  AND2X2 AND2X2_4969 ( .A(_abc_17692_n12063), .B(_abc_17692_n11933), .Y(_abc_17692_n12064) );
  AND2X2 AND2X2_497 ( .A(_abc_17692_n1824), .B(_abc_17692_n1819), .Y(_abc_17692_n1825) );
  AND2X2 AND2X2_4970 ( .A(_abc_17692_n12067), .B(_abc_17692_n12068), .Y(_abc_17692_n12069) );
  AND2X2 AND2X2_4971 ( .A(_abc_17692_n12070), .B(workunit2_26_), .Y(_abc_17692_n12071) );
  AND2X2 AND2X2_4972 ( .A(_abc_17692_n12069), .B(_abc_17692_n7128), .Y(_abc_17692_n12072) );
  AND2X2 AND2X2_4973 ( .A(_abc_17692_n12066), .B(_abc_17692_n12073), .Y(_abc_17692_n12074) );
  AND2X2 AND2X2_4974 ( .A(_abc_17692_n12065), .B(_abc_17692_n12075), .Y(_abc_17692_n12076) );
  AND2X2 AND2X2_4975 ( .A(_abc_17692_n12080), .B(_abc_17692_n12079), .Y(_abc_17692_n12081) );
  AND2X2 AND2X2_4976 ( .A(_abc_17692_n12081), .B(workunit1_26_), .Y(_abc_17692_n12082) );
  AND2X2 AND2X2_4977 ( .A(_abc_17692_n12083), .B(_abc_17692_n12084), .Y(_abc_17692_n12085) );
  AND2X2 AND2X2_4978 ( .A(_abc_17692_n12060), .B(_abc_17692_n12085), .Y(_abc_17692_n12087) );
  AND2X2 AND2X2_4979 ( .A(_abc_17692_n12088), .B(_abc_17692_n1877_bF_buf7), .Y(_abc_17692_n12089) );
  AND2X2 AND2X2_498 ( .A(_abc_17692_n1826), .B(_abc_17692_n1823), .Y(_abc_17692_n1827) );
  AND2X2 AND2X2_4980 ( .A(_abc_17692_n12089), .B(_abc_17692_n12086), .Y(_abc_17692_n12090) );
  AND2X2 AND2X2_4981 ( .A(_abc_17692_n7168), .B(_abc_17692_n12077), .Y(_abc_17692_n12091) );
  AND2X2 AND2X2_4982 ( .A(_abc_17692_n7166), .B(_abc_17692_n12078), .Y(_abc_17692_n12092) );
  AND2X2 AND2X2_4983 ( .A(_abc_17692_n12095), .B(_abc_17692_n12096), .Y(_abc_17692_n12097) );
  AND2X2 AND2X2_4984 ( .A(_abc_17692_n11806), .B(_abc_17692_n12100), .Y(_abc_17692_n12101) );
  AND2X2 AND2X2_4985 ( .A(_abc_17692_n12105), .B(_abc_17692_n1830_bF_buf7), .Y(_abc_17692_n12106) );
  AND2X2 AND2X2_4986 ( .A(_abc_17692_n12106), .B(_abc_17692_n12104), .Y(_abc_17692_n12107) );
  AND2X2 AND2X2_4987 ( .A(_abc_17692_n12108), .B(_abc_17692_n12109), .Y(_abc_17692_n12110) );
  AND2X2 AND2X2_4988 ( .A(_abc_17692_n12111), .B(_abc_17692_n6065), .Y(_abc_17692_n12112) );
  AND2X2 AND2X2_4989 ( .A(_abc_17692_n12110), .B(workunit1_26_), .Y(_abc_17692_n12113) );
  AND2X2 AND2X2_499 ( .A(selectslice_0_), .B(selectslice_1_), .Y(_abc_17692_n1830) );
  AND2X2 AND2X2_4990 ( .A(_abc_17692_n11966), .B(_abc_17692_n11969), .Y(_abc_17692_n12117) );
  AND2X2 AND2X2_4991 ( .A(_abc_17692_n11967), .B(_abc_17692_n11816), .Y(_abc_17692_n12120) );
  AND2X2 AND2X2_4992 ( .A(_abc_17692_n11827), .B(_abc_17692_n12120), .Y(_abc_17692_n12121) );
  AND2X2 AND2X2_4993 ( .A(_abc_17692_n12122), .B(_abc_17692_n12115), .Y(_abc_17692_n12123) );
  AND2X2 AND2X2_4994 ( .A(_abc_17692_n12125), .B(_abc_17692_n1846_bF_buf7), .Y(_abc_17692_n12126) );
  AND2X2 AND2X2_4995 ( .A(_abc_17692_n12126), .B(_abc_17692_n12124), .Y(_abc_17692_n12127) );
  AND2X2 AND2X2_4996 ( .A(_abc_17692_n12131), .B(_abc_17692_n12001), .Y(_abc_17692_n12132) );
  AND2X2 AND2X2_4997 ( .A(_abc_17692_n12007), .B(_abc_17692_n11741), .Y(_abc_17692_n12133) );
  AND2X2 AND2X2_4998 ( .A(_abc_17692_n11756), .B(_abc_17692_n12133), .Y(_abc_17692_n12134) );
  AND2X2 AND2X2_4999 ( .A(_abc_17692_n12136), .B(_abc_17692_n12137), .Y(_abc_17692_n12138) );
  AND2X2 AND2X2_5 ( .A(_abc_17692_n632), .B(delta_2_), .Y(delta_2__FF_INPUT) );
  AND2X2 AND2X2_50 ( .A(_abc_17692_n755), .B(_abc_17692_n754), .Y(data_out2_9__FF_INPUT) );
  AND2X2 AND2X2_500 ( .A(_abc_17692_n1832), .B(_abc_17692_n1830_bF_buf10), .Y(_abc_17692_n1833) );
  AND2X2 AND2X2_5000 ( .A(_abc_17692_n12141), .B(_abc_17692_n12139), .Y(_abc_17692_n12142) );
  AND2X2 AND2X2_5001 ( .A(_abc_17692_n12135), .B(_abc_17692_n12143), .Y(_abc_17692_n12144) );
  AND2X2 AND2X2_5002 ( .A(_abc_17692_n12145), .B(_abc_17692_n12146), .Y(_abc_17692_n12147) );
  AND2X2 AND2X2_5003 ( .A(_abc_17692_n12148), .B(state_10_bF_buf4), .Y(_abc_17692_n12149) );
  AND2X2 AND2X2_5004 ( .A(_abc_17692_n12149), .B(_abc_17692_n12130), .Y(_abc_17692_n12150) );
  AND2X2 AND2X2_5005 ( .A(_abc_17692_n11999), .B(workunit1_25_), .Y(_abc_17692_n12151) );
  AND2X2 AND2X2_5006 ( .A(_abc_17692_n12012), .B(_abc_17692_n11738), .Y(_abc_17692_n12152) );
  AND2X2 AND2X2_5007 ( .A(_abc_17692_n12012), .B(_abc_17692_n11838), .Y(_abc_17692_n12154) );
  AND2X2 AND2X2_5008 ( .A(_abc_17692_n11849), .B(_abc_17692_n12154), .Y(_abc_17692_n12155) );
  AND2X2 AND2X2_5009 ( .A(_abc_17692_n12156), .B(_abc_17692_n12142), .Y(_abc_17692_n12157) );
  AND2X2 AND2X2_501 ( .A(_abc_17692_n1833), .B(_abc_17692_n1829), .Y(_abc_17692_n1834) );
  AND2X2 AND2X2_5010 ( .A(_abc_17692_n12159), .B(_abc_17692_n1863_bF_buf6), .Y(_abc_17692_n12160) );
  AND2X2 AND2X2_5011 ( .A(_abc_17692_n12160), .B(_abc_17692_n12158), .Y(_abc_17692_n12161) );
  AND2X2 AND2X2_5012 ( .A(_abc_17692_n11946), .B(workunit1_25_), .Y(_abc_17692_n12163) );
  AND2X2 AND2X2_5013 ( .A(_abc_17692_n12165), .B(_abc_17692_n12164), .Y(_abc_17692_n12166) );
  AND2X2 AND2X2_5014 ( .A(_abc_17692_n11949), .B(_abc_17692_n11768), .Y(_abc_17692_n12168) );
  AND2X2 AND2X2_5015 ( .A(_abc_17692_n11871), .B(_abc_17692_n12168), .Y(_abc_17692_n12169) );
  AND2X2 AND2X2_5016 ( .A(_abc_17692_n12170), .B(_abc_17692_n12162), .Y(_abc_17692_n12171) );
  AND2X2 AND2X2_5017 ( .A(_abc_17692_n12173), .B(_abc_17692_n1877_bF_buf6), .Y(_abc_17692_n12174) );
  AND2X2 AND2X2_5018 ( .A(_abc_17692_n12174), .B(_abc_17692_n12172), .Y(_abc_17692_n12175) );
  AND2X2 AND2X2_5019 ( .A(_abc_17692_n11965), .B(workunit1_25_), .Y(_abc_17692_n12176) );
  AND2X2 AND2X2_502 ( .A(sum_0_), .B(\key_in[32] ), .Y(_abc_17692_n1835) );
  AND2X2 AND2X2_5020 ( .A(_abc_17692_n12178), .B(_abc_17692_n12177), .Y(_abc_17692_n12179) );
  AND2X2 AND2X2_5021 ( .A(_abc_17692_n11892), .B(_abc_17692_n12182), .Y(_abc_17692_n12183) );
  AND2X2 AND2X2_5022 ( .A(_abc_17692_n12184), .B(_abc_17692_n12114), .Y(_abc_17692_n12186) );
  AND2X2 AND2X2_5023 ( .A(_abc_17692_n12187), .B(_abc_17692_n1846_bF_buf6), .Y(_abc_17692_n12188) );
  AND2X2 AND2X2_5024 ( .A(_abc_17692_n12188), .B(_abc_17692_n12185), .Y(_abc_17692_n12189) );
  AND2X2 AND2X2_5025 ( .A(_abc_17692_n11985), .B(_abc_17692_n11911), .Y(_abc_17692_n12190) );
  AND2X2 AND2X2_5026 ( .A(_abc_17692_n11985), .B(_abc_17692_n11789), .Y(_abc_17692_n12193) );
  AND2X2 AND2X2_5027 ( .A(_abc_17692_n11979), .B(workunit1_25_), .Y(_abc_17692_n12194) );
  AND2X2 AND2X2_5028 ( .A(_abc_17692_n12192), .B(_abc_17692_n12196), .Y(_abc_17692_n12197) );
  AND2X2 AND2X2_5029 ( .A(_abc_17692_n12200), .B(_abc_17692_n1830_bF_buf6), .Y(_abc_17692_n12201) );
  AND2X2 AND2X2_503 ( .A(_abc_17692_n1836), .B(_abc_17692_n1837), .Y(_abc_17692_n1838) );
  AND2X2 AND2X2_5030 ( .A(_abc_17692_n12201), .B(_abc_17692_n12198), .Y(_abc_17692_n12202) );
  AND2X2 AND2X2_5031 ( .A(_abc_17692_n12205), .B(state_14_bF_buf4), .Y(_abc_17692_n12206) );
  AND2X2 AND2X2_5032 ( .A(_abc_17692_n8383_bF_buf3), .B(workunit1_26_), .Y(_abc_17692_n12207) );
  AND2X2 AND2X2_5033 ( .A(state_8_bF_buf1), .B(\data_in1[26] ), .Y(_abc_17692_n12208) );
  AND2X2 AND2X2_5034 ( .A(workunit2_23_), .B(workunit2_27_), .Y(_abc_17692_n12213) );
  AND2X2 AND2X2_5035 ( .A(_abc_17692_n6505), .B(_abc_17692_n7385), .Y(_abc_17692_n12215) );
  AND2X2 AND2X2_5036 ( .A(_abc_17692_n12216), .B(_abc_17692_n12214), .Y(_abc_17692_n12217) );
  AND2X2 AND2X2_5037 ( .A(_abc_17692_n12212), .B(_abc_17692_n12218), .Y(_abc_17692_n12219) );
  AND2X2 AND2X2_5038 ( .A(_abc_17692_n12220), .B(_abc_17692_n12221), .Y(_abc_17692_n12222) );
  AND2X2 AND2X2_5039 ( .A(_abc_17692_n12223), .B(_abc_17692_n12225), .Y(_abc_17692_n12226) );
  AND2X2 AND2X2_504 ( .A(_abc_17692_n1839), .B(_abc_17692_n1819), .Y(_abc_17692_n1840) );
  AND2X2 AND2X2_5040 ( .A(_abc_17692_n12229), .B(_abc_17692_n12228), .Y(_abc_17692_n12230) );
  AND2X2 AND2X2_5041 ( .A(_abc_17692_n12227), .B(_abc_17692_n12231), .Y(_abc_17692_n12232) );
  AND2X2 AND2X2_5042 ( .A(_abc_17692_n12236), .B(_abc_17692_n12232), .Y(_abc_17692_n12237) );
  AND2X2 AND2X2_5043 ( .A(_abc_17692_n12230), .B(_abc_17692_n6242), .Y(_abc_17692_n12238) );
  AND2X2 AND2X2_5044 ( .A(_abc_17692_n12226), .B(workunit1_27_), .Y(_abc_17692_n12239) );
  AND2X2 AND2X2_5045 ( .A(_abc_17692_n12235), .B(_abc_17692_n12240), .Y(_abc_17692_n12241) );
  AND2X2 AND2X2_5046 ( .A(_abc_17692_n12244), .B(_abc_17692_n12245), .Y(_abc_17692_n12246) );
  AND2X2 AND2X2_5047 ( .A(_abc_17692_n12246), .B(_abc_17692_n6242), .Y(_abc_17692_n12247) );
  AND2X2 AND2X2_5048 ( .A(_abc_17692_n12248), .B(_abc_17692_n12249), .Y(_abc_17692_n12250) );
  AND2X2 AND2X2_5049 ( .A(_abc_17692_n12250), .B(workunit1_27_), .Y(_abc_17692_n12251) );
  AND2X2 AND2X2_505 ( .A(_abc_17692_n1826), .B(_abc_17692_n1838), .Y(_abc_17692_n1841) );
  AND2X2 AND2X2_5050 ( .A(_abc_17692_n12094), .B(workunit1_26_), .Y(_abc_17692_n12254) );
  AND2X2 AND2X2_5051 ( .A(_abc_17692_n12105), .B(_abc_17692_n12255), .Y(_abc_17692_n12256) );
  AND2X2 AND2X2_5052 ( .A(_abc_17692_n12259), .B(_abc_17692_n1830_bF_buf5), .Y(_abc_17692_n12260) );
  AND2X2 AND2X2_5053 ( .A(_abc_17692_n12260), .B(_abc_17692_n12258), .Y(_abc_17692_n12261) );
  AND2X2 AND2X2_5054 ( .A(_abc_17692_n12262), .B(_abc_17692_n12263), .Y(_abc_17692_n12264) );
  AND2X2 AND2X2_5055 ( .A(_abc_17692_n12267), .B(_abc_17692_n12266), .Y(_abc_17692_n12268) );
  AND2X2 AND2X2_5056 ( .A(_abc_17692_n12265), .B(_abc_17692_n12269), .Y(_abc_17692_n12270) );
  AND2X2 AND2X2_5057 ( .A(_abc_17692_n12088), .B(_abc_17692_n12083), .Y(_abc_17692_n12271) );
  AND2X2 AND2X2_5058 ( .A(_abc_17692_n12275), .B(_abc_17692_n1877_bF_buf5), .Y(_abc_17692_n12276) );
  AND2X2 AND2X2_5059 ( .A(_abc_17692_n12276), .B(_abc_17692_n12273), .Y(_abc_17692_n12277) );
  AND2X2 AND2X2_506 ( .A(_abc_17692_n1845), .B(selectslice_1_), .Y(_abc_17692_n1846) );
  AND2X2 AND2X2_5060 ( .A(_abc_17692_n12278), .B(_abc_17692_n12279), .Y(_abc_17692_n12280) );
  AND2X2 AND2X2_5061 ( .A(_abc_17692_n12280), .B(_abc_17692_n6242), .Y(_abc_17692_n12281) );
  AND2X2 AND2X2_5062 ( .A(_abc_17692_n12282), .B(_abc_17692_n12283), .Y(_abc_17692_n12284) );
  AND2X2 AND2X2_5063 ( .A(_abc_17692_n12284), .B(workunit1_27_), .Y(_abc_17692_n12285) );
  AND2X2 AND2X2_5064 ( .A(_abc_17692_n12290), .B(_abc_17692_n12291), .Y(_abc_17692_n12292) );
  AND2X2 AND2X2_5065 ( .A(_abc_17692_n12293), .B(_abc_17692_n1846_bF_buf5), .Y(_abc_17692_n12294) );
  AND2X2 AND2X2_5066 ( .A(_abc_17692_n12294), .B(_abc_17692_n12289), .Y(_abc_17692_n12295) );
  AND2X2 AND2X2_5067 ( .A(_abc_17692_n12298), .B(state_10_bF_buf3), .Y(_abc_17692_n12299) );
  AND2X2 AND2X2_5068 ( .A(_abc_17692_n12299), .B(_abc_17692_n12243), .Y(_abc_17692_n12300) );
  AND2X2 AND2X2_5069 ( .A(_abc_17692_n12158), .B(_abc_17692_n12139), .Y(_abc_17692_n12301) );
  AND2X2 AND2X2_507 ( .A(_abc_17692_n1847), .B(_abc_17692_n1846_bF_buf10), .Y(_abc_17692_n1848) );
  AND2X2 AND2X2_5070 ( .A(_abc_17692_n12304), .B(_abc_17692_n1863_bF_buf4), .Y(_abc_17692_n12305) );
  AND2X2 AND2X2_5071 ( .A(_abc_17692_n12305), .B(_abc_17692_n12303), .Y(_abc_17692_n12306) );
  AND2X2 AND2X2_5072 ( .A(_abc_17692_n12307), .B(workunit1_26_), .Y(_abc_17692_n12308) );
  AND2X2 AND2X2_5073 ( .A(_abc_17692_n12172), .B(_abc_17692_n12309), .Y(_abc_17692_n12310) );
  AND2X2 AND2X2_5074 ( .A(_abc_17692_n12313), .B(_abc_17692_n1877_bF_buf4), .Y(_abc_17692_n12314) );
  AND2X2 AND2X2_5075 ( .A(_abc_17692_n12314), .B(_abc_17692_n12312), .Y(_abc_17692_n12315) );
  AND2X2 AND2X2_5076 ( .A(_abc_17692_n12111), .B(workunit1_26_), .Y(_abc_17692_n12316) );
  AND2X2 AND2X2_5077 ( .A(_abc_17692_n12187), .B(_abc_17692_n12317), .Y(_abc_17692_n12318) );
  AND2X2 AND2X2_5078 ( .A(_abc_17692_n12321), .B(_abc_17692_n1846_bF_buf4), .Y(_abc_17692_n12322) );
  AND2X2 AND2X2_5079 ( .A(_abc_17692_n12322), .B(_abc_17692_n12320), .Y(_abc_17692_n12323) );
  AND2X2 AND2X2_508 ( .A(_abc_17692_n1848), .B(_abc_17692_n1844), .Y(_abc_17692_n1849) );
  AND2X2 AND2X2_5080 ( .A(_abc_17692_n12198), .B(_abc_17692_n12095), .Y(_abc_17692_n12324) );
  AND2X2 AND2X2_5081 ( .A(_abc_17692_n12327), .B(_abc_17692_n1830_bF_buf4), .Y(_abc_17692_n12328) );
  AND2X2 AND2X2_5082 ( .A(_abc_17692_n12328), .B(_abc_17692_n12326), .Y(_abc_17692_n12329) );
  AND2X2 AND2X2_5083 ( .A(_abc_17692_n12332), .B(state_14_bF_buf3), .Y(_abc_17692_n12333) );
  AND2X2 AND2X2_5084 ( .A(_abc_17692_n8383_bF_buf2), .B(workunit1_27_), .Y(_abc_17692_n12334) );
  AND2X2 AND2X2_5085 ( .A(state_8_bF_buf0), .B(\data_in1[27] ), .Y(_abc_17692_n12335) );
  AND2X2 AND2X2_5086 ( .A(workunit2_24_), .B(workunit2_28_), .Y(_abc_17692_n12339) );
  AND2X2 AND2X2_5087 ( .A(_abc_17692_n6657_1), .B(_abc_17692_n7535), .Y(_abc_17692_n12340) );
  AND2X2 AND2X2_5088 ( .A(_abc_17692_n12343), .B(_abc_17692_n12216), .Y(_abc_17692_n12344) );
  AND2X2 AND2X2_5089 ( .A(_abc_17692_n12345), .B(_abc_17692_n12341), .Y(_abc_17692_n12346) );
  AND2X2 AND2X2_509 ( .A(sum_0_), .B(\key_in[96] ), .Y(_abc_17692_n1851) );
  AND2X2 AND2X2_5090 ( .A(_abc_17692_n12344), .B(_abc_17692_n12347), .Y(_abc_17692_n12348) );
  AND2X2 AND2X2_5091 ( .A(_abc_17692_n12351), .B(_abc_17692_n12352), .Y(_abc_17692_n12353) );
  AND2X2 AND2X2_5092 ( .A(_abc_17692_n12355), .B(_abc_17692_n12356), .Y(_abc_17692_n12357) );
  AND2X2 AND2X2_5093 ( .A(_abc_17692_n12232), .B(_abc_17692_n12143), .Y(_abc_17692_n12359) );
  AND2X2 AND2X2_5094 ( .A(_abc_17692_n12359), .B(_abc_17692_n12133), .Y(_abc_17692_n12360) );
  AND2X2 AND2X2_5095 ( .A(_abc_17692_n12359), .B(_abc_17692_n12132), .Y(_abc_17692_n12363) );
  AND2X2 AND2X2_5096 ( .A(_abc_17692_n12364), .B(_abc_17692_n12227), .Y(_abc_17692_n12365) );
  AND2X2 AND2X2_5097 ( .A(_abc_17692_n12362), .B(_abc_17692_n12367), .Y(_abc_17692_n12368) );
  AND2X2 AND2X2_5098 ( .A(_abc_17692_n12369), .B(_abc_17692_n12358), .Y(_abc_17692_n12371) );
  AND2X2 AND2X2_5099 ( .A(_abc_17692_n12372), .B(_abc_17692_n12370), .Y(_abc_17692_n12373) );
  AND2X2 AND2X2_51 ( .A(_abc_17692_n758), .B(_abc_17692_n757), .Y(data_out2_10__FF_INPUT) );
  AND2X2 AND2X2_510 ( .A(_abc_17692_n1852_1), .B(_abc_17692_n1853), .Y(_abc_17692_n1854) );
  AND2X2 AND2X2_5100 ( .A(_abc_17692_n12375), .B(_abc_17692_n12376), .Y(_abc_17692_n12377) );
  AND2X2 AND2X2_5101 ( .A(_abc_17692_n12377), .B(workunit1_28_), .Y(_abc_17692_n12378) );
  AND2X2 AND2X2_5102 ( .A(_abc_17692_n12379), .B(_abc_17692_n12380), .Y(_abc_17692_n12381) );
  AND2X2 AND2X2_5103 ( .A(_abc_17692_n12270), .B(_abc_17692_n12085), .Y(_abc_17692_n12383) );
  AND2X2 AND2X2_5104 ( .A(_abc_17692_n12383), .B(_abc_17692_n12055), .Y(_abc_17692_n12384) );
  AND2X2 AND2X2_5105 ( .A(_abc_17692_n11780), .B(_abc_17692_n12384), .Y(_abc_17692_n12385) );
  AND2X2 AND2X2_5106 ( .A(_abc_17692_n12059), .B(_abc_17692_n12383), .Y(_abc_17692_n12386) );
  AND2X2 AND2X2_5107 ( .A(_abc_17692_n12265), .B(_abc_17692_n12082), .Y(_abc_17692_n12388) );
  AND2X2 AND2X2_5108 ( .A(_abc_17692_n12391), .B(_abc_17692_n12382), .Y(_abc_17692_n12392) );
  AND2X2 AND2X2_5109 ( .A(_abc_17692_n12394), .B(_abc_17692_n1877_bF_buf3), .Y(_abc_17692_n12395) );
  AND2X2 AND2X2_511 ( .A(_abc_17692_n1855_1), .B(_abc_17692_n1819), .Y(_abc_17692_n1856) );
  AND2X2 AND2X2_5110 ( .A(_abc_17692_n12395), .B(_abc_17692_n12393), .Y(_abc_17692_n12396) );
  AND2X2 AND2X2_5111 ( .A(_abc_17692_n12397), .B(_abc_17692_n12398), .Y(_abc_17692_n12399) );
  AND2X2 AND2X2_5112 ( .A(_abc_17692_n12401), .B(_abc_17692_n12402), .Y(_abc_17692_n12403) );
  AND2X2 AND2X2_5113 ( .A(_abc_17692_n11990), .B(_abc_17692_n11792), .Y(_abc_17692_n12405) );
  AND2X2 AND2X2_5114 ( .A(_abc_17692_n12253), .B(_abc_17692_n12098), .Y(_abc_17692_n12406) );
  AND2X2 AND2X2_5115 ( .A(_abc_17692_n12406), .B(_abc_17692_n12405), .Y(_abc_17692_n12407) );
  AND2X2 AND2X2_5116 ( .A(_abc_17692_n11804), .B(_abc_17692_n12407), .Y(_abc_17692_n12408) );
  AND2X2 AND2X2_5117 ( .A(_abc_17692_n12406), .B(_abc_17692_n12410), .Y(_abc_17692_n12411) );
  AND2X2 AND2X2_5118 ( .A(_abc_17692_n12253), .B(_abc_17692_n12254), .Y(_abc_17692_n12412) );
  AND2X2 AND2X2_5119 ( .A(_abc_17692_n12415), .B(_abc_17692_n12404), .Y(_abc_17692_n12417) );
  AND2X2 AND2X2_512 ( .A(_abc_17692_n1826), .B(_abc_17692_n1854), .Y(_abc_17692_n1857) );
  AND2X2 AND2X2_5120 ( .A(_abc_17692_n12418), .B(_abc_17692_n1830_bF_buf3), .Y(_abc_17692_n12419) );
  AND2X2 AND2X2_5121 ( .A(_abc_17692_n12419), .B(_abc_17692_n12416), .Y(_abc_17692_n12420) );
  AND2X2 AND2X2_5122 ( .A(_abc_17692_n12421), .B(_abc_17692_n12422), .Y(_abc_17692_n12423) );
  AND2X2 AND2X2_5123 ( .A(_abc_17692_n12425), .B(_abc_17692_n12426), .Y(_abc_17692_n12427) );
  AND2X2 AND2X2_5124 ( .A(_abc_17692_n12434), .B(_abc_17692_n12290), .Y(_abc_17692_n12435) );
  AND2X2 AND2X2_5125 ( .A(_abc_17692_n12433), .B(_abc_17692_n12436), .Y(_abc_17692_n12437) );
  AND2X2 AND2X2_5126 ( .A(_abc_17692_n12432), .B(_abc_17692_n12437), .Y(_abc_17692_n12438) );
  AND2X2 AND2X2_5127 ( .A(_abc_17692_n12439), .B(_abc_17692_n12428), .Y(_abc_17692_n12440) );
  AND2X2 AND2X2_5128 ( .A(_abc_17692_n12442), .B(_abc_17692_n1846_bF_buf3), .Y(_abc_17692_n12443) );
  AND2X2 AND2X2_5129 ( .A(_abc_17692_n12443), .B(_abc_17692_n12441), .Y(_abc_17692_n12444) );
  AND2X2 AND2X2_513 ( .A(_abc_17692_n1859), .B(workunit2_0_), .Y(_abc_17692_n1860) );
  AND2X2 AND2X2_5130 ( .A(_abc_17692_n12447), .B(state_10_bF_buf2), .Y(_abc_17692_n12448) );
  AND2X2 AND2X2_5131 ( .A(_abc_17692_n12374), .B(_abc_17692_n12448), .Y(_abc_17692_n12449) );
  AND2X2 AND2X2_5132 ( .A(_abc_17692_n12240), .B(_abc_17692_n12142), .Y(_abc_17692_n12450) );
  AND2X2 AND2X2_5133 ( .A(_abc_17692_n12450), .B(_abc_17692_n12154), .Y(_abc_17692_n12451) );
  AND2X2 AND2X2_5134 ( .A(_abc_17692_n11849), .B(_abc_17692_n12451), .Y(_abc_17692_n12452) );
  AND2X2 AND2X2_5135 ( .A(_abc_17692_n12450), .B(_abc_17692_n12153), .Y(_abc_17692_n12453) );
  AND2X2 AND2X2_5136 ( .A(_abc_17692_n12230), .B(workunit1_27_), .Y(_abc_17692_n12454) );
  AND2X2 AND2X2_5137 ( .A(_abc_17692_n12240), .B(_abc_17692_n12455), .Y(_abc_17692_n12456) );
  AND2X2 AND2X2_5138 ( .A(_abc_17692_n12459), .B(_abc_17692_n12357), .Y(_abc_17692_n12460) );
  AND2X2 AND2X2_5139 ( .A(_abc_17692_n12462), .B(_abc_17692_n1863_bF_buf2), .Y(_abc_17692_n12463) );
  AND2X2 AND2X2_514 ( .A(_abc_17692_n1845), .B(_abc_17692_n1862), .Y(_abc_17692_n1863) );
  AND2X2 AND2X2_5140 ( .A(_abc_17692_n12463), .B(_abc_17692_n12461), .Y(_abc_17692_n12464) );
  AND2X2 AND2X2_5141 ( .A(_abc_17692_n12268), .B(workunit1_27_), .Y(_abc_17692_n12470) );
  AND2X2 AND2X2_5142 ( .A(_abc_17692_n12472), .B(_abc_17692_n12471), .Y(_abc_17692_n12473) );
  AND2X2 AND2X2_5143 ( .A(_abc_17692_n12469), .B(_abc_17692_n12473), .Y(_abc_17692_n12474) );
  AND2X2 AND2X2_5144 ( .A(_abc_17692_n12468), .B(_abc_17692_n12474), .Y(_abc_17692_n12475) );
  AND2X2 AND2X2_5145 ( .A(_abc_17692_n12476), .B(_abc_17692_n12381), .Y(_abc_17692_n12477) );
  AND2X2 AND2X2_5146 ( .A(_abc_17692_n12479), .B(_abc_17692_n1877_bF_buf2), .Y(_abc_17692_n12480) );
  AND2X2 AND2X2_5147 ( .A(_abc_17692_n12480), .B(_abc_17692_n12478), .Y(_abc_17692_n12481) );
  AND2X2 AND2X2_5148 ( .A(_abc_17692_n12280), .B(workunit1_27_), .Y(_abc_17692_n12486) );
  AND2X2 AND2X2_5149 ( .A(_abc_17692_n12488), .B(_abc_17692_n12487), .Y(_abc_17692_n12489) );
  AND2X2 AND2X2_515 ( .A(_abc_17692_n1864), .B(_abc_17692_n1863_bF_buf10), .Y(_abc_17692_n1865) );
  AND2X2 AND2X2_5150 ( .A(_abc_17692_n12485), .B(_abc_17692_n12489), .Y(_abc_17692_n12490) );
  AND2X2 AND2X2_5151 ( .A(_abc_17692_n12484), .B(_abc_17692_n12490), .Y(_abc_17692_n12491) );
  AND2X2 AND2X2_5152 ( .A(_abc_17692_n12492), .B(_abc_17692_n12427), .Y(_abc_17692_n12494) );
  AND2X2 AND2X2_5153 ( .A(_abc_17692_n12495), .B(_abc_17692_n1846_bF_buf2), .Y(_abc_17692_n12496) );
  AND2X2 AND2X2_5154 ( .A(_abc_17692_n12496), .B(_abc_17692_n12493), .Y(_abc_17692_n12497) );
  AND2X2 AND2X2_5155 ( .A(_abc_17692_n12252), .B(_abc_17692_n12097), .Y(_abc_17692_n12498) );
  AND2X2 AND2X2_5156 ( .A(_abc_17692_n12498), .B(_abc_17692_n12190), .Y(_abc_17692_n12499) );
  AND2X2 AND2X2_5157 ( .A(_abc_17692_n11908), .B(_abc_17692_n12499), .Y(_abc_17692_n12500) );
  AND2X2 AND2X2_5158 ( .A(_abc_17692_n12498), .B(_abc_17692_n12195), .Y(_abc_17692_n12501) );
  AND2X2 AND2X2_5159 ( .A(_abc_17692_n12246), .B(workunit1_27_), .Y(_abc_17692_n12502) );
  AND2X2 AND2X2_516 ( .A(_abc_17692_n1865), .B(_abc_17692_n1861), .Y(_abc_17692_n1866) );
  AND2X2 AND2X2_5160 ( .A(_abc_17692_n12252), .B(_abc_17692_n12503), .Y(_abc_17692_n12504) );
  AND2X2 AND2X2_5161 ( .A(_abc_17692_n12507), .B(_abc_17692_n12403), .Y(_abc_17692_n12508) );
  AND2X2 AND2X2_5162 ( .A(_abc_17692_n12510), .B(_abc_17692_n1830_bF_buf2), .Y(_abc_17692_n12511) );
  AND2X2 AND2X2_5163 ( .A(_abc_17692_n12511), .B(_abc_17692_n12509), .Y(_abc_17692_n12512) );
  AND2X2 AND2X2_5164 ( .A(_abc_17692_n12515), .B(state_14_bF_buf2), .Y(_abc_17692_n12516) );
  AND2X2 AND2X2_5165 ( .A(_abc_17692_n8383_bF_buf1), .B(workunit1_28_), .Y(_abc_17692_n12517) );
  AND2X2 AND2X2_5166 ( .A(state_8_bF_buf9), .B(\data_in1[28] ), .Y(_abc_17692_n12518) );
  AND2X2 AND2X2_5167 ( .A(workunit2_25_), .B(workunit2_29_), .Y(_abc_17692_n12523) );
  AND2X2 AND2X2_5168 ( .A(_abc_17692_n6952), .B(_abc_17692_n7812), .Y(_abc_17692_n12525) );
  AND2X2 AND2X2_5169 ( .A(_abc_17692_n12526), .B(_abc_17692_n12524), .Y(_abc_17692_n12527) );
  AND2X2 AND2X2_517 ( .A(sum_0_), .B(\key_in[64] ), .Y(_abc_17692_n1867_1) );
  AND2X2 AND2X2_5170 ( .A(_abc_17692_n12522), .B(_abc_17692_n12528), .Y(_abc_17692_n12529) );
  AND2X2 AND2X2_5171 ( .A(_abc_17692_n12530), .B(_abc_17692_n12531), .Y(_abc_17692_n12532) );
  AND2X2 AND2X2_5172 ( .A(_abc_17692_n12533), .B(_abc_17692_n12535), .Y(_abc_17692_n12536) );
  AND2X2 AND2X2_5173 ( .A(_abc_17692_n12536), .B(_abc_17692_n6659_1), .Y(_abc_17692_n12537) );
  AND2X2 AND2X2_5174 ( .A(_abc_17692_n12539), .B(_abc_17692_n12538), .Y(_abc_17692_n12540) );
  AND2X2 AND2X2_5175 ( .A(_abc_17692_n12540), .B(workunit1_29_), .Y(_abc_17692_n12541) );
  AND2X2 AND2X2_5176 ( .A(_abc_17692_n12372), .B(_abc_17692_n12543), .Y(_abc_17692_n12544) );
  AND2X2 AND2X2_5177 ( .A(_abc_17692_n12545), .B(_abc_17692_n12542), .Y(_abc_17692_n12546) );
  AND2X2 AND2X2_5178 ( .A(_abc_17692_n12547), .B(_abc_17692_n12548), .Y(_abc_17692_n12549) );
  AND2X2 AND2X2_5179 ( .A(_abc_17692_n12544), .B(_abc_17692_n12549), .Y(_abc_17692_n12550) );
  AND2X2 AND2X2_518 ( .A(_abc_17692_n1868), .B(_abc_17692_n1869), .Y(_abc_17692_n1870) );
  AND2X2 AND2X2_5180 ( .A(_abc_17692_n12554), .B(_abc_17692_n12553), .Y(_abc_17692_n12555) );
  AND2X2 AND2X2_5181 ( .A(_abc_17692_n12557), .B(_abc_17692_n12558), .Y(_abc_17692_n12559) );
  AND2X2 AND2X2_5182 ( .A(_abc_17692_n12556), .B(_abc_17692_n12560), .Y(_abc_17692_n12561) );
  AND2X2 AND2X2_5183 ( .A(_abc_17692_n12563), .B(workunit1_28_), .Y(_abc_17692_n12564) );
  AND2X2 AND2X2_5184 ( .A(_abc_17692_n12568), .B(_abc_17692_n1877_bF_buf1), .Y(_abc_17692_n12569) );
  AND2X2 AND2X2_5185 ( .A(_abc_17692_n12569), .B(_abc_17692_n12567), .Y(_abc_17692_n12570) );
  AND2X2 AND2X2_5186 ( .A(_abc_17692_n12571), .B(_abc_17692_n12572), .Y(_abc_17692_n12573) );
  AND2X2 AND2X2_5187 ( .A(_abc_17692_n12573), .B(_abc_17692_n6659_1), .Y(_abc_17692_n12574) );
  AND2X2 AND2X2_5188 ( .A(_abc_17692_n12576), .B(_abc_17692_n12575), .Y(_abc_17692_n12577) );
  AND2X2 AND2X2_5189 ( .A(_abc_17692_n12577), .B(workunit1_29_), .Y(_abc_17692_n12578) );
  AND2X2 AND2X2_519 ( .A(_abc_17692_n1871), .B(_abc_17692_n1819), .Y(_abc_17692_n1872) );
  AND2X2 AND2X2_5190 ( .A(_abc_17692_n12400), .B(workunit1_28_), .Y(_abc_17692_n12580) );
  AND2X2 AND2X2_5191 ( .A(_abc_17692_n12418), .B(_abc_17692_n12581), .Y(_abc_17692_n12582) );
  AND2X2 AND2X2_5192 ( .A(_abc_17692_n12586), .B(_abc_17692_n1830_bF_buf1), .Y(_abc_17692_n12587) );
  AND2X2 AND2X2_5193 ( .A(_abc_17692_n12587), .B(_abc_17692_n12583), .Y(_abc_17692_n12588) );
  AND2X2 AND2X2_5194 ( .A(_abc_17692_n12589), .B(_abc_17692_n12590), .Y(_abc_17692_n12591) );
  AND2X2 AND2X2_5195 ( .A(_abc_17692_n12591), .B(_abc_17692_n6659_1), .Y(_abc_17692_n12592) );
  AND2X2 AND2X2_5196 ( .A(_abc_17692_n12594), .B(_abc_17692_n12593), .Y(_abc_17692_n12595) );
  AND2X2 AND2X2_5197 ( .A(_abc_17692_n12595), .B(workunit1_29_), .Y(_abc_17692_n12596) );
  AND2X2 AND2X2_5198 ( .A(_abc_17692_n12603), .B(_abc_17692_n12604), .Y(_abc_17692_n12605) );
  AND2X2 AND2X2_5199 ( .A(_abc_17692_n12606), .B(_abc_17692_n1846_bF_buf1), .Y(_abc_17692_n12607) );
  AND2X2 AND2X2_52 ( .A(_abc_17692_n761), .B(_abc_17692_n760), .Y(data_out2_11__FF_INPUT) );
  AND2X2 AND2X2_520 ( .A(_abc_17692_n1826), .B(_abc_17692_n1870), .Y(_abc_17692_n1873) );
  AND2X2 AND2X2_5200 ( .A(_abc_17692_n12607), .B(_abc_17692_n12602), .Y(_abc_17692_n12608) );
  AND2X2 AND2X2_5201 ( .A(_abc_17692_n12611), .B(state_10_bF_buf1), .Y(_abc_17692_n12612) );
  AND2X2 AND2X2_5202 ( .A(_abc_17692_n12552), .B(_abc_17692_n12612), .Y(_abc_17692_n12613) );
  AND2X2 AND2X2_5203 ( .A(_abc_17692_n12461), .B(_abc_17692_n12355), .Y(_abc_17692_n12614) );
  AND2X2 AND2X2_5204 ( .A(_abc_17692_n12616), .B(_abc_17692_n12617), .Y(_abc_17692_n12618) );
  AND2X2 AND2X2_5205 ( .A(_abc_17692_n12618), .B(_abc_17692_n1863_bF_buf0), .Y(_abc_17692_n12619) );
  AND2X2 AND2X2_5206 ( .A(_abc_17692_n12478), .B(_abc_17692_n12379), .Y(_abc_17692_n12620) );
  AND2X2 AND2X2_5207 ( .A(_abc_17692_n12623), .B(_abc_17692_n1877_bF_buf0), .Y(_abc_17692_n12624) );
  AND2X2 AND2X2_5208 ( .A(_abc_17692_n12624), .B(_abc_17692_n12622), .Y(_abc_17692_n12625) );
  AND2X2 AND2X2_5209 ( .A(_abc_17692_n12509), .B(_abc_17692_n12401), .Y(_abc_17692_n12626) );
  AND2X2 AND2X2_521 ( .A(_abc_17692_n1862), .B(selectslice_0_), .Y(_abc_17692_n1877) );
  AND2X2 AND2X2_5210 ( .A(_abc_17692_n12629), .B(_abc_17692_n1830_bF_buf0), .Y(_abc_17692_n12630) );
  AND2X2 AND2X2_5211 ( .A(_abc_17692_n12630), .B(_abc_17692_n12627), .Y(_abc_17692_n12631) );
  AND2X2 AND2X2_5212 ( .A(_abc_17692_n12495), .B(_abc_17692_n12425), .Y(_abc_17692_n12632) );
  AND2X2 AND2X2_5213 ( .A(_abc_17692_n12635), .B(_abc_17692_n1846_bF_buf0), .Y(_abc_17692_n12636) );
  AND2X2 AND2X2_5214 ( .A(_abc_17692_n12636), .B(_abc_17692_n12634), .Y(_abc_17692_n12637) );
  AND2X2 AND2X2_5215 ( .A(_abc_17692_n12640), .B(state_14_bF_buf1), .Y(_abc_17692_n12641) );
  AND2X2 AND2X2_5216 ( .A(_abc_17692_n8383_bF_buf0), .B(workunit1_29_), .Y(_abc_17692_n12642) );
  AND2X2 AND2X2_5217 ( .A(state_8_bF_buf8), .B(\data_in1[29] ), .Y(_abc_17692_n12643) );
  AND2X2 AND2X2_5218 ( .A(workunit2_26_), .B(workunit2_30_), .Y(_abc_17692_n12648) );
  AND2X2 AND2X2_5219 ( .A(_abc_17692_n7128), .B(_abc_17692_n7968), .Y(_abc_17692_n12649) );
  AND2X2 AND2X2_522 ( .A(_abc_17692_n1875), .B(workunit2_0_), .Y(_abc_17692_n1878) );
  AND2X2 AND2X2_5220 ( .A(_abc_17692_n12652), .B(_abc_17692_n12526), .Y(_abc_17692_n12653) );
  AND2X2 AND2X2_5221 ( .A(_abc_17692_n12653), .B(_abc_17692_n12651), .Y(_abc_17692_n12654) );
  AND2X2 AND2X2_5222 ( .A(_abc_17692_n12655), .B(_abc_17692_n12656), .Y(_abc_17692_n12657) );
  AND2X2 AND2X2_5223 ( .A(_abc_17692_n12658), .B(_abc_17692_n12660), .Y(_abc_17692_n12661) );
  AND2X2 AND2X2_5224 ( .A(_abc_17692_n12664), .B(_abc_17692_n12663), .Y(_abc_17692_n12665) );
  AND2X2 AND2X2_5225 ( .A(_abc_17692_n12662), .B(_abc_17692_n12666), .Y(_abc_17692_n12667) );
  AND2X2 AND2X2_5226 ( .A(_abc_17692_n12584), .B(_abc_17692_n12404), .Y(_abc_17692_n12669) );
  AND2X2 AND2X2_5227 ( .A(_abc_17692_n12415), .B(_abc_17692_n12669), .Y(_abc_17692_n12670) );
  AND2X2 AND2X2_5228 ( .A(_abc_17692_n12584), .B(_abc_17692_n12580), .Y(_abc_17692_n12671) );
  AND2X2 AND2X2_5229 ( .A(_abc_17692_n12673), .B(_abc_17692_n12668), .Y(_abc_17692_n12675) );
  AND2X2 AND2X2_523 ( .A(_abc_17692_n1879), .B(_abc_17692_n1877_bF_buf10), .Y(_abc_17692_n1880) );
  AND2X2 AND2X2_5230 ( .A(_abc_17692_n12676), .B(_abc_17692_n1830_bF_buf10), .Y(_abc_17692_n12677) );
  AND2X2 AND2X2_5231 ( .A(_abc_17692_n12677), .B(_abc_17692_n12674), .Y(_abc_17692_n12678) );
  AND2X2 AND2X2_5232 ( .A(_abc_17692_n8023), .B(_abc_17692_n12659), .Y(_abc_17692_n12679) );
  AND2X2 AND2X2_5233 ( .A(_abc_17692_n8024), .B(_abc_17692_n12657), .Y(_abc_17692_n12680) );
  AND2X2 AND2X2_5234 ( .A(_abc_17692_n12683), .B(_abc_17692_n12684), .Y(_abc_17692_n12685) );
  AND2X2 AND2X2_5235 ( .A(_abc_17692_n12561), .B(_abc_17692_n12382), .Y(_abc_17692_n12686) );
  AND2X2 AND2X2_5236 ( .A(_abc_17692_n12391), .B(_abc_17692_n12686), .Y(_abc_17692_n12687) );
  AND2X2 AND2X2_5237 ( .A(_abc_17692_n12561), .B(_abc_17692_n12564), .Y(_abc_17692_n12689) );
  AND2X2 AND2X2_5238 ( .A(_abc_17692_n12691), .B(_abc_17692_n12685), .Y(_abc_17692_n12692) );
  AND2X2 AND2X2_5239 ( .A(_abc_17692_n12694), .B(_abc_17692_n1877_bF_buf10), .Y(_abc_17692_n12695) );
  AND2X2 AND2X2_524 ( .A(_abc_17692_n1880), .B(_abc_17692_n1876), .Y(_abc_17692_n1881) );
  AND2X2 AND2X2_5240 ( .A(_abc_17692_n12695), .B(_abc_17692_n12693), .Y(_abc_17692_n12696) );
  AND2X2 AND2X2_5241 ( .A(_abc_17692_n12697), .B(_abc_17692_n12698), .Y(_abc_17692_n12699) );
  AND2X2 AND2X2_5242 ( .A(_abc_17692_n12702), .B(_abc_17692_n12701), .Y(_abc_17692_n12703) );
  AND2X2 AND2X2_5243 ( .A(_abc_17692_n12700), .B(_abc_17692_n12704), .Y(_abc_17692_n12705) );
  AND2X2 AND2X2_5244 ( .A(_abc_17692_n12708), .B(_abc_17692_n12604), .Y(_abc_17692_n12709) );
  AND2X2 AND2X2_5245 ( .A(_abc_17692_n12707), .B(_abc_17692_n12709), .Y(_abc_17692_n12710) );
  AND2X2 AND2X2_5246 ( .A(_abc_17692_n12713), .B(_abc_17692_n12714), .Y(_abc_17692_n12715) );
  AND2X2 AND2X2_5247 ( .A(_abc_17692_n12716), .B(_abc_17692_n1846_bF_buf10), .Y(_abc_17692_n12717) );
  AND2X2 AND2X2_5248 ( .A(_abc_17692_n12717), .B(_abc_17692_n12712), .Y(_abc_17692_n12718) );
  AND2X2 AND2X2_5249 ( .A(_abc_17692_n12723), .B(_abc_17692_n12722), .Y(_abc_17692_n12724) );
  AND2X2 AND2X2_525 ( .A(_abc_17692_n1883), .B(_abc_17692_n714_1), .Y(_abc_17692_n1884_1) );
  AND2X2 AND2X2_5250 ( .A(_abc_17692_n12726), .B(_abc_17692_n12727), .Y(_abc_17692_n12728) );
  AND2X2 AND2X2_5251 ( .A(_abc_17692_n12549), .B(_abc_17692_n12358), .Y(_abc_17692_n12729) );
  AND2X2 AND2X2_5252 ( .A(_abc_17692_n12548), .B(_abc_17692_n12543), .Y(_abc_17692_n12732) );
  AND2X2 AND2X2_5253 ( .A(_abc_17692_n12731), .B(_abc_17692_n12733), .Y(_abc_17692_n12734) );
  AND2X2 AND2X2_5254 ( .A(_abc_17692_n12738), .B(_abc_17692_n12737), .Y(_abc_17692_n12739) );
  AND2X2 AND2X2_5255 ( .A(_abc_17692_n12736), .B(_abc_17692_n12740), .Y(_abc_17692_n12741) );
  AND2X2 AND2X2_5256 ( .A(_abc_17692_n12742), .B(state_10_bF_buf0), .Y(_abc_17692_n12743) );
  AND2X2 AND2X2_5257 ( .A(_abc_17692_n12743), .B(_abc_17692_n12721), .Y(_abc_17692_n12744) );
  AND2X2 AND2X2_5258 ( .A(_abc_17692_n12747), .B(_abc_17692_n12748), .Y(_abc_17692_n12749) );
  AND2X2 AND2X2_5259 ( .A(_abc_17692_n12745), .B(_abc_17692_n12749), .Y(_abc_17692_n12750) );
  AND2X2 AND2X2_526 ( .A(_abc_17692_n715_1), .B(_abc_17692_n632), .Y(_abc_17692_n1885) );
  AND2X2 AND2X2_5260 ( .A(_abc_17692_n12757), .B(_abc_17692_n12756), .Y(_abc_17692_n12758) );
  AND2X2 AND2X2_5261 ( .A(_abc_17692_n12755), .B(_abc_17692_n12758), .Y(_abc_17692_n12759) );
  AND2X2 AND2X2_5262 ( .A(_abc_17692_n12753), .B(_abc_17692_n12759), .Y(_abc_17692_n12760) );
  AND2X2 AND2X2_5263 ( .A(_abc_17692_n12764), .B(_abc_17692_n12760), .Y(_abc_17692_n12765) );
  AND2X2 AND2X2_5264 ( .A(_abc_17692_n12771), .B(_abc_17692_n12770), .Y(_abc_17692_n12772) );
  AND2X2 AND2X2_5265 ( .A(_abc_17692_n12775), .B(_abc_17692_n12774), .Y(_abc_17692_n12776) );
  AND2X2 AND2X2_5266 ( .A(_abc_17692_n12773), .B(_abc_17692_n12776), .Y(_abc_17692_n12777) );
  AND2X2 AND2X2_5267 ( .A(_abc_17692_n12769), .B(_abc_17692_n12777), .Y(_abc_17692_n12778) );
  AND2X2 AND2X2_5268 ( .A(_abc_17692_n12536), .B(workunit1_29_), .Y(_abc_17692_n12781) );
  AND2X2 AND2X2_5269 ( .A(_abc_17692_n12783), .B(_abc_17692_n12782), .Y(_abc_17692_n12784) );
  AND2X2 AND2X2_527 ( .A(_abc_17692_n1885_bF_buf4), .B(workunit2_0_), .Y(_abc_17692_n1886) );
  AND2X2 AND2X2_5270 ( .A(_abc_17692_n12780), .B(_abc_17692_n12784), .Y(_abc_17692_n12785) );
  AND2X2 AND2X2_5271 ( .A(_abc_17692_n12542), .B(_abc_17692_n12357), .Y(_abc_17692_n12787) );
  AND2X2 AND2X2_5272 ( .A(_abc_17692_n12459), .B(_abc_17692_n12787), .Y(_abc_17692_n12788) );
  AND2X2 AND2X2_5273 ( .A(_abc_17692_n12542), .B(_abc_17692_n12789), .Y(_abc_17692_n12790) );
  AND2X2 AND2X2_5274 ( .A(_abc_17692_n12793), .B(_abc_17692_n1863_bF_buf9), .Y(_abc_17692_n12794) );
  AND2X2 AND2X2_5275 ( .A(_abc_17692_n12794), .B(_abc_17692_n12786), .Y(_abc_17692_n12795) );
  AND2X2 AND2X2_5276 ( .A(_abc_17692_n12559), .B(workunit1_29_), .Y(_abc_17692_n12799) );
  AND2X2 AND2X2_5277 ( .A(_abc_17692_n12801), .B(_abc_17692_n12800), .Y(_abc_17692_n12802) );
  AND2X2 AND2X2_5278 ( .A(_abc_17692_n12798), .B(_abc_17692_n12802), .Y(_abc_17692_n12803) );
  AND2X2 AND2X2_5279 ( .A(_abc_17692_n12806), .B(_abc_17692_n1877_bF_buf9), .Y(_abc_17692_n12807) );
  AND2X2 AND2X2_528 ( .A(state_8_bF_buf9), .B(\data_in2[0] ), .Y(_abc_17692_n1887) );
  AND2X2 AND2X2_5280 ( .A(_abc_17692_n12807), .B(_abc_17692_n12805), .Y(_abc_17692_n12808) );
  AND2X2 AND2X2_5281 ( .A(_abc_17692_n12591), .B(workunit1_29_), .Y(_abc_17692_n12811) );
  AND2X2 AND2X2_5282 ( .A(_abc_17692_n12813), .B(_abc_17692_n12812), .Y(_abc_17692_n12814) );
  AND2X2 AND2X2_5283 ( .A(_abc_17692_n12810), .B(_abc_17692_n12814), .Y(_abc_17692_n12815) );
  AND2X2 AND2X2_5284 ( .A(_abc_17692_n12818), .B(_abc_17692_n1846_bF_buf9), .Y(_abc_17692_n12819) );
  AND2X2 AND2X2_5285 ( .A(_abc_17692_n12819), .B(_abc_17692_n12816), .Y(_abc_17692_n12820) );
  AND2X2 AND2X2_5286 ( .A(_abc_17692_n12579), .B(_abc_17692_n12403), .Y(_abc_17692_n12821) );
  AND2X2 AND2X2_5287 ( .A(_abc_17692_n12507), .B(_abc_17692_n12821), .Y(_abc_17692_n12822) );
  AND2X2 AND2X2_5288 ( .A(_abc_17692_n12573), .B(workunit1_29_), .Y(_abc_17692_n12823) );
  AND2X2 AND2X2_5289 ( .A(_abc_17692_n12579), .B(_abc_17692_n12824), .Y(_abc_17692_n12825) );
  AND2X2 AND2X2_529 ( .A(workunit1_1_bF_buf2), .B(workunit1_6_), .Y(_abc_17692_n1891) );
  AND2X2 AND2X2_5290 ( .A(_abc_17692_n12827), .B(_abc_17692_n12667), .Y(_abc_17692_n12828) );
  AND2X2 AND2X2_5291 ( .A(_abc_17692_n12830), .B(_abc_17692_n1830_bF_buf9), .Y(_abc_17692_n12831) );
  AND2X2 AND2X2_5292 ( .A(_abc_17692_n12831), .B(_abc_17692_n12829), .Y(_abc_17692_n12832) );
  AND2X2 AND2X2_5293 ( .A(_abc_17692_n12835), .B(state_14_bF_buf0), .Y(_abc_17692_n12836) );
  AND2X2 AND2X2_5294 ( .A(_abc_17692_n8383_bF_buf4), .B(workunit1_30_), .Y(_abc_17692_n12837) );
  AND2X2 AND2X2_5295 ( .A(state_8_bF_buf7), .B(\data_in1[30] ), .Y(_abc_17692_n12838) );
  AND2X2 AND2X2_5296 ( .A(_abc_17692_n12740), .B(_abc_17692_n12726), .Y(_abc_17692_n12842) );
  AND2X2 AND2X2_5297 ( .A(_abc_17692_n8202), .B(workunit2_27_), .Y(_abc_17692_n12845) );
  AND2X2 AND2X2_5298 ( .A(_abc_17692_n7385), .B(workunit2_31_), .Y(_abc_17692_n12846) );
  AND2X2 AND2X2_5299 ( .A(_abc_17692_n12844), .B(_abc_17692_n12847), .Y(_abc_17692_n12848) );
  AND2X2 AND2X2_53 ( .A(_abc_17692_n764), .B(_abc_17692_n763), .Y(data_out2_12__FF_INPUT) );
  AND2X2 AND2X2_530 ( .A(_abc_17692_n1896), .B(_abc_17692_n1892), .Y(_abc_17692_n1897) );
  AND2X2 AND2X2_5300 ( .A(_abc_17692_n12849), .B(_abc_17692_n12850), .Y(_abc_17692_n12851) );
  AND2X2 AND2X2_5301 ( .A(_abc_17692_n12852), .B(_abc_17692_n7135), .Y(_abc_17692_n12853) );
  AND2X2 AND2X2_5302 ( .A(_abc_17692_n12854), .B(_abc_17692_n12855), .Y(_abc_17692_n12856) );
  AND2X2 AND2X2_5303 ( .A(_abc_17692_n8217), .B(_abc_17692_n12857), .Y(_abc_17692_n12858) );
  AND2X2 AND2X2_5304 ( .A(_abc_17692_n8201), .B(_abc_17692_n12856), .Y(_abc_17692_n12859) );
  AND2X2 AND2X2_5305 ( .A(_abc_17692_n12843), .B(_abc_17692_n12860), .Y(_abc_17692_n12861) );
  AND2X2 AND2X2_5306 ( .A(_abc_17692_n12842), .B(_abc_17692_n12862), .Y(_abc_17692_n12863) );
  AND2X2 AND2X2_5307 ( .A(_abc_17692_n12870), .B(_abc_17692_n12869), .Y(_abc_17692_n12871) );
  AND2X2 AND2X2_5308 ( .A(_abc_17692_n12874), .B(_abc_17692_n1877_bF_buf8), .Y(_abc_17692_n12875) );
  AND2X2 AND2X2_5309 ( .A(_abc_17692_n12875), .B(_abc_17692_n12873), .Y(_abc_17692_n12876) );
  AND2X2 AND2X2_531 ( .A(_abc_17692_n1895), .B(_abc_17692_n1898), .Y(_abc_17692_n1899) );
  AND2X2 AND2X2_5310 ( .A(_abc_17692_n12661), .B(workunit1_30_), .Y(_abc_17692_n12877) );
  AND2X2 AND2X2_5311 ( .A(_abc_17692_n12880), .B(_abc_17692_n12881), .Y(_abc_17692_n12882) );
  AND2X2 AND2X2_5312 ( .A(_abc_17692_n12885), .B(_abc_17692_n1830_bF_buf8), .Y(_abc_17692_n12886) );
  AND2X2 AND2X2_5313 ( .A(_abc_17692_n12886), .B(_abc_17692_n12883), .Y(_abc_17692_n12887) );
  AND2X2 AND2X2_5314 ( .A(_abc_17692_n12716), .B(_abc_17692_n12704), .Y(_abc_17692_n12888) );
  AND2X2 AND2X2_5315 ( .A(_abc_17692_n12891), .B(_abc_17692_n12890), .Y(_abc_17692_n12892) );
  AND2X2 AND2X2_5316 ( .A(_abc_17692_n12895), .B(_abc_17692_n1846_bF_buf8), .Y(_abc_17692_n12896) );
  AND2X2 AND2X2_5317 ( .A(_abc_17692_n12896), .B(_abc_17692_n12893), .Y(_abc_17692_n12897) );
  AND2X2 AND2X2_5318 ( .A(_abc_17692_n12900), .B(state_10_bF_buf4), .Y(_abc_17692_n12901) );
  AND2X2 AND2X2_5319 ( .A(_abc_17692_n12901), .B(_abc_17692_n12865), .Y(_abc_17692_n12902) );
  AND2X2 AND2X2_532 ( .A(sum_1_), .B(\key_in[65] ), .Y(_abc_17692_n1900) );
  AND2X2 AND2X2_5320 ( .A(_abc_17692_n12792), .B(_abc_17692_n12739), .Y(_abc_17692_n12904) );
  AND2X2 AND2X2_5321 ( .A(_abc_17692_n12786), .B(_abc_17692_n12737), .Y(_abc_17692_n12907) );
  AND2X2 AND2X2_5322 ( .A(_abc_17692_n12906), .B(_abc_17692_n12908), .Y(_abc_17692_n12909) );
  AND2X2 AND2X2_5323 ( .A(_abc_17692_n12909), .B(_abc_17692_n1863_bF_buf7), .Y(_abc_17692_n12910) );
  AND2X2 AND2X2_5324 ( .A(_abc_17692_n12681), .B(workunit1_30_), .Y(_abc_17692_n12911) );
  AND2X2 AND2X2_5325 ( .A(_abc_17692_n12806), .B(_abc_17692_n12912), .Y(_abc_17692_n12913) );
  AND2X2 AND2X2_5326 ( .A(_abc_17692_n12916), .B(_abc_17692_n1877_bF_buf7), .Y(_abc_17692_n12917) );
  AND2X2 AND2X2_5327 ( .A(_abc_17692_n12917), .B(_abc_17692_n12915), .Y(_abc_17692_n12918) );
  AND2X2 AND2X2_5328 ( .A(_abc_17692_n12816), .B(_abc_17692_n12713), .Y(_abc_17692_n12919) );
  AND2X2 AND2X2_5329 ( .A(_abc_17692_n12922), .B(_abc_17692_n1846_bF_buf7), .Y(_abc_17692_n12923) );
  AND2X2 AND2X2_533 ( .A(_abc_17692_n1901_1), .B(_abc_17692_n1902), .Y(_abc_17692_n1903) );
  AND2X2 AND2X2_5330 ( .A(_abc_17692_n12923), .B(_abc_17692_n12921), .Y(_abc_17692_n12924) );
  AND2X2 AND2X2_5331 ( .A(_abc_17692_n12929), .B(_abc_17692_n1830_bF_buf7), .Y(_abc_17692_n12930) );
  AND2X2 AND2X2_5332 ( .A(_abc_17692_n12930), .B(_abc_17692_n12928), .Y(_abc_17692_n12931) );
  AND2X2 AND2X2_5333 ( .A(_abc_17692_n12934), .B(state_14_bF_buf4), .Y(_abc_17692_n12935) );
  AND2X2 AND2X2_5334 ( .A(_abc_17692_n8383_bF_buf3), .B(workunit1_31_), .Y(_abc_17692_n12936) );
  AND2X2 AND2X2_5335 ( .A(state_8_bF_buf6), .B(\data_in1[31] ), .Y(_abc_17692_n12937) );
  AND2X2 AND2X2_5336 ( .A(_abc_17692_n12941), .B(_abc_17692_n12943), .Y(_abc_17692_n12944) );
  AND2X2 AND2X2_5337 ( .A(_abc_17692_n12944), .B(selectslice_0_), .Y(_abc_17692_n12945) );
  AND2X2 AND2X2_5338 ( .A(_abc_17692_n12942), .B(sum_11_), .Y(_abc_17692_n12946) );
  AND2X2 AND2X2_5339 ( .A(_abc_17692_n709), .B(sum_0_), .Y(_abc_17692_n12947) );
  AND2X2 AND2X2_534 ( .A(_abc_17692_n1903), .B(_abc_17692_n1867_1), .Y(_abc_17692_n1904) );
  AND2X2 AND2X2_5340 ( .A(_abc_17692_n12944), .B(selectslice_1_), .Y(_abc_17692_n12950) );
  AND2X2 AND2X2_5341 ( .A(_abc_17692_n12942), .B(sum_12_), .Y(_abc_17692_n12951) );
  AND2X2 AND2X2_5342 ( .A(_abc_17692_n709), .B(sum_1_), .Y(_abc_17692_n12952) );
  AND2X2 AND2X2_5343 ( .A(_abc_17692_n12955), .B(state_2_), .Y(_abc_10892_n6074) );
  AND2X2 AND2X2_5344 ( .A(while_flag), .B(state_13_), .Y(_abc_10892_n7323) );
  AND2X2 AND2X2_5345 ( .A(modereg), .B(state_2_), .Y(_abc_10892_n7419) );
  AND2X2 AND2X2_535 ( .A(_abc_17692_n1906), .B(_abc_17692_n1868), .Y(_abc_17692_n1907) );
  AND2X2 AND2X2_536 ( .A(_abc_17692_n1899), .B(_abc_17692_n1908), .Y(_abc_17692_n1909) );
  AND2X2 AND2X2_537 ( .A(_abc_17692_n1897), .B(_abc_17692_n1815_1), .Y(_abc_17692_n1910) );
  AND2X2 AND2X2_538 ( .A(_abc_17692_n1894), .B(_abc_17692_n1890), .Y(_abc_17692_n1911) );
  AND2X2 AND2X2_539 ( .A(_abc_17692_n1913), .B(_abc_17692_n1914), .Y(_abc_17692_n1915) );
  AND2X2 AND2X2_54 ( .A(_abc_17692_n767), .B(_abc_17692_n766_1), .Y(data_out2_13__FF_INPUT) );
  AND2X2 AND2X2_540 ( .A(_abc_17692_n1912), .B(_abc_17692_n1915), .Y(_abc_17692_n1916) );
  AND2X2 AND2X2_541 ( .A(_abc_17692_n1917), .B(workunit2_1_bF_buf2), .Y(_abc_17692_n1918) );
  AND2X2 AND2X2_542 ( .A(_abc_17692_n1920), .B(_abc_17692_n1921), .Y(_abc_17692_n1922) );
  AND2X2 AND2X2_543 ( .A(_abc_17692_n1922), .B(_abc_17692_n1919_1), .Y(_abc_17692_n1923) );
  AND2X2 AND2X2_544 ( .A(_abc_17692_n1875), .B(_abc_17692_n1814), .Y(_abc_17692_n1925) );
  AND2X2 AND2X2_545 ( .A(_abc_17692_n1924), .B(_abc_17692_n1926), .Y(_abc_17692_n1928) );
  AND2X2 AND2X2_546 ( .A(_abc_17692_n1929), .B(_abc_17692_n1877_bF_buf9), .Y(_abc_17692_n1930) );
  AND2X2 AND2X2_547 ( .A(_abc_17692_n1930), .B(_abc_17692_n1927), .Y(_abc_17692_n1931) );
  AND2X2 AND2X2_548 ( .A(_abc_17692_n1831), .B(_abc_17692_n1814), .Y(_abc_17692_n1932) );
  AND2X2 AND2X2_549 ( .A(sum_1_), .B(\key_in[1] ), .Y(_abc_17692_n1934) );
  AND2X2 AND2X2_55 ( .A(_abc_17692_n770), .B(_abc_17692_n769), .Y(data_out2_14__FF_INPUT) );
  AND2X2 AND2X2_550 ( .A(_abc_17692_n1935), .B(_abc_17692_n1936), .Y(_abc_17692_n1937) );
  AND2X2 AND2X2_551 ( .A(_abc_17692_n1937), .B(_abc_17692_n1820), .Y(_abc_17692_n1938) );
  AND2X2 AND2X2_552 ( .A(_abc_17692_n1940), .B(_abc_17692_n1821), .Y(_abc_17692_n1941) );
  AND2X2 AND2X2_553 ( .A(_abc_17692_n1899), .B(_abc_17692_n1942), .Y(_abc_17692_n1943) );
  AND2X2 AND2X2_554 ( .A(_abc_17692_n1944), .B(_abc_17692_n1945), .Y(_abc_17692_n1946) );
  AND2X2 AND2X2_555 ( .A(_abc_17692_n1912), .B(_abc_17692_n1946), .Y(_abc_17692_n1947) );
  AND2X2 AND2X2_556 ( .A(_abc_17692_n1948), .B(workunit2_1_bF_buf0), .Y(_abc_17692_n1949) );
  AND2X2 AND2X2_557 ( .A(_abc_17692_n1950), .B(_abc_17692_n1951), .Y(_abc_17692_n1952) );
  AND2X2 AND2X2_558 ( .A(_abc_17692_n1952), .B(_abc_17692_n1919_1), .Y(_abc_17692_n1953) );
  AND2X2 AND2X2_559 ( .A(_abc_17692_n1956), .B(_abc_17692_n1957), .Y(_abc_17692_n1958) );
  AND2X2 AND2X2_56 ( .A(_abc_17692_n773), .B(_abc_17692_n772), .Y(data_out2_15__FF_INPUT) );
  AND2X2 AND2X2_560 ( .A(_abc_17692_n1959), .B(_abc_17692_n1830_bF_buf9), .Y(_abc_17692_n1960) );
  AND2X2 AND2X2_561 ( .A(_abc_17692_n1960), .B(_abc_17692_n1955), .Y(_abc_17692_n1961) );
  AND2X2 AND2X2_562 ( .A(_abc_17692_n1843), .B(_abc_17692_n1814), .Y(_abc_17692_n1962) );
  AND2X2 AND2X2_563 ( .A(sum_1_), .B(\key_in[33] ), .Y(_abc_17692_n1964) );
  AND2X2 AND2X2_564 ( .A(_abc_17692_n1965), .B(_abc_17692_n1966), .Y(_abc_17692_n1967) );
  AND2X2 AND2X2_565 ( .A(_abc_17692_n1967), .B(_abc_17692_n1835), .Y(_abc_17692_n1968) );
  AND2X2 AND2X2_566 ( .A(_abc_17692_n1969), .B(_abc_17692_n1970), .Y(_abc_17692_n1971_1) );
  AND2X2 AND2X2_567 ( .A(_abc_17692_n1972), .B(_abc_17692_n1836), .Y(_abc_17692_n1973) );
  AND2X2 AND2X2_568 ( .A(_abc_17692_n1976), .B(_abc_17692_n1977), .Y(_abc_17692_n1978) );
  AND2X2 AND2X2_569 ( .A(_abc_17692_n1975), .B(_abc_17692_n1979), .Y(_abc_17692_n1980) );
  AND2X2 AND2X2_57 ( .A(_abc_17692_n776), .B(_abc_17692_n775), .Y(data_out2_16__FF_INPUT) );
  AND2X2 AND2X2_570 ( .A(_abc_17692_n1980), .B(workunit2_1_bF_buf2), .Y(_abc_17692_n1981_1) );
  AND2X2 AND2X2_571 ( .A(_abc_17692_n1982), .B(_abc_17692_n1983), .Y(_abc_17692_n1984) );
  AND2X2 AND2X2_572 ( .A(_abc_17692_n1984), .B(_abc_17692_n1919_1), .Y(_abc_17692_n1985) );
  AND2X2 AND2X2_573 ( .A(_abc_17692_n1986), .B(_abc_17692_n1963), .Y(_abc_17692_n1987) );
  AND2X2 AND2X2_574 ( .A(_abc_17692_n1989), .B(_abc_17692_n1846_bF_buf9), .Y(_abc_17692_n1990) );
  AND2X2 AND2X2_575 ( .A(_abc_17692_n1990), .B(_abc_17692_n1988), .Y(_abc_17692_n1991) );
  AND2X2 AND2X2_576 ( .A(_abc_17692_n1859), .B(_abc_17692_n1814), .Y(_abc_17692_n1994) );
  AND2X2 AND2X2_577 ( .A(sum_1_), .B(\key_in[97] ), .Y(_abc_17692_n1995) );
  AND2X2 AND2X2_578 ( .A(_abc_17692_n1996), .B(_abc_17692_n1997), .Y(_abc_17692_n1998) );
  AND2X2 AND2X2_579 ( .A(_abc_17692_n1998), .B(_abc_17692_n1851), .Y(_abc_17692_n1999) );
  AND2X2 AND2X2_58 ( .A(_abc_17692_n779), .B(_abc_17692_n778), .Y(data_out2_17__FF_INPUT) );
  AND2X2 AND2X2_580 ( .A(_abc_17692_n2000), .B(_abc_17692_n2001), .Y(_abc_17692_n2002) );
  AND2X2 AND2X2_581 ( .A(_abc_17692_n2005), .B(_abc_17692_n1852_1), .Y(_abc_17692_n2006) );
  AND2X2 AND2X2_582 ( .A(_abc_17692_n2003), .B(_abc_17692_n2008), .Y(_abc_17692_n2009) );
  AND2X2 AND2X2_583 ( .A(_abc_17692_n1899), .B(_abc_17692_n2007), .Y(_abc_17692_n2011) );
  AND2X2 AND2X2_584 ( .A(_abc_17692_n2002), .B(_abc_17692_n1912), .Y(_abc_17692_n2012) );
  AND2X2 AND2X2_585 ( .A(_abc_17692_n2010), .B(_abc_17692_n2014), .Y(_abc_17692_n2015) );
  AND2X2 AND2X2_586 ( .A(_abc_17692_n2013), .B(workunit2_1_bF_buf0), .Y(_abc_17692_n2018) );
  AND2X2 AND2X2_587 ( .A(_abc_17692_n2009), .B(_abc_17692_n1919_1), .Y(_abc_17692_n2019) );
  AND2X2 AND2X2_588 ( .A(_abc_17692_n2021), .B(_abc_17692_n1863_bF_buf9), .Y(_abc_17692_n2022) );
  AND2X2 AND2X2_589 ( .A(_abc_17692_n2022), .B(_abc_17692_n2016_1), .Y(_abc_17692_n2023) );
  AND2X2 AND2X2_59 ( .A(_abc_17692_n782), .B(_abc_17692_n781), .Y(data_out2_18__FF_INPUT) );
  AND2X2 AND2X2_590 ( .A(_abc_17692_n2024), .B(state_6_bF_buf3), .Y(_abc_17692_n2025) );
  AND2X2 AND2X2_591 ( .A(_abc_17692_n2026), .B(_abc_17692_n2027), .Y(_abc_17692_n2028) );
  AND2X2 AND2X2_592 ( .A(_abc_17692_n2030), .B(_abc_17692_n1877_bF_buf8), .Y(_abc_17692_n2031) );
  AND2X2 AND2X2_593 ( .A(_abc_17692_n2031), .B(_abc_17692_n2029), .Y(_abc_17692_n2032) );
  AND2X2 AND2X2_594 ( .A(_abc_17692_n1958), .B(_abc_17692_n2033), .Y(_abc_17692_n2034) );
  AND2X2 AND2X2_595 ( .A(_abc_17692_n2036), .B(_abc_17692_n1830_bF_buf8), .Y(_abc_17692_n2037) );
  AND2X2 AND2X2_596 ( .A(_abc_17692_n2037), .B(_abc_17692_n2035), .Y(_abc_17692_n2038) );
  AND2X2 AND2X2_597 ( .A(_abc_17692_n2041), .B(_abc_17692_n1863_bF_buf8), .Y(_abc_17692_n2042) );
  AND2X2 AND2X2_598 ( .A(_abc_17692_n2042), .B(_abc_17692_n2040), .Y(_abc_17692_n2043) );
  AND2X2 AND2X2_599 ( .A(_abc_17692_n2046), .B(_abc_17692_n2047), .Y(_abc_17692_n2048) );
  AND2X2 AND2X2_6 ( .A(_abc_17692_n632), .B(delta_6_), .Y(delta_6__FF_INPUT) );
  AND2X2 AND2X2_60 ( .A(_abc_17692_n785), .B(_abc_17692_n784), .Y(data_out2_19__FF_INPUT) );
  AND2X2 AND2X2_600 ( .A(_abc_17692_n2049_1), .B(_abc_17692_n1846_bF_buf8), .Y(_abc_17692_n2050) );
  AND2X2 AND2X2_601 ( .A(_abc_17692_n2050), .B(_abc_17692_n2044), .Y(_abc_17692_n2051) );
  AND2X2 AND2X2_602 ( .A(_abc_17692_n2053), .B(state_7_bF_buf2), .Y(_abc_17692_n2054) );
  AND2X2 AND2X2_603 ( .A(_abc_17692_n1885_bF_buf3), .B(workunit2_1_bF_buf1), .Y(_abc_17692_n2055) );
  AND2X2 AND2X2_604 ( .A(state_8_bF_buf8), .B(\data_in2[1] ), .Y(_abc_17692_n2056) );
  AND2X2 AND2X2_605 ( .A(workunit1_2_), .B(workunit1_7_), .Y(_abc_17692_n2061) );
  AND2X2 AND2X2_606 ( .A(_abc_17692_n2062_1), .B(_abc_17692_n2063), .Y(_abc_17692_n2064) );
  AND2X2 AND2X2_607 ( .A(_abc_17692_n2060), .B(_abc_17692_n2066), .Y(_abc_17692_n2067) );
  AND2X2 AND2X2_608 ( .A(_abc_17692_n1895), .B(_abc_17692_n1896), .Y(_abc_17692_n2068) );
  AND2X2 AND2X2_609 ( .A(_abc_17692_n2068), .B(_abc_17692_n2065), .Y(_abc_17692_n2069) );
  AND2X2 AND2X2_61 ( .A(_abc_17692_n788), .B(_abc_17692_n787), .Y(data_out2_20__FF_INPUT) );
  AND2X2 AND2X2_610 ( .A(_abc_17692_n1913), .B(_abc_17692_n1901_1), .Y(_abc_17692_n2071) );
  AND2X2 AND2X2_611 ( .A(sum_2_), .B(\key_in[66] ), .Y(_abc_17692_n2072) );
  AND2X2 AND2X2_612 ( .A(_abc_17692_n2073), .B(_abc_17692_n2074), .Y(_abc_17692_n2075) );
  AND2X2 AND2X2_613 ( .A(_abc_17692_n2077), .B(_abc_17692_n2079), .Y(_abc_17692_n2080) );
  AND2X2 AND2X2_614 ( .A(_abc_17692_n2082), .B(_abc_17692_n2083), .Y(_abc_17692_n2084) );
  AND2X2 AND2X2_615 ( .A(_abc_17692_n2078), .B(_abc_17692_n2075), .Y(_abc_17692_n2085) );
  AND2X2 AND2X2_616 ( .A(_abc_17692_n2071), .B(_abc_17692_n2076), .Y(_abc_17692_n2086) );
  AND2X2 AND2X2_617 ( .A(_abc_17692_n2081), .B(_abc_17692_n2088), .Y(_abc_17692_n2089) );
  AND2X2 AND2X2_618 ( .A(_abc_17692_n2084), .B(_abc_17692_n2087_1), .Y(_abc_17692_n2092) );
  AND2X2 AND2X2_619 ( .A(_abc_17692_n2070), .B(_abc_17692_n2080), .Y(_abc_17692_n2093) );
  AND2X2 AND2X2_62 ( .A(_abc_17692_n791), .B(_abc_17692_n790), .Y(data_out2_21__FF_INPUT) );
  AND2X2 AND2X2_620 ( .A(_abc_17692_n2090), .B(_abc_17692_n2095), .Y(_abc_17692_n2096) );
  AND2X2 AND2X2_621 ( .A(_abc_17692_n1922), .B(workunit2_1_bF_buf0), .Y(_abc_17692_n2097) );
  AND2X2 AND2X2_622 ( .A(_abc_17692_n2098), .B(_abc_17692_n2096), .Y(_abc_17692_n2099) );
  AND2X2 AND2X2_623 ( .A(_abc_17692_n2101), .B(_abc_17692_n1877_bF_buf7), .Y(_abc_17692_n2102) );
  AND2X2 AND2X2_624 ( .A(_abc_17692_n2102), .B(_abc_17692_n2100), .Y(_abc_17692_n2103) );
  AND2X2 AND2X2_625 ( .A(sum_2_), .B(\key_in[34] ), .Y(_abc_17692_n2105) );
  AND2X2 AND2X2_626 ( .A(_abc_17692_n2106), .B(_abc_17692_n2107), .Y(_abc_17692_n2108) );
  AND2X2 AND2X2_627 ( .A(_abc_17692_n2104), .B(_abc_17692_n2108), .Y(_abc_17692_n2109) );
  AND2X2 AND2X2_628 ( .A(_abc_17692_n1976), .B(_abc_17692_n1965), .Y(_abc_17692_n2110) );
  AND2X2 AND2X2_629 ( .A(_abc_17692_n2110), .B(_abc_17692_n2111), .Y(_abc_17692_n2112_1) );
  AND2X2 AND2X2_63 ( .A(_abc_17692_n794), .B(_abc_17692_n793), .Y(data_out2_22__FF_INPUT) );
  AND2X2 AND2X2_630 ( .A(_abc_17692_n2115), .B(_abc_17692_n2116), .Y(_abc_17692_n2117) );
  AND2X2 AND2X2_631 ( .A(_abc_17692_n2114), .B(_abc_17692_n2118), .Y(_abc_17692_n2119) );
  AND2X2 AND2X2_632 ( .A(_abc_17692_n2121), .B(_abc_17692_n2122), .Y(_abc_17692_n2123) );
  AND2X2 AND2X2_633 ( .A(_abc_17692_n2120), .B(_abc_17692_n2124), .Y(_abc_17692_n2125) );
  AND2X2 AND2X2_634 ( .A(_abc_17692_n1984), .B(workunit2_1_bF_buf3), .Y(_abc_17692_n2126) );
  AND2X2 AND2X2_635 ( .A(_abc_17692_n2127), .B(_abc_17692_n2125), .Y(_abc_17692_n2128) );
  AND2X2 AND2X2_636 ( .A(_abc_17692_n2130), .B(_abc_17692_n1846_bF_buf7), .Y(_abc_17692_n2131) );
  AND2X2 AND2X2_637 ( .A(_abc_17692_n2131), .B(_abc_17692_n2129), .Y(_abc_17692_n2132) );
  AND2X2 AND2X2_638 ( .A(sum_2_), .B(\key_in[2] ), .Y(_abc_17692_n2134) );
  AND2X2 AND2X2_639 ( .A(_abc_17692_n2135), .B(_abc_17692_n2136), .Y(_abc_17692_n2137_1) );
  AND2X2 AND2X2_64 ( .A(_abc_17692_n797), .B(_abc_17692_n796), .Y(data_out2_23__FF_INPUT) );
  AND2X2 AND2X2_640 ( .A(_abc_17692_n2133), .B(_abc_17692_n2137_1), .Y(_abc_17692_n2138) );
  AND2X2 AND2X2_641 ( .A(_abc_17692_n2139), .B(_abc_17692_n2140), .Y(_abc_17692_n2141) );
  AND2X2 AND2X2_642 ( .A(_abc_17692_n1944), .B(_abc_17692_n1935), .Y(_abc_17692_n2143) );
  AND2X2 AND2X2_643 ( .A(_abc_17692_n2143), .B(_abc_17692_n2144), .Y(_abc_17692_n2145) );
  AND2X2 AND2X2_644 ( .A(_abc_17692_n2142), .B(_abc_17692_n2147), .Y(_abc_17692_n2148) );
  AND2X2 AND2X2_645 ( .A(_abc_17692_n2084), .B(_abc_17692_n2146), .Y(_abc_17692_n2150) );
  AND2X2 AND2X2_646 ( .A(_abc_17692_n2141), .B(_abc_17692_n2070), .Y(_abc_17692_n2151) );
  AND2X2 AND2X2_647 ( .A(_abc_17692_n2149), .B(_abc_17692_n2153), .Y(_abc_17692_n2154) );
  AND2X2 AND2X2_648 ( .A(_abc_17692_n1952), .B(workunit2_1_bF_buf2), .Y(_abc_17692_n2155) );
  AND2X2 AND2X2_649 ( .A(_abc_17692_n1959), .B(_abc_17692_n2156), .Y(_abc_17692_n2157) );
  AND2X2 AND2X2_65 ( .A(_abc_17692_n800), .B(_abc_17692_n799_1), .Y(data_out2_24__FF_INPUT) );
  AND2X2 AND2X2_650 ( .A(_abc_17692_n2159), .B(_abc_17692_n2160), .Y(_abc_17692_n2161) );
  AND2X2 AND2X2_651 ( .A(_abc_17692_n1954), .B(_abc_17692_n1933), .Y(_abc_17692_n2162) );
  AND2X2 AND2X2_652 ( .A(_abc_17692_n2164), .B(_abc_17692_n1830_bF_buf7), .Y(_abc_17692_n2165) );
  AND2X2 AND2X2_653 ( .A(_abc_17692_n2165), .B(_abc_17692_n2158), .Y(_abc_17692_n2166) );
  AND2X2 AND2X2_654 ( .A(sum_2_), .B(\key_in[98] ), .Y(_abc_17692_n2170) );
  AND2X2 AND2X2_655 ( .A(_abc_17692_n2171), .B(_abc_17692_n2172), .Y(_abc_17692_n2173) );
  AND2X2 AND2X2_656 ( .A(_abc_17692_n2169), .B(_abc_17692_n2173), .Y(_abc_17692_n2174) );
  AND2X2 AND2X2_657 ( .A(_abc_17692_n2175), .B(_abc_17692_n2176), .Y(_abc_17692_n2177) );
  AND2X2 AND2X2_658 ( .A(_abc_17692_n2000), .B(_abc_17692_n1996), .Y(_abc_17692_n2179) );
  AND2X2 AND2X2_659 ( .A(_abc_17692_n2179), .B(_abc_17692_n2180), .Y(_abc_17692_n2181) );
  AND2X2 AND2X2_66 ( .A(_abc_17692_n803), .B(_abc_17692_n802), .Y(data_out2_25__FF_INPUT) );
  AND2X2 AND2X2_660 ( .A(_abc_17692_n2178), .B(_abc_17692_n2183), .Y(_abc_17692_n2184) );
  AND2X2 AND2X2_661 ( .A(_abc_17692_n2186), .B(_abc_17692_n2187), .Y(_abc_17692_n2188) );
  AND2X2 AND2X2_662 ( .A(_abc_17692_n2185), .B(_abc_17692_n2189), .Y(_abc_17692_n2190) );
  AND2X2 AND2X2_663 ( .A(_abc_17692_n2009), .B(workunit2_1_bF_buf1), .Y(_abc_17692_n2191) );
  AND2X2 AND2X2_664 ( .A(_abc_17692_n2016_1), .B(_abc_17692_n2192), .Y(_abc_17692_n2193) );
  AND2X2 AND2X2_665 ( .A(_abc_17692_n2195), .B(_abc_17692_n2196), .Y(_abc_17692_n2197) );
  AND2X2 AND2X2_666 ( .A(_abc_17692_n2199), .B(_abc_17692_n1863_bF_buf7), .Y(_abc_17692_n2200) );
  AND2X2 AND2X2_667 ( .A(_abc_17692_n2200), .B(_abc_17692_n2194), .Y(_abc_17692_n2201) );
  AND2X2 AND2X2_668 ( .A(_abc_17692_n2202), .B(state_6_bF_buf2), .Y(_abc_17692_n2203) );
  AND2X2 AND2X2_669 ( .A(_abc_17692_n2204), .B(_abc_17692_n2205), .Y(_abc_17692_n2206) );
  AND2X2 AND2X2_67 ( .A(_abc_17692_n806), .B(_abc_17692_n805), .Y(data_out2_26__FF_INPUT) );
  AND2X2 AND2X2_670 ( .A(_abc_17692_n2028), .B(_abc_17692_n1878), .Y(_abc_17692_n2207) );
  AND2X2 AND2X2_671 ( .A(_abc_17692_n2030), .B(_abc_17692_n2026), .Y(_abc_17692_n2210) );
  AND2X2 AND2X2_672 ( .A(_abc_17692_n2211_1), .B(_abc_17692_n1877_bF_buf6), .Y(_abc_17692_n2212) );
  AND2X2 AND2X2_673 ( .A(_abc_17692_n2212), .B(_abc_17692_n2209), .Y(_abc_17692_n2213) );
  AND2X2 AND2X2_674 ( .A(_abc_17692_n2154), .B(_abc_17692_n2214_1), .Y(_abc_17692_n2215) );
  AND2X2 AND2X2_675 ( .A(_abc_17692_n2217), .B(_abc_17692_n1830_bF_buf6), .Y(_abc_17692_n2218) );
  AND2X2 AND2X2_676 ( .A(_abc_17692_n2218), .B(_abc_17692_n2216), .Y(_abc_17692_n2219) );
  AND2X2 AND2X2_677 ( .A(_abc_17692_n2040), .B(_abc_17692_n2010), .Y(_abc_17692_n2221) );
  AND2X2 AND2X2_678 ( .A(_abc_17692_n2015), .B(_abc_17692_n1860), .Y(_abc_17692_n2223) );
  AND2X2 AND2X2_679 ( .A(_abc_17692_n2225), .B(_abc_17692_n1863_bF_buf6), .Y(_abc_17692_n2226_1) );
  AND2X2 AND2X2_68 ( .A(_abc_17692_n809), .B(_abc_17692_n808), .Y(data_out2_27__FF_INPUT) );
  AND2X2 AND2X2_680 ( .A(_abc_17692_n2226_1), .B(_abc_17692_n2222), .Y(_abc_17692_n2227) );
  AND2X2 AND2X2_681 ( .A(_abc_17692_n2044), .B(_abc_17692_n2046), .Y(_abc_17692_n2228) );
  AND2X2 AND2X2_682 ( .A(_abc_17692_n2230), .B(_abc_17692_n2231), .Y(_abc_17692_n2232) );
  AND2X2 AND2X2_683 ( .A(_abc_17692_n2048), .B(_abc_17692_n2045), .Y(_abc_17692_n2233) );
  AND2X2 AND2X2_684 ( .A(_abc_17692_n2235), .B(_abc_17692_n1846_bF_buf6), .Y(_abc_17692_n2236) );
  AND2X2 AND2X2_685 ( .A(_abc_17692_n2236), .B(_abc_17692_n2229), .Y(_abc_17692_n2237) );
  AND2X2 AND2X2_686 ( .A(_abc_17692_n2239), .B(state_7_bF_buf1), .Y(_abc_17692_n2240) );
  AND2X2 AND2X2_687 ( .A(_abc_17692_n1885_bF_buf2), .B(workunit2_2_), .Y(_abc_17692_n2241) );
  AND2X2 AND2X2_688 ( .A(state_8_bF_buf7), .B(\data_in2[2] ), .Y(_abc_17692_n2242_1) );
  AND2X2 AND2X2_689 ( .A(workunit1_3_), .B(workunit1_8_bF_buf2), .Y(_abc_17692_n2248) );
  AND2X2 AND2X2_69 ( .A(_abc_17692_n812), .B(_abc_17692_n811), .Y(data_out2_28__FF_INPUT) );
  AND2X2 AND2X2_690 ( .A(_abc_17692_n2249), .B(_abc_17692_n2250), .Y(_abc_17692_n2251) );
  AND2X2 AND2X2_691 ( .A(_abc_17692_n2082), .B(_abc_17692_n2254), .Y(_abc_17692_n2255) );
  AND2X2 AND2X2_692 ( .A(_abc_17692_n2257_1), .B(_abc_17692_n2253), .Y(_abc_17692_n2258) );
  AND2X2 AND2X2_693 ( .A(sum_3_), .B(\key_in[35] ), .Y(_abc_17692_n2260) );
  AND2X2 AND2X2_694 ( .A(_abc_17692_n2261), .B(_abc_17692_n2262), .Y(_abc_17692_n2263) );
  AND2X2 AND2X2_695 ( .A(_abc_17692_n2115), .B(_abc_17692_n2106), .Y(_abc_17692_n2266) );
  AND2X2 AND2X2_696 ( .A(_abc_17692_n2267), .B(_abc_17692_n2265), .Y(_abc_17692_n2268) );
  AND2X2 AND2X2_697 ( .A(_abc_17692_n2255), .B(_abc_17692_n2256), .Y(_abc_17692_n2270) );
  AND2X2 AND2X2_698 ( .A(_abc_17692_n2247), .B(_abc_17692_n2252), .Y(_abc_17692_n2271) );
  AND2X2 AND2X2_699 ( .A(_abc_17692_n2266), .B(_abc_17692_n2263), .Y(_abc_17692_n2273) );
  AND2X2 AND2X2_7 ( .A(_abc_17692_n632), .B(delta_9_), .Y(delta_9__FF_INPUT) );
  AND2X2 AND2X2_70 ( .A(_abc_17692_n815_1), .B(_abc_17692_n814_1), .Y(data_out2_29__FF_INPUT) );
  AND2X2 AND2X2_700 ( .A(_abc_17692_n2259), .B(_abc_17692_n2264), .Y(_abc_17692_n2274) );
  AND2X2 AND2X2_701 ( .A(_abc_17692_n2269), .B(_abc_17692_n2276), .Y(_abc_17692_n2277) );
  AND2X2 AND2X2_702 ( .A(_abc_17692_n2279), .B(_abc_17692_n2280), .Y(_abc_17692_n2281) );
  AND2X2 AND2X2_703 ( .A(_abc_17692_n2278_1), .B(_abc_17692_n2282), .Y(_abc_17692_n2283) );
  AND2X2 AND2X2_704 ( .A(_abc_17692_n2129), .B(_abc_17692_n2120), .Y(_abc_17692_n2284) );
  AND2X2 AND2X2_705 ( .A(_abc_17692_n2287), .B(_abc_17692_n2288), .Y(_abc_17692_n2289) );
  AND2X2 AND2X2_706 ( .A(_abc_17692_n2290), .B(_abc_17692_n1846_bF_buf5), .Y(_abc_17692_n2291) );
  AND2X2 AND2X2_707 ( .A(_abc_17692_n2291), .B(_abc_17692_n2286), .Y(_abc_17692_n2292) );
  AND2X2 AND2X2_708 ( .A(sum_3_), .B(\key_in[67] ), .Y(_abc_17692_n2294) );
  AND2X2 AND2X2_709 ( .A(_abc_17692_n2295), .B(_abc_17692_n2296), .Y(_abc_17692_n2297) );
  AND2X2 AND2X2_71 ( .A(_abc_17692_n818), .B(_abc_17692_n817), .Y(data_out2_30__FF_INPUT) );
  AND2X2 AND2X2_710 ( .A(_abc_17692_n2077), .B(_abc_17692_n2073), .Y(_abc_17692_n2300) );
  AND2X2 AND2X2_711 ( .A(_abc_17692_n2301), .B(_abc_17692_n2299), .Y(_abc_17692_n2302) );
  AND2X2 AND2X2_712 ( .A(_abc_17692_n2300), .B(_abc_17692_n2297), .Y(_abc_17692_n2304) );
  AND2X2 AND2X2_713 ( .A(_abc_17692_n2293), .B(_abc_17692_n2298), .Y(_abc_17692_n2305) );
  AND2X2 AND2X2_714 ( .A(_abc_17692_n2303), .B(_abc_17692_n2307), .Y(_abc_17692_n2308) );
  AND2X2 AND2X2_715 ( .A(_abc_17692_n2272), .B(_abc_17692_n2306), .Y(_abc_17692_n2310) );
  AND2X2 AND2X2_716 ( .A(_abc_17692_n2258), .B(_abc_17692_n2302), .Y(_abc_17692_n2311) );
  AND2X2 AND2X2_717 ( .A(_abc_17692_n2309), .B(_abc_17692_n2313), .Y(_abc_17692_n2314) );
  AND2X2 AND2X2_718 ( .A(_abc_17692_n2316), .B(_abc_17692_n2314), .Y(_abc_17692_n2317) );
  AND2X2 AND2X2_719 ( .A(_abc_17692_n2319), .B(_abc_17692_n1877_bF_buf5), .Y(_abc_17692_n2320) );
  AND2X2 AND2X2_72 ( .A(_abc_17692_n821), .B(_abc_17692_n820), .Y(data_out2_31__FF_INPUT) );
  AND2X2 AND2X2_720 ( .A(_abc_17692_n2320), .B(_abc_17692_n2318), .Y(_abc_17692_n2321) );
  AND2X2 AND2X2_721 ( .A(_abc_17692_n2139), .B(_abc_17692_n2135), .Y(_abc_17692_n2322) );
  AND2X2 AND2X2_722 ( .A(sum_3_), .B(\key_in[3] ), .Y(_abc_17692_n2323) );
  AND2X2 AND2X2_723 ( .A(_abc_17692_n2324), .B(_abc_17692_n2325), .Y(_abc_17692_n2326_1) );
  AND2X2 AND2X2_724 ( .A(_abc_17692_n2322), .B(_abc_17692_n2326_1), .Y(_abc_17692_n2327) );
  AND2X2 AND2X2_725 ( .A(_abc_17692_n2328), .B(_abc_17692_n2329_1), .Y(_abc_17692_n2330) );
  AND2X2 AND2X2_726 ( .A(_abc_17692_n2334), .B(_abc_17692_n2333), .Y(_abc_17692_n2335) );
  AND2X2 AND2X2_727 ( .A(_abc_17692_n2332), .B(_abc_17692_n2336), .Y(_abc_17692_n2337) );
  AND2X2 AND2X2_728 ( .A(_abc_17692_n2339), .B(_abc_17692_n2340_1), .Y(_abc_17692_n2341) );
  AND2X2 AND2X2_729 ( .A(_abc_17692_n2338), .B(_abc_17692_n2342), .Y(_abc_17692_n2343) );
  AND2X2 AND2X2_73 ( .A(_abc_17692_n824), .B(_abc_17692_n823), .Y(data_out1_0__FF_INPUT) );
  AND2X2 AND2X2_730 ( .A(_abc_17692_n2158), .B(_abc_17692_n2159), .Y(_abc_17692_n2344) );
  AND2X2 AND2X2_731 ( .A(_abc_17692_n2346), .B(_abc_17692_n2347), .Y(_abc_17692_n2348) );
  AND2X2 AND2X2_732 ( .A(_abc_17692_n2163), .B(_abc_17692_n2161), .Y(_abc_17692_n2350) );
  AND2X2 AND2X2_733 ( .A(_abc_17692_n2352), .B(_abc_17692_n1830_bF_buf5), .Y(_abc_17692_n2353) );
  AND2X2 AND2X2_734 ( .A(_abc_17692_n2353), .B(_abc_17692_n2345), .Y(_abc_17692_n2354) );
  AND2X2 AND2X2_735 ( .A(sum_3_), .B(\key_in[99] ), .Y(_abc_17692_n2358) );
  AND2X2 AND2X2_736 ( .A(_abc_17692_n2359), .B(_abc_17692_n2360), .Y(_abc_17692_n2361_1) );
  AND2X2 AND2X2_737 ( .A(_abc_17692_n2357), .B(_abc_17692_n2361_1), .Y(_abc_17692_n2362) );
  AND2X2 AND2X2_738 ( .A(_abc_17692_n2175), .B(_abc_17692_n2171), .Y(_abc_17692_n2363) );
  AND2X2 AND2X2_739 ( .A(_abc_17692_n2363), .B(_abc_17692_n2364), .Y(_abc_17692_n2365) );
  AND2X2 AND2X2_74 ( .A(_abc_17692_n827), .B(_abc_17692_n826), .Y(data_out1_1__FF_INPUT) );
  AND2X2 AND2X2_740 ( .A(_abc_17692_n2368), .B(_abc_17692_n2369), .Y(_abc_17692_n2370) );
  AND2X2 AND2X2_741 ( .A(_abc_17692_n2367), .B(_abc_17692_n2371), .Y(_abc_17692_n2372) );
  AND2X2 AND2X2_742 ( .A(_abc_17692_n2374), .B(_abc_17692_n2375), .Y(_abc_17692_n2376) );
  AND2X2 AND2X2_743 ( .A(_abc_17692_n2373), .B(_abc_17692_n2377), .Y(_abc_17692_n2378) );
  AND2X2 AND2X2_744 ( .A(_abc_17692_n2194), .B(_abc_17692_n2195), .Y(_abc_17692_n2379) );
  AND2X2 AND2X2_745 ( .A(_abc_17692_n2382), .B(_abc_17692_n2383), .Y(_abc_17692_n2384) );
  AND2X2 AND2X2_746 ( .A(_abc_17692_n2385), .B(_abc_17692_n1863_bF_buf5), .Y(_abc_17692_n2386) );
  AND2X2 AND2X2_747 ( .A(_abc_17692_n2386), .B(_abc_17692_n2381), .Y(_abc_17692_n2387) );
  AND2X2 AND2X2_748 ( .A(_abc_17692_n2388), .B(state_6_bF_buf1), .Y(_abc_17692_n2389) );
  AND2X2 AND2X2_749 ( .A(_abc_17692_n2390), .B(_abc_17692_n2391), .Y(_abc_17692_n2392) );
  AND2X2 AND2X2_75 ( .A(_abc_17692_n830), .B(_abc_17692_n829), .Y(data_out1_2__FF_INPUT) );
  AND2X2 AND2X2_750 ( .A(_abc_17692_n2206), .B(_abc_17692_n2208), .Y(_abc_17692_n2394) );
  AND2X2 AND2X2_751 ( .A(_abc_17692_n2211_1), .B(_abc_17692_n2204), .Y(_abc_17692_n2397) );
  AND2X2 AND2X2_752 ( .A(_abc_17692_n2398), .B(_abc_17692_n1877_bF_buf4), .Y(_abc_17692_n2399_1) );
  AND2X2 AND2X2_753 ( .A(_abc_17692_n2399_1), .B(_abc_17692_n2396), .Y(_abc_17692_n2400) );
  AND2X2 AND2X2_754 ( .A(_abc_17692_n2402), .B(_abc_17692_n2343), .Y(_abc_17692_n2403) );
  AND2X2 AND2X2_755 ( .A(_abc_17692_n2405), .B(_abc_17692_n1830_bF_buf4), .Y(_abc_17692_n2406) );
  AND2X2 AND2X2_756 ( .A(_abc_17692_n2406), .B(_abc_17692_n2404), .Y(_abc_17692_n2407) );
  AND2X2 AND2X2_757 ( .A(_abc_17692_n2222), .B(_abc_17692_n2185), .Y(_abc_17692_n2409) );
  AND2X2 AND2X2_758 ( .A(_abc_17692_n2190), .B(_abc_17692_n2224), .Y(_abc_17692_n2412) );
  AND2X2 AND2X2_759 ( .A(_abc_17692_n2414), .B(_abc_17692_n1863_bF_buf4), .Y(_abc_17692_n2415) );
  AND2X2 AND2X2_76 ( .A(_abc_17692_n833), .B(_abc_17692_n832), .Y(data_out1_3__FF_INPUT) );
  AND2X2 AND2X2_760 ( .A(_abc_17692_n2415), .B(_abc_17692_n2410), .Y(_abc_17692_n2416) );
  AND2X2 AND2X2_761 ( .A(_abc_17692_n2229), .B(_abc_17692_n2230), .Y(_abc_17692_n2417) );
  AND2X2 AND2X2_762 ( .A(_abc_17692_n2232), .B(_abc_17692_n2234), .Y(_abc_17692_n2420) );
  AND2X2 AND2X2_763 ( .A(_abc_17692_n2422), .B(_abc_17692_n1846_bF_buf4), .Y(_abc_17692_n2423) );
  AND2X2 AND2X2_764 ( .A(_abc_17692_n2423), .B(_abc_17692_n2418), .Y(_abc_17692_n2424) );
  AND2X2 AND2X2_765 ( .A(_abc_17692_n2426), .B(state_7_bF_buf0), .Y(_abc_17692_n2427) );
  AND2X2 AND2X2_766 ( .A(_abc_17692_n1885_bF_buf1), .B(workunit2_3_), .Y(_abc_17692_n2428) );
  AND2X2 AND2X2_767 ( .A(state_8_bF_buf6), .B(\data_in2[3] ), .Y(_abc_17692_n2429) );
  AND2X2 AND2X2_768 ( .A(_abc_17692_n2434), .B(_abc_17692_n2436), .Y(_abc_17692_n2437) );
  AND2X2 AND2X2_769 ( .A(_abc_17692_n2435), .B(workunit1_0_), .Y(_abc_17692_n2439) );
  AND2X2 AND2X2_77 ( .A(_abc_17692_n836_1), .B(_abc_17692_n835), .Y(data_out1_4__FF_INPUT) );
  AND2X2 AND2X2_770 ( .A(_abc_17692_n1816), .B(workunit1_9_), .Y(_abc_17692_n2440) );
  AND2X2 AND2X2_771 ( .A(_abc_17692_n2442), .B(_abc_17692_n2438), .Y(_abc_17692_n2443) );
  AND2X2 AND2X2_772 ( .A(_abc_17692_n2256), .B(_abc_17692_n2061), .Y(_abc_17692_n2444) );
  AND2X2 AND2X2_773 ( .A(_abc_17692_n2066), .B(_abc_17692_n2256), .Y(_abc_17692_n2446) );
  AND2X2 AND2X2_774 ( .A(_abc_17692_n2060), .B(_abc_17692_n2446), .Y(_abc_17692_n2447) );
  AND2X2 AND2X2_775 ( .A(_abc_17692_n2448), .B(_abc_17692_n2443), .Y(_abc_17692_n2449) );
  AND2X2 AND2X2_776 ( .A(_abc_17692_n2441), .B(workunit1_4_), .Y(_abc_17692_n2450) );
  AND2X2 AND2X2_777 ( .A(_abc_17692_n2437), .B(_abc_17692_n2433), .Y(_abc_17692_n2451) );
  AND2X2 AND2X2_778 ( .A(_abc_17692_n2455), .B(_abc_17692_n2453), .Y(_abc_17692_n2456) );
  AND2X2 AND2X2_779 ( .A(_abc_17692_n2456), .B(_abc_17692_n2452), .Y(_abc_17692_n2457) );
  AND2X2 AND2X2_78 ( .A(_abc_17692_n839), .B(_abc_17692_n838), .Y(data_out1_5__FF_INPUT) );
  AND2X2 AND2X2_780 ( .A(_abc_17692_n2326_1), .B(_abc_17692_n2134), .Y(_abc_17692_n2460) );
  AND2X2 AND2X2_781 ( .A(_abc_17692_n2137_1), .B(_abc_17692_n2326_1), .Y(_abc_17692_n2462_1) );
  AND2X2 AND2X2_782 ( .A(_abc_17692_n2133), .B(_abc_17692_n2462_1), .Y(_abc_17692_n2463) );
  AND2X2 AND2X2_783 ( .A(sum_4_), .B(\key_in[4] ), .Y(_abc_17692_n2465) );
  AND2X2 AND2X2_784 ( .A(_abc_17692_n2466), .B(_abc_17692_n2467), .Y(_abc_17692_n2468) );
  AND2X2 AND2X2_785 ( .A(_abc_17692_n2464), .B(_abc_17692_n2468), .Y(_abc_17692_n2469_1) );
  AND2X2 AND2X2_786 ( .A(_abc_17692_n2472), .B(_abc_17692_n2470), .Y(_abc_17692_n2473) );
  AND2X2 AND2X2_787 ( .A(_abc_17692_n2473), .B(_abc_17692_n2474), .Y(_abc_17692_n2475) );
  AND2X2 AND2X2_788 ( .A(_abc_17692_n2459_1), .B(_abc_17692_n2476), .Y(_abc_17692_n2477) );
  AND2X2 AND2X2_789 ( .A(_abc_17692_n2478), .B(_abc_17692_n2458), .Y(_abc_17692_n2479_1) );
  AND2X2 AND2X2_79 ( .A(_abc_17692_n842), .B(_abc_17692_n841), .Y(data_out1_6__FF_INPUT) );
  AND2X2 AND2X2_790 ( .A(_abc_17692_n2480), .B(workunit2_4_), .Y(_abc_17692_n2481) );
  AND2X2 AND2X2_791 ( .A(_abc_17692_n2483), .B(_abc_17692_n2482), .Y(_abc_17692_n2484) );
  AND2X2 AND2X2_792 ( .A(_abc_17692_n2345), .B(_abc_17692_n2346), .Y(_abc_17692_n2487) );
  AND2X2 AND2X2_793 ( .A(_abc_17692_n2351), .B(_abc_17692_n2348), .Y(_abc_17692_n2490_1) );
  AND2X2 AND2X2_794 ( .A(_abc_17692_n2492), .B(_abc_17692_n1830_bF_buf3), .Y(_abc_17692_n2493) );
  AND2X2 AND2X2_795 ( .A(_abc_17692_n2493), .B(_abc_17692_n2488), .Y(_abc_17692_n2494) );
  AND2X2 AND2X2_796 ( .A(sum_4_), .B(\key_in[68] ), .Y(_abc_17692_n2495) );
  AND2X2 AND2X2_797 ( .A(_abc_17692_n2496), .B(_abc_17692_n2497), .Y(_abc_17692_n2498) );
  AND2X2 AND2X2_798 ( .A(_abc_17692_n2297), .B(_abc_17692_n2072), .Y(_abc_17692_n2499) );
  AND2X2 AND2X2_799 ( .A(_abc_17692_n2075), .B(_abc_17692_n2297), .Y(_abc_17692_n2501) );
  AND2X2 AND2X2_8 ( .A(_abc_17692_n632), .B(delta_10_), .Y(delta_10__FF_INPUT) );
  AND2X2 AND2X2_80 ( .A(_abc_17692_n845), .B(_abc_17692_n844), .Y(data_out1_7__FF_INPUT) );
  AND2X2 AND2X2_800 ( .A(_abc_17692_n2078), .B(_abc_17692_n2501), .Y(_abc_17692_n2502) );
  AND2X2 AND2X2_801 ( .A(_abc_17692_n2503), .B(_abc_17692_n2498), .Y(_abc_17692_n2504) );
  AND2X2 AND2X2_802 ( .A(_abc_17692_n2506), .B(_abc_17692_n2505), .Y(_abc_17692_n2507) );
  AND2X2 AND2X2_803 ( .A(_abc_17692_n2508), .B(_abc_17692_n2458), .Y(_abc_17692_n2509) );
  AND2X2 AND2X2_804 ( .A(_abc_17692_n2510), .B(_abc_17692_n2459_1), .Y(_abc_17692_n2511) );
  AND2X2 AND2X2_805 ( .A(_abc_17692_n2515), .B(_abc_17692_n2513), .Y(_abc_17692_n2516) );
  AND2X2 AND2X2_806 ( .A(_abc_17692_n2519), .B(_abc_17692_n2517), .Y(_abc_17692_n2521) );
  AND2X2 AND2X2_807 ( .A(_abc_17692_n2522), .B(_abc_17692_n1877_bF_buf3), .Y(_abc_17692_n2523) );
  AND2X2 AND2X2_808 ( .A(_abc_17692_n2523), .B(_abc_17692_n2520), .Y(_abc_17692_n2524) );
  AND2X2 AND2X2_809 ( .A(_abc_17692_n2263), .B(_abc_17692_n2105), .Y(_abc_17692_n2525) );
  AND2X2 AND2X2_81 ( .A(_abc_17692_n848), .B(_abc_17692_n847), .Y(data_out1_8__FF_INPUT) );
  AND2X2 AND2X2_810 ( .A(_abc_17692_n2108), .B(_abc_17692_n2263), .Y(_abc_17692_n2527) );
  AND2X2 AND2X2_811 ( .A(_abc_17692_n2104), .B(_abc_17692_n2527), .Y(_abc_17692_n2528) );
  AND2X2 AND2X2_812 ( .A(sum_4_), .B(\key_in[36] ), .Y(_abc_17692_n2530) );
  AND2X2 AND2X2_813 ( .A(_abc_17692_n2531), .B(_abc_17692_n2532), .Y(_abc_17692_n2533) );
  AND2X2 AND2X2_814 ( .A(_abc_17692_n2529), .B(_abc_17692_n2533), .Y(_abc_17692_n2534) );
  AND2X2 AND2X2_815 ( .A(_abc_17692_n2537), .B(_abc_17692_n2535_1), .Y(_abc_17692_n2538_1) );
  AND2X2 AND2X2_816 ( .A(_abc_17692_n2538_1), .B(_abc_17692_n2539), .Y(_abc_17692_n2540) );
  AND2X2 AND2X2_817 ( .A(_abc_17692_n2459_1), .B(_abc_17692_n2541), .Y(_abc_17692_n2542) );
  AND2X2 AND2X2_818 ( .A(_abc_17692_n2543), .B(_abc_17692_n2458), .Y(_abc_17692_n2544) );
  AND2X2 AND2X2_819 ( .A(_abc_17692_n2545), .B(workunit2_4_), .Y(_abc_17692_n2546) );
  AND2X2 AND2X2_82 ( .A(_abc_17692_n851_1), .B(_abc_17692_n850_1), .Y(data_out1_9__FF_INPUT) );
  AND2X2 AND2X2_820 ( .A(_abc_17692_n2547), .B(_abc_17692_n2482), .Y(_abc_17692_n2548) );
  AND2X2 AND2X2_821 ( .A(_abc_17692_n2290), .B(_abc_17692_n2278_1), .Y(_abc_17692_n2550) );
  AND2X2 AND2X2_822 ( .A(_abc_17692_n2551), .B(_abc_17692_n2549), .Y(_abc_17692_n2552_1) );
  AND2X2 AND2X2_823 ( .A(_abc_17692_n2554), .B(_abc_17692_n1846_bF_buf3), .Y(_abc_17692_n2555) );
  AND2X2 AND2X2_824 ( .A(_abc_17692_n2555), .B(_abc_17692_n2553), .Y(_abc_17692_n2556) );
  AND2X2 AND2X2_825 ( .A(sum_4_), .B(\key_in[100] ), .Y(_abc_17692_n2560) );
  AND2X2 AND2X2_826 ( .A(_abc_17692_n2561), .B(_abc_17692_n2562), .Y(_abc_17692_n2563) );
  AND2X2 AND2X2_827 ( .A(_abc_17692_n2559), .B(_abc_17692_n2563), .Y(_abc_17692_n2564) );
  AND2X2 AND2X2_828 ( .A(_abc_17692_n2565), .B(_abc_17692_n2566), .Y(_abc_17692_n2567) );
  AND2X2 AND2X2_829 ( .A(_abc_17692_n2368), .B(_abc_17692_n2359), .Y(_abc_17692_n2569) );
  AND2X2 AND2X2_83 ( .A(_abc_17692_n854), .B(_abc_17692_n853), .Y(data_out1_10__FF_INPUT) );
  AND2X2 AND2X2_830 ( .A(_abc_17692_n2569), .B(_abc_17692_n2570), .Y(_abc_17692_n2571) );
  AND2X2 AND2X2_831 ( .A(_abc_17692_n2568), .B(_abc_17692_n2573), .Y(_abc_17692_n2574) );
  AND2X2 AND2X2_832 ( .A(_abc_17692_n2576), .B(_abc_17692_n2577), .Y(_abc_17692_n2578) );
  AND2X2 AND2X2_833 ( .A(_abc_17692_n2579), .B(_abc_17692_n2575), .Y(_abc_17692_n2580) );
  AND2X2 AND2X2_834 ( .A(_abc_17692_n2385), .B(_abc_17692_n2373), .Y(_abc_17692_n2581_1) );
  AND2X2 AND2X2_835 ( .A(_abc_17692_n2583), .B(_abc_17692_n2584), .Y(_abc_17692_n2585) );
  AND2X2 AND2X2_836 ( .A(_abc_17692_n2587), .B(_abc_17692_n1863_bF_buf3), .Y(_abc_17692_n2588) );
  AND2X2 AND2X2_837 ( .A(_abc_17692_n2588), .B(_abc_17692_n2582), .Y(_abc_17692_n2589) );
  AND2X2 AND2X2_838 ( .A(_abc_17692_n2590), .B(state_6_bF_buf0), .Y(_abc_17692_n2591) );
  AND2X2 AND2X2_839 ( .A(_abc_17692_n2395), .B(_abc_17692_n2392), .Y(_abc_17692_n2593) );
  AND2X2 AND2X2_84 ( .A(_abc_17692_n857), .B(_abc_17692_n856), .Y(data_out1_11__FF_INPUT) );
  AND2X2 AND2X2_840 ( .A(_abc_17692_n2398), .B(_abc_17692_n2390), .Y(_abc_17692_n2596) );
  AND2X2 AND2X2_841 ( .A(_abc_17692_n2597), .B(_abc_17692_n1877_bF_buf2), .Y(_abc_17692_n2598) );
  AND2X2 AND2X2_842 ( .A(_abc_17692_n2598), .B(_abc_17692_n2595), .Y(_abc_17692_n2599) );
  AND2X2 AND2X2_843 ( .A(_abc_17692_n2601), .B(_abc_17692_n2486), .Y(_abc_17692_n2602) );
  AND2X2 AND2X2_844 ( .A(_abc_17692_n2604), .B(_abc_17692_n1830_bF_buf2), .Y(_abc_17692_n2605) );
  AND2X2 AND2X2_845 ( .A(_abc_17692_n2605), .B(_abc_17692_n2603), .Y(_abc_17692_n2606) );
  AND2X2 AND2X2_846 ( .A(_abc_17692_n2410), .B(_abc_17692_n2382), .Y(_abc_17692_n2608_1) );
  AND2X2 AND2X2_847 ( .A(_abc_17692_n2413), .B(_abc_17692_n2384), .Y(_abc_17692_n2611) );
  AND2X2 AND2X2_848 ( .A(_abc_17692_n2613), .B(_abc_17692_n1863_bF_buf2), .Y(_abc_17692_n2614) );
  AND2X2 AND2X2_849 ( .A(_abc_17692_n2614), .B(_abc_17692_n2609), .Y(_abc_17692_n2615) );
  AND2X2 AND2X2_85 ( .A(_abc_17692_n860), .B(_abc_17692_n859), .Y(data_out1_12__FF_INPUT) );
  AND2X2 AND2X2_850 ( .A(_abc_17692_n2418), .B(_abc_17692_n2287), .Y(_abc_17692_n2616) );
  AND2X2 AND2X2_851 ( .A(_abc_17692_n2421), .B(_abc_17692_n2289), .Y(_abc_17692_n2620) );
  AND2X2 AND2X2_852 ( .A(_abc_17692_n2622), .B(_abc_17692_n1846_bF_buf2), .Y(_abc_17692_n2623) );
  AND2X2 AND2X2_853 ( .A(_abc_17692_n2623), .B(_abc_17692_n2617), .Y(_abc_17692_n2624) );
  AND2X2 AND2X2_854 ( .A(_abc_17692_n2626), .B(state_7_bF_buf4), .Y(_abc_17692_n2627) );
  AND2X2 AND2X2_855 ( .A(_abc_17692_n1885_bF_buf0), .B(workunit2_4_), .Y(_abc_17692_n2628) );
  AND2X2 AND2X2_856 ( .A(state_8_bF_buf5), .B(\data_in2[4] ), .Y(_abc_17692_n2629) );
  AND2X2 AND2X2_857 ( .A(_abc_17692_n2634_1), .B(_abc_17692_n2438), .Y(_abc_17692_n2635) );
  AND2X2 AND2X2_858 ( .A(workunit1_1_bF_buf0), .B(workunit1_10_), .Y(_abc_17692_n2636) );
  AND2X2 AND2X2_859 ( .A(_abc_17692_n2637), .B(_abc_17692_n2638), .Y(_abc_17692_n2639) );
  AND2X2 AND2X2_86 ( .A(_abc_17692_n863), .B(_abc_17692_n862), .Y(data_out1_13__FF_INPUT) );
  AND2X2 AND2X2_860 ( .A(_abc_17692_n2642), .B(_abc_17692_n2643), .Y(_abc_17692_n2644) );
  AND2X2 AND2X2_861 ( .A(_abc_17692_n2641), .B(_abc_17692_n2645), .Y(_abc_17692_n2646) );
  AND2X2 AND2X2_862 ( .A(_abc_17692_n2635), .B(_abc_17692_n2646), .Y(_abc_17692_n2647) );
  AND2X2 AND2X2_863 ( .A(_abc_17692_n2644), .B(workunit1_5_), .Y(_abc_17692_n2649) );
  AND2X2 AND2X2_864 ( .A(_abc_17692_n2640), .B(_abc_17692_n1817), .Y(_abc_17692_n2650) );
  AND2X2 AND2X2_865 ( .A(_abc_17692_n2648), .B(_abc_17692_n2651), .Y(_abc_17692_n2652) );
  AND2X2 AND2X2_866 ( .A(sum_5_), .B(\key_in[69] ), .Y(_abc_17692_n2655) );
  AND2X2 AND2X2_867 ( .A(_abc_17692_n2656), .B(_abc_17692_n2657), .Y(_abc_17692_n2658) );
  AND2X2 AND2X2_868 ( .A(_abc_17692_n2654), .B(_abc_17692_n2659), .Y(_abc_17692_n2661) );
  AND2X2 AND2X2_869 ( .A(_abc_17692_n2662), .B(_abc_17692_n2660), .Y(_abc_17692_n2663) );
  AND2X2 AND2X2_87 ( .A(_abc_17692_n866), .B(_abc_17692_n865), .Y(data_out1_14__FF_INPUT) );
  AND2X2 AND2X2_870 ( .A(_abc_17692_n2664), .B(_abc_17692_n2653), .Y(_abc_17692_n2665) );
  AND2X2 AND2X2_871 ( .A(_abc_17692_n2667), .B(_abc_17692_n2666), .Y(_abc_17692_n2668) );
  AND2X2 AND2X2_872 ( .A(_abc_17692_n2663), .B(_abc_17692_n2668), .Y(_abc_17692_n2669) );
  AND2X2 AND2X2_873 ( .A(_abc_17692_n2672), .B(_abc_17692_n2673), .Y(_abc_17692_n2674) );
  AND2X2 AND2X2_874 ( .A(_abc_17692_n2677), .B(_abc_17692_n2674), .Y(_abc_17692_n2678) );
  AND2X2 AND2X2_875 ( .A(_abc_17692_n2680), .B(_abc_17692_n1877_bF_buf1), .Y(_abc_17692_n2681) );
  AND2X2 AND2X2_876 ( .A(_abc_17692_n2681), .B(_abc_17692_n2679), .Y(_abc_17692_n2682) );
  AND2X2 AND2X2_877 ( .A(sum_5_), .B(\key_in[5] ), .Y(_abc_17692_n2684) );
  AND2X2 AND2X2_878 ( .A(_abc_17692_n1024), .B(_abc_17692_n2685), .Y(_abc_17692_n2686) );
  AND2X2 AND2X2_879 ( .A(_abc_17692_n2683), .B(_abc_17692_n2687), .Y(_abc_17692_n2689) );
  AND2X2 AND2X2_88 ( .A(_abc_17692_n869), .B(_abc_17692_n868), .Y(data_out1_15__FF_INPUT) );
  AND2X2 AND2X2_880 ( .A(_abc_17692_n2690), .B(_abc_17692_n2688), .Y(_abc_17692_n2691) );
  AND2X2 AND2X2_881 ( .A(_abc_17692_n2694), .B(_abc_17692_n2692), .Y(_abc_17692_n2695) );
  AND2X2 AND2X2_882 ( .A(_abc_17692_n2698), .B(_abc_17692_n2696), .Y(_abc_17692_n2699) );
  AND2X2 AND2X2_883 ( .A(_abc_17692_n2483), .B(workunit2_4_), .Y(_abc_17692_n2701) );
  AND2X2 AND2X2_884 ( .A(_abc_17692_n2488), .B(_abc_17692_n2702), .Y(_abc_17692_n2703) );
  AND2X2 AND2X2_885 ( .A(_abc_17692_n2491), .B(_abc_17692_n2485), .Y(_abc_17692_n2705) );
  AND2X2 AND2X2_886 ( .A(_abc_17692_n2707), .B(_abc_17692_n1830_bF_buf1), .Y(_abc_17692_n2708) );
  AND2X2 AND2X2_887 ( .A(_abc_17692_n2708), .B(_abc_17692_n2704), .Y(_abc_17692_n2709) );
  AND2X2 AND2X2_888 ( .A(_abc_17692_n2710), .B(_abc_17692_n2531), .Y(_abc_17692_n2711) );
  AND2X2 AND2X2_889 ( .A(sum_5_), .B(\key_in[37] ), .Y(_abc_17692_n2712) );
  AND2X2 AND2X2_89 ( .A(_abc_17692_n872), .B(_abc_17692_n871), .Y(data_out1_16__FF_INPUT) );
  AND2X2 AND2X2_890 ( .A(_abc_17692_n1024), .B(_abc_17692_n2713_1), .Y(_abc_17692_n2714) );
  AND2X2 AND2X2_891 ( .A(_abc_17692_n2711), .B(_abc_17692_n2716_1), .Y(_abc_17692_n2717) );
  AND2X2 AND2X2_892 ( .A(_abc_17692_n2718), .B(_abc_17692_n2715), .Y(_abc_17692_n2719) );
  AND2X2 AND2X2_893 ( .A(_abc_17692_n2723_1), .B(_abc_17692_n2722), .Y(_abc_17692_n2724) );
  AND2X2 AND2X2_894 ( .A(_abc_17692_n2721), .B(_abc_17692_n2725), .Y(_abc_17692_n2726) );
  AND2X2 AND2X2_895 ( .A(_abc_17692_n2728), .B(_abc_17692_n2729), .Y(_abc_17692_n2730) );
  AND2X2 AND2X2_896 ( .A(_abc_17692_n2727), .B(_abc_17692_n2731), .Y(_abc_17692_n2732) );
  AND2X2 AND2X2_897 ( .A(_abc_17692_n2547), .B(workunit2_4_), .Y(_abc_17692_n2734_1) );
  AND2X2 AND2X2_898 ( .A(_abc_17692_n2735), .B(_abc_17692_n2733), .Y(_abc_17692_n2737) );
  AND2X2 AND2X2_899 ( .A(_abc_17692_n2738), .B(_abc_17692_n1846_bF_buf1), .Y(_abc_17692_n2739) );
  AND2X2 AND2X2_9 ( .A(_abc_17692_n632), .B(delta_15_), .Y(delta_15__FF_INPUT) );
  AND2X2 AND2X2_90 ( .A(_abc_17692_n875_1), .B(_abc_17692_n874), .Y(data_out1_17__FF_INPUT) );
  AND2X2 AND2X2_900 ( .A(_abc_17692_n2739), .B(_abc_17692_n2736), .Y(_abc_17692_n2740) );
  AND2X2 AND2X2_901 ( .A(_abc_17692_n2565), .B(_abc_17692_n2561), .Y(_abc_17692_n2743) );
  AND2X2 AND2X2_902 ( .A(sum_5_), .B(\key_in[101] ), .Y(_abc_17692_n2744) );
  AND2X2 AND2X2_903 ( .A(_abc_17692_n2745_1), .B(_abc_17692_n2746), .Y(_abc_17692_n2747) );
  AND2X2 AND2X2_904 ( .A(_abc_17692_n2743), .B(_abc_17692_n2747), .Y(_abc_17692_n2748) );
  AND2X2 AND2X2_905 ( .A(_abc_17692_n2749), .B(_abc_17692_n2750), .Y(_abc_17692_n2751) );
  AND2X2 AND2X2_906 ( .A(_abc_17692_n2755), .B(_abc_17692_n2754), .Y(_abc_17692_n2756) );
  AND2X2 AND2X2_907 ( .A(_abc_17692_n2753), .B(_abc_17692_n2757_1), .Y(_abc_17692_n2758) );
  AND2X2 AND2X2_908 ( .A(_abc_17692_n2760), .B(_abc_17692_n2761), .Y(_abc_17692_n2762) );
  AND2X2 AND2X2_909 ( .A(_abc_17692_n2759), .B(_abc_17692_n2763), .Y(_abc_17692_n2764) );
  AND2X2 AND2X2_91 ( .A(_abc_17692_n878), .B(_abc_17692_n877), .Y(data_out1_18__FF_INPUT) );
  AND2X2 AND2X2_910 ( .A(_abc_17692_n2582), .B(_abc_17692_n2583), .Y(_abc_17692_n2765) );
  AND2X2 AND2X2_911 ( .A(_abc_17692_n2767), .B(_abc_17692_n2768), .Y(_abc_17692_n2769) );
  AND2X2 AND2X2_912 ( .A(_abc_17692_n2771), .B(_abc_17692_n1863_bF_buf1), .Y(_abc_17692_n2772) );
  AND2X2 AND2X2_913 ( .A(_abc_17692_n2772), .B(_abc_17692_n2766), .Y(_abc_17692_n2773) );
  AND2X2 AND2X2_914 ( .A(_abc_17692_n2774), .B(state_6_bF_buf4), .Y(_abc_17692_n2775) );
  AND2X2 AND2X2_915 ( .A(_abc_17692_n2594), .B(_abc_17692_n2516), .Y(_abc_17692_n2778) );
  AND2X2 AND2X2_916 ( .A(_abc_17692_n2597), .B(_abc_17692_n2513), .Y(_abc_17692_n2781) );
  AND2X2 AND2X2_917 ( .A(_abc_17692_n2782), .B(_abc_17692_n1877_bF_buf0), .Y(_abc_17692_n2783) );
  AND2X2 AND2X2_918 ( .A(_abc_17692_n2783), .B(_abc_17692_n2780), .Y(_abc_17692_n2784) );
  AND2X2 AND2X2_919 ( .A(_abc_17692_n2785), .B(_abc_17692_n2700), .Y(_abc_17692_n2786) );
  AND2X2 AND2X2_92 ( .A(_abc_17692_n881), .B(_abc_17692_n880), .Y(data_out1_19__FF_INPUT) );
  AND2X2 AND2X2_920 ( .A(_abc_17692_n2788), .B(_abc_17692_n1830_bF_buf0), .Y(_abc_17692_n2789) );
  AND2X2 AND2X2_921 ( .A(_abc_17692_n2789), .B(_abc_17692_n2787), .Y(_abc_17692_n2790) );
  AND2X2 AND2X2_922 ( .A(_abc_17692_n2609), .B(_abc_17692_n2575), .Y(_abc_17692_n2792) );
  AND2X2 AND2X2_923 ( .A(_abc_17692_n2612), .B(_abc_17692_n2580), .Y(_abc_17692_n2795) );
  AND2X2 AND2X2_924 ( .A(_abc_17692_n2797_1), .B(_abc_17692_n1863_bF_buf0), .Y(_abc_17692_n2798) );
  AND2X2 AND2X2_925 ( .A(_abc_17692_n2798), .B(_abc_17692_n2793), .Y(_abc_17692_n2799) );
  AND2X2 AND2X2_926 ( .A(_abc_17692_n2617), .B(_abc_17692_n2800_1), .Y(_abc_17692_n2801) );
  AND2X2 AND2X2_927 ( .A(_abc_17692_n2621), .B(_abc_17692_n2618), .Y(_abc_17692_n2803) );
  AND2X2 AND2X2_928 ( .A(_abc_17692_n2805), .B(_abc_17692_n1846_bF_buf0), .Y(_abc_17692_n2806) );
  AND2X2 AND2X2_929 ( .A(_abc_17692_n2806), .B(_abc_17692_n2802), .Y(_abc_17692_n2807) );
  AND2X2 AND2X2_93 ( .A(_abc_17692_n884), .B(_abc_17692_n883), .Y(data_out1_20__FF_INPUT) );
  AND2X2 AND2X2_930 ( .A(_abc_17692_n2809), .B(state_7_bF_buf3), .Y(_abc_17692_n2810) );
  AND2X2 AND2X2_931 ( .A(_abc_17692_n1885_bF_buf4), .B(workunit2_5_), .Y(_abc_17692_n2811) );
  AND2X2 AND2X2_932 ( .A(state_8_bF_buf4), .B(\data_in2[5] ), .Y(_abc_17692_n2812_1) );
  AND2X2 AND2X2_933 ( .A(_abc_17692_n2443), .B(_abc_17692_n2646), .Y(_abc_17692_n2816) );
  AND2X2 AND2X2_934 ( .A(_abc_17692_n2448), .B(_abc_17692_n2816), .Y(_abc_17692_n2817) );
  AND2X2 AND2X2_935 ( .A(_abc_17692_n2818), .B(_abc_17692_n2645), .Y(_abc_17692_n2819) );
  AND2X2 AND2X2_936 ( .A(workunit1_2_), .B(workunit1_11_bF_buf2), .Y(_abc_17692_n2822) );
  AND2X2 AND2X2_937 ( .A(_abc_17692_n2062_1), .B(_abc_17692_n2823), .Y(_abc_17692_n2824) );
  AND2X2 AND2X2_938 ( .A(_abc_17692_n2827), .B(_abc_17692_n2828), .Y(_abc_17692_n2829) );
  AND2X2 AND2X2_939 ( .A(_abc_17692_n2826), .B(_abc_17692_n2830_1), .Y(_abc_17692_n2831) );
  AND2X2 AND2X2_94 ( .A(_abc_17692_n887), .B(_abc_17692_n886), .Y(data_out1_21__FF_INPUT) );
  AND2X2 AND2X2_940 ( .A(_abc_17692_n2820), .B(_abc_17692_n2831), .Y(_abc_17692_n2832) );
  AND2X2 AND2X2_941 ( .A(_abc_17692_n2834), .B(_abc_17692_n2641), .Y(_abc_17692_n2835) );
  AND2X2 AND2X2_942 ( .A(_abc_17692_n2833), .B(_abc_17692_n2835), .Y(_abc_17692_n2836) );
  AND2X2 AND2X2_943 ( .A(_abc_17692_n2829), .B(workunit1_6_), .Y(_abc_17692_n2837) );
  AND2X2 AND2X2_944 ( .A(_abc_17692_n2825), .B(_abc_17692_n2821), .Y(_abc_17692_n2838) );
  AND2X2 AND2X2_945 ( .A(_abc_17692_n2836), .B(_abc_17692_n2839), .Y(_abc_17692_n2840) );
  AND2X2 AND2X2_946 ( .A(_abc_17692_n2498), .B(_abc_17692_n2658), .Y(_abc_17692_n2843) );
  AND2X2 AND2X2_947 ( .A(_abc_17692_n2503), .B(_abc_17692_n2843), .Y(_abc_17692_n2844) );
  AND2X2 AND2X2_948 ( .A(_abc_17692_n2845), .B(_abc_17692_n2656), .Y(_abc_17692_n2846) );
  AND2X2 AND2X2_949 ( .A(sum_6_), .B(\key_in[70] ), .Y(_abc_17692_n2849_1) );
  AND2X2 AND2X2_95 ( .A(_abc_17692_n890_1), .B(_abc_17692_n889_1), .Y(data_out1_22__FF_INPUT) );
  AND2X2 AND2X2_950 ( .A(_abc_17692_n2850), .B(_abc_17692_n2851), .Y(_abc_17692_n2852) );
  AND2X2 AND2X2_951 ( .A(_abc_17692_n2848), .B(_abc_17692_n2852), .Y(_abc_17692_n2853) );
  AND2X2 AND2X2_952 ( .A(_abc_17692_n2854), .B(_abc_17692_n2855), .Y(_abc_17692_n2856) );
  AND2X2 AND2X2_953 ( .A(_abc_17692_n2857), .B(_abc_17692_n2842), .Y(_abc_17692_n2858) );
  AND2X2 AND2X2_954 ( .A(_abc_17692_n2856), .B(_abc_17692_n2841), .Y(_abc_17692_n2859) );
  AND2X2 AND2X2_955 ( .A(_abc_17692_n2860), .B(workunit2_6_), .Y(_abc_17692_n2861) );
  AND2X2 AND2X2_956 ( .A(_abc_17692_n2863), .B(_abc_17692_n2862), .Y(_abc_17692_n2864) );
  AND2X2 AND2X2_957 ( .A(_abc_17692_n2867_1), .B(_abc_17692_n2865), .Y(_abc_17692_n2869) );
  AND2X2 AND2X2_958 ( .A(_abc_17692_n2870), .B(_abc_17692_n1877_bF_buf10), .Y(_abc_17692_n2871) );
  AND2X2 AND2X2_959 ( .A(_abc_17692_n2871), .B(_abc_17692_n2868), .Y(_abc_17692_n2872) );
  AND2X2 AND2X2_96 ( .A(_abc_17692_n893), .B(_abc_17692_n892), .Y(data_out1_23__FF_INPUT) );
  AND2X2 AND2X2_960 ( .A(_abc_17692_n2464), .B(_abc_17692_n2874), .Y(_abc_17692_n2875) );
  AND2X2 AND2X2_961 ( .A(_abc_17692_n2877), .B(_abc_17692_n2876), .Y(_abc_17692_n2878) );
  AND2X2 AND2X2_962 ( .A(sum_6_), .B(\key_in[6] ), .Y(_abc_17692_n2880) );
  AND2X2 AND2X2_963 ( .A(_abc_17692_n2881), .B(_abc_17692_n2882), .Y(_abc_17692_n2883) );
  AND2X2 AND2X2_964 ( .A(_abc_17692_n2879), .B(_abc_17692_n2883), .Y(_abc_17692_n2884) );
  AND2X2 AND2X2_965 ( .A(_abc_17692_n2885), .B(_abc_17692_n2886), .Y(_abc_17692_n2887) );
  AND2X2 AND2X2_966 ( .A(_abc_17692_n2842), .B(_abc_17692_n2888), .Y(_abc_17692_n2889) );
  AND2X2 AND2X2_967 ( .A(_abc_17692_n2890), .B(_abc_17692_n2841), .Y(_abc_17692_n2891) );
  AND2X2 AND2X2_968 ( .A(_abc_17692_n2892), .B(workunit2_6_), .Y(_abc_17692_n2893) );
  AND2X2 AND2X2_969 ( .A(_abc_17692_n2894), .B(_abc_17692_n2895), .Y(_abc_17692_n2896) );
  AND2X2 AND2X2_97 ( .A(_abc_17692_n896), .B(_abc_17692_n895), .Y(data_out1_24__FF_INPUT) );
  AND2X2 AND2X2_970 ( .A(_abc_17692_n2704), .B(_abc_17692_n2696), .Y(_abc_17692_n2897) );
  AND2X2 AND2X2_971 ( .A(_abc_17692_n2706), .B(_abc_17692_n2699), .Y(_abc_17692_n2901) );
  AND2X2 AND2X2_972 ( .A(_abc_17692_n2903), .B(_abc_17692_n1830_bF_buf10), .Y(_abc_17692_n2904) );
  AND2X2 AND2X2_973 ( .A(_abc_17692_n2904), .B(_abc_17692_n2898), .Y(_abc_17692_n2905) );
  AND2X2 AND2X2_974 ( .A(_abc_17692_n2716_1), .B(_abc_17692_n2533), .Y(_abc_17692_n2906) );
  AND2X2 AND2X2_975 ( .A(_abc_17692_n2529), .B(_abc_17692_n2906), .Y(_abc_17692_n2907) );
  AND2X2 AND2X2_976 ( .A(_abc_17692_n2909), .B(_abc_17692_n2908), .Y(_abc_17692_n2910) );
  AND2X2 AND2X2_977 ( .A(sum_6_), .B(\key_in[38] ), .Y(_abc_17692_n2912) );
  AND2X2 AND2X2_978 ( .A(_abc_17692_n2913), .B(_abc_17692_n2914), .Y(_abc_17692_n2915) );
  AND2X2 AND2X2_979 ( .A(_abc_17692_n2911), .B(_abc_17692_n2915), .Y(_abc_17692_n2916_1) );
  AND2X2 AND2X2_98 ( .A(_abc_17692_n899), .B(_abc_17692_n898), .Y(data_out1_25__FF_INPUT) );
  AND2X2 AND2X2_980 ( .A(_abc_17692_n2918), .B(_abc_17692_n2919_1), .Y(_abc_17692_n2920) );
  AND2X2 AND2X2_981 ( .A(_abc_17692_n2920), .B(_abc_17692_n2921), .Y(_abc_17692_n2922) );
  AND2X2 AND2X2_982 ( .A(_abc_17692_n2842), .B(_abc_17692_n2923), .Y(_abc_17692_n2924) );
  AND2X2 AND2X2_983 ( .A(_abc_17692_n2925), .B(_abc_17692_n2841), .Y(_abc_17692_n2926_1) );
  AND2X2 AND2X2_984 ( .A(_abc_17692_n2929), .B(_abc_17692_n2930), .Y(_abc_17692_n2931) );
  AND2X2 AND2X2_985 ( .A(_abc_17692_n2726), .B(workunit2_5_), .Y(_abc_17692_n2935) );
  AND2X2 AND2X2_986 ( .A(_abc_17692_n2938_1), .B(_abc_17692_n2936), .Y(_abc_17692_n2939) );
  AND2X2 AND2X2_987 ( .A(_abc_17692_n2934), .B(_abc_17692_n2939), .Y(_abc_17692_n2940) );
  AND2X2 AND2X2_988 ( .A(_abc_17692_n2941), .B(_abc_17692_n2932), .Y(_abc_17692_n2943) );
  AND2X2 AND2X2_989 ( .A(_abc_17692_n2944), .B(_abc_17692_n1846_bF_buf10), .Y(_abc_17692_n2945) );
  AND2X2 AND2X2_99 ( .A(_abc_17692_n902), .B(_abc_17692_n901), .Y(data_out1_26__FF_INPUT) );
  AND2X2 AND2X2_990 ( .A(_abc_17692_n2945), .B(_abc_17692_n2942), .Y(_abc_17692_n2946) );
  AND2X2 AND2X2_991 ( .A(_abc_17692_n2563), .B(_abc_17692_n2747), .Y(_abc_17692_n2949_1) );
  AND2X2 AND2X2_992 ( .A(_abc_17692_n2559), .B(_abc_17692_n2949_1), .Y(_abc_17692_n2950) );
  AND2X2 AND2X2_993 ( .A(_abc_17692_n2951), .B(_abc_17692_n2745_1), .Y(_abc_17692_n2952) );
  AND2X2 AND2X2_994 ( .A(sum_6_), .B(\key_in[102] ), .Y(_abc_17692_n2955) );
  AND2X2 AND2X2_995 ( .A(_abc_17692_n2956), .B(_abc_17692_n2957), .Y(_abc_17692_n2958) );
  AND2X2 AND2X2_996 ( .A(_abc_17692_n2954), .B(_abc_17692_n2958), .Y(_abc_17692_n2959) );
  AND2X2 AND2X2_997 ( .A(_abc_17692_n2960_1), .B(_abc_17692_n2961), .Y(_abc_17692_n2962) );
  AND2X2 AND2X2_998 ( .A(_abc_17692_n2963), .B(_abc_17692_n2842), .Y(_abc_17692_n2964) );
  AND2X2 AND2X2_999 ( .A(_abc_17692_n2962), .B(_abc_17692_n2841), .Y(_abc_17692_n2965) );
  BUFX2 BUFX2_1 ( .A(workunit2_12_), .Y(workunit2_12_bF_buf3) );
  BUFX2 BUFX2_10 ( .A(clock), .Y(clock_bF_buf12) );
  BUFX2 BUFX2_100 ( .A(_abc_17692_n1877), .Y(_abc_17692_n1877_bF_buf0) );
  BUFX2 BUFX2_101 ( .A(workunit1_14_), .Y(workunit1_14_bF_buf3) );
  BUFX2 BUFX2_102 ( .A(workunit1_14_), .Y(workunit1_14_bF_buf2) );
  BUFX2 BUFX2_103 ( .A(workunit1_14_), .Y(workunit1_14_bF_buf1) );
  BUFX2 BUFX2_104 ( .A(workunit1_14_), .Y(workunit1_14_bF_buf0) );
  BUFX2 BUFX2_105 ( .A(_abc_17692_n1846), .Y(_abc_17692_n1846_bF_buf10) );
  BUFX2 BUFX2_106 ( .A(_abc_17692_n1846), .Y(_abc_17692_n1846_bF_buf9) );
  BUFX2 BUFX2_107 ( .A(_abc_17692_n1846), .Y(_abc_17692_n1846_bF_buf8) );
  BUFX2 BUFX2_108 ( .A(_abc_17692_n1846), .Y(_abc_17692_n1846_bF_buf7) );
  BUFX2 BUFX2_109 ( .A(_abc_17692_n1846), .Y(_abc_17692_n1846_bF_buf6) );
  BUFX2 BUFX2_11 ( .A(clock), .Y(clock_bF_buf11) );
  BUFX2 BUFX2_110 ( .A(_abc_17692_n1846), .Y(_abc_17692_n1846_bF_buf5) );
  BUFX2 BUFX2_111 ( .A(_abc_17692_n1846), .Y(_abc_17692_n1846_bF_buf4) );
  BUFX2 BUFX2_112 ( .A(_abc_17692_n1846), .Y(_abc_17692_n1846_bF_buf3) );
  BUFX2 BUFX2_113 ( .A(_abc_17692_n1846), .Y(_abc_17692_n1846_bF_buf2) );
  BUFX2 BUFX2_114 ( .A(_abc_17692_n1846), .Y(_abc_17692_n1846_bF_buf1) );
  BUFX2 BUFX2_115 ( .A(_abc_17692_n1846), .Y(_abc_17692_n1846_bF_buf0) );
  BUFX2 BUFX2_116 ( .A(workunit1_11_), .Y(workunit1_11_bF_buf3) );
  BUFX2 BUFX2_117 ( .A(workunit1_11_), .Y(workunit1_11_bF_buf2) );
  BUFX2 BUFX2_118 ( .A(workunit1_11_), .Y(workunit1_11_bF_buf1) );
  BUFX2 BUFX2_119 ( .A(workunit1_11_), .Y(workunit1_11_bF_buf0) );
  BUFX2 BUFX2_12 ( .A(clock), .Y(clock_bF_buf10) );
  BUFX2 BUFX2_120 ( .A(workunit2_8_), .Y(workunit2_8_bF_buf3) );
  BUFX2 BUFX2_121 ( .A(workunit2_8_), .Y(workunit2_8_bF_buf2) );
  BUFX2 BUFX2_122 ( .A(workunit2_8_), .Y(workunit2_8_bF_buf1) );
  BUFX2 BUFX2_123 ( .A(workunit2_8_), .Y(workunit2_8_bF_buf0) );
  BUFX2 BUFX2_124 ( .A(workunit1_8_), .Y(workunit1_8_bF_buf3) );
  BUFX2 BUFX2_125 ( .A(workunit1_8_), .Y(workunit1_8_bF_buf2) );
  BUFX2 BUFX2_126 ( .A(workunit1_8_), .Y(workunit1_8_bF_buf1) );
  BUFX2 BUFX2_127 ( .A(workunit1_8_), .Y(workunit1_8_bF_buf0) );
  BUFX2 BUFX2_128 ( .A(workunit2_16_), .Y(workunit2_16_bF_buf3) );
  BUFX2 BUFX2_129 ( .A(workunit2_16_), .Y(workunit2_16_bF_buf2) );
  BUFX2 BUFX2_13 ( .A(clock), .Y(clock_bF_buf9) );
  BUFX2 BUFX2_130 ( .A(workunit2_16_), .Y(workunit2_16_bF_buf1) );
  BUFX2 BUFX2_131 ( .A(workunit2_16_), .Y(workunit2_16_bF_buf0) );
  BUFX2 BUFX2_132 ( .A(workunit2_10_), .Y(workunit2_10_bF_buf3) );
  BUFX2 BUFX2_133 ( .A(workunit2_10_), .Y(workunit2_10_bF_buf2) );
  BUFX2 BUFX2_134 ( .A(workunit2_10_), .Y(workunit2_10_bF_buf1) );
  BUFX2 BUFX2_135 ( .A(workunit2_10_), .Y(workunit2_10_bF_buf0) );
  BUFX2 BUFX2_136 ( .A(state_10_), .Y(state_10_bF_buf4) );
  BUFX2 BUFX2_137 ( .A(state_10_), .Y(state_10_bF_buf3) );
  BUFX2 BUFX2_138 ( .A(state_10_), .Y(state_10_bF_buf2) );
  BUFX2 BUFX2_139 ( .A(state_10_), .Y(state_10_bF_buf1) );
  BUFX2 BUFX2_14 ( .A(clock), .Y(clock_bF_buf8) );
  BUFX2 BUFX2_140 ( .A(state_10_), .Y(state_10_bF_buf0) );
  BUFX2 BUFX2_141 ( .A(state_8_), .Y(state_8_bF_buf9) );
  BUFX2 BUFX2_142 ( .A(state_8_), .Y(state_8_bF_buf8) );
  BUFX2 BUFX2_143 ( .A(state_8_), .Y(state_8_bF_buf7) );
  BUFX2 BUFX2_144 ( .A(state_8_), .Y(state_8_bF_buf6) );
  BUFX2 BUFX2_145 ( .A(state_8_), .Y(state_8_bF_buf5) );
  BUFX2 BUFX2_146 ( .A(state_8_), .Y(state_8_bF_buf4) );
  BUFX2 BUFX2_147 ( .A(state_8_), .Y(state_8_bF_buf3) );
  BUFX2 BUFX2_148 ( .A(state_8_), .Y(state_8_bF_buf2) );
  BUFX2 BUFX2_149 ( .A(state_8_), .Y(state_8_bF_buf1) );
  BUFX2 BUFX2_15 ( .A(clock), .Y(clock_bF_buf7) );
  BUFX2 BUFX2_150 ( .A(state_8_), .Y(state_8_bF_buf0) );
  BUFX2 BUFX2_151 ( .A(_abc_17692_n4047), .Y(_abc_17692_n4047_bF_buf4) );
  BUFX2 BUFX2_152 ( .A(_abc_17692_n4047), .Y(_abc_17692_n4047_bF_buf3) );
  BUFX2 BUFX2_153 ( .A(_abc_17692_n4047), .Y(_abc_17692_n4047_bF_buf2) );
  BUFX2 BUFX2_154 ( .A(_abc_17692_n4047), .Y(_abc_17692_n4047_bF_buf1) );
  BUFX2 BUFX2_155 ( .A(_abc_17692_n4047), .Y(_abc_17692_n4047_bF_buf0) );
  BUFX2 BUFX2_156 ( .A(workunit1_16_), .Y(workunit1_16_bF_buf3) );
  BUFX2 BUFX2_157 ( .A(workunit1_16_), .Y(workunit1_16_bF_buf2) );
  BUFX2 BUFX2_158 ( .A(workunit1_16_), .Y(workunit1_16_bF_buf1) );
  BUFX2 BUFX2_159 ( .A(workunit1_16_), .Y(workunit1_16_bF_buf0) );
  BUFX2 BUFX2_16 ( .A(clock), .Y(clock_bF_buf6) );
  BUFX2 BUFX2_160 ( .A(_abc_17692_n1863), .Y(_abc_17692_n1863_bF_buf10) );
  BUFX2 BUFX2_161 ( .A(_abc_17692_n1863), .Y(_abc_17692_n1863_bF_buf9) );
  BUFX2 BUFX2_162 ( .A(_abc_17692_n1863), .Y(_abc_17692_n1863_bF_buf8) );
  BUFX2 BUFX2_163 ( .A(_abc_17692_n1863), .Y(_abc_17692_n1863_bF_buf7) );
  BUFX2 BUFX2_164 ( .A(_abc_17692_n1863), .Y(_abc_17692_n1863_bF_buf6) );
  BUFX2 BUFX2_165 ( .A(_abc_17692_n1863), .Y(_abc_17692_n1863_bF_buf5) );
  BUFX2 BUFX2_166 ( .A(_abc_17692_n1863), .Y(_abc_17692_n1863_bF_buf4) );
  BUFX2 BUFX2_167 ( .A(_abc_17692_n1863), .Y(_abc_17692_n1863_bF_buf3) );
  BUFX2 BUFX2_168 ( .A(_abc_17692_n1863), .Y(_abc_17692_n1863_bF_buf2) );
  BUFX2 BUFX2_169 ( .A(_abc_17692_n1863), .Y(_abc_17692_n1863_bF_buf1) );
  BUFX2 BUFX2_17 ( .A(clock), .Y(clock_bF_buf5) );
  BUFX2 BUFX2_170 ( .A(_abc_17692_n1863), .Y(_abc_17692_n1863_bF_buf0) );
  BUFX2 BUFX2_171 ( .A(workunit1_13_), .Y(workunit1_13_bF_buf3) );
  BUFX2 BUFX2_172 ( .A(workunit1_13_), .Y(workunit1_13_bF_buf2) );
  BUFX2 BUFX2_173 ( .A(workunit1_13_), .Y(workunit1_13_bF_buf1) );
  BUFX2 BUFX2_174 ( .A(workunit1_13_), .Y(workunit1_13_bF_buf0) );
  BUFX2 BUFX2_175 ( .A(_abc_17692_n1830), .Y(_abc_17692_n1830_bF_buf10) );
  BUFX2 BUFX2_176 ( .A(_abc_17692_n1830), .Y(_abc_17692_n1830_bF_buf9) );
  BUFX2 BUFX2_177 ( .A(_abc_17692_n1830), .Y(_abc_17692_n1830_bF_buf8) );
  BUFX2 BUFX2_178 ( .A(_abc_17692_n1830), .Y(_abc_17692_n1830_bF_buf7) );
  BUFX2 BUFX2_179 ( .A(_abc_17692_n1830), .Y(_abc_17692_n1830_bF_buf6) );
  BUFX2 BUFX2_18 ( .A(clock), .Y(clock_bF_buf4) );
  BUFX2 BUFX2_180 ( .A(_abc_17692_n1830), .Y(_abc_17692_n1830_bF_buf5) );
  BUFX2 BUFX2_181 ( .A(_abc_17692_n1830), .Y(_abc_17692_n1830_bF_buf4) );
  BUFX2 BUFX2_182 ( .A(_abc_17692_n1830), .Y(_abc_17692_n1830_bF_buf3) );
  BUFX2 BUFX2_183 ( .A(_abc_17692_n1830), .Y(_abc_17692_n1830_bF_buf2) );
  BUFX2 BUFX2_184 ( .A(_abc_17692_n1830), .Y(_abc_17692_n1830_bF_buf1) );
  BUFX2 BUFX2_185 ( .A(_abc_17692_n1830), .Y(_abc_17692_n1830_bF_buf0) );
  BUFX2 BUFX2_186 ( .A(workunit2_1_), .Y(workunit2_1_bF_buf3) );
  BUFX2 BUFX2_187 ( .A(workunit2_1_), .Y(workunit2_1_bF_buf2) );
  BUFX2 BUFX2_188 ( .A(workunit2_1_), .Y(workunit2_1_bF_buf1) );
  BUFX2 BUFX2_189 ( .A(workunit2_1_), .Y(workunit2_1_bF_buf0) );
  BUFX2 BUFX2_19 ( .A(clock), .Y(clock_bF_buf3) );
  BUFX2 BUFX2_190 ( .A(_abc_17692_n8383), .Y(_abc_17692_n8383_bF_buf4) );
  BUFX2 BUFX2_191 ( .A(_abc_17692_n8383), .Y(_abc_17692_n8383_bF_buf3) );
  BUFX2 BUFX2_192 ( .A(_abc_17692_n8383), .Y(_abc_17692_n8383_bF_buf2) );
  BUFX2 BUFX2_193 ( .A(_abc_17692_n8383), .Y(_abc_17692_n8383_bF_buf1) );
  BUFX2 BUFX2_194 ( .A(_abc_17692_n8383), .Y(_abc_17692_n8383_bF_buf0) );
  BUFX2 BUFX2_195 ( .A(state_15_), .Y(state_15_bF_buf4) );
  BUFX2 BUFX2_196 ( .A(state_15_), .Y(state_15_bF_buf3) );
  BUFX2 BUFX2_197 ( .A(state_15_), .Y(state_15_bF_buf2) );
  BUFX2 BUFX2_198 ( .A(state_15_), .Y(state_15_bF_buf1) );
  BUFX2 BUFX2_199 ( .A(state_15_), .Y(state_15_bF_buf0) );
  BUFX2 BUFX2_2 ( .A(workunit2_12_), .Y(workunit2_12_bF_buf2) );
  BUFX2 BUFX2_20 ( .A(clock), .Y(clock_bF_buf2) );
  BUFX2 BUFX2_200 ( .A(1'b0), .Y(all_done) );
  BUFX2 BUFX2_201 ( .A(_auto_iopadmap_cc_313_execute_30032_0_), .Y(\data_out1[0] ) );
  BUFX2 BUFX2_202 ( .A(_auto_iopadmap_cc_313_execute_30032_1_), .Y(\data_out1[1] ) );
  BUFX2 BUFX2_203 ( .A(_auto_iopadmap_cc_313_execute_30032_2_), .Y(\data_out1[2] ) );
  BUFX2 BUFX2_204 ( .A(_auto_iopadmap_cc_313_execute_30032_3_), .Y(\data_out1[3] ) );
  BUFX2 BUFX2_205 ( .A(_auto_iopadmap_cc_313_execute_30032_4_), .Y(\data_out1[4] ) );
  BUFX2 BUFX2_206 ( .A(_auto_iopadmap_cc_313_execute_30032_5_), .Y(\data_out1[5] ) );
  BUFX2 BUFX2_207 ( .A(_auto_iopadmap_cc_313_execute_30032_6_), .Y(\data_out1[6] ) );
  BUFX2 BUFX2_208 ( .A(_auto_iopadmap_cc_313_execute_30032_7_), .Y(\data_out1[7] ) );
  BUFX2 BUFX2_209 ( .A(_auto_iopadmap_cc_313_execute_30032_8_), .Y(\data_out1[8] ) );
  BUFX2 BUFX2_21 ( .A(clock), .Y(clock_bF_buf1) );
  BUFX2 BUFX2_210 ( .A(_auto_iopadmap_cc_313_execute_30032_9_), .Y(\data_out1[9] ) );
  BUFX2 BUFX2_211 ( .A(_auto_iopadmap_cc_313_execute_30032_10_), .Y(\data_out1[10] ) );
  BUFX2 BUFX2_212 ( .A(_auto_iopadmap_cc_313_execute_30032_11_), .Y(\data_out1[11] ) );
  BUFX2 BUFX2_213 ( .A(_auto_iopadmap_cc_313_execute_30032_12_), .Y(\data_out1[12] ) );
  BUFX2 BUFX2_214 ( .A(_auto_iopadmap_cc_313_execute_30032_13_), .Y(\data_out1[13] ) );
  BUFX2 BUFX2_215 ( .A(_auto_iopadmap_cc_313_execute_30032_14_), .Y(\data_out1[14] ) );
  BUFX2 BUFX2_216 ( .A(_auto_iopadmap_cc_313_execute_30032_15_), .Y(\data_out1[15] ) );
  BUFX2 BUFX2_217 ( .A(_auto_iopadmap_cc_313_execute_30032_16_), .Y(\data_out1[16] ) );
  BUFX2 BUFX2_218 ( .A(_auto_iopadmap_cc_313_execute_30032_17_), .Y(\data_out1[17] ) );
  BUFX2 BUFX2_219 ( .A(_auto_iopadmap_cc_313_execute_30032_18_), .Y(\data_out1[18] ) );
  BUFX2 BUFX2_22 ( .A(clock), .Y(clock_bF_buf0) );
  BUFX2 BUFX2_220 ( .A(_auto_iopadmap_cc_313_execute_30032_19_), .Y(\data_out1[19] ) );
  BUFX2 BUFX2_221 ( .A(_auto_iopadmap_cc_313_execute_30032_20_), .Y(\data_out1[20] ) );
  BUFX2 BUFX2_222 ( .A(_auto_iopadmap_cc_313_execute_30032_21_), .Y(\data_out1[21] ) );
  BUFX2 BUFX2_223 ( .A(_auto_iopadmap_cc_313_execute_30032_22_), .Y(\data_out1[22] ) );
  BUFX2 BUFX2_224 ( .A(_auto_iopadmap_cc_313_execute_30032_23_), .Y(\data_out1[23] ) );
  BUFX2 BUFX2_225 ( .A(_auto_iopadmap_cc_313_execute_30032_24_), .Y(\data_out1[24] ) );
  BUFX2 BUFX2_226 ( .A(_auto_iopadmap_cc_313_execute_30032_25_), .Y(\data_out1[25] ) );
  BUFX2 BUFX2_227 ( .A(_auto_iopadmap_cc_313_execute_30032_26_), .Y(\data_out1[26] ) );
  BUFX2 BUFX2_228 ( .A(_auto_iopadmap_cc_313_execute_30032_27_), .Y(\data_out1[27] ) );
  BUFX2 BUFX2_229 ( .A(_auto_iopadmap_cc_313_execute_30032_28_), .Y(\data_out1[28] ) );
  BUFX2 BUFX2_23 ( .A(state_7_), .Y(state_7_bF_buf4) );
  BUFX2 BUFX2_230 ( .A(_auto_iopadmap_cc_313_execute_30032_29_), .Y(\data_out1[29] ) );
  BUFX2 BUFX2_231 ( .A(_auto_iopadmap_cc_313_execute_30032_30_), .Y(\data_out1[30] ) );
  BUFX2 BUFX2_232 ( .A(_auto_iopadmap_cc_313_execute_30032_31_), .Y(\data_out1[31] ) );
  BUFX2 BUFX2_233 ( .A(_auto_iopadmap_cc_313_execute_30065_0_), .Y(\data_out2[0] ) );
  BUFX2 BUFX2_234 ( .A(_auto_iopadmap_cc_313_execute_30065_1_), .Y(\data_out2[1] ) );
  BUFX2 BUFX2_235 ( .A(_auto_iopadmap_cc_313_execute_30065_2_), .Y(\data_out2[2] ) );
  BUFX2 BUFX2_236 ( .A(_auto_iopadmap_cc_313_execute_30065_3_), .Y(\data_out2[3] ) );
  BUFX2 BUFX2_237 ( .A(_auto_iopadmap_cc_313_execute_30065_4_), .Y(\data_out2[4] ) );
  BUFX2 BUFX2_238 ( .A(_auto_iopadmap_cc_313_execute_30065_5_), .Y(\data_out2[5] ) );
  BUFX2 BUFX2_239 ( .A(_auto_iopadmap_cc_313_execute_30065_6_), .Y(\data_out2[6] ) );
  BUFX2 BUFX2_24 ( .A(state_7_), .Y(state_7_bF_buf3) );
  BUFX2 BUFX2_240 ( .A(_auto_iopadmap_cc_313_execute_30065_7_), .Y(\data_out2[7] ) );
  BUFX2 BUFX2_241 ( .A(_auto_iopadmap_cc_313_execute_30065_8_), .Y(\data_out2[8] ) );
  BUFX2 BUFX2_242 ( .A(_auto_iopadmap_cc_313_execute_30065_9_), .Y(\data_out2[9] ) );
  BUFX2 BUFX2_243 ( .A(_auto_iopadmap_cc_313_execute_30065_10_), .Y(\data_out2[10] ) );
  BUFX2 BUFX2_244 ( .A(_auto_iopadmap_cc_313_execute_30065_11_), .Y(\data_out2[11] ) );
  BUFX2 BUFX2_245 ( .A(_auto_iopadmap_cc_313_execute_30065_12_), .Y(\data_out2[12] ) );
  BUFX2 BUFX2_246 ( .A(_auto_iopadmap_cc_313_execute_30065_13_), .Y(\data_out2[13] ) );
  BUFX2 BUFX2_247 ( .A(_auto_iopadmap_cc_313_execute_30065_14_), .Y(\data_out2[14] ) );
  BUFX2 BUFX2_248 ( .A(_auto_iopadmap_cc_313_execute_30065_15_), .Y(\data_out2[15] ) );
  BUFX2 BUFX2_249 ( .A(_auto_iopadmap_cc_313_execute_30065_16_), .Y(\data_out2[16] ) );
  BUFX2 BUFX2_25 ( .A(state_7_), .Y(state_7_bF_buf2) );
  BUFX2 BUFX2_250 ( .A(_auto_iopadmap_cc_313_execute_30065_17_), .Y(\data_out2[17] ) );
  BUFX2 BUFX2_251 ( .A(_auto_iopadmap_cc_313_execute_30065_18_), .Y(\data_out2[18] ) );
  BUFX2 BUFX2_252 ( .A(_auto_iopadmap_cc_313_execute_30065_19_), .Y(\data_out2[19] ) );
  BUFX2 BUFX2_253 ( .A(_auto_iopadmap_cc_313_execute_30065_20_), .Y(\data_out2[20] ) );
  BUFX2 BUFX2_254 ( .A(_auto_iopadmap_cc_313_execute_30065_21_), .Y(\data_out2[21] ) );
  BUFX2 BUFX2_255 ( .A(_auto_iopadmap_cc_313_execute_30065_22_), .Y(\data_out2[22] ) );
  BUFX2 BUFX2_256 ( .A(_auto_iopadmap_cc_313_execute_30065_23_), .Y(\data_out2[23] ) );
  BUFX2 BUFX2_257 ( .A(_auto_iopadmap_cc_313_execute_30065_24_), .Y(\data_out2[24] ) );
  BUFX2 BUFX2_258 ( .A(_auto_iopadmap_cc_313_execute_30065_25_), .Y(\data_out2[25] ) );
  BUFX2 BUFX2_259 ( .A(_auto_iopadmap_cc_313_execute_30065_26_), .Y(\data_out2[26] ) );
  BUFX2 BUFX2_26 ( .A(state_7_), .Y(state_7_bF_buf1) );
  BUFX2 BUFX2_260 ( .A(_auto_iopadmap_cc_313_execute_30065_27_), .Y(\data_out2[27] ) );
  BUFX2 BUFX2_261 ( .A(_auto_iopadmap_cc_313_execute_30065_28_), .Y(\data_out2[28] ) );
  BUFX2 BUFX2_262 ( .A(_auto_iopadmap_cc_313_execute_30065_29_), .Y(\data_out2[29] ) );
  BUFX2 BUFX2_263 ( .A(_auto_iopadmap_cc_313_execute_30065_30_), .Y(\data_out2[30] ) );
  BUFX2 BUFX2_264 ( .A(_auto_iopadmap_cc_313_execute_30065_31_), .Y(\data_out2[31] ) );
  BUFX2 BUFX2_27 ( .A(state_7_), .Y(state_7_bF_buf0) );
  BUFX2 BUFX2_28 ( .A(_abc_17692_n1885), .Y(_abc_17692_n1885_bF_buf4) );
  BUFX2 BUFX2_29 ( .A(_abc_17692_n1885), .Y(_abc_17692_n1885_bF_buf3) );
  BUFX2 BUFX2_3 ( .A(workunit2_12_), .Y(workunit2_12_bF_buf1) );
  BUFX2 BUFX2_30 ( .A(_abc_17692_n1885), .Y(_abc_17692_n1885_bF_buf2) );
  BUFX2 BUFX2_31 ( .A(_abc_17692_n1885), .Y(_abc_17692_n1885_bF_buf1) );
  BUFX2 BUFX2_32 ( .A(_abc_17692_n1885), .Y(_abc_17692_n1885_bF_buf0) );
  BUFX2 BUFX2_33 ( .A(workunit1_12_), .Y(workunit1_12_bF_buf3) );
  BUFX2 BUFX2_34 ( .A(workunit1_12_), .Y(workunit1_12_bF_buf2) );
  BUFX2 BUFX2_35 ( .A(workunit1_12_), .Y(workunit1_12_bF_buf1) );
  BUFX2 BUFX2_36 ( .A(workunit1_12_), .Y(workunit1_12_bF_buf0) );
  BUFX2 BUFX2_37 ( .A(_abc_17692_n722), .Y(_abc_17692_n722_bF_buf3) );
  BUFX2 BUFX2_38 ( .A(_abc_17692_n722), .Y(_abc_17692_n722_bF_buf2) );
  BUFX2 BUFX2_39 ( .A(_abc_17692_n722), .Y(_abc_17692_n722_bF_buf1) );
  BUFX2 BUFX2_4 ( .A(workunit2_12_), .Y(workunit2_12_bF_buf0) );
  BUFX2 BUFX2_40 ( .A(_abc_17692_n722), .Y(_abc_17692_n722_bF_buf0) );
  BUFX2 BUFX2_41 ( .A(_abc_17692_n725), .Y(_abc_17692_n725_bF_buf7) );
  BUFX2 BUFX2_42 ( .A(_abc_17692_n725), .Y(_abc_17692_n725_bF_buf6) );
  BUFX2 BUFX2_43 ( .A(_abc_17692_n725), .Y(_abc_17692_n725_bF_buf5) );
  BUFX2 BUFX2_44 ( .A(_abc_17692_n725), .Y(_abc_17692_n725_bF_buf4) );
  BUFX2 BUFX2_45 ( .A(_abc_17692_n725), .Y(_abc_17692_n725_bF_buf3) );
  BUFX2 BUFX2_46 ( .A(_abc_17692_n725), .Y(_abc_17692_n725_bF_buf2) );
  BUFX2 BUFX2_47 ( .A(_abc_17692_n725), .Y(_abc_17692_n725_bF_buf1) );
  BUFX2 BUFX2_48 ( .A(_abc_17692_n725), .Y(_abc_17692_n725_bF_buf0) );
  BUFX2 BUFX2_49 ( .A(_abc_17692_n727), .Y(_abc_17692_n727_bF_buf7) );
  BUFX2 BUFX2_5 ( .A(workunit1_1_), .Y(workunit1_1_bF_buf3) );
  BUFX2 BUFX2_50 ( .A(_abc_17692_n727), .Y(_abc_17692_n727_bF_buf6) );
  BUFX2 BUFX2_51 ( .A(_abc_17692_n727), .Y(_abc_17692_n727_bF_buf5) );
  BUFX2 BUFX2_52 ( .A(_abc_17692_n727), .Y(_abc_17692_n727_bF_buf4) );
  BUFX2 BUFX2_53 ( .A(_abc_17692_n727), .Y(_abc_17692_n727_bF_buf3) );
  BUFX2 BUFX2_54 ( .A(_abc_17692_n727), .Y(_abc_17692_n727_bF_buf2) );
  BUFX2 BUFX2_55 ( .A(_abc_17692_n727), .Y(_abc_17692_n727_bF_buf1) );
  BUFX2 BUFX2_56 ( .A(_abc_17692_n727), .Y(_abc_17692_n727_bF_buf0) );
  BUFX2 BUFX2_57 ( .A(workunit2_14_), .Y(workunit2_14_bF_buf3) );
  BUFX2 BUFX2_58 ( .A(workunit2_14_), .Y(workunit2_14_bF_buf2) );
  BUFX2 BUFX2_59 ( .A(workunit2_14_), .Y(workunit2_14_bF_buf1) );
  BUFX2 BUFX2_6 ( .A(workunit1_1_), .Y(workunit1_1_bF_buf2) );
  BUFX2 BUFX2_60 ( .A(workunit2_14_), .Y(workunit2_14_bF_buf0) );
  BUFX2 BUFX2_61 ( .A(state_14_), .Y(state_14_bF_buf4) );
  BUFX2 BUFX2_62 ( .A(state_14_), .Y(state_14_bF_buf3) );
  BUFX2 BUFX2_63 ( .A(state_14_), .Y(state_14_bF_buf2) );
  BUFX2 BUFX2_64 ( .A(state_14_), .Y(state_14_bF_buf1) );
  BUFX2 BUFX2_65 ( .A(state_14_), .Y(state_14_bF_buf0) );
  BUFX2 BUFX2_66 ( .A(state_6_), .Y(state_6_bF_buf4) );
  BUFX2 BUFX2_67 ( .A(state_6_), .Y(state_6_bF_buf3) );
  BUFX2 BUFX2_68 ( .A(state_6_), .Y(state_6_bF_buf2) );
  BUFX2 BUFX2_69 ( .A(state_6_), .Y(state_6_bF_buf1) );
  BUFX2 BUFX2_7 ( .A(workunit1_1_), .Y(workunit1_1_bF_buf1) );
  BUFX2 BUFX2_70 ( .A(state_6_), .Y(state_6_bF_buf0) );
  BUFX2 BUFX2_71 ( .A(_abc_17692_n6660), .Y(_abc_17692_n6660_bF_buf13) );
  BUFX2 BUFX2_72 ( .A(_abc_17692_n6660), .Y(_abc_17692_n6660_bF_buf12) );
  BUFX2 BUFX2_73 ( .A(_abc_17692_n6660), .Y(_abc_17692_n6660_bF_buf11) );
  BUFX2 BUFX2_74 ( .A(_abc_17692_n6660), .Y(_abc_17692_n6660_bF_buf10) );
  BUFX2 BUFX2_75 ( .A(_abc_17692_n6660), .Y(_abc_17692_n6660_bF_buf9) );
  BUFX2 BUFX2_76 ( .A(_abc_17692_n6660), .Y(_abc_17692_n6660_bF_buf8) );
  BUFX2 BUFX2_77 ( .A(_abc_17692_n6660), .Y(_abc_17692_n6660_bF_buf7) );
  BUFX2 BUFX2_78 ( .A(_abc_17692_n6660), .Y(_abc_17692_n6660_bF_buf6) );
  BUFX2 BUFX2_79 ( .A(_abc_17692_n6660), .Y(_abc_17692_n6660_bF_buf5) );
  BUFX2 BUFX2_8 ( .A(workunit1_1_), .Y(workunit1_1_bF_buf0) );
  BUFX2 BUFX2_80 ( .A(_abc_17692_n6660), .Y(_abc_17692_n6660_bF_buf4) );
  BUFX2 BUFX2_81 ( .A(_abc_17692_n6660), .Y(_abc_17692_n6660_bF_buf3) );
  BUFX2 BUFX2_82 ( .A(_abc_17692_n6660), .Y(_abc_17692_n6660_bF_buf2) );
  BUFX2 BUFX2_83 ( .A(_abc_17692_n6660), .Y(_abc_17692_n6660_bF_buf1) );
  BUFX2 BUFX2_84 ( .A(_abc_17692_n6660), .Y(_abc_17692_n6660_bF_buf0) );
  BUFX2 BUFX2_85 ( .A(state_3_), .Y(state_3_bF_buf4) );
  BUFX2 BUFX2_86 ( .A(state_3_), .Y(state_3_bF_buf3) );
  BUFX2 BUFX2_87 ( .A(state_3_), .Y(state_3_bF_buf2) );
  BUFX2 BUFX2_88 ( .A(state_3_), .Y(state_3_bF_buf1) );
  BUFX2 BUFX2_89 ( .A(state_3_), .Y(state_3_bF_buf0) );
  BUFX2 BUFX2_9 ( .A(clock), .Y(clock_bF_buf13) );
  BUFX2 BUFX2_90 ( .A(_abc_17692_n1877), .Y(_abc_17692_n1877_bF_buf10) );
  BUFX2 BUFX2_91 ( .A(_abc_17692_n1877), .Y(_abc_17692_n1877_bF_buf9) );
  BUFX2 BUFX2_92 ( .A(_abc_17692_n1877), .Y(_abc_17692_n1877_bF_buf8) );
  BUFX2 BUFX2_93 ( .A(_abc_17692_n1877), .Y(_abc_17692_n1877_bF_buf7) );
  BUFX2 BUFX2_94 ( .A(_abc_17692_n1877), .Y(_abc_17692_n1877_bF_buf6) );
  BUFX2 BUFX2_95 ( .A(_abc_17692_n1877), .Y(_abc_17692_n1877_bF_buf5) );
  BUFX2 BUFX2_96 ( .A(_abc_17692_n1877), .Y(_abc_17692_n1877_bF_buf4) );
  BUFX2 BUFX2_97 ( .A(_abc_17692_n1877), .Y(_abc_17692_n1877_bF_buf3) );
  BUFX2 BUFX2_98 ( .A(_abc_17692_n1877), .Y(_abc_17692_n1877_bF_buf2) );
  BUFX2 BUFX2_99 ( .A(_abc_17692_n1877), .Y(_abc_17692_n1877_bF_buf1) );
  DFFSR DFFSR_1 ( .CLK(clock_bF_buf13), .D(data_out1_0__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30032_0_), .R(_abc_17692_n6660_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_10 ( .CLK(clock_bF_buf4), .D(data_out1_9__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30032_9_), .R(_abc_17692_n6660_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_100 ( .CLK(clock_bF_buf12), .D(sum_23__FF_INPUT), .Q(sum_23_), .R(_abc_17692_n6660_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_101 ( .CLK(clock_bF_buf11), .D(sum_24__FF_INPUT), .Q(sum_24_), .R(_abc_17692_n6660_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_102 ( .CLK(clock_bF_buf10), .D(sum_25__FF_INPUT), .Q(sum_25_), .R(_abc_17692_n6660_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_103 ( .CLK(clock_bF_buf9), .D(sum_26__FF_INPUT), .Q(sum_26_), .R(_abc_17692_n6660_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_104 ( .CLK(clock_bF_buf8), .D(sum_27__FF_INPUT), .Q(sum_27_), .R(_abc_17692_n6660_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_105 ( .CLK(clock_bF_buf7), .D(sum_28__FF_INPUT), .Q(sum_28_), .R(_abc_17692_n6660_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_106 ( .CLK(clock_bF_buf6), .D(sum_29__FF_INPUT), .Q(sum_29_), .R(_abc_17692_n6660_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_107 ( .CLK(clock_bF_buf5), .D(sum_30__FF_INPUT), .Q(sum_30_), .R(_abc_17692_n6660_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_108 ( .CLK(clock_bF_buf4), .D(sum_31__FF_INPUT), .Q(sum_31_), .R(_abc_17692_n6660_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_109 ( .CLK(clock_bF_buf3), .D(workunit1_0__FF_INPUT), .Q(workunit1_0_), .R(_abc_17692_n6660_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_11 ( .CLK(clock_bF_buf3), .D(data_out1_10__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30032_10_), .R(_abc_17692_n6660_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_110 ( .CLK(clock_bF_buf2), .D(workunit1_1__FF_INPUT), .Q(workunit1_1_), .R(_abc_17692_n6660_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_111 ( .CLK(clock_bF_buf1), .D(workunit1_2__FF_INPUT), .Q(workunit1_2_), .R(_abc_17692_n6660_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_112 ( .CLK(clock_bF_buf0), .D(workunit1_3__FF_INPUT), .Q(workunit1_3_), .R(_abc_17692_n6660_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_113 ( .CLK(clock_bF_buf13), .D(workunit1_4__FF_INPUT), .Q(workunit1_4_), .R(_abc_17692_n6660_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_114 ( .CLK(clock_bF_buf12), .D(workunit1_5__FF_INPUT), .Q(workunit1_5_), .R(_abc_17692_n6660_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_115 ( .CLK(clock_bF_buf11), .D(workunit1_6__FF_INPUT), .Q(workunit1_6_), .R(_abc_17692_n6660_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_116 ( .CLK(clock_bF_buf10), .D(workunit1_7__FF_INPUT), .Q(workunit1_7_), .R(_abc_17692_n6660_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_117 ( .CLK(clock_bF_buf9), .D(workunit1_8__FF_INPUT), .Q(workunit1_8_), .R(_abc_17692_n6660_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_118 ( .CLK(clock_bF_buf8), .D(workunit1_9__FF_INPUT), .Q(workunit1_9_), .R(_abc_17692_n6660_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_119 ( .CLK(clock_bF_buf7), .D(workunit1_10__FF_INPUT), .Q(workunit1_10_), .R(_abc_17692_n6660_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_12 ( .CLK(clock_bF_buf2), .D(data_out1_11__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30032_11_), .R(_abc_17692_n6660_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_120 ( .CLK(clock_bF_buf6), .D(workunit1_11__FF_INPUT), .Q(workunit1_11_), .R(_abc_17692_n6660_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_121 ( .CLK(clock_bF_buf5), .D(workunit1_12__FF_INPUT), .Q(workunit1_12_), .R(_abc_17692_n6660_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_122 ( .CLK(clock_bF_buf4), .D(workunit1_13__FF_INPUT), .Q(workunit1_13_), .R(_abc_17692_n6660_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_123 ( .CLK(clock_bF_buf3), .D(workunit1_14__FF_INPUT), .Q(workunit1_14_), .R(_abc_17692_n6660_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_124 ( .CLK(clock_bF_buf2), .D(workunit1_15__FF_INPUT), .Q(workunit1_15_), .R(_abc_17692_n6660_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_125 ( .CLK(clock_bF_buf1), .D(workunit1_16__FF_INPUT), .Q(workunit1_16_), .R(_abc_17692_n6660_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_126 ( .CLK(clock_bF_buf0), .D(workunit1_17__FF_INPUT), .Q(workunit1_17_), .R(_abc_17692_n6660_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_127 ( .CLK(clock_bF_buf13), .D(workunit1_18__FF_INPUT), .Q(workunit1_18_), .R(_abc_17692_n6660_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_128 ( .CLK(clock_bF_buf12), .D(workunit1_19__FF_INPUT), .Q(workunit1_19_), .R(_abc_17692_n6660_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_129 ( .CLK(clock_bF_buf11), .D(workunit1_20__FF_INPUT), .Q(workunit1_20_), .R(_abc_17692_n6660_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_13 ( .CLK(clock_bF_buf1), .D(data_out1_12__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30032_12_), .R(_abc_17692_n6660_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_130 ( .CLK(clock_bF_buf10), .D(workunit1_21__FF_INPUT), .Q(workunit1_21_), .R(_abc_17692_n6660_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_131 ( .CLK(clock_bF_buf9), .D(workunit1_22__FF_INPUT), .Q(workunit1_22_), .R(_abc_17692_n6660_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_132 ( .CLK(clock_bF_buf8), .D(workunit1_23__FF_INPUT), .Q(workunit1_23_), .R(_abc_17692_n6660_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_133 ( .CLK(clock_bF_buf7), .D(workunit1_24__FF_INPUT), .Q(workunit1_24_), .R(_abc_17692_n6660_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_134 ( .CLK(clock_bF_buf6), .D(workunit1_25__FF_INPUT), .Q(workunit1_25_), .R(_abc_17692_n6660_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_135 ( .CLK(clock_bF_buf5), .D(workunit1_26__FF_INPUT), .Q(workunit1_26_), .R(_abc_17692_n6660_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_136 ( .CLK(clock_bF_buf4), .D(workunit1_27__FF_INPUT), .Q(workunit1_27_), .R(_abc_17692_n6660_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_137 ( .CLK(clock_bF_buf3), .D(workunit1_28__FF_INPUT), .Q(workunit1_28_), .R(_abc_17692_n6660_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_138 ( .CLK(clock_bF_buf2), .D(workunit1_29__FF_INPUT), .Q(workunit1_29_), .R(_abc_17692_n6660_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_139 ( .CLK(clock_bF_buf1), .D(workunit1_30__FF_INPUT), .Q(workunit1_30_), .R(_abc_17692_n6660_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_14 ( .CLK(clock_bF_buf0), .D(data_out1_13__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30032_13_), .R(_abc_17692_n6660_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_140 ( .CLK(clock_bF_buf0), .D(workunit1_31__FF_INPUT), .Q(workunit1_31_), .R(_abc_17692_n6660_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_141 ( .CLK(clock_bF_buf13), .D(workunit2_0__FF_INPUT), .Q(workunit2_0_), .R(_abc_17692_n6660_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_142 ( .CLK(clock_bF_buf12), .D(workunit2_1__FF_INPUT), .Q(workunit2_1_), .R(_abc_17692_n6660_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_143 ( .CLK(clock_bF_buf11), .D(workunit2_2__FF_INPUT), .Q(workunit2_2_), .R(_abc_17692_n6660_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_144 ( .CLK(clock_bF_buf10), .D(workunit2_3__FF_INPUT), .Q(workunit2_3_), .R(_abc_17692_n6660_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_145 ( .CLK(clock_bF_buf9), .D(workunit2_4__FF_INPUT), .Q(workunit2_4_), .R(_abc_17692_n6660_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_146 ( .CLK(clock_bF_buf8), .D(workunit2_5__FF_INPUT), .Q(workunit2_5_), .R(_abc_17692_n6660_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_147 ( .CLK(clock_bF_buf7), .D(workunit2_6__FF_INPUT), .Q(workunit2_6_), .R(_abc_17692_n6660_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_148 ( .CLK(clock_bF_buf6), .D(workunit2_7__FF_INPUT), .Q(workunit2_7_), .R(_abc_17692_n6660_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_149 ( .CLK(clock_bF_buf5), .D(workunit2_8__FF_INPUT), .Q(workunit2_8_), .R(_abc_17692_n6660_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_15 ( .CLK(clock_bF_buf13), .D(data_out1_14__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30032_14_), .R(_abc_17692_n6660_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_150 ( .CLK(clock_bF_buf4), .D(workunit2_9__FF_INPUT), .Q(workunit2_9_), .R(_abc_17692_n6660_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_151 ( .CLK(clock_bF_buf3), .D(workunit2_10__FF_INPUT), .Q(workunit2_10_), .R(_abc_17692_n6660_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_152 ( .CLK(clock_bF_buf2), .D(workunit2_11__FF_INPUT), .Q(workunit2_11_), .R(_abc_17692_n6660_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_153 ( .CLK(clock_bF_buf1), .D(workunit2_12__FF_INPUT), .Q(workunit2_12_), .R(_abc_17692_n6660_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_154 ( .CLK(clock_bF_buf0), .D(workunit2_13__FF_INPUT), .Q(workunit2_13_), .R(_abc_17692_n6660_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_155 ( .CLK(clock_bF_buf13), .D(workunit2_14__FF_INPUT), .Q(workunit2_14_), .R(_abc_17692_n6660_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_156 ( .CLK(clock_bF_buf12), .D(workunit2_15__FF_INPUT), .Q(workunit2_15_), .R(_abc_17692_n6660_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_157 ( .CLK(clock_bF_buf11), .D(workunit2_16__FF_INPUT), .Q(workunit2_16_), .R(_abc_17692_n6660_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_158 ( .CLK(clock_bF_buf10), .D(workunit2_17__FF_INPUT), .Q(workunit2_17_), .R(_abc_17692_n6660_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_159 ( .CLK(clock_bF_buf9), .D(workunit2_18__FF_INPUT), .Q(workunit2_18_), .R(_abc_17692_n6660_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_16 ( .CLK(clock_bF_buf12), .D(data_out1_15__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30032_15_), .R(_abc_17692_n6660_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_160 ( .CLK(clock_bF_buf8), .D(workunit2_19__FF_INPUT), .Q(workunit2_19_), .R(_abc_17692_n6660_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_161 ( .CLK(clock_bF_buf7), .D(workunit2_20__FF_INPUT), .Q(workunit2_20_), .R(_abc_17692_n6660_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_162 ( .CLK(clock_bF_buf6), .D(workunit2_21__FF_INPUT), .Q(workunit2_21_), .R(_abc_17692_n6660_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_163 ( .CLK(clock_bF_buf5), .D(workunit2_22__FF_INPUT), .Q(workunit2_22_), .R(_abc_17692_n6660_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_164 ( .CLK(clock_bF_buf4), .D(workunit2_23__FF_INPUT), .Q(workunit2_23_), .R(_abc_17692_n6660_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_165 ( .CLK(clock_bF_buf3), .D(workunit2_24__FF_INPUT), .Q(workunit2_24_), .R(_abc_17692_n6660_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_166 ( .CLK(clock_bF_buf2), .D(workunit2_25__FF_INPUT), .Q(workunit2_25_), .R(_abc_17692_n6660_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_167 ( .CLK(clock_bF_buf1), .D(workunit2_26__FF_INPUT), .Q(workunit2_26_), .R(_abc_17692_n6660_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_168 ( .CLK(clock_bF_buf0), .D(workunit2_27__FF_INPUT), .Q(workunit2_27_), .R(_abc_17692_n6660_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_169 ( .CLK(clock_bF_buf13), .D(workunit2_28__FF_INPUT), .Q(workunit2_28_), .R(_abc_17692_n6660_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_17 ( .CLK(clock_bF_buf11), .D(data_out1_16__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30032_16_), .R(_abc_17692_n6660_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_170 ( .CLK(clock_bF_buf12), .D(workunit2_29__FF_INPUT), .Q(workunit2_29_), .R(_abc_17692_n6660_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_171 ( .CLK(clock_bF_buf11), .D(workunit2_30__FF_INPUT), .Q(workunit2_30_), .R(_abc_17692_n6660_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_172 ( .CLK(clock_bF_buf10), .D(workunit2_31__FF_INPUT), .Q(workunit2_31_), .R(_abc_17692_n6660_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_173 ( .CLK(clock_bF_buf9), .D(delta_0__FF_INPUT), .Q(delta_0_), .R(_abc_17692_n6660_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_174 ( .CLK(clock_bF_buf8), .D(delta_1__FF_INPUT), .Q(delta_1_), .R(_abc_17692_n6660_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_175 ( .CLK(clock_bF_buf7), .D(delta_2__FF_INPUT), .Q(delta_2_), .R(_abc_17692_n6660_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_176 ( .CLK(clock_bF_buf6), .D(delta_3__FF_INPUT), .Q(delta_3_), .R(_abc_17692_n6660_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_177 ( .CLK(clock_bF_buf5), .D(delta_4__FF_INPUT), .Q(delta_4_), .R(_abc_17692_n6660_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_178 ( .CLK(clock_bF_buf4), .D(delta_5__FF_INPUT), .Q(delta_5_), .R(_abc_17692_n6660_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_179 ( .CLK(clock_bF_buf3), .D(delta_6__FF_INPUT), .Q(delta_6_), .R(_abc_17692_n6660_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_18 ( .CLK(clock_bF_buf10), .D(data_out1_17__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30032_17_), .R(_abc_17692_n6660_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_180 ( .CLK(clock_bF_buf2), .D(delta_7__FF_INPUT), .Q(delta_7_), .R(_abc_17692_n6660_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_181 ( .CLK(clock_bF_buf1), .D(delta_8__FF_INPUT), .Q(delta_8_), .R(_abc_17692_n6660_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_182 ( .CLK(clock_bF_buf0), .D(delta_9__FF_INPUT), .Q(delta_9_), .R(_abc_17692_n6660_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_183 ( .CLK(clock_bF_buf13), .D(delta_10__FF_INPUT), .Q(delta_10_), .R(_abc_17692_n6660_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_184 ( .CLK(clock_bF_buf12), .D(delta_11__FF_INPUT), .Q(delta_11_), .R(_abc_17692_n6660_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_185 ( .CLK(clock_bF_buf11), .D(delta_12__FF_INPUT), .Q(delta_12_), .R(_abc_17692_n6660_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_186 ( .CLK(clock_bF_buf10), .D(delta_13__FF_INPUT), .Q(delta_13_), .R(_abc_17692_n6660_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_187 ( .CLK(clock_bF_buf9), .D(delta_14__FF_INPUT), .Q(delta_14_), .R(_abc_17692_n6660_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_188 ( .CLK(clock_bF_buf8), .D(delta_15__FF_INPUT), .Q(delta_15_), .R(_abc_17692_n6660_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_189 ( .CLK(clock_bF_buf7), .D(delta_16__FF_INPUT), .Q(delta_16_), .R(_abc_17692_n6660_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_19 ( .CLK(clock_bF_buf9), .D(data_out1_18__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30032_18_), .R(_abc_17692_n6660_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_190 ( .CLK(clock_bF_buf6), .D(delta_17__FF_INPUT), .Q(delta_17_), .R(_abc_17692_n6660_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_191 ( .CLK(clock_bF_buf5), .D(delta_18__FF_INPUT), .Q(delta_18_), .R(_abc_17692_n6660_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_192 ( .CLK(clock_bF_buf4), .D(delta_19__FF_INPUT), .Q(delta_19_), .R(_abc_17692_n6660_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_193 ( .CLK(clock_bF_buf3), .D(delta_20__FF_INPUT), .Q(delta_20_), .R(_abc_17692_n6660_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_194 ( .CLK(clock_bF_buf2), .D(delta_21__FF_INPUT), .Q(delta_21_), .R(_abc_17692_n6660_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_195 ( .CLK(clock_bF_buf1), .D(delta_22__FF_INPUT), .Q(delta_22_), .R(_abc_17692_n6660_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_196 ( .CLK(clock_bF_buf0), .D(delta_23__FF_INPUT), .Q(delta_23_), .R(_abc_17692_n6660_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_197 ( .CLK(clock_bF_buf13), .D(delta_24__FF_INPUT), .Q(delta_24_), .R(_abc_17692_n6660_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_198 ( .CLK(clock_bF_buf12), .D(delta_25__FF_INPUT), .Q(delta_25_), .R(_abc_17692_n6660_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_199 ( .CLK(clock_bF_buf11), .D(delta_26__FF_INPUT), .Q(delta_26_), .R(_abc_17692_n6660_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_2 ( .CLK(clock_bF_buf12), .D(data_out1_1__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30032_1_), .R(_abc_17692_n6660_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_20 ( .CLK(clock_bF_buf8), .D(data_out1_19__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30032_19_), .R(_abc_17692_n6660_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_200 ( .CLK(clock_bF_buf10), .D(delta_27__FF_INPUT), .Q(delta_27_), .R(_abc_17692_n6660_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_201 ( .CLK(clock_bF_buf9), .D(delta_28__FF_INPUT), .Q(delta_28_), .R(_abc_17692_n6660_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_202 ( .CLK(clock_bF_buf8), .D(delta_29__FF_INPUT), .Q(delta_29_), .R(_abc_17692_n6660_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_203 ( .CLK(clock_bF_buf7), .D(delta_30__FF_INPUT), .Q(delta_30_), .R(_abc_17692_n6660_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_204 ( .CLK(clock_bF_buf6), .D(delta_31__FF_INPUT), .Q(delta_31_), .R(_abc_17692_n6660_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_205 ( .CLK(clock_bF_buf5), .D(1'b0), .Q(state_0_), .R(1'b1), .S(_abc_17692_n6660_bF_buf5) );
  DFFSR DFFSR_206 ( .CLK(clock_bF_buf4), .D(state_15_bF_buf2), .Q(state_1_), .R(_abc_17692_n6660_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_207 ( .CLK(clock_bF_buf3), .D(_abc_10892_n7323), .Q(state_2_), .R(_abc_17692_n6660_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_208 ( .CLK(clock_bF_buf2), .D(state_14_bF_buf3), .Q(state_3_), .R(_abc_17692_n6660_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_209 ( .CLK(clock_bF_buf1), .D(_abc_10892_n1125), .Q(state_4_), .R(_abc_17692_n6660_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_21 ( .CLK(clock_bF_buf7), .D(data_out1_20__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30032_20_), .R(_abc_17692_n6660_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_210 ( .CLK(clock_bF_buf0), .D(_abc_10892_n7419), .Q(state_5_), .R(_abc_17692_n6660_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_211 ( .CLK(clock_bF_buf13), .D(state_11_), .Q(state_6_), .R(_abc_17692_n6660_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_212 ( .CLK(clock_bF_buf12), .D(_abc_10892_n1037), .Q(state_7_), .R(_abc_17692_n6660_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_213 ( .CLK(clock_bF_buf11), .D(state_0_), .Q(state_8_), .R(_abc_17692_n6660_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_214 ( .CLK(clock_bF_buf10), .D(state_1_), .Q(state_10_), .R(_abc_17692_n6660_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_215 ( .CLK(clock_bF_buf9), .D(_abc_10892_n6074), .Q(state_11_), .R(_abc_17692_n6660_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_216 ( .CLK(clock_bF_buf8), .D(state_3_bF_buf2), .Q(state_12_), .R(_abc_17692_n6660_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_217 ( .CLK(clock_bF_buf7), .D(state_4_), .Q(state_13_), .R(_abc_17692_n6660_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_218 ( .CLK(clock_bF_buf6), .D(state_5_), .Q(state_14_), .R(_abc_17692_n6660_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_219 ( .CLK(clock_bF_buf5), .D(state_6_bF_buf2), .Q(state_15_), .R(_abc_17692_n6660_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_22 ( .CLK(clock_bF_buf6), .D(data_out1_21__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30032_21_), .R(_abc_17692_n6660_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_23 ( .CLK(clock_bF_buf5), .D(data_out1_22__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30032_22_), .R(_abc_17692_n6660_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_24 ( .CLK(clock_bF_buf4), .D(data_out1_23__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30032_23_), .R(_abc_17692_n6660_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_25 ( .CLK(clock_bF_buf3), .D(data_out1_24__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30032_24_), .R(_abc_17692_n6660_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_26 ( .CLK(clock_bF_buf2), .D(data_out1_25__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30032_25_), .R(_abc_17692_n6660_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_27 ( .CLK(clock_bF_buf1), .D(data_out1_26__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30032_26_), .R(_abc_17692_n6660_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_28 ( .CLK(clock_bF_buf0), .D(data_out1_27__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30032_27_), .R(_abc_17692_n6660_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_29 ( .CLK(clock_bF_buf13), .D(data_out1_28__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30032_28_), .R(_abc_17692_n6660_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_3 ( .CLK(clock_bF_buf11), .D(data_out1_2__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30032_2_), .R(_abc_17692_n6660_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_30 ( .CLK(clock_bF_buf12), .D(data_out1_29__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30032_29_), .R(_abc_17692_n6660_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_31 ( .CLK(clock_bF_buf11), .D(data_out1_30__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30032_30_), .R(_abc_17692_n6660_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_32 ( .CLK(clock_bF_buf10), .D(data_out1_31__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30032_31_), .R(_abc_17692_n6660_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_33 ( .CLK(clock_bF_buf9), .D(data_out2_0__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30065_0_), .R(_abc_17692_n6660_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_34 ( .CLK(clock_bF_buf8), .D(data_out2_1__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30065_1_), .R(_abc_17692_n6660_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_35 ( .CLK(clock_bF_buf7), .D(data_out2_2__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30065_2_), .R(_abc_17692_n6660_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_36 ( .CLK(clock_bF_buf6), .D(data_out2_3__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30065_3_), .R(_abc_17692_n6660_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_37 ( .CLK(clock_bF_buf5), .D(data_out2_4__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30065_4_), .R(_abc_17692_n6660_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_38 ( .CLK(clock_bF_buf4), .D(data_out2_5__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30065_5_), .R(_abc_17692_n6660_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_39 ( .CLK(clock_bF_buf3), .D(data_out2_6__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30065_6_), .R(_abc_17692_n6660_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_4 ( .CLK(clock_bF_buf10), .D(data_out1_3__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30032_3_), .R(_abc_17692_n6660_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_40 ( .CLK(clock_bF_buf2), .D(data_out2_7__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30065_7_), .R(_abc_17692_n6660_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_41 ( .CLK(clock_bF_buf1), .D(data_out2_8__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30065_8_), .R(_abc_17692_n6660_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_42 ( .CLK(clock_bF_buf0), .D(data_out2_9__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30065_9_), .R(_abc_17692_n6660_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_43 ( .CLK(clock_bF_buf13), .D(data_out2_10__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30065_10_), .R(_abc_17692_n6660_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_44 ( .CLK(clock_bF_buf12), .D(data_out2_11__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30065_11_), .R(_abc_17692_n6660_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_45 ( .CLK(clock_bF_buf11), .D(data_out2_12__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30065_12_), .R(_abc_17692_n6660_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_46 ( .CLK(clock_bF_buf10), .D(data_out2_13__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30065_13_), .R(_abc_17692_n6660_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_47 ( .CLK(clock_bF_buf9), .D(data_out2_14__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30065_14_), .R(_abc_17692_n6660_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_48 ( .CLK(clock_bF_buf8), .D(data_out2_15__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30065_15_), .R(_abc_17692_n6660_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_49 ( .CLK(clock_bF_buf7), .D(data_out2_16__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30065_16_), .R(_abc_17692_n6660_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_5 ( .CLK(clock_bF_buf9), .D(data_out1_4__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30032_4_), .R(_abc_17692_n6660_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_50 ( .CLK(clock_bF_buf6), .D(data_out2_17__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30065_17_), .R(_abc_17692_n6660_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_51 ( .CLK(clock_bF_buf5), .D(data_out2_18__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30065_18_), .R(_abc_17692_n6660_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_52 ( .CLK(clock_bF_buf4), .D(data_out2_19__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30065_19_), .R(_abc_17692_n6660_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_53 ( .CLK(clock_bF_buf3), .D(data_out2_20__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30065_20_), .R(_abc_17692_n6660_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_54 ( .CLK(clock_bF_buf2), .D(data_out2_21__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30065_21_), .R(_abc_17692_n6660_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_55 ( .CLK(clock_bF_buf1), .D(data_out2_22__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30065_22_), .R(_abc_17692_n6660_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_56 ( .CLK(clock_bF_buf0), .D(data_out2_23__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30065_23_), .R(_abc_17692_n6660_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_57 ( .CLK(clock_bF_buf13), .D(data_out2_24__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30065_24_), .R(_abc_17692_n6660_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_58 ( .CLK(clock_bF_buf12), .D(data_out2_25__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30065_25_), .R(_abc_17692_n6660_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_59 ( .CLK(clock_bF_buf11), .D(data_out2_26__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30065_26_), .R(_abc_17692_n6660_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_6 ( .CLK(clock_bF_buf8), .D(data_out1_5__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30032_5_), .R(_abc_17692_n6660_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_60 ( .CLK(clock_bF_buf10), .D(data_out2_27__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30065_27_), .R(_abc_17692_n6660_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_61 ( .CLK(clock_bF_buf9), .D(data_out2_28__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30065_28_), .R(_abc_17692_n6660_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_62 ( .CLK(clock_bF_buf8), .D(data_out2_29__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30065_29_), .R(_abc_17692_n6660_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_63 ( .CLK(clock_bF_buf7), .D(data_out2_30__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30065_30_), .R(_abc_17692_n6660_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_64 ( .CLK(clock_bF_buf6), .D(data_out2_31__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30065_31_), .R(_abc_17692_n6660_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_65 ( .CLK(clock_bF_buf5), .D(while_flag_FF_INPUT), .Q(while_flag), .R(_abc_17692_n6660_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_66 ( .CLK(clock_bF_buf4), .D(modereg_FF_INPUT), .Q(modereg), .R(_abc_17692_n6660_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_67 ( .CLK(clock_bF_buf3), .D(selectslice_0__FF_INPUT), .Q(selectslice_0_), .R(_abc_17692_n6660_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_68 ( .CLK(clock_bF_buf2), .D(selectslice_1__FF_INPUT), .Q(selectslice_1_), .R(_abc_17692_n6660_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_69 ( .CLK(clock_bF_buf1), .D(x_0__FF_INPUT), .Q(x_0_), .R(_abc_17692_n6660_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_7 ( .CLK(clock_bF_buf7), .D(data_out1_6__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30032_6_), .R(_abc_17692_n6660_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_70 ( .CLK(clock_bF_buf0), .D(x_1__FF_INPUT), .Q(x_1_), .R(_abc_17692_n6660_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_71 ( .CLK(clock_bF_buf13), .D(x_2__FF_INPUT), .Q(x_2_), .R(_abc_17692_n6660_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_72 ( .CLK(clock_bF_buf12), .D(x_3__FF_INPUT), .Q(x_3_), .R(_abc_17692_n6660_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_73 ( .CLK(clock_bF_buf11), .D(x_4__FF_INPUT), .Q(x_4_), .R(_abc_17692_n6660_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_74 ( .CLK(clock_bF_buf10), .D(x_5__FF_INPUT), .Q(x_5_), .R(_abc_17692_n6660_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_75 ( .CLK(clock_bF_buf9), .D(x_6__FF_INPUT), .Q(x_6_), .R(_abc_17692_n6660_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_76 ( .CLK(clock_bF_buf8), .D(x_7__FF_INPUT), .Q(x_7_), .R(_abc_17692_n6660_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_77 ( .CLK(clock_bF_buf7), .D(sum_0__FF_INPUT), .Q(sum_0_), .R(_abc_17692_n6660_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_78 ( .CLK(clock_bF_buf6), .D(sum_1__FF_INPUT), .Q(sum_1_), .R(_abc_17692_n6660_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_79 ( .CLK(clock_bF_buf5), .D(sum_2__FF_INPUT), .Q(sum_2_), .R(_abc_17692_n6660_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_8 ( .CLK(clock_bF_buf6), .D(data_out1_7__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30032_7_), .R(_abc_17692_n6660_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_80 ( .CLK(clock_bF_buf4), .D(sum_3__FF_INPUT), .Q(sum_3_), .R(_abc_17692_n6660_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_81 ( .CLK(clock_bF_buf3), .D(sum_4__FF_INPUT), .Q(sum_4_), .R(_abc_17692_n6660_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_82 ( .CLK(clock_bF_buf2), .D(sum_5__FF_INPUT), .Q(sum_5_), .R(_abc_17692_n6660_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_83 ( .CLK(clock_bF_buf1), .D(sum_6__FF_INPUT), .Q(sum_6_), .R(_abc_17692_n6660_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_84 ( .CLK(clock_bF_buf0), .D(sum_7__FF_INPUT), .Q(sum_7_), .R(_abc_17692_n6660_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_85 ( .CLK(clock_bF_buf13), .D(sum_8__FF_INPUT), .Q(sum_8_), .R(_abc_17692_n6660_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_86 ( .CLK(clock_bF_buf12), .D(sum_9__FF_INPUT), .Q(sum_9_), .R(_abc_17692_n6660_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_87 ( .CLK(clock_bF_buf11), .D(sum_10__FF_INPUT), .Q(sum_10_), .R(_abc_17692_n6660_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_88 ( .CLK(clock_bF_buf10), .D(sum_11__FF_INPUT), .Q(sum_11_), .R(_abc_17692_n6660_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_89 ( .CLK(clock_bF_buf9), .D(sum_12__FF_INPUT), .Q(sum_12_), .R(_abc_17692_n6660_bF_buf9), .S(1'b1) );
  DFFSR DFFSR_9 ( .CLK(clock_bF_buf5), .D(data_out1_8__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_30032_8_), .R(_abc_17692_n6660_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_90 ( .CLK(clock_bF_buf8), .D(sum_13__FF_INPUT), .Q(sum_13_), .R(_abc_17692_n6660_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_91 ( .CLK(clock_bF_buf7), .D(sum_14__FF_INPUT), .Q(sum_14_), .R(_abc_17692_n6660_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_92 ( .CLK(clock_bF_buf6), .D(sum_15__FF_INPUT), .Q(sum_15_), .R(_abc_17692_n6660_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_93 ( .CLK(clock_bF_buf5), .D(sum_16__FF_INPUT), .Q(sum_16_), .R(_abc_17692_n6660_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_94 ( .CLK(clock_bF_buf4), .D(sum_17__FF_INPUT), .Q(sum_17_), .R(_abc_17692_n6660_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_95 ( .CLK(clock_bF_buf3), .D(sum_18__FF_INPUT), .Q(sum_18_), .R(_abc_17692_n6660_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_96 ( .CLK(clock_bF_buf2), .D(sum_19__FF_INPUT), .Q(sum_19_), .R(_abc_17692_n6660_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_97 ( .CLK(clock_bF_buf1), .D(sum_20__FF_INPUT), .Q(sum_20_), .R(_abc_17692_n6660_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_98 ( .CLK(clock_bF_buf0), .D(sum_21__FF_INPUT), .Q(sum_21_), .R(_abc_17692_n6660_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_99 ( .CLK(clock_bF_buf13), .D(sum_22__FF_INPUT), .Q(sum_22_), .R(_abc_17692_n6660_bF_buf13), .S(1'b1) );
  INVX1 INVX1_1 ( .A(while_flag), .Y(_abc_17692_n623) );
  INVX1 INVX1_10 ( .A(_abc_17692_n688), .Y(_abc_17692_n689) );
  INVX1 INVX1_100 ( .A(_abc_17692_n1216), .Y(_abc_17692_n1217) );
  INVX1 INVX1_1000 ( .A(_abc_17692_n5521), .Y(_abc_17692_n5522) );
  INVX1 INVX1_1001 ( .A(_abc_17692_n5525), .Y(_abc_17692_n5526) );
  INVX1 INVX1_1002 ( .A(_abc_17692_n5529), .Y(_abc_17692_n5530) );
  INVX1 INVX1_1003 ( .A(_abc_17692_n5531), .Y(_abc_17692_n5532) );
  INVX1 INVX1_1004 ( .A(_abc_17692_n5534), .Y(_abc_17692_n5535) );
  INVX1 INVX1_1005 ( .A(_abc_17692_n5539), .Y(_abc_17692_n5540) );
  INVX1 INVX1_1006 ( .A(_abc_17692_n5551), .Y(_abc_17692_n5552) );
  INVX1 INVX1_1007 ( .A(_abc_17692_n5419), .Y(_abc_17692_n5556) );
  INVX1 INVX1_1008 ( .A(_abc_17692_n5559), .Y(_abc_17692_n5560) );
  INVX1 INVX1_1009 ( .A(_abc_17692_n5569), .Y(_abc_17692_n5570) );
  INVX1 INVX1_101 ( .A(_abc_17692_n1219), .Y(_abc_17692_n1220) );
  INVX1 INVX1_1010 ( .A(_abc_17692_n5293), .Y(_abc_17692_n5574) );
  INVX1 INVX1_1011 ( .A(_abc_17692_n5576), .Y(_abc_17692_n5577) );
  INVX1 INVX1_1012 ( .A(_abc_17692_n5581), .Y(_abc_17692_n5582) );
  INVX1 INVX1_1013 ( .A(_abc_17692_n5595), .Y(_abc_17692_n5596) );
  INVX1 INVX1_1014 ( .A(_abc_17692_n5600), .Y(_abc_17692_n5601) );
  INVX1 INVX1_1015 ( .A(_abc_17692_n5602), .Y(_abc_17692_n5603) );
  INVX1 INVX1_1016 ( .A(_abc_17692_n5604), .Y(_abc_17692_n5605) );
  INVX1 INVX1_1017 ( .A(_abc_17692_n5606), .Y(_abc_17692_n5608_1) );
  INVX1 INVX1_1018 ( .A(_abc_17692_n5613), .Y(_abc_17692_n5614) );
  INVX1 INVX1_1019 ( .A(_abc_17692_n5617), .Y(_abc_17692_n5618) );
  INVX1 INVX1_102 ( .A(_abc_17692_n1226), .Y(_abc_17692_n1227) );
  INVX1 INVX1_1020 ( .A(_abc_17692_n5620), .Y(_abc_17692_n5622) );
  INVX1 INVX1_1021 ( .A(_abc_17692_n5624), .Y(_abc_17692_n5627) );
  INVX1 INVX1_1022 ( .A(_abc_17692_n5415), .Y(_abc_17692_n5630) );
  INVX1 INVX1_1023 ( .A(_abc_17692_n5629), .Y(_abc_17692_n5634) );
  INVX1 INVX1_1024 ( .A(_abc_17692_n5632), .Y(_abc_17692_n5635) );
  INVX1 INVX1_1025 ( .A(_abc_17692_n5639), .Y(_abc_17692_n5640) );
  INVX1 INVX1_1026 ( .A(_abc_17692_n5641), .Y(_abc_17692_n5642) );
  INVX1 INVX1_1027 ( .A(_abc_17692_n5645), .Y(_abc_17692_n5646) );
  INVX1 INVX1_1028 ( .A(_abc_17692_n5647), .Y(_abc_17692_n5650) );
  INVX1 INVX1_1029 ( .A(_abc_17692_n5660), .Y(_abc_17692_n5661) );
  INVX1 INVX1_103 ( .A(_abc_17692_n1231), .Y(_abc_17692_n1232) );
  INVX1 INVX1_1030 ( .A(_abc_17692_n5662), .Y(_abc_17692_n5667) );
  INVX1 INVX1_1031 ( .A(_abc_17692_n5671), .Y(_abc_17692_n5672) );
  INVX1 INVX1_1032 ( .A(_abc_17692_n5673), .Y(_abc_17692_n5674) );
  INVX1 INVX1_1033 ( .A(_abc_17692_n5678), .Y(_abc_17692_n5679) );
  INVX1 INVX1_1034 ( .A(_abc_17692_n5677), .Y(_abc_17692_n5682) );
  INVX1 INVX1_1035 ( .A(_abc_17692_n5692_1), .Y(_abc_17692_n5693) );
  INVX1 INVX1_1036 ( .A(_abc_17692_n5691), .Y(_abc_17692_n5695_1) );
  INVX1 INVX1_1037 ( .A(_abc_17692_n5699), .Y(_abc_17692_n5700) );
  INVX1 INVX1_1038 ( .A(_abc_17692_n5701), .Y(_abc_17692_n5702) );
  INVX1 INVX1_1039 ( .A(_abc_17692_n5706), .Y(_abc_17692_n5707) );
  INVX1 INVX1_104 ( .A(_abc_17692_n1233), .Y(_abc_17692_n1234) );
  INVX1 INVX1_1040 ( .A(_abc_17692_n5705), .Y(_abc_17692_n5710) );
  INVX1 INVX1_1041 ( .A(_abc_17692_n5719), .Y(_abc_17692_n5720) );
  INVX1 INVX1_1042 ( .A(_abc_17692_n5721), .Y(_abc_17692_n5723) );
  INVX1 INVX1_1043 ( .A(_abc_17692_n5528), .Y(_abc_17692_n5731) );
  INVX1 INVX1_1044 ( .A(_abc_17692_n5732), .Y(_abc_17692_n5733) );
  INVX1 INVX1_1045 ( .A(_abc_17692_n5738), .Y(_abc_17692_n5739) );
  INVX1 INVX1_1046 ( .A(_abc_17692_n5745_1), .Y(_abc_17692_n5746) );
  INVX1 INVX1_1047 ( .A(_abc_17692_n5751), .Y(_abc_17692_n5752) );
  INVX1 INVX1_1048 ( .A(_abc_17692_n5753), .Y(_abc_17692_n5754) );
  INVX1 INVX1_1049 ( .A(_abc_17692_n5773), .Y(_abc_17692_n5774) );
  INVX1 INVX1_105 ( .A(_abc_17692_n1235), .Y(_abc_17692_n1236) );
  INVX1 INVX1_1050 ( .A(_abc_17692_n5382), .Y(_abc_17692_n5775) );
  INVX1 INVX1_1051 ( .A(_abc_17692_n5778), .Y(_abc_17692_n5779) );
  INVX1 INVX1_1052 ( .A(_abc_17692_n5784), .Y(_abc_17692_n5785) );
  INVX1 INVX1_1053 ( .A(_abc_17692_n5788), .Y(_abc_17692_n5789) );
  INVX1 INVX1_1054 ( .A(_abc_17692_n5771), .Y(_abc_17692_n5791) );
  INVX1 INVX1_1055 ( .A(_abc_17692_n5804), .Y(_abc_17692_n5805) );
  INVX1 INVX1_1056 ( .A(_abc_17692_n5798), .Y(_abc_17692_n5809) );
  INVX1 INVX1_1057 ( .A(_abc_17692_n5802), .Y(_abc_17692_n5810) );
  INVX1 INVX1_1058 ( .A(_abc_17692_n5807), .Y(_abc_17692_n5812) );
  INVX1 INVX1_1059 ( .A(_abc_17692_n5814), .Y(_abc_17692_n5815) );
  INVX1 INVX1_106 ( .A(_abc_17692_n1244), .Y(_abc_17692_n1245) );
  INVX1 INVX1_1060 ( .A(_abc_17692_n5819), .Y(_abc_17692_n5820) );
  INVX1 INVX1_1061 ( .A(_abc_17692_n5823), .Y(_abc_17692_n5824) );
  INVX1 INVX1_1062 ( .A(_abc_17692_n5826), .Y(_abc_17692_n5827) );
  INVX1 INVX1_1063 ( .A(_abc_17692_n5829), .Y(_abc_17692_n5830) );
  INVX1 INVX1_1064 ( .A(_abc_17692_n5833), .Y(_abc_17692_n5834) );
  INVX1 INVX1_1065 ( .A(_abc_17692_n5836), .Y(_abc_17692_n5837) );
  INVX1 INVX1_1066 ( .A(_abc_17692_n5838), .Y(_abc_17692_n5839) );
  INVX1 INVX1_1067 ( .A(_abc_17692_n5851), .Y(_abc_17692_n5852) );
  INVX1 INVX1_1068 ( .A(_abc_17692_n5850), .Y(_abc_17692_n5856) );
  INVX1 INVX1_1069 ( .A(_abc_17692_n5854), .Y(_abc_17692_n5857) );
  INVX1 INVX1_107 ( .A(delta_13_), .Y(_abc_17692_n1246) );
  INVX1 INVX1_1070 ( .A(_abc_17692_n5859), .Y(_abc_17692_n5860) );
  INVX1 INVX1_1071 ( .A(_abc_17692_n5864), .Y(_abc_17692_n5865) );
  INVX1 INVX1_1072 ( .A(_abc_17692_n5868), .Y(_abc_17692_n5869) );
  INVX1 INVX1_1073 ( .A(_abc_17692_n5873), .Y(_abc_17692_n5874) );
  INVX1 INVX1_1074 ( .A(_abc_17692_n5877), .Y(_abc_17692_n5878) );
  INVX1 INVX1_1075 ( .A(_abc_17692_n5879), .Y(_abc_17692_n5880) );
  INVX1 INVX1_1076 ( .A(_abc_17692_n5881), .Y(_abc_17692_n5882) );
  INVX1 INVX1_1077 ( .A(_abc_17692_n5894), .Y(_abc_17692_n5895) );
  INVX1 INVX1_1078 ( .A(_abc_17692_n5887), .Y(_abc_17692_n5899) );
  INVX1 INVX1_1079 ( .A(_abc_17692_n5892), .Y(_abc_17692_n5901) );
  INVX1 INVX1_108 ( .A(sum_13_), .Y(_abc_17692_n1247) );
  INVX1 INVX1_1080 ( .A(_abc_17692_n5897), .Y(_abc_17692_n5903_1) );
  INVX1 INVX1_1081 ( .A(_abc_17692_n5905), .Y(_abc_17692_n5906) );
  INVX1 INVX1_1082 ( .A(_abc_17692_n5909), .Y(_abc_17692_n5910) );
  INVX1 INVX1_1083 ( .A(_abc_17692_n5914), .Y(_abc_17692_n5915) );
  INVX1 INVX1_1084 ( .A(_abc_17692_n5917), .Y(_abc_17692_n5918) );
  INVX1 INVX1_1085 ( .A(_abc_17692_n5919), .Y(_abc_17692_n5920) );
  INVX1 INVX1_1086 ( .A(_abc_17692_n5923), .Y(_abc_17692_n5924) );
  INVX1 INVX1_1087 ( .A(_abc_17692_n5913), .Y(_abc_17692_n5928) );
  INVX1 INVX1_1088 ( .A(_abc_17692_n5926), .Y(_abc_17692_n5929) );
  INVX1 INVX1_1089 ( .A(_abc_17692_n5941), .Y(_abc_17692_n5942) );
  INVX1 INVX1_109 ( .A(_abc_17692_n1248), .Y(_abc_17692_n1249) );
  INVX1 INVX1_1090 ( .A(_abc_17692_n5934), .Y(_abc_17692_n5946) );
  INVX1 INVX1_1091 ( .A(_abc_17692_n5939), .Y(_abc_17692_n5948) );
  INVX1 INVX1_1092 ( .A(_abc_17692_n5944), .Y(_abc_17692_n5950) );
  INVX1 INVX1_1093 ( .A(_abc_17692_n5952), .Y(_abc_17692_n5953) );
  INVX1 INVX1_1094 ( .A(_abc_17692_n5956), .Y(_abc_17692_n5957) );
  INVX1 INVX1_1095 ( .A(_abc_17692_n5963), .Y(_abc_17692_n5964) );
  INVX1 INVX1_1096 ( .A(_abc_17692_n5961), .Y(_abc_17692_n5968) );
  INVX1 INVX1_1097 ( .A(_abc_17692_n5969), .Y(_abc_17692_n5970) );
  INVX1 INVX1_1098 ( .A(_abc_17692_n5960), .Y(_abc_17692_n5974) );
  INVX1 INVX1_1099 ( .A(_abc_17692_n5972), .Y(_abc_17692_n5975) );
  INVX1 INVX1_11 ( .A(_abc_17692_n692_1), .Y(_abc_17692_n693_1) );
  INVX1 INVX1_110 ( .A(_abc_17692_n1204), .Y(_abc_17692_n1252) );
  INVX1 INVX1_1100 ( .A(_abc_17692_n5987), .Y(_abc_17692_n5988) );
  INVX1 INVX1_1101 ( .A(_abc_17692_n5994), .Y(_abc_17692_n5995) );
  INVX1 INVX1_1102 ( .A(_abc_17692_n5867), .Y(_abc_17692_n5998) );
  INVX1 INVX1_1103 ( .A(_abc_17692_n5625), .Y(_abc_17692_n6003) );
  INVX1 INVX1_1104 ( .A(_abc_17692_n5631), .Y(_abc_17692_n6004) );
  INVX1 INVX1_1105 ( .A(_abc_17692_n6001), .Y(_abc_17692_n6009) );
  INVX1 INVX1_1106 ( .A(_abc_17692_n6010), .Y(_abc_17692_n6011) );
  INVX1 INVX1_1107 ( .A(_abc_17692_n6013), .Y(_abc_17692_n6014) );
  INVX1 INVX1_1108 ( .A(_abc_17692_n6015), .Y(_abc_17692_n6016) );
  INVX1 INVX1_1109 ( .A(_abc_17692_n5686), .Y(_abc_17692_n6022) );
  INVX1 INVX1_111 ( .A(_abc_17692_n1253), .Y(_abc_17692_n1255) );
  INVX1 INVX1_1110 ( .A(_abc_17692_n5449), .Y(_abc_17692_n6023) );
  INVX1 INVX1_1111 ( .A(_abc_17692_n6026), .Y(_abc_17692_n6027) );
  INVX1 INVX1_1112 ( .A(_abc_17692_n6029), .Y(_abc_17692_n6030) );
  INVX1 INVX1_1113 ( .A(_abc_17692_n6031), .Y(_abc_17692_n6032) );
  INVX1 INVX1_1114 ( .A(_abc_17692_n6034), .Y(_abc_17692_n6035) );
  INVX1 INVX1_1115 ( .A(_abc_17692_n5714), .Y(_abc_17692_n6040) );
  INVX1 INVX1_1116 ( .A(_abc_17692_n5487), .Y(_abc_17692_n6041_1) );
  INVX1 INVX1_1117 ( .A(_abc_17692_n6048), .Y(_abc_17692_n6049) );
  INVX1 INVX1_1118 ( .A(_abc_17692_n6062), .Y(_abc_17692_n6063) );
  INVX1 INVX1_1119 ( .A(_abc_17692_n6067), .Y(_abc_17692_n6068) );
  INVX1 INVX1_112 ( .A(_abc_17692_n1263), .Y(_abc_17692_n1264) );
  INVX1 INVX1_1120 ( .A(_abc_17692_n6069), .Y(_abc_17692_n6070) );
  INVX1 INVX1_1121 ( .A(_abc_17692_n6071), .Y(_abc_17692_n6072) );
  INVX1 INVX1_1122 ( .A(_abc_17692_n6074), .Y(_abc_17692_n6075) );
  INVX1 INVX1_1123 ( .A(_abc_17692_n6078), .Y(_abc_17692_n6079) );
  INVX1 INVX1_1124 ( .A(_abc_17692_n6080), .Y(_abc_17692_n6081) );
  INVX1 INVX1_1125 ( .A(_abc_17692_n6083), .Y(_abc_17692_n6085) );
  INVX1 INVX1_1126 ( .A(_abc_17692_n6087), .Y(_abc_17692_n6088) );
  INVX1 INVX1_1127 ( .A(_abc_17692_n6076), .Y(_abc_17692_n6090) );
  INVX1 INVX1_1128 ( .A(_abc_17692_n6093), .Y(_abc_17692_n6096) );
  INVX1 INVX1_1129 ( .A(_abc_17692_n6099), .Y(_abc_17692_n6100) );
  INVX1 INVX1_113 ( .A(_abc_17692_n1265), .Y(_abc_17692_n1266) );
  INVX1 INVX1_1130 ( .A(_abc_17692_n6098), .Y(_abc_17692_n6102) );
  INVX1 INVX1_1131 ( .A(_abc_17692_n6107), .Y(_abc_17692_n6108) );
  INVX1 INVX1_1132 ( .A(_abc_17692_n6110), .Y(_abc_17692_n6111) );
  INVX1 INVX1_1133 ( .A(_abc_17692_n6113), .Y(_abc_17692_n6114) );
  INVX1 INVX1_1134 ( .A(_abc_17692_n6115), .Y(_abc_17692_n6116) );
  INVX1 INVX1_1135 ( .A(_abc_17692_n6119), .Y(_abc_17692_n6120) );
  INVX1 INVX1_1136 ( .A(_abc_17692_n5912), .Y(_abc_17692_n6124) );
  INVX1 INVX1_1137 ( .A(_abc_17692_n6125), .Y(_abc_17692_n6126) );
  INVX1 INVX1_1138 ( .A(_abc_17692_n6121), .Y(_abc_17692_n6128) );
  INVX1 INVX1_1139 ( .A(_abc_17692_n6122), .Y(_abc_17692_n6129) );
  INVX1 INVX1_114 ( .A(sum_14_), .Y(_abc_17692_n1274) );
  INVX1 INVX1_1140 ( .A(_abc_17692_n6134), .Y(_abc_17692_n6135) );
  INVX1 INVX1_1141 ( .A(_abc_17692_n6136), .Y(_abc_17692_n6137) );
  INVX1 INVX1_1142 ( .A(_abc_17692_n6140), .Y(_abc_17692_n6141) );
  INVX1 INVX1_1143 ( .A(_abc_17692_n6143), .Y(_abc_17692_n6144) );
  INVX1 INVX1_1144 ( .A(_abc_17692_n6153), .Y(_abc_17692_n6154) );
  INVX1 INVX1_1145 ( .A(_abc_17692_n5959), .Y(_abc_17692_n6155) );
  INVX1 INVX1_1146 ( .A(_abc_17692_n6156), .Y(_abc_17692_n6157) );
  INVX1 INVX1_1147 ( .A(_abc_17692_n6166_1), .Y(_abc_17692_n6167) );
  INVX1 INVX1_1148 ( .A(_abc_17692_n6169_1), .Y(_abc_17692_n6170) );
  INVX1 INVX1_1149 ( .A(_abc_17692_n6172), .Y(_abc_17692_n6173) );
  INVX1 INVX1_115 ( .A(_abc_17692_n1276), .Y(_abc_17692_n1277) );
  INVX1 INVX1_1150 ( .A(_abc_17692_n6174), .Y(_abc_17692_n6176) );
  INVX1 INVX1_1151 ( .A(_abc_17692_n6179), .Y(_abc_17692_n6180) );
  INVX1 INVX1_1152 ( .A(_abc_17692_n6178), .Y(_abc_17692_n6181) );
  INVX1 INVX1_1153 ( .A(_abc_17692_n6182), .Y(_abc_17692_n6183) );
  INVX1 INVX1_1154 ( .A(_abc_17692_n5822), .Y(_abc_17692_n6185) );
  INVX1 INVX1_1155 ( .A(_abc_17692_n6186), .Y(_abc_17692_n6187) );
  INVX1 INVX1_1156 ( .A(_abc_17692_n6184), .Y(_abc_17692_n6189) );
  INVX1 INVX1_1157 ( .A(_abc_17692_n6195), .Y(_abc_17692_n6196) );
  INVX1 INVX1_1158 ( .A(_abc_17692_n6197), .Y(_abc_17692_n6199) );
  INVX1 INVX1_1159 ( .A(_abc_17692_n5863), .Y(_abc_17692_n6203) );
  INVX1 INVX1_116 ( .A(_abc_17692_n1282), .Y(_abc_17692_n1283) );
  INVX1 INVX1_1160 ( .A(_abc_17692_n6204), .Y(_abc_17692_n6205) );
  INVX1 INVX1_1161 ( .A(_abc_17692_n6206), .Y(_abc_17692_n6208) );
  INVX1 INVX1_1162 ( .A(_abc_17692_n6212), .Y(_abc_17692_n6213) );
  INVX1 INVX1_1163 ( .A(_abc_17692_n6214), .Y(_abc_17692_n6216) );
  INVX1 INVX1_1164 ( .A(_abc_17692_n6221), .Y(_abc_17692_n6223) );
  INVX1 INVX1_1165 ( .A(_abc_17692_n6244), .Y(_abc_17692_n6245) );
  INVX1 INVX1_1166 ( .A(_abc_17692_n6248), .Y(_abc_17692_n6249) );
  INVX1 INVX1_1167 ( .A(_abc_17692_n6236), .Y(_abc_17692_n6251) );
  INVX1 INVX1_1168 ( .A(_abc_17692_n6239), .Y(_abc_17692_n6253) );
  INVX1 INVX1_1169 ( .A(_abc_17692_n6258), .Y(_abc_17692_n6259) );
  INVX1 INVX1_117 ( .A(_abc_17692_n1285), .Y(_abc_17692_n1286) );
  INVX1 INVX1_1170 ( .A(_abc_17692_n6082), .Y(_abc_17692_n6260) );
  INVX1 INVX1_1171 ( .A(_abc_17692_n6263), .Y(_abc_17692_n6264) );
  INVX1 INVX1_1172 ( .A(_abc_17692_n6265), .Y(_abc_17692_n6266) );
  INVX1 INVX1_1173 ( .A(_abc_17692_n6268), .Y(_abc_17692_n6270) );
  INVX1 INVX1_1174 ( .A(_abc_17692_n6272), .Y(_abc_17692_n6273) );
  INVX1 INVX1_1175 ( .A(_abc_17692_n6256), .Y(_abc_17692_n6275) );
  INVX1 INVX1_1176 ( .A(_abc_17692_n6278), .Y(_abc_17692_n6279) );
  INVX1 INVX1_1177 ( .A(_abc_17692_n6288), .Y(_abc_17692_n6289) );
  INVX1 INVX1_1178 ( .A(_abc_17692_n6109), .Y(_abc_17692_n6296) );
  INVX1 INVX1_1179 ( .A(_abc_17692_n6298), .Y(_abc_17692_n6299) );
  INVX1 INVX1_118 ( .A(_abc_17692_n1278), .Y(_abc_17692_n1290) );
  INVX1 INVX1_1180 ( .A(_abc_17692_n6301), .Y(_abc_17692_n6302) );
  INVX1 INVX1_1181 ( .A(_abc_17692_n6294), .Y(_abc_17692_n6306) );
  INVX1 INVX1_1182 ( .A(_abc_17692_n6304), .Y(_abc_17692_n6309) );
  INVX1 INVX1_1183 ( .A(_abc_17692_n6311), .Y(_abc_17692_n6313) );
  INVX1 INVX1_1184 ( .A(_abc_17692_n6315), .Y(_abc_17692_n6316_1) );
  INVX1 INVX1_1185 ( .A(_abc_17692_n6319_1), .Y(_abc_17692_n6320) );
  INVX1 INVX1_1186 ( .A(_abc_17692_n6327), .Y(_abc_17692_n6328) );
  INVX1 INVX1_1187 ( .A(_abc_17692_n6138), .Y(_abc_17692_n6334) );
  INVX1 INVX1_1188 ( .A(_abc_17692_n6336), .Y(_abc_17692_n6337) );
  INVX1 INVX1_1189 ( .A(_abc_17692_n6339), .Y(_abc_17692_n6340) );
  INVX1 INVX1_119 ( .A(_abc_17692_n1292), .Y(_abc_17692_n1293) );
  INVX1 INVX1_1190 ( .A(_abc_17692_n6332), .Y(_abc_17692_n6344) );
  INVX1 INVX1_1191 ( .A(_abc_17692_n6342), .Y(_abc_17692_n6347) );
  INVX1 INVX1_1192 ( .A(_abc_17692_n6349), .Y(_abc_17692_n6350) );
  INVX1 INVX1_1193 ( .A(_abc_17692_n6353), .Y(_abc_17692_n6354) );
  INVX1 INVX1_1194 ( .A(_abc_17692_n6357), .Y(_abc_17692_n6358) );
  INVX1 INVX1_1195 ( .A(_abc_17692_n6359), .Y(_abc_17692_n6360) );
  INVX1 INVX1_1196 ( .A(_abc_17692_n6365), .Y(_abc_17692_n6366) );
  INVX1 INVX1_1197 ( .A(_abc_17692_n6168), .Y(_abc_17692_n6375) );
  INVX1 INVX1_1198 ( .A(_abc_17692_n6377), .Y(_abc_17692_n6378) );
  INVX1 INVX1_1199 ( .A(_abc_17692_n6380), .Y(_abc_17692_n6381) );
  INVX1 INVX1_12 ( .A(_abc_17692_n696), .Y(_abc_17692_n697) );
  INVX1 INVX1_120 ( .A(_abc_17692_n1294), .Y(_abc_17692_n1295) );
  INVX1 INVX1_1200 ( .A(_abc_17692_n6374_1), .Y(_abc_17692_n6385) );
  INVX1 INVX1_1201 ( .A(_abc_17692_n6383), .Y(_abc_17692_n6387) );
  INVX1 INVX1_1202 ( .A(_abc_17692_n6389), .Y(_abc_17692_n6391) );
  INVX1 INVX1_1203 ( .A(_abc_17692_n6393), .Y(_abc_17692_n6394) );
  INVX1 INVX1_1204 ( .A(_abc_17692_n6405), .Y(_abc_17692_n6406) );
  INVX1 INVX1_1205 ( .A(_abc_17692_n6414), .Y(_abc_17692_n6416) );
  INVX1 INVX1_1206 ( .A(_abc_17692_n6281), .Y(_abc_17692_n6420) );
  INVX1 INVX1_1207 ( .A(_abc_17692_n6421), .Y(_abc_17692_n6422) );
  INVX1 INVX1_1208 ( .A(_abc_17692_n6094), .Y(_abc_17692_n6424) );
  INVX1 INVX1_1209 ( .A(_abc_17692_n6426), .Y(_abc_17692_n6427) );
  INVX1 INVX1_121 ( .A(_abc_17692_n1296), .Y(_abc_17692_n1297) );
  INVX1 INVX1_1210 ( .A(_abc_17692_n6429), .Y(_abc_17692_n6430) );
  INVX1 INVX1_1211 ( .A(_abc_17692_n6148), .Y(_abc_17692_n6434) );
  INVX1 INVX1_1212 ( .A(_abc_17692_n6436), .Y(_abc_17692_n6437) );
  INVX1 INVX1_1213 ( .A(_abc_17692_n6438), .Y(_abc_17692_n6439) );
  INVX1 INVX1_1214 ( .A(_abc_17692_n6441), .Y(_abc_17692_n6443) );
  INVX1 INVX1_1215 ( .A(_abc_17692_n6452), .Y(_abc_17692_n6453) );
  INVX1 INVX1_1216 ( .A(_abc_17692_n6470), .Y(_abc_17692_n6471) );
  INVX1 INVX1_1217 ( .A(_abc_17692_n6472), .Y(_abc_17692_n6473) );
  INVX1 INVX1_1218 ( .A(_abc_17692_n6474), .Y(_abc_17692_n6475) );
  INVX1 INVX1_1219 ( .A(_abc_17692_n6476), .Y(_abc_17692_n6477) );
  INVX1 INVX1_122 ( .A(sum_15_), .Y(_abc_17692_n1303) );
  INVX1 INVX1_1220 ( .A(_abc_17692_n6246), .Y(_abc_17692_n6479) );
  INVX1 INVX1_1221 ( .A(_abc_17692_n6486), .Y(_abc_17692_n6487) );
  INVX1 INVX1_1222 ( .A(_abc_17692_n6490), .Y(_abc_17692_n6491) );
  INVX1 INVX1_1223 ( .A(_abc_17692_n6485), .Y(_abc_17692_n6498) );
  INVX1 INVX1_1224 ( .A(_abc_17692_n6489), .Y(_abc_17692_n6499) );
  INVX1 INVX1_1225 ( .A(_abc_17692_n6511), .Y(_abc_17692_n6512) );
  INVX1 INVX1_1226 ( .A(_abc_17692_n6510), .Y(_abc_17692_n6514) );
  INVX1 INVX1_1227 ( .A(_abc_17692_n6520), .Y(_abc_17692_n6521) );
  INVX1 INVX1_1228 ( .A(_abc_17692_n6523_1), .Y(_abc_17692_n6526_1) );
  INVX1 INVX1_1229 ( .A(_abc_17692_n6540), .Y(_abc_17692_n6541) );
  INVX1 INVX1_123 ( .A(_abc_17692_n1304), .Y(_abc_17692_n1305) );
  INVX1 INVX1_1230 ( .A(_abc_17692_n6356), .Y(_abc_17692_n6542) );
  INVX1 INVX1_1231 ( .A(_abc_17692_n6543), .Y(_abc_17692_n6544) );
  INVX1 INVX1_1232 ( .A(_abc_17692_n6551), .Y(_abc_17692_n6552) );
  INVX1 INVX1_1233 ( .A(_abc_17692_n6554), .Y(_abc_17692_n6557) );
  INVX1 INVX1_1234 ( .A(_abc_17692_n6571), .Y(_abc_17692_n6572) );
  INVX1 INVX1_1235 ( .A(_abc_17692_n6573), .Y(_abc_17692_n6574) );
  INVX1 INVX1_1236 ( .A(_abc_17692_n6575), .Y(_abc_17692_n6576) );
  INVX1 INVX1_1237 ( .A(_abc_17692_n6584), .Y(_abc_17692_n6585) );
  INVX1 INVX1_1238 ( .A(_abc_17692_n6587), .Y(_abc_17692_n6588) );
  INVX1 INVX1_1239 ( .A(_abc_17692_n6590), .Y(_abc_17692_n6591) );
  INVX1 INVX1_124 ( .A(_abc_17692_n1308_1), .Y(_abc_17692_n1309) );
  INVX1 INVX1_1240 ( .A(_abc_17692_n6384), .Y(_abc_17692_n6594) );
  INVX1 INVX1_1241 ( .A(_abc_17692_n6606), .Y(_abc_17692_n6607) );
  INVX1 INVX1_1242 ( .A(_abc_17692_n6608), .Y(_abc_17692_n6609) );
  INVX1 INVX1_1243 ( .A(_abc_17692_n6619), .Y(_abc_17692_n6620) );
  INVX1 INVX1_1244 ( .A(_abc_17692_n6277), .Y(_abc_17692_n6625) );
  INVX1 INVX1_1245 ( .A(_abc_17692_n6627), .Y(_abc_17692_n6629) );
  INVX1 INVX1_1246 ( .A(_abc_17692_n6633), .Y(_abc_17692_n6634) );
  INVX1 INVX1_1247 ( .A(_abc_17692_n6635), .Y(_abc_17692_n6636) );
  INVX1 INVX1_1248 ( .A(_abc_17692_n6317), .Y(_abc_17692_n6641) );
  INVX1 INVX1_1249 ( .A(_abc_17692_n6642), .Y(_abc_17692_n6643) );
  INVX1 INVX1_125 ( .A(_abc_17692_n1310), .Y(_abc_17692_n1313) );
  INVX1 INVX1_1250 ( .A(_abc_17692_n6661), .Y(_abc_17692_n6662) );
  INVX1 INVX1_1251 ( .A(_abc_17692_n6665), .Y(_abc_17692_n6666) );
  INVX1 INVX1_1252 ( .A(_abc_17692_n6668), .Y(_abc_17692_n6669) );
  INVX1 INVX1_1253 ( .A(_abc_17692_n6672), .Y(_abc_17692_n6673) );
  INVX1 INVX1_1254 ( .A(_abc_17692_n6671), .Y(_abc_17692_n6677) );
  INVX1 INVX1_1255 ( .A(_abc_17692_n6682), .Y(_abc_17692_n6683) );
  INVX1 INVX1_1256 ( .A(_abc_17692_n6687), .Y(_abc_17692_n6688) );
  INVX1 INVX1_1257 ( .A(_abc_17692_n6689), .Y(_abc_17692_n6690) );
  INVX1 INVX1_1258 ( .A(_abc_17692_n6685), .Y(_abc_17692_n6696) );
  INVX1 INVX1_1259 ( .A(_abc_17692_n6694), .Y(_abc_17692_n6697) );
  INVX1 INVX1_126 ( .A(_abc_17692_n1318), .Y(_abc_17692_n1319) );
  INVX1 INVX1_1260 ( .A(_abc_17692_n6699), .Y(_abc_17692_n6700) );
  INVX1 INVX1_1261 ( .A(_abc_17692_n6704), .Y(_abc_17692_n6705) );
  INVX1 INVX1_1262 ( .A(_abc_17692_n6708), .Y(_abc_17692_n6709) );
  INVX1 INVX1_1263 ( .A(_abc_17692_n6715), .Y(_abc_17692_n6716) );
  INVX1 INVX1_1264 ( .A(_abc_17692_n6717), .Y(_abc_17692_n6718) );
  INVX1 INVX1_1265 ( .A(_abc_17692_n6720), .Y(_abc_17692_n6721) );
  INVX1 INVX1_1266 ( .A(_abc_17692_n6722), .Y(_abc_17692_n6723) );
  INVX1 INVX1_1267 ( .A(_abc_17692_n6727), .Y(_abc_17692_n6728) );
  INVX1 INVX1_1268 ( .A(_abc_17692_n6732), .Y(_abc_17692_n6733) );
  INVX1 INVX1_1269 ( .A(_abc_17692_n6734), .Y(_abc_17692_n6735) );
  INVX1 INVX1_127 ( .A(delta_16_), .Y(_abc_17692_n1327) );
  INVX1 INVX1_1270 ( .A(_abc_17692_n6730), .Y(_abc_17692_n6741) );
  INVX1 INVX1_1271 ( .A(_abc_17692_n6738), .Y(_abc_17692_n6743) );
  INVX1 INVX1_1272 ( .A(_abc_17692_n6746), .Y(_abc_17692_n6747) );
  INVX1 INVX1_1273 ( .A(_abc_17692_n6750), .Y(_abc_17692_n6751) );
  INVX1 INVX1_1274 ( .A(_abc_17692_n6754), .Y(_abc_17692_n6755) );
  INVX1 INVX1_1275 ( .A(_abc_17692_n6757), .Y(_abc_17692_n6758) );
  INVX1 INVX1_1276 ( .A(_abc_17692_n6765), .Y(_abc_17692_n6766) );
  INVX1 INVX1_1277 ( .A(_abc_17692_n6768), .Y(_abc_17692_n6769) );
  INVX1 INVX1_1278 ( .A(_abc_17692_n6771), .Y(_abc_17692_n6772) );
  INVX1 INVX1_1279 ( .A(_abc_17692_n6775), .Y(_abc_17692_n6776) );
  INVX1 INVX1_128 ( .A(sum_16_), .Y(_abc_17692_n1328) );
  INVX1 INVX1_1280 ( .A(_abc_17692_n6780), .Y(_abc_17692_n6781) );
  INVX1 INVX1_1281 ( .A(_abc_17692_n6785), .Y(_abc_17692_n6786) );
  INVX1 INVX1_1282 ( .A(_abc_17692_n6787), .Y(_abc_17692_n6788) );
  INVX1 INVX1_1283 ( .A(_abc_17692_n6778), .Y(_abc_17692_n6790) );
  INVX1 INVX1_1284 ( .A(_abc_17692_n6792), .Y(_abc_17692_n6793) );
  INVX1 INVX1_1285 ( .A(_abc_17692_n6796), .Y(_abc_17692_n6797) );
  INVX1 INVX1_1286 ( .A(_abc_17692_n6802), .Y(_abc_17692_n6804) );
  INVX1 INVX1_1287 ( .A(_abc_17692_n6806), .Y(_abc_17692_n6807) );
  INVX1 INVX1_1288 ( .A(_abc_17692_n6810), .Y(_abc_17692_n6811) );
  INVX1 INVX1_1289 ( .A(_abc_17692_n6813), .Y(_abc_17692_n6814) );
  INVX1 INVX1_129 ( .A(_abc_17692_n1330), .Y(_abc_17692_n1331_1) );
  INVX1 INVX1_1290 ( .A(_abc_17692_n6816), .Y(_abc_17692_n6817) );
  INVX1 INVX1_1291 ( .A(_abc_17692_n6821), .Y(_abc_17692_n6822) );
  INVX1 INVX1_1292 ( .A(_abc_17692_n6826), .Y(_abc_17692_n6827) );
  INVX1 INVX1_1293 ( .A(_abc_17692_n6828), .Y(_abc_17692_n6829) );
  INVX1 INVX1_1294 ( .A(_abc_17692_n6824), .Y(_abc_17692_n6835) );
  INVX1 INVX1_1295 ( .A(_abc_17692_n6832), .Y(_abc_17692_n6837) );
  INVX1 INVX1_1296 ( .A(_abc_17692_n6840), .Y(_abc_17692_n6841) );
  INVX1 INVX1_1297 ( .A(_abc_17692_n6844), .Y(_abc_17692_n6845) );
  INVX1 INVX1_1298 ( .A(_abc_17692_n6848), .Y(_abc_17692_n6849) );
  INVX1 INVX1_1299 ( .A(_abc_17692_n6855), .Y(_abc_17692_n6856) );
  INVX1 INVX1_13 ( .A(state_4_), .Y(_abc_17692_n699) );
  INVX1 INVX1_130 ( .A(_abc_17692_n1332), .Y(_abc_17692_n1333) );
  INVX1 INVX1_1300 ( .A(_abc_17692_n6861), .Y(_abc_17692_n6862) );
  INVX1 INVX1_1301 ( .A(_abc_17692_n6863), .Y(_abc_17692_n6864) );
  INVX1 INVX1_1302 ( .A(_abc_17692_n6412), .Y(_abc_17692_n6877) );
  INVX1 INVX1_1303 ( .A(_abc_17692_n6881), .Y(_abc_17692_n6882) );
  INVX1 INVX1_1304 ( .A(_abc_17692_n6888), .Y(_abc_17692_n6889) );
  INVX1 INVX1_1305 ( .A(_abc_17692_n6509), .Y(_abc_17692_n6897) );
  INVX1 INVX1_1306 ( .A(_abc_17692_n6899), .Y(_abc_17692_n6900) );
  INVX1 INVX1_1307 ( .A(_abc_17692_n6800), .Y(_abc_17692_n6905) );
  INVX1 INVX1_1308 ( .A(_abc_17692_n6903), .Y(_abc_17692_n6906) );
  INVX1 INVX1_1309 ( .A(_abc_17692_n6535), .Y(_abc_17692_n6914) );
  INVX1 INVX1_131 ( .A(_abc_17692_n1337), .Y(_abc_17692_n1338) );
  INVX1 INVX1_1310 ( .A(_abc_17692_n6922), .Y(_abc_17692_n6923) );
  INVX1 INVX1_1311 ( .A(_abc_17692_n6566), .Y(_abc_17692_n6930) );
  INVX1 INVX1_1312 ( .A(_abc_17692_n6938), .Y(_abc_17692_n6939) );
  INVX1 INVX1_1313 ( .A(_abc_17692_n6953), .Y(_abc_17692_n6954) );
  INVX1 INVX1_1314 ( .A(_abc_17692_n6958), .Y(_abc_17692_n6959) );
  INVX1 INVX1_1315 ( .A(_abc_17692_n6960), .Y(_abc_17692_n6961) );
  INVX1 INVX1_1316 ( .A(_abc_17692_n6962), .Y(_abc_17692_n6963) );
  INVX1 INVX1_1317 ( .A(_abc_17692_n6965), .Y(_abc_17692_n6966) );
  INVX1 INVX1_1318 ( .A(_abc_17692_n6969), .Y(_abc_17692_n6970) );
  INVX1 INVX1_1319 ( .A(_abc_17692_n6971), .Y(_abc_17692_n6972) );
  INVX1 INVX1_132 ( .A(_abc_17692_n1341), .Y(_abc_17692_n1342) );
  INVX1 INVX1_1320 ( .A(_abc_17692_n6976), .Y(_abc_17692_n6977) );
  INVX1 INVX1_1321 ( .A(_abc_17692_n6967), .Y(_abc_17692_n6980) );
  INVX1 INVX1_1322 ( .A(_abc_17692_n6975), .Y(_abc_17692_n6982) );
  INVX1 INVX1_1323 ( .A(_abc_17692_n6987), .Y(_abc_17692_n6988) );
  INVX1 INVX1_1324 ( .A(_abc_17692_n6707), .Y(_abc_17692_n6990) );
  INVX1 INVX1_1325 ( .A(_abc_17692_n6991), .Y(_abc_17692_n6992) );
  INVX1 INVX1_1326 ( .A(_abc_17692_n6989), .Y(_abc_17692_n6994) );
  INVX1 INVX1_1327 ( .A(_abc_17692_n6999), .Y(_abc_17692_n7000) );
  INVX1 INVX1_1328 ( .A(_abc_17692_n7002), .Y(_abc_17692_n7003) );
  INVX1 INVX1_1329 ( .A(_abc_17692_n7005), .Y(_abc_17692_n7006) );
  INVX1 INVX1_133 ( .A(_abc_17692_n1344), .Y(_abc_17692_n1345) );
  INVX1 INVX1_1330 ( .A(_abc_17692_n7004), .Y(_abc_17692_n7009) );
  INVX1 INVX1_1331 ( .A(_abc_17692_n7012), .Y(_abc_17692_n7014) );
  INVX1 INVX1_1332 ( .A(_abc_17692_n7016), .Y(_abc_17692_n7017) );
  INVX1 INVX1_1333 ( .A(_abc_17692_n7018), .Y(_abc_17692_n7019) );
  INVX1 INVX1_1334 ( .A(_abc_17692_n7020), .Y(_abc_17692_n7022) );
  INVX1 INVX1_1335 ( .A(_abc_17692_n7026), .Y(_abc_17692_n7027) );
  INVX1 INVX1_1336 ( .A(_abc_17692_n7028), .Y(_abc_17692_n7029) );
  INVX1 INVX1_1337 ( .A(_abc_17692_n7032), .Y(_abc_17692_n7033) );
  INVX1 INVX1_1338 ( .A(_abc_17692_n7034), .Y(_abc_17692_n7037) );
  INVX1 INVX1_1339 ( .A(_abc_17692_n7041), .Y(_abc_17692_n7042) );
  INVX1 INVX1_134 ( .A(_abc_17692_n1230), .Y(_abc_17692_n1352) );
  INVX1 INVX1_1340 ( .A(_abc_17692_n7040), .Y(_abc_17692_n7043) );
  INVX1 INVX1_1341 ( .A(_abc_17692_n7044), .Y(_abc_17692_n7045) );
  INVX1 INVX1_1342 ( .A(_abc_17692_n7046), .Y(_abc_17692_n7047) );
  INVX1 INVX1_1343 ( .A(_abc_17692_n6753), .Y(_abc_17692_n7048) );
  INVX1 INVX1_1344 ( .A(_abc_17692_n7049), .Y(_abc_17692_n7050) );
  INVX1 INVX1_1345 ( .A(_abc_17692_n7055), .Y(_abc_17692_n7056) );
  INVX1 INVX1_1346 ( .A(_abc_17692_n7057), .Y(_abc_17692_n7058) );
  INVX1 INVX1_1347 ( .A(_abc_17692_n7061), .Y(_abc_17692_n7062) );
  INVX1 INVX1_1348 ( .A(_abc_17692_n7064), .Y(_abc_17692_n7065) );
  INVX1 INVX1_1349 ( .A(_abc_17692_n7074), .Y(_abc_17692_n7075) );
  INVX1 INVX1_135 ( .A(_abc_17692_n1355_1), .Y(_abc_17692_n1356) );
  INVX1 INVX1_1350 ( .A(_abc_17692_n6847), .Y(_abc_17692_n7076) );
  INVX1 INVX1_1351 ( .A(_abc_17692_n7077), .Y(_abc_17692_n7078) );
  INVX1 INVX1_1352 ( .A(_abc_17692_n7088), .Y(_abc_17692_n7089) );
  INVX1 INVX1_1353 ( .A(_abc_17692_n7090), .Y(_abc_17692_n7091) );
  INVX1 INVX1_1354 ( .A(_abc_17692_n6798), .Y(_abc_17692_n7096) );
  INVX1 INVX1_1355 ( .A(_abc_17692_n7097), .Y(_abc_17692_n7098) );
  INVX1 INVX1_1356 ( .A(_abc_17692_n7103), .Y(_abc_17692_n7104) );
  INVX1 INVX1_1357 ( .A(_abc_17692_n7105), .Y(_abc_17692_n7106) );
  INVX1 INVX1_1358 ( .A(_abc_17692_n7111), .Y(_abc_17692_n7112) );
  INVX1 INVX1_1359 ( .A(_abc_17692_n7113), .Y(_abc_17692_n7115) );
  INVX1 INVX1_136 ( .A(_abc_17692_n1360), .Y(_abc_17692_n1361) );
  INVX1 INVX1_1360 ( .A(workunit1_31_), .Y(_abc_17692_n7135) );
  INVX1 INVX1_1361 ( .A(_abc_17692_n7137), .Y(_abc_17692_n7138) );
  INVX1 INVX1_1362 ( .A(_abc_17692_n7141), .Y(_abc_17692_n7142) );
  INVX1 INVX1_1363 ( .A(_abc_17692_n7129), .Y(_abc_17692_n7144) );
  INVX1 INVX1_1364 ( .A(_abc_17692_n7132), .Y(_abc_17692_n7146) );
  INVX1 INVX1_1365 ( .A(_abc_17692_n7149), .Y(_abc_17692_n7150) );
  INVX1 INVX1_1366 ( .A(_abc_17692_n7156), .Y(_abc_17692_n7157) );
  INVX1 INVX1_1367 ( .A(_abc_17692_n7152), .Y(_abc_17692_n7161) );
  INVX1 INVX1_1368 ( .A(_abc_17692_n7154), .Y(_abc_17692_n7162) );
  INVX1 INVX1_1369 ( .A(_abc_17692_n7159), .Y(_abc_17692_n7164) );
  INVX1 INVX1_137 ( .A(_abc_17692_n1369), .Y(_abc_17692_n1370) );
  INVX1 INVX1_1370 ( .A(_abc_17692_n7166), .Y(_abc_17692_n7168) );
  INVX1 INVX1_1371 ( .A(_abc_17692_n7170), .Y(_abc_17692_n7171) );
  INVX1 INVX1_1372 ( .A(_abc_17692_n7174), .Y(_abc_17692_n7175) );
  INVX1 INVX1_1373 ( .A(_abc_17692_n7176), .Y(_abc_17692_n7177) );
  INVX1 INVX1_1374 ( .A(_abc_17692_n7179), .Y(_abc_17692_n7180) );
  INVX1 INVX1_1375 ( .A(_abc_17692_n7181), .Y(_abc_17692_n7182) );
  INVX1 INVX1_1376 ( .A(_abc_17692_n7186), .Y(_abc_17692_n7187) );
  INVX1 INVX1_1377 ( .A(_abc_17692_n7190), .Y(_abc_17692_n7191) );
  INVX1 INVX1_1378 ( .A(_abc_17692_n7194), .Y(_abc_17692_n7195) );
  INVX1 INVX1_1379 ( .A(_abc_17692_n7196), .Y(_abc_17692_n7197) );
  INVX1 INVX1_138 ( .A(delta_17_), .Y(_abc_17692_n1371) );
  INVX1 INVX1_1380 ( .A(_abc_17692_n7198), .Y(_abc_17692_n7199) );
  INVX1 INVX1_1381 ( .A(_abc_17692_n7201), .Y(_abc_17692_n7203) );
  INVX1 INVX1_1382 ( .A(_abc_17692_n7205), .Y(_abc_17692_n7206) );
  INVX1 INVX1_1383 ( .A(_abc_17692_n7210), .Y(_abc_17692_n7211) );
  INVX1 INVX1_1384 ( .A(_abc_17692_n7220), .Y(_abc_17692_n7221) );
  INVX1 INVX1_1385 ( .A(_abc_17692_n7230), .Y(_abc_17692_n7231) );
  INVX1 INVX1_1386 ( .A(_abc_17692_n7234), .Y(_abc_17692_n7235) );
  INVX1 INVX1_1387 ( .A(_abc_17692_n7237), .Y(_abc_17692_n7239) );
  INVX1 INVX1_1388 ( .A(_abc_17692_n7241), .Y(_abc_17692_n7243) );
  INVX1 INVX1_1389 ( .A(_abc_17692_n7245), .Y(_abc_17692_n7246) );
  INVX1 INVX1_139 ( .A(sum_17_), .Y(_abc_17692_n1372) );
  INVX1 INVX1_1390 ( .A(_abc_17692_n7247), .Y(_abc_17692_n7248) );
  INVX1 INVX1_1391 ( .A(_abc_17692_n7253), .Y(_abc_17692_n7254) );
  INVX1 INVX1_1392 ( .A(_abc_17692_n7267), .Y(_abc_17692_n7268) );
  INVX1 INVX1_1393 ( .A(_abc_17692_n7271), .Y(_abc_17692_n7272) );
  INVX1 INVX1_1394 ( .A(_abc_17692_n7274), .Y(_abc_17692_n7276) );
  INVX1 INVX1_1395 ( .A(_abc_17692_n7278), .Y(_abc_17692_n7280) );
  INVX1 INVX1_1396 ( .A(_abc_17692_n7285), .Y(_abc_17692_n7286) );
  INVX1 INVX1_1397 ( .A(_abc_17692_n7287), .Y(_abc_17692_n7288) );
  INVX1 INVX1_1398 ( .A(_abc_17692_n7282), .Y(_abc_17692_n7292) );
  INVX1 INVX1_1399 ( .A(_abc_17692_n7290), .Y(_abc_17692_n7293) );
  INVX1 INVX1_14 ( .A(x_5_), .Y(_abc_17692_n700) );
  INVX1 INVX1_140 ( .A(_abc_17692_n1373), .Y(_abc_17692_n1374) );
  INVX1 INVX1_1400 ( .A(_abc_17692_n7300), .Y(_abc_17692_n7301) );
  INVX1 INVX1_1401 ( .A(_abc_17692_n7305), .Y(_abc_17692_n7306) );
  INVX1 INVX1_1402 ( .A(_abc_17692_n7213), .Y(_abc_17692_n7310) );
  INVX1 INVX1_1403 ( .A(_abc_17692_n7311), .Y(_abc_17692_n7312) );
  INVX1 INVX1_1404 ( .A(_abc_17692_n7313), .Y(_abc_17692_n7314) );
  INVX1 INVX1_1405 ( .A(_abc_17692_n7315), .Y(_abc_17692_n7316) );
  INVX1 INVX1_1406 ( .A(_abc_17692_n7319), .Y(_abc_17692_n7320) );
  INVX1 INVX1_1407 ( .A(_abc_17692_n7069), .Y(_abc_17692_n7324) );
  INVX1 INVX1_1408 ( .A(_abc_17692_n7330), .Y(_abc_17692_n7331) );
  INVX1 INVX1_1409 ( .A(_abc_17692_n7340), .Y(_abc_17692_n7341) );
  INVX1 INVX1_141 ( .A(_abc_17692_n1326), .Y(_abc_17692_n1376) );
  INVX1 INVX1_1410 ( .A(_abc_17692_n7139), .Y(_abc_17692_n7354) );
  INVX1 INVX1_1411 ( .A(_abc_17692_n7359), .Y(_abc_17692_n7360) );
  INVX1 INVX1_1412 ( .A(_abc_17692_n7366), .Y(_abc_17692_n7367) );
  INVX1 INVX1_1413 ( .A(_abc_17692_n7369), .Y(_abc_17692_n7370) );
  INVX1 INVX1_1414 ( .A(_abc_17692_n7372), .Y(_abc_17692_n7373) );
  INVX1 INVX1_1415 ( .A(_abc_17692_n7365), .Y(_abc_17692_n7379) );
  INVX1 INVX1_1416 ( .A(_abc_17692_n7279), .Y(_abc_17692_n7391) );
  INVX1 INVX1_1417 ( .A(_abc_17692_n7392), .Y(_abc_17692_n7393) );
  INVX1 INVX1_1418 ( .A(_abc_17692_n7403), .Y(_abc_17692_n7404) );
  INVX1 INVX1_1419 ( .A(_abc_17692_n7407), .Y(_abc_17692_n7408) );
  INVX1 INVX1_142 ( .A(_abc_17692_n1377), .Y(_abc_17692_n1378) );
  INVX1 INVX1_1420 ( .A(_abc_17692_n7402), .Y(_abc_17692_n7412) );
  INVX1 INVX1_1421 ( .A(_abc_17692_n7406), .Y(_abc_17692_n7413) );
  INVX1 INVX1_1422 ( .A(_abc_17692_n7423), .Y(_abc_17692_n7424) );
  INVX1 INVX1_1423 ( .A(_abc_17692_n7209), .Y(_abc_17692_n7425) );
  INVX1 INVX1_1424 ( .A(_abc_17692_n7426), .Y(_abc_17692_n7427) );
  INVX1 INVX1_1425 ( .A(_abc_17692_n7428), .Y(_abc_17692_n7429) );
  INVX1 INVX1_1426 ( .A(_abc_17692_n7435), .Y(_abc_17692_n7436) );
  INVX1 INVX1_1427 ( .A(_abc_17692_n7438), .Y(_abc_17692_n7441) );
  INVX1 INVX1_1428 ( .A(_abc_17692_n7442), .Y(_abc_17692_n7446) );
  INVX1 INVX1_1429 ( .A(_abc_17692_n7456), .Y(_abc_17692_n7457) );
  INVX1 INVX1_143 ( .A(_abc_17692_n1375), .Y(_abc_17692_n1380) );
  INVX1 INVX1_1430 ( .A(_abc_17692_n7455), .Y(_abc_17692_n7459) );
  INVX1 INVX1_1431 ( .A(_abc_17692_n7160), .Y(_abc_17692_n7463) );
  INVX1 INVX1_1432 ( .A(_abc_17692_n7465), .Y(_abc_17692_n7466) );
  INVX1 INVX1_1433 ( .A(_abc_17692_n7468), .Y(_abc_17692_n7471) );
  INVX1 INVX1_1434 ( .A(_abc_17692_n7472), .Y(_abc_17692_n7476) );
  INVX1 INVX1_1435 ( .A(_abc_17692_n7485), .Y(_abc_17692_n7486) );
  INVX1 INVX1_1436 ( .A(_abc_17692_n7487), .Y(_abc_17692_n7489) );
  INVX1 INVX1_1437 ( .A(_abc_17692_n7498), .Y(_abc_17692_n7499) );
  INVX1 INVX1_1438 ( .A(_abc_17692_n7504), .Y(_abc_17692_n7505) );
  INVX1 INVX1_1439 ( .A(_abc_17692_n7511), .Y(_abc_17692_n7512) );
  INVX1 INVX1_144 ( .A(_abc_17692_n1387), .Y(_abc_17692_n1388) );
  INVX1 INVX1_1440 ( .A(_abc_17692_n7517), .Y(_abc_17692_n7518) );
  INVX1 INVX1_1441 ( .A(_abc_17692_n7519), .Y(_abc_17692_n7520) );
  INVX1 INVX1_1442 ( .A(_abc_17692_n7545), .Y(_abc_17692_n7546) );
  INVX1 INVX1_1443 ( .A(_abc_17692_n7547), .Y(_abc_17692_n7548) );
  INVX1 INVX1_1444 ( .A(_abc_17692_n7551), .Y(_abc_17692_n7552) );
  INVX1 INVX1_1445 ( .A(_abc_17692_n7555), .Y(_abc_17692_n7556) );
  INVX1 INVX1_1446 ( .A(_abc_17692_n7554), .Y(_abc_17692_n7560) );
  INVX1 INVX1_1447 ( .A(_abc_17692_n7558), .Y(_abc_17692_n7561) );
  INVX1 INVX1_1448 ( .A(_abc_17692_n7550), .Y(_abc_17692_n7565) );
  INVX1 INVX1_1449 ( .A(_abc_17692_n7563), .Y(_abc_17692_n7566) );
  INVX1 INVX1_145 ( .A(_abc_17692_n1389_1), .Y(_abc_17692_n1390) );
  INVX1 INVX1_1450 ( .A(_abc_17692_n7568), .Y(_abc_17692_n7570) );
  INVX1 INVX1_1451 ( .A(_abc_17692_n7574), .Y(_abc_17692_n7575) );
  INVX1 INVX1_1452 ( .A(_abc_17692_n7577), .Y(_abc_17692_n7578) );
  INVX1 INVX1_1453 ( .A(_abc_17692_n7579), .Y(_abc_17692_n7580) );
  INVX1 INVX1_1454 ( .A(_abc_17692_n7584), .Y(_abc_17692_n7585) );
  INVX1 INVX1_1455 ( .A(_abc_17692_n7572), .Y(_abc_17692_n7587) );
  INVX1 INVX1_1456 ( .A(_abc_17692_n7591), .Y(_abc_17692_n7592) );
  INVX1 INVX1_1457 ( .A(_abc_17692_n7595), .Y(_abc_17692_n7596) );
  INVX1 INVX1_1458 ( .A(_abc_17692_n7594), .Y(_abc_17692_n7600) );
  INVX1 INVX1_1459 ( .A(_abc_17692_n7598), .Y(_abc_17692_n7601) );
  INVX1 INVX1_146 ( .A(delta_18_), .Y(_abc_17692_n1399) );
  INVX1 INVX1_1460 ( .A(_abc_17692_n7603), .Y(_abc_17692_n7605) );
  INVX1 INVX1_1461 ( .A(_abc_17692_n7607), .Y(_abc_17692_n7608) );
  INVX1 INVX1_1462 ( .A(_abc_17692_n7611), .Y(_abc_17692_n7612) );
  INVX1 INVX1_1463 ( .A(_abc_17692_n7614), .Y(_abc_17692_n7615) );
  INVX1 INVX1_1464 ( .A(_abc_17692_n7613), .Y(_abc_17692_n7617) );
  INVX1 INVX1_1465 ( .A(_abc_17692_n7621), .Y(_abc_17692_n7622) );
  INVX1 INVX1_1466 ( .A(_abc_17692_n7624), .Y(_abc_17692_n7625) );
  INVX1 INVX1_1467 ( .A(_abc_17692_n7627), .Y(_abc_17692_n7628) );
  INVX1 INVX1_1468 ( .A(_abc_17692_n7631), .Y(_abc_17692_n7632) );
  INVX1 INVX1_1469 ( .A(_abc_17692_n7405), .Y(_abc_17692_n7635) );
  INVX1 INVX1_147 ( .A(sum_18_), .Y(_abc_17692_n1400) );
  INVX1 INVX1_1470 ( .A(_abc_17692_n7638), .Y(_abc_17692_n7639) );
  INVX1 INVX1_1471 ( .A(_abc_17692_n7634), .Y(_abc_17692_n7641) );
  INVX1 INVX1_1472 ( .A(_abc_17692_n7643), .Y(_abc_17692_n7644) );
  INVX1 INVX1_1473 ( .A(_abc_17692_n7648), .Y(_abc_17692_n7649) );
  INVX1 INVX1_1474 ( .A(_abc_17692_n7217), .Y(_abc_17692_n7652) );
  INVX1 INVX1_1475 ( .A(_abc_17692_n7654), .Y(_abc_17692_n7655) );
  INVX1 INVX1_1476 ( .A(_abc_17692_n7216), .Y(_abc_17692_n7657) );
  INVX1 INVX1_1477 ( .A(_abc_17692_n7661), .Y(_abc_17692_n7662) );
  INVX1 INVX1_1478 ( .A(_abc_17692_n7663), .Y(_abc_17692_n7664) );
  INVX1 INVX1_1479 ( .A(_abc_17692_n7666), .Y(_abc_17692_n7667) );
  INVX1 INVX1_148 ( .A(_abc_17692_n1402), .Y(_abc_17692_n1403_1) );
  INVX1 INVX1_1480 ( .A(_abc_17692_n7671), .Y(_abc_17692_n7672) );
  INVX1 INVX1_1481 ( .A(_abc_17692_n7675), .Y(_abc_17692_n7676) );
  INVX1 INVX1_1482 ( .A(_abc_17692_n7674), .Y(_abc_17692_n7680) );
  INVX1 INVX1_1483 ( .A(_abc_17692_n7678), .Y(_abc_17692_n7681) );
  INVX1 INVX1_1484 ( .A(_abc_17692_n7683), .Y(_abc_17692_n7685) );
  INVX1 INVX1_1485 ( .A(_abc_17692_n7687), .Y(_abc_17692_n7688) );
  INVX1 INVX1_1486 ( .A(_abc_17692_n7691), .Y(_abc_17692_n7692) );
  INVX1 INVX1_1487 ( .A(_abc_17692_n7697), .Y(_abc_17692_n7698) );
  INVX1 INVX1_1488 ( .A(_abc_17692_n7702), .Y(_abc_17692_n7703) );
  INVX1 INVX1_1489 ( .A(_abc_17692_n7704), .Y(_abc_17692_n7705) );
  INVX1 INVX1_149 ( .A(_abc_17692_n1404), .Y(_abc_17692_n1405) );
  INVX1 INVX1_1490 ( .A(_abc_17692_n7723), .Y(_abc_17692_n7724) );
  INVX1 INVX1_1491 ( .A(_abc_17692_n7651), .Y(_abc_17692_n7727) );
  INVX1 INVX1_1492 ( .A(_abc_17692_n7422), .Y(_abc_17692_n7732) );
  INVX1 INVX1_1493 ( .A(_abc_17692_n7734), .Y(_abc_17692_n7735) );
  INVX1 INVX1_1494 ( .A(_abc_17692_n7737), .Y(_abc_17692_n7738) );
  INVX1 INVX1_1495 ( .A(_abc_17692_n7739), .Y(_abc_17692_n7740) );
  INVX1 INVX1_1496 ( .A(_abc_17692_n7242), .Y(_abc_17692_n7748) );
  INVX1 INVX1_1497 ( .A(_abc_17692_n7450), .Y(_abc_17692_n7749) );
  INVX1 INVX1_1498 ( .A(_abc_17692_n7755), .Y(_abc_17692_n7756) );
  INVX1 INVX1_1499 ( .A(_abc_17692_n7480), .Y(_abc_17692_n7763) );
  INVX1 INVX1_15 ( .A(x_6_), .Y(_abc_17692_n701) );
  INVX1 INVX1_150 ( .A(_abc_17692_n1409), .Y(_abc_17692_n1410) );
  INVX1 INVX1_1500 ( .A(_abc_17692_n7172), .Y(_abc_17692_n7764) );
  INVX1 INVX1_1501 ( .A(_abc_17692_n7769), .Y(_abc_17692_n7770) );
  INVX1 INVX1_1502 ( .A(_abc_17692_n7784), .Y(_abc_17692_n7785) );
  INVX1 INVX1_1503 ( .A(_abc_17692_n7786), .Y(_abc_17692_n7787) );
  INVX1 INVX1_1504 ( .A(_abc_17692_n7790), .Y(_abc_17692_n7791) );
  INVX1 INVX1_1505 ( .A(_abc_17692_n7795), .Y(_abc_17692_n7796) );
  INVX1 INVX1_1506 ( .A(_abc_17692_n7798), .Y(_abc_17692_n7799) );
  INVX1 INVX1_1507 ( .A(_abc_17692_n7800), .Y(_abc_17692_n7801) );
  INVX1 INVX1_1508 ( .A(_abc_17692_n7794), .Y(_abc_17692_n7806) );
  INVX1 INVX1_1509 ( .A(_abc_17692_n7817), .Y(_abc_17692_n7818) );
  INVX1 INVX1_151 ( .A(_abc_17692_n1412), .Y(_abc_17692_n1413) );
  INVX1 INVX1_1510 ( .A(_abc_17692_n7819), .Y(_abc_17692_n7821) );
  INVX1 INVX1_1511 ( .A(_abc_17692_n7825), .Y(_abc_17692_n7826) );
  INVX1 INVX1_1512 ( .A(_abc_17692_n7827), .Y(_abc_17692_n7828) );
  INVX1 INVX1_1513 ( .A(_abc_17692_n7830), .Y(_abc_17692_n7831) );
  INVX1 INVX1_1514 ( .A(_abc_17692_n7833), .Y(_abc_17692_n7837) );
  INVX1 INVX1_1515 ( .A(_abc_17692_n7846), .Y(_abc_17692_n7847) );
  INVX1 INVX1_1516 ( .A(_abc_17692_n7848), .Y(_abc_17692_n7849) );
  INVX1 INVX1_1517 ( .A(_abc_17692_n7850), .Y(_abc_17692_n7851) );
  INVX1 INVX1_1518 ( .A(_abc_17692_n7856), .Y(_abc_17692_n7857) );
  INVX1 INVX1_1519 ( .A(_abc_17692_n7858), .Y(_abc_17692_n7859) );
  INVX1 INVX1_152 ( .A(_abc_17692_n1416), .Y(_abc_17692_n1417) );
  INVX1 INVX1_1520 ( .A(_abc_17692_n7861), .Y(_abc_17692_n7862) );
  INVX1 INVX1_1521 ( .A(_abc_17692_n7864), .Y(_abc_17692_n7868) );
  INVX1 INVX1_1522 ( .A(_abc_17692_n7878), .Y(_abc_17692_n7879) );
  INVX1 INVX1_1523 ( .A(_abc_17692_n7877), .Y(_abc_17692_n7882) );
  INVX1 INVX1_1524 ( .A(_abc_17692_n7880), .Y(_abc_17692_n7883) );
  INVX1 INVX1_1525 ( .A(_abc_17692_n7891), .Y(_abc_17692_n7892) );
  INVX1 INVX1_1526 ( .A(_abc_17692_n7895), .Y(_abc_17692_n7896) );
  INVX1 INVX1_1527 ( .A(_abc_17692_n7897), .Y(_abc_17692_n7900) );
  INVX1 INVX1_1528 ( .A(_abc_17692_n7910), .Y(_abc_17692_n7911) );
  INVX1 INVX1_1529 ( .A(_abc_17692_n7647), .Y(_abc_17692_n7921) );
  INVX1 INVX1_153 ( .A(_abc_17692_n1419), .Y(_abc_17692_n1420) );
  INVX1 INVX1_1530 ( .A(_abc_17692_n7923), .Y(_abc_17692_n7925) );
  INVX1 INVX1_1531 ( .A(_abc_17692_n7929), .Y(_abc_17692_n7930) );
  INVX1 INVX1_1532 ( .A(_abc_17692_n7931), .Y(_abc_17692_n7932) );
  INVX1 INVX1_1533 ( .A(_abc_17692_n7609), .Y(_abc_17692_n7937) );
  INVX1 INVX1_1534 ( .A(_abc_17692_n7938), .Y(_abc_17692_n7939) );
  INVX1 INVX1_1535 ( .A(_abc_17692_n7689), .Y(_abc_17692_n7944) );
  INVX1 INVX1_1536 ( .A(_abc_17692_n7945), .Y(_abc_17692_n7946) );
  INVX1 INVX1_1537 ( .A(_abc_17692_n7964), .Y(_abc_17692_n7965) );
  INVX1 INVX1_1538 ( .A(_abc_17692_n7966), .Y(_abc_17692_n7967) );
  INVX1 INVX1_1539 ( .A(_abc_17692_n7971), .Y(_abc_17692_n7972) );
  INVX1 INVX1_154 ( .A(_abc_17692_n1421_1), .Y(_abc_17692_n1422) );
  INVX1 INVX1_1540 ( .A(_abc_17692_n7975), .Y(_abc_17692_n7976) );
  INVX1 INVX1_1541 ( .A(_abc_17692_n7979), .Y(_abc_17692_n7980) );
  INVX1 INVX1_1542 ( .A(_abc_17692_n7982), .Y(_abc_17692_n7983) );
  INVX1 INVX1_1543 ( .A(_abc_17692_n7829), .Y(_abc_17692_n7984) );
  INVX1 INVX1_1544 ( .A(_abc_17692_n7987), .Y(_abc_17692_n7988) );
  INVX1 INVX1_1545 ( .A(_abc_17692_n7991), .Y(_abc_17692_n7992) );
  INVX1 INVX1_1546 ( .A(_abc_17692_n7993), .Y(_abc_17692_n7996) );
  INVX1 INVX1_1547 ( .A(_abc_17692_n7999), .Y(_abc_17692_n8000) );
  INVX1 INVX1_1548 ( .A(_abc_17692_n7978), .Y(_abc_17692_n8011) );
  INVX1 INVX1_1549 ( .A(_abc_17692_n8012), .Y(_abc_17692_n8013) );
  INVX1 INVX1_155 ( .A(_abc_17692_n1430), .Y(_abc_17692_n1431) );
  INVX1 INVX1_1550 ( .A(_abc_17692_n8015), .Y(_abc_17692_n8016) );
  INVX1 INVX1_1551 ( .A(_abc_17692_n7797), .Y(_abc_17692_n8017) );
  INVX1 INVX1_1552 ( .A(_abc_17692_n8020), .Y(_abc_17692_n8021) );
  INVX1 INVX1_1553 ( .A(_abc_17692_n8023), .Y(_abc_17692_n8024) );
  INVX1 INVX1_1554 ( .A(_abc_17692_n8027), .Y(_abc_17692_n8029) );
  INVX1 INVX1_1555 ( .A(_abc_17692_n8033), .Y(_abc_17692_n8034) );
  INVX1 INVX1_1556 ( .A(_abc_17692_n8039), .Y(_abc_17692_n8040) );
  INVX1 INVX1_1557 ( .A(_abc_17692_n8043), .Y(_abc_17692_n8044) );
  INVX1 INVX1_1558 ( .A(_abc_17692_n8045), .Y(_abc_17692_n8046) );
  INVX1 INVX1_1559 ( .A(_abc_17692_n8048), .Y(_abc_17692_n8049) );
  INVX1 INVX1_156 ( .A(delta_19_), .Y(_abc_17692_n1432) );
  INVX1 INVX1_1560 ( .A(_abc_17692_n7860), .Y(_abc_17692_n8050) );
  INVX1 INVX1_1561 ( .A(_abc_17692_n8053), .Y(_abc_17692_n8054) );
  INVX1 INVX1_1562 ( .A(_abc_17692_n8066), .Y(_abc_17692_n8067) );
  INVX1 INVX1_1563 ( .A(_abc_17692_n8075), .Y(_abc_17692_n8076) );
  INVX1 INVX1_1564 ( .A(_abc_17692_n8078), .Y(_abc_17692_n8079) );
  INVX1 INVX1_1565 ( .A(_abc_17692_n8082), .Y(_abc_17692_n8083) );
  INVX1 INVX1_1566 ( .A(_abc_17692_n8084), .Y(_abc_17692_n8085) );
  INVX1 INVX1_1567 ( .A(_abc_17692_n8087), .Y(_abc_17692_n8088) );
  INVX1 INVX1_1568 ( .A(_abc_17692_n8090), .Y(_abc_17692_n8091) );
  INVX1 INVX1_1569 ( .A(_abc_17692_n8094), .Y(_abc_17692_n8096) );
  INVX1 INVX1_157 ( .A(sum_19_), .Y(_abc_17692_n1433) );
  INVX1 INVX1_1570 ( .A(_abc_17692_n8098), .Y(_abc_17692_n8099) );
  INVX1 INVX1_1571 ( .A(_abc_17692_n8115), .Y(_abc_17692_n8116) );
  INVX1 INVX1_1572 ( .A(_abc_17692_n6876), .Y(_abc_17692_n8119) );
  INVX1 INVX1_1573 ( .A(_abc_17692_n6879), .Y(_abc_17692_n8120) );
  INVX1 INVX1_1574 ( .A(_abc_17692_n5139), .Y(_abc_17692_n8123) );
  INVX1 INVX1_1575 ( .A(_abc_17692_n5990), .Y(_abc_17692_n8124) );
  INVX1 INVX1_1576 ( .A(_abc_17692_n6873), .Y(_abc_17692_n8125) );
  INVX1 INVX1_1577 ( .A(_abc_17692_n7302), .Y(_abc_17692_n8131) );
  INVX1 INVX1_1578 ( .A(_abc_17692_n7719), .Y(_abc_17692_n8136) );
  INVX1 INVX1_1579 ( .A(_abc_17692_n8031), .Y(_abc_17692_n8145) );
  INVX1 INVX1_158 ( .A(_abc_17692_n1434), .Y(_abc_17692_n1435) );
  INVX1 INVX1_1580 ( .A(_abc_17692_n7816), .Y(_abc_17692_n8148) );
  INVX1 INVX1_1581 ( .A(_abc_17692_n8150), .Y(_abc_17692_n8151) );
  INVX1 INVX1_1582 ( .A(_abc_17692_n8152), .Y(_abc_17692_n8153) );
  INVX1 INVX1_1583 ( .A(_abc_17692_n7872), .Y(_abc_17692_n8160) );
  INVX1 INVX1_1584 ( .A(_abc_17692_n8164), .Y(_abc_17692_n8165) );
  INVX1 INVX1_1585 ( .A(_abc_17692_n7841), .Y(_abc_17692_n8171) );
  INVX1 INVX1_1586 ( .A(_abc_17692_n8175), .Y(_abc_17692_n8176) );
  INVX1 INVX1_1587 ( .A(_abc_17692_n8189), .Y(_abc_17692_n8190) );
  INVX1 INVX1_1588 ( .A(_abc_17692_n8093), .Y(_abc_17692_n8191) );
  INVX1 INVX1_1589 ( .A(\key_in[127] ), .Y(_abc_17692_n8194) );
  INVX1 INVX1_159 ( .A(_abc_17692_n1436), .Y(_abc_17692_n1437) );
  INVX1 INVX1_1590 ( .A(_abc_17692_n8196), .Y(_abc_17692_n8197) );
  INVX1 INVX1_1591 ( .A(_abc_17692_n8198), .Y(_abc_17692_n8199) );
  INVX1 INVX1_1592 ( .A(workunit2_31_), .Y(_abc_17692_n8202) );
  INVX1 INVX1_1593 ( .A(_abc_17692_n8203), .Y(_abc_17692_n8204) );
  INVX1 INVX1_1594 ( .A(_abc_17692_n8208), .Y(_abc_17692_n8209) );
  INVX1 INVX1_1595 ( .A(_abc_17692_n8213), .Y(_abc_17692_n8214) );
  INVX1 INVX1_1596 ( .A(_abc_17692_n8201), .Y(_abc_17692_n8217) );
  INVX1 INVX1_1597 ( .A(_abc_17692_n8220), .Y(_abc_17692_n8221) );
  INVX1 INVX1_1598 ( .A(_abc_17692_n8030), .Y(_abc_17692_n8226) );
  INVX1 INVX1_1599 ( .A(_abc_17692_n8227), .Y(_abc_17692_n8228) );
  INVX1 INVX1_16 ( .A(x_7_), .Y(_abc_17692_n702) );
  INVX1 INVX1_160 ( .A(_abc_17692_n1438), .Y(_abc_17692_n1439) );
  INVX1 INVX1_1600 ( .A(\key_in[95] ), .Y(_abc_17692_n8231) );
  INVX1 INVX1_1601 ( .A(_abc_17692_n8233), .Y(_abc_17692_n8234) );
  INVX1 INVX1_1602 ( .A(_abc_17692_n8235), .Y(_abc_17692_n8236) );
  INVX1 INVX1_1603 ( .A(_abc_17692_n8238), .Y(_abc_17692_n8240) );
  INVX1 INVX1_1604 ( .A(_abc_17692_n8242), .Y(_abc_17692_n8243) );
  INVX1 INVX1_1605 ( .A(_abc_17692_n8248), .Y(_abc_17692_n8249) );
  INVX1 INVX1_1606 ( .A(_abc_17692_n8250), .Y(_abc_17692_n8251) );
  INVX1 INVX1_1607 ( .A(\key_in[31] ), .Y(_abc_17692_n8254) );
  INVX1 INVX1_1608 ( .A(_abc_17692_n8256), .Y(_abc_17692_n8257) );
  INVX1 INVX1_1609 ( .A(_abc_17692_n8258), .Y(_abc_17692_n8259) );
  INVX1 INVX1_161 ( .A(_abc_17692_n1444), .Y(_abc_17692_n1445) );
  INVX1 INVX1_1610 ( .A(_abc_17692_n8261), .Y(_abc_17692_n8263) );
  INVX1 INVX1_1611 ( .A(_abc_17692_n8265), .Y(_abc_17692_n8266) );
  INVX1 INVX1_1612 ( .A(_abc_17692_n8271), .Y(_abc_17692_n8272) );
  INVX1 INVX1_1613 ( .A(_abc_17692_n8273), .Y(_abc_17692_n8274) );
  INVX1 INVX1_1614 ( .A(\key_in[63] ), .Y(_abc_17692_n8277) );
  INVX1 INVX1_1615 ( .A(_abc_17692_n8279), .Y(_abc_17692_n8280) );
  INVX1 INVX1_1616 ( .A(_abc_17692_n8281), .Y(_abc_17692_n8282) );
  INVX1 INVX1_1617 ( .A(_abc_17692_n8284), .Y(_abc_17692_n8286) );
  INVX1 INVX1_1618 ( .A(_abc_17692_n8288), .Y(_abc_17692_n8289) );
  INVX1 INVX1_1619 ( .A(_abc_17692_n8104), .Y(_abc_17692_n8301) );
  INVX1 INVX1_162 ( .A(_abc_17692_n1446), .Y(_abc_17692_n1447) );
  INVX1 INVX1_1620 ( .A(_abc_17692_n8307), .Y(_abc_17692_n8308) );
  INVX1 INVX1_1621 ( .A(_abc_17692_n8309), .Y(_abc_17692_n8310) );
  INVX1 INVX1_1622 ( .A(_abc_17692_n8061), .Y(_abc_17692_n8315) );
  INVX1 INVX1_1623 ( .A(_abc_17692_n8316), .Y(_abc_17692_n8317) );
  INVX1 INVX1_1624 ( .A(_abc_17692_n7995), .Y(_abc_17692_n8322) );
  INVX1 INVX1_1625 ( .A(_abc_17692_n8323), .Y(_abc_17692_n8324) );
  INVX1 INVX1_1626 ( .A(_abc_17692_n713), .Y(_abc_17692_n8338) );
  INVX1 INVX1_1627 ( .A(_abc_17692_n8341), .Y(_abc_17692_n8343) );
  INVX1 INVX1_1628 ( .A(_abc_17692_n8345), .Y(_abc_17692_n8346) );
  INVX1 INVX1_1629 ( .A(_abc_17692_n8347), .Y(_abc_17692_n8348) );
  INVX1 INVX1_163 ( .A(sum_20_), .Y(_abc_17692_n1456) );
  INVX1 INVX1_1630 ( .A(_abc_17692_n8354), .Y(_abc_17692_n8355) );
  INVX1 INVX1_1631 ( .A(_abc_17692_n8357), .Y(_abc_17692_n8358) );
  INVX1 INVX1_1632 ( .A(_abc_17692_n8364), .Y(_abc_17692_n8365) );
  INVX1 INVX1_1633 ( .A(_abc_17692_n8366), .Y(_abc_17692_n8367) );
  INVX1 INVX1_1634 ( .A(_abc_17692_n8373), .Y(_abc_17692_n8374) );
  INVX1 INVX1_1635 ( .A(_abc_17692_n8376), .Y(_abc_17692_n8377) );
  INVX1 INVX1_1636 ( .A(_abc_17692_n8388), .Y(_abc_17692_n8389) );
  INVX1 INVX1_1637 ( .A(_abc_17692_n8390), .Y(_abc_17692_n8391) );
  INVX1 INVX1_1638 ( .A(_abc_17692_n8339), .Y(_abc_17692_n8395) );
  INVX1 INVX1_1639 ( .A(_abc_17692_n8406), .Y(_abc_17692_n8407) );
  INVX1 INVX1_164 ( .A(_abc_17692_n1458), .Y(_abc_17692_n1459_1) );
  INVX1 INVX1_1640 ( .A(_abc_17692_n8409), .Y(_abc_17692_n8410) );
  INVX1 INVX1_1641 ( .A(_abc_17692_n8411), .Y(_abc_17692_n8412) );
  INVX1 INVX1_1642 ( .A(_abc_17692_n8425), .Y(_abc_17692_n8426) );
  INVX1 INVX1_1643 ( .A(_abc_17692_n8428), .Y(_abc_17692_n8429) );
  INVX1 INVX1_1644 ( .A(_abc_17692_n8432), .Y(_abc_17692_n8433) );
  INVX1 INVX1_1645 ( .A(_abc_17692_n8437), .Y(_abc_17692_n8438) );
  INVX1 INVX1_1646 ( .A(_abc_17692_n8440), .Y(_abc_17692_n8441) );
  INVX1 INVX1_1647 ( .A(_abc_17692_n8448), .Y(_abc_17692_n8449) );
  INVX1 INVX1_1648 ( .A(_abc_17692_n8451), .Y(_abc_17692_n8452) );
  INVX1 INVX1_1649 ( .A(_abc_17692_n8458), .Y(_abc_17692_n8459) );
  INVX1 INVX1_165 ( .A(_abc_17692_n1461), .Y(_abc_17692_n1462) );
  INVX1 INVX1_1650 ( .A(_abc_17692_n8460), .Y(_abc_17692_n8461) );
  INVX1 INVX1_1651 ( .A(_abc_17692_n8424), .Y(_abc_17692_n8467) );
  INVX1 INVX1_1652 ( .A(_abc_17692_n8472), .Y(_abc_17692_n8473) );
  INVX1 INVX1_1653 ( .A(_abc_17692_n8478), .Y(_abc_17692_n8479) );
  INVX1 INVX1_1654 ( .A(_abc_17692_n8483), .Y(_abc_17692_n8484) );
  INVX1 INVX1_1655 ( .A(_abc_17692_n8499), .Y(_abc_17692_n8502) );
  INVX1 INVX1_1656 ( .A(_abc_17692_n8519), .Y(_abc_17692_n8520) );
  INVX1 INVX1_1657 ( .A(_abc_17692_n8524), .Y(_abc_17692_n8525) );
  INVX1 INVX1_1658 ( .A(_abc_17692_n8526), .Y(_abc_17692_n8527) );
  INVX1 INVX1_1659 ( .A(_abc_17692_n8532), .Y(_abc_17692_n8533) );
  INVX1 INVX1_166 ( .A(_abc_17692_n1465), .Y(_abc_17692_n1466) );
  INVX1 INVX1_1660 ( .A(_abc_17692_n8434), .Y(_abc_17692_n8534) );
  INVX1 INVX1_1661 ( .A(_abc_17692_n8435), .Y(_abc_17692_n8535) );
  INVX1 INVX1_1662 ( .A(_abc_17692_n8537), .Y(_abc_17692_n8538) );
  INVX1 INVX1_1663 ( .A(_abc_17692_n8539), .Y(_abc_17692_n8540) );
  INVX1 INVX1_1664 ( .A(_abc_17692_n8548), .Y(_abc_17692_n8549) );
  INVX1 INVX1_1665 ( .A(_abc_17692_n8551), .Y(_abc_17692_n8552) );
  INVX1 INVX1_1666 ( .A(_abc_17692_n8405), .Y(_abc_17692_n8553) );
  INVX1 INVX1_1667 ( .A(_abc_17692_n8556), .Y(_abc_17692_n8557) );
  INVX1 INVX1_1668 ( .A(_abc_17692_n8571), .Y(_abc_17692_n8572) );
  INVX1 INVX1_1669 ( .A(_abc_17692_n8575), .Y(_abc_17692_n8576) );
  INVX1 INVX1_167 ( .A(_abc_17692_n1469), .Y(_abc_17692_n1470) );
  INVX1 INVX1_1670 ( .A(_abc_17692_n8516), .Y(_abc_17692_n8582) );
  INVX1 INVX1_1671 ( .A(_abc_17692_n8419), .Y(_abc_17692_n8583) );
  INVX1 INVX1_1672 ( .A(_abc_17692_n8584), .Y(_abc_17692_n8585) );
  INVX1 INVX1_1673 ( .A(_abc_17692_n8591), .Y(_abc_17692_n8592) );
  INVX1 INVX1_1674 ( .A(_abc_17692_n8454), .Y(_abc_17692_n8597) );
  INVX1 INVX1_1675 ( .A(_abc_17692_n8599), .Y(_abc_17692_n8600) );
  INVX1 INVX1_1676 ( .A(_abc_17692_n8605), .Y(_abc_17692_n8606) );
  INVX1 INVX1_1677 ( .A(_abc_17692_n8497), .Y(_abc_17692_n8621) );
  INVX1 INVX1_1678 ( .A(_abc_17692_n8620), .Y(_abc_17692_n8624) );
  INVX1 INVX1_1679 ( .A(_abc_17692_n8626), .Y(_abc_17692_n8630) );
  INVX1 INVX1_168 ( .A(_abc_17692_n1472), .Y(_abc_17692_n1473) );
  INVX1 INVX1_1680 ( .A(_abc_17692_n8515), .Y(_abc_17692_n8640) );
  INVX1 INVX1_1681 ( .A(_abc_17692_n8642), .Y(_abc_17692_n8643) );
  INVX1 INVX1_1682 ( .A(_abc_17692_n8655), .Y(_abc_17692_n8656) );
  INVX1 INVX1_1683 ( .A(_abc_17692_n8657), .Y(_abc_17692_n8658) );
  INVX1 INVX1_1684 ( .A(_abc_17692_n8659), .Y(_abc_17692_n8660) );
  INVX1 INVX1_1685 ( .A(_abc_17692_n8667), .Y(_abc_17692_n8668) );
  INVX1 INVX1_1686 ( .A(_abc_17692_n8672), .Y(_abc_17692_n8673) );
  INVX1 INVX1_1687 ( .A(_abc_17692_n8675), .Y(_abc_17692_n8676) );
  INVX1 INVX1_1688 ( .A(_abc_17692_n8690), .Y(_abc_17692_n8691) );
  INVX1 INVX1_1689 ( .A(_abc_17692_n8693), .Y(_abc_17692_n8694) );
  INVX1 INVX1_169 ( .A(_abc_17692_n1460), .Y(_abc_17692_n1477) );
  INVX1 INVX1_1690 ( .A(_abc_17692_n8696), .Y(_abc_17692_n8697) );
  INVX1 INVX1_1691 ( .A(_abc_17692_n8639), .Y(_abc_17692_n8702) );
  INVX1 INVX1_1692 ( .A(_abc_17692_n8704), .Y(_abc_17692_n8705) );
  INVX1 INVX1_1693 ( .A(_abc_17692_n8714), .Y(_abc_17692_n8715) );
  INVX1 INVX1_1694 ( .A(_abc_17692_n8566), .Y(_abc_17692_n8720) );
  INVX1 INVX1_1695 ( .A(_abc_17692_n8722), .Y(_abc_17692_n8723) );
  INVX1 INVX1_1696 ( .A(_abc_17692_n8529), .Y(_abc_17692_n8727) );
  INVX1 INVX1_1697 ( .A(_abc_17692_n8729), .Y(_abc_17692_n8730) );
  INVX1 INVX1_1698 ( .A(_abc_17692_n8751), .Y(_abc_17692_n8752) );
  INVX1 INVX1_1699 ( .A(_abc_17692_n8755), .Y(_abc_17692_n8762) );
  INVX1 INVX1_17 ( .A(_abc_17692_n710), .Y(_abc_17692_n711) );
  INVX1 INVX1_170 ( .A(_abc_17692_n1418), .Y(_abc_17692_n1480) );
  INVX1 INVX1_1700 ( .A(_abc_17692_n8769), .Y(_abc_17692_n8771) );
  INVX1 INVX1_1701 ( .A(_abc_17692_n8669), .Y(_abc_17692_n8774) );
  INVX1 INVX1_1702 ( .A(_abc_17692_n8776), .Y(_abc_17692_n8777) );
  INVX1 INVX1_1703 ( .A(_abc_17692_n8783), .Y(_abc_17692_n8784) );
  INVX1 INVX1_1704 ( .A(_abc_17692_n8634), .Y(_abc_17692_n8788) );
  INVX1 INVX1_1705 ( .A(_abc_17692_n8791), .Y(_abc_17692_n8792) );
  INVX1 INVX1_1706 ( .A(_abc_17692_n8797), .Y(_abc_17692_n8799) );
  INVX1 INVX1_1707 ( .A(_abc_17692_n8802), .Y(_abc_17692_n8803) );
  INVX1 INVX1_1708 ( .A(_abc_17692_n8804), .Y(_abc_17692_n8805) );
  INVX1 INVX1_1709 ( .A(_abc_17692_n8806), .Y(_abc_17692_n8807) );
  INVX1 INVX1_171 ( .A(_abc_17692_n1487), .Y(_abc_17692_n1488) );
  INVX1 INVX1_1710 ( .A(_abc_17692_n8821), .Y(_abc_17692_n8822) );
  INVX1 INVX1_1711 ( .A(_abc_17692_n8823), .Y(_abc_17692_n8824) );
  INVX1 INVX1_1712 ( .A(_abc_17692_n8826), .Y(_abc_17692_n8827) );
  INVX1 INVX1_1713 ( .A(_abc_17692_n8787), .Y(_abc_17692_n8833) );
  INVX1 INVX1_1714 ( .A(_abc_17692_n8835), .Y(_abc_17692_n8836) );
  INVX1 INVX1_1715 ( .A(_abc_17692_n8773), .Y(_abc_17692_n8841) );
  INVX1 INVX1_1716 ( .A(_abc_17692_n8710), .Y(_abc_17692_n8842) );
  INVX1 INVX1_1717 ( .A(_abc_17692_n8844), .Y(_abc_17692_n8845) );
  INVX1 INVX1_1718 ( .A(_abc_17692_n8685), .Y(_abc_17692_n8850) );
  INVX1 INVX1_1719 ( .A(_abc_17692_n8852), .Y(_abc_17692_n8853) );
  INVX1 INVX1_172 ( .A(_abc_17692_n1494), .Y(_abc_17692_n1495) );
  INVX1 INVX1_1720 ( .A(_abc_17692_n8801), .Y(_abc_17692_n8857) );
  INVX1 INVX1_1721 ( .A(_abc_17692_n8650), .Y(_abc_17692_n8858) );
  INVX1 INVX1_1722 ( .A(_abc_17692_n8860), .Y(_abc_17692_n8861) );
  INVX1 INVX1_1723 ( .A(_abc_17692_n8875), .Y(_abc_17692_n8879) );
  INVX1 INVX1_1724 ( .A(_abc_17692_n8889), .Y(_abc_17692_n8893) );
  INVX1 INVX1_1725 ( .A(_abc_17692_n8896), .Y(_abc_17692_n8897) );
  INVX1 INVX1_1726 ( .A(_abc_17692_n8786), .Y(_abc_17692_n8901) );
  INVX1 INVX1_1727 ( .A(_abc_17692_n8903), .Y(_abc_17692_n8904) );
  INVX1 INVX1_1728 ( .A(_abc_17692_n8910), .Y(_abc_17692_n8911) );
  INVX1 INVX1_1729 ( .A(_abc_17692_n8912), .Y(_abc_17692_n8913) );
  INVX1 INVX1_173 ( .A(delta_21_), .Y(_abc_17692_n1496) );
  INVX1 INVX1_1730 ( .A(_abc_17692_n8918), .Y(_abc_17692_n8919) );
  INVX1 INVX1_1731 ( .A(_abc_17692_n8931), .Y(_abc_17692_n8932) );
  INVX1 INVX1_1732 ( .A(_abc_17692_n8936), .Y(_abc_17692_n8937) );
  INVX1 INVX1_1733 ( .A(_abc_17692_n8950), .Y(_abc_17692_n8951) );
  INVX1 INVX1_1734 ( .A(_abc_17692_n8952), .Y(_abc_17692_n8953) );
  INVX1 INVX1_1735 ( .A(_abc_17692_n8955), .Y(_abc_17692_n8956) );
  INVX1 INVX1_1736 ( .A(_abc_17692_n8900), .Y(_abc_17692_n8962) );
  INVX1 INVX1_1737 ( .A(_abc_17692_n8963), .Y(_abc_17692_n8964) );
  INVX1 INVX1_1738 ( .A(_abc_17692_n8965), .Y(_abc_17692_n8966) );
  INVX1 INVX1_1739 ( .A(_abc_17692_n8915), .Y(_abc_17692_n8971) );
  INVX1 INVX1_174 ( .A(sum_21_), .Y(_abc_17692_n1497) );
  INVX1 INVX1_1740 ( .A(_abc_17692_n8973), .Y(_abc_17692_n8974) );
  INVX1 INVX1_1741 ( .A(_abc_17692_n8816), .Y(_abc_17692_n8979) );
  INVX1 INVX1_1742 ( .A(_abc_17692_n8981), .Y(_abc_17692_n8982) );
  INVX1 INVX1_1743 ( .A(_abc_17692_n8987), .Y(_abc_17692_n8988) );
  INVX1 INVX1_1744 ( .A(_abc_17692_n9005), .Y(_abc_17692_n9006) );
  INVX1 INVX1_1745 ( .A(_abc_17692_n9024), .Y(_abc_17692_n9026) );
  INVX1 INVX1_1746 ( .A(_abc_17692_n9028), .Y(_abc_17692_n9030) );
  INVX1 INVX1_1747 ( .A(_abc_17692_n9034), .Y(_abc_17692_n9035) );
  INVX1 INVX1_1748 ( .A(_abc_17692_n9041), .Y(_abc_17692_n9043) );
  INVX1 INVX1_1749 ( .A(_abc_17692_n8898), .Y(_abc_17692_n9046) );
  INVX1 INVX1_175 ( .A(_abc_17692_n1498), .Y(_abc_17692_n1499) );
  INVX1 INVX1_1750 ( .A(_abc_17692_n9049), .Y(_abc_17692_n9050) );
  INVX1 INVX1_1751 ( .A(_abc_17692_n9055), .Y(_abc_17692_n9056) );
  INVX1 INVX1_1752 ( .A(_abc_17692_n9059), .Y(_abc_17692_n9060) );
  INVX1 INVX1_1753 ( .A(_abc_17692_n9063), .Y(_abc_17692_n9064) );
  INVX1 INVX1_1754 ( .A(_abc_17692_n8933), .Y(_abc_17692_n9065) );
  INVX1 INVX1_1755 ( .A(_abc_17692_n9068), .Y(_abc_17692_n9069) );
  INVX1 INVX1_1756 ( .A(_abc_17692_n9071), .Y(_abc_17692_n9072) );
  INVX1 INVX1_1757 ( .A(_abc_17692_n9079), .Y(_abc_17692_n9081) );
  INVX1 INVX1_1758 ( .A(_abc_17692_n9084), .Y(_abc_17692_n9085) );
  INVX1 INVX1_1759 ( .A(_abc_17692_n9088), .Y(_abc_17692_n9089) );
  INVX1 INVX1_176 ( .A(_abc_17692_n1501), .Y(_abc_17692_n1502) );
  INVX1 INVX1_1760 ( .A(_abc_17692_n9032), .Y(_abc_17692_n9094) );
  INVX1 INVX1_1761 ( .A(_abc_17692_n9095), .Y(_abc_17692_n9096) );
  INVX1 INVX1_1762 ( .A(_abc_17692_n9098), .Y(_abc_17692_n9099) );
  INVX1 INVX1_1763 ( .A(_abc_17692_n8926), .Y(_abc_17692_n9103) );
  INVX1 INVX1_1764 ( .A(_abc_17692_n9106), .Y(_abc_17692_n9107) );
  INVX1 INVX1_1765 ( .A(_abc_17692_n9083), .Y(_abc_17692_n9111) );
  INVX1 INVX1_1766 ( .A(_abc_17692_n8945), .Y(_abc_17692_n9112) );
  INVX1 INVX1_1767 ( .A(_abc_17692_n9114), .Y(_abc_17692_n9115) );
  INVX1 INVX1_1768 ( .A(_abc_17692_n9119), .Y(_abc_17692_n9120) );
  INVX1 INVX1_1769 ( .A(_abc_17692_n9045), .Y(_abc_17692_n9123) );
  INVX1 INVX1_177 ( .A(_abc_17692_n1503), .Y(_abc_17692_n1504) );
  INVX1 INVX1_1770 ( .A(_abc_17692_n9121), .Y(_abc_17692_n9124) );
  INVX1 INVX1_1771 ( .A(_abc_17692_n9138), .Y(_abc_17692_n9139) );
  INVX1 INVX1_1772 ( .A(_abc_17692_n9166), .Y(_abc_17692_n9167) );
  INVX1 INVX1_1773 ( .A(_abc_17692_n9057), .Y(_abc_17692_n9168) );
  INVX1 INVX1_1774 ( .A(_abc_17692_n9169), .Y(_abc_17692_n9170) );
  INVX1 INVX1_1775 ( .A(_abc_17692_n9177), .Y(_abc_17692_n9178) );
  INVX1 INVX1_1776 ( .A(_abc_17692_n9184), .Y(_abc_17692_n9185) );
  INVX1 INVX1_1777 ( .A(_abc_17692_n9192), .Y(_abc_17692_n9193) );
  INVX1 INVX1_1778 ( .A(_abc_17692_n9199), .Y(_abc_17692_n9200) );
  INVX1 INVX1_1779 ( .A(_abc_17692_n9201), .Y(_abc_17692_n9202) );
  INVX1 INVX1_178 ( .A(_abc_17692_n1500), .Y(_abc_17692_n1506) );
  INVX1 INVX1_1780 ( .A(_abc_17692_n9210), .Y(_abc_17692_n9211) );
  INVX1 INVX1_1781 ( .A(_abc_17692_n9214), .Y(_abc_17692_n9215) );
  INVX1 INVX1_1782 ( .A(_abc_17692_n9080), .Y(_abc_17692_n9216) );
  INVX1 INVX1_1783 ( .A(_abc_17692_n9219), .Y(_abc_17692_n9220) );
  INVX1 INVX1_1784 ( .A(_abc_17692_n9029), .Y(_abc_17692_n9225) );
  INVX1 INVX1_1785 ( .A(_abc_17692_n9194), .Y(_abc_17692_n9228) );
  INVX1 INVX1_1786 ( .A(_abc_17692_n9195), .Y(_abc_17692_n9229) );
  INVX1 INVX1_1787 ( .A(_abc_17692_n9226), .Y(_abc_17692_n9231) );
  INVX1 INVX1_1788 ( .A(_abc_17692_n9235), .Y(_abc_17692_n9236) );
  INVX1 INVX1_1789 ( .A(_abc_17692_n9237), .Y(_abc_17692_n9238) );
  INVX1 INVX1_179 ( .A(_abc_17692_n1513), .Y(_abc_17692_n1514) );
  INVX1 INVX1_1790 ( .A(_abc_17692_n9244), .Y(_abc_17692_n9245) );
  INVX1 INVX1_1791 ( .A(_abc_17692_n9248), .Y(_abc_17692_n9249) );
  INVX1 INVX1_1792 ( .A(_abc_17692_n9122), .Y(_abc_17692_n9252) );
  INVX1 INVX1_1793 ( .A(_abc_17692_n9181), .Y(_abc_17692_n9253) );
  INVX1 INVX1_1794 ( .A(_abc_17692_n9042), .Y(_abc_17692_n9257) );
  INVX1 INVX1_1795 ( .A(_abc_17692_n9275), .Y(_abc_17692_n9276) );
  INVX1 INVX1_1796 ( .A(_abc_17692_n9287), .Y(_abc_17692_n9288) );
  INVX1 INVX1_1797 ( .A(_abc_17692_n9302), .Y(_abc_17692_n9303) );
  INVX1 INVX1_1798 ( .A(_abc_17692_n9305), .Y(_abc_17692_n9306) );
  INVX1 INVX1_1799 ( .A(_abc_17692_n9307), .Y(_abc_17692_n9308) );
  INVX1 INVX1_18 ( .A(state_14_bF_buf4), .Y(_abc_17692_n712) );
  INVX1 INVX1_180 ( .A(_abc_17692_n1515), .Y(_abc_17692_n1516) );
  INVX1 INVX1_1800 ( .A(_abc_17692_n9315), .Y(_abc_17692_n9316) );
  INVX1 INVX1_1801 ( .A(_abc_17692_n9319), .Y(_abc_17692_n9320) );
  INVX1 INVX1_1802 ( .A(_abc_17692_n9324), .Y(_abc_17692_n9325) );
  INVX1 INVX1_1803 ( .A(_abc_17692_n9331), .Y(_abc_17692_n9332) );
  INVX1 INVX1_1804 ( .A(_abc_17692_n9339), .Y(_abc_17692_n9340) );
  INVX1 INVX1_1805 ( .A(_abc_17692_n9346), .Y(_abc_17692_n9347) );
  INVX1 INVX1_1806 ( .A(_abc_17692_n9351), .Y(_abc_17692_n9352) );
  INVX1 INVX1_1807 ( .A(_abc_17692_n9356), .Y(_abc_17692_n9357) );
  INVX1 INVX1_1808 ( .A(_abc_17692_n9359), .Y(_abc_17692_n9360) );
  INVX1 INVX1_1809 ( .A(_abc_17692_n9371), .Y(_abc_17692_n9372) );
  INVX1 INVX1_181 ( .A(delta_22_), .Y(_abc_17692_n1525) );
  INVX1 INVX1_1810 ( .A(_abc_17692_n9179), .Y(_abc_17692_n9375) );
  INVX1 INVX1_1811 ( .A(_abc_17692_n9377), .Y(_abc_17692_n9378) );
  INVX1 INVX1_1812 ( .A(_abc_17692_n9379), .Y(_abc_17692_n9380) );
  INVX1 INVX1_1813 ( .A(_abc_17692_n9349), .Y(_abc_17692_n9384) );
  INVX1 INVX1_1814 ( .A(_abc_17692_n9161), .Y(_abc_17692_n9385) );
  INVX1 INVX1_1815 ( .A(_abc_17692_n9392), .Y(_abc_17692_n9393) );
  INVX1 INVX1_1816 ( .A(_abc_17692_n9334), .Y(_abc_17692_n9396) );
  INVX1 INVX1_1817 ( .A(_abc_17692_n9399), .Y(_abc_17692_n9400) );
  INVX1 INVX1_1818 ( .A(_abc_17692_n9403), .Y(_abc_17692_n9404) );
  INVX1 INVX1_1819 ( .A(_abc_17692_n9318), .Y(_abc_17692_n9417) );
  INVX1 INVX1_182 ( .A(sum_22_), .Y(_abc_17692_n1526_1) );
  INVX1 INVX1_1820 ( .A(_abc_17692_n9419), .Y(_abc_17692_n9420) );
  INVX1 INVX1_1821 ( .A(_abc_17692_n9421), .Y(_abc_17692_n9422) );
  INVX1 INVX1_1822 ( .A(_abc_17692_n9423), .Y(_abc_17692_n9426) );
  INVX1 INVX1_1823 ( .A(_abc_17692_n9429), .Y(_abc_17692_n9430) );
  INVX1 INVX1_1824 ( .A(_abc_17692_n9437), .Y(_abc_17692_n9439) );
  INVX1 INVX1_1825 ( .A(_abc_17692_n9418), .Y(_abc_17692_n9443) );
  INVX1 INVX1_1826 ( .A(_abc_17692_n9441), .Y(_abc_17692_n9444) );
  INVX1 INVX1_1827 ( .A(_abc_17692_n9448), .Y(_abc_17692_n9449) );
  INVX1 INVX1_1828 ( .A(_abc_17692_n9458), .Y(_abc_17692_n9459) );
  INVX1 INVX1_1829 ( .A(_abc_17692_n9464), .Y(_abc_17692_n9465) );
  INVX1 INVX1_183 ( .A(_abc_17692_n1528), .Y(_abc_17692_n1529) );
  INVX1 INVX1_1830 ( .A(_abc_17692_n9469), .Y(_abc_17692_n9470) );
  INVX1 INVX1_1831 ( .A(_abc_17692_n9472), .Y(_abc_17692_n9473) );
  INVX1 INVX1_1832 ( .A(_abc_17692_n9484), .Y(_abc_17692_n9485) );
  INVX1 INVX1_1833 ( .A(_abc_17692_n9483), .Y(_abc_17692_n9486) );
  INVX1 INVX1_1834 ( .A(_abc_17692_n9487), .Y(_abc_17692_n9488) );
  INVX1 INVX1_1835 ( .A(_abc_17692_n9489), .Y(_abc_17692_n9490) );
  INVX1 INVX1_1836 ( .A(_abc_17692_n9480), .Y(_abc_17692_n9492) );
  INVX1 INVX1_1837 ( .A(_abc_17692_n9301), .Y(_abc_17692_n9498) );
  INVX1 INVX1_1838 ( .A(_abc_17692_n9499), .Y(_abc_17692_n9500) );
  INVX1 INVX1_1839 ( .A(_abc_17692_n9501), .Y(_abc_17692_n9502) );
  INVX1 INVX1_184 ( .A(_abc_17692_n1531), .Y(_abc_17692_n1532) );
  INVX1 INVX1_1840 ( .A(_abc_17692_n9507), .Y(_abc_17692_n9508) );
  INVX1 INVX1_1841 ( .A(_abc_17692_n9509), .Y(_abc_17692_n9510) );
  INVX1 INVX1_1842 ( .A(_abc_17692_n9330), .Y(_abc_17692_n9515) );
  INVX1 INVX1_1843 ( .A(_abc_17692_n9516), .Y(_abc_17692_n9517) );
  INVX1 INVX1_1844 ( .A(_abc_17692_n9518), .Y(_abc_17692_n9520) );
  INVX1 INVX1_1845 ( .A(_abc_17692_n9345), .Y(_abc_17692_n9524) );
  INVX1 INVX1_1846 ( .A(_abc_17692_n9525), .Y(_abc_17692_n9526) );
  INVX1 INVX1_1847 ( .A(_abc_17692_n9527), .Y(_abc_17692_n9528) );
  INVX1 INVX1_1848 ( .A(_abc_17692_n9425), .Y(_abc_17692_n9544) );
  INVX1 INVX1_1849 ( .A(_abc_17692_n9542), .Y(_abc_17692_n9559) );
  INVX1 INVX1_185 ( .A(_abc_17692_n1537), .Y(_abc_17692_n1538_1) );
  INVX1 INVX1_1850 ( .A(_abc_17692_n9428), .Y(_abc_17692_n9561) );
  INVX1 INVX1_1851 ( .A(_abc_17692_n9569), .Y(_abc_17692_n9571) );
  INVX1 INVX1_1852 ( .A(_abc_17692_n9573), .Y(_abc_17692_n9574) );
  INVX1 INVX1_1853 ( .A(_abc_17692_n9577), .Y(_abc_17692_n9578) );
  INVX1 INVX1_1854 ( .A(_abc_17692_n9581), .Y(_abc_17692_n9582) );
  INVX1 INVX1_1855 ( .A(_abc_17692_n9584), .Y(_abc_17692_n9585) );
  INVX1 INVX1_1856 ( .A(_abc_17692_n9586), .Y(_abc_17692_n9587) );
  INVX1 INVX1_1857 ( .A(_abc_17692_n9588), .Y(_abc_17692_n9589) );
  INVX1 INVX1_1858 ( .A(_abc_17692_n9595), .Y(_abc_17692_n9597) );
  INVX1 INVX1_1859 ( .A(_abc_17692_n9599), .Y(_abc_17692_n9600) );
  INVX1 INVX1_186 ( .A(_abc_17692_n1542), .Y(_abc_17692_n1543) );
  INVX1 INVX1_1860 ( .A(_abc_17692_n9607), .Y(_abc_17692_n9608) );
  INVX1 INVX1_1861 ( .A(_abc_17692_n9614), .Y(_abc_17692_n9615) );
  INVX1 INVX1_1862 ( .A(_abc_17692_n9618), .Y(_abc_17692_n9619) );
  INVX1 INVX1_1863 ( .A(_abc_17692_n9337), .Y(_abc_17692_n9620) );
  INVX1 INVX1_1864 ( .A(_abc_17692_n9621), .Y(_abc_17692_n9622) );
  INVX1 INVX1_1865 ( .A(_abc_17692_n9468), .Y(_abc_17692_n9624) );
  INVX1 INVX1_1866 ( .A(_abc_17692_n9627), .Y(_abc_17692_n9628) );
  INVX1 INVX1_1867 ( .A(_abc_17692_n9629), .Y(_abc_17692_n9630) );
  INVX1 INVX1_1868 ( .A(_abc_17692_n9631), .Y(_abc_17692_n9632) );
  INVX1 INVX1_1869 ( .A(_abc_17692_n9638), .Y(_abc_17692_n9639) );
  INVX1 INVX1_187 ( .A(_abc_17692_n1544), .Y(_abc_17692_n1545) );
  INVX1 INVX1_1870 ( .A(_abc_17692_n9642), .Y(_abc_17692_n9643) );
  INVX1 INVX1_1871 ( .A(_abc_17692_n9646), .Y(_abc_17692_n9647) );
  INVX1 INVX1_1872 ( .A(_abc_17692_n9650), .Y(_abc_17692_n9651) );
  INVX1 INVX1_1873 ( .A(_abc_17692_n9652), .Y(_abc_17692_n9653) );
  INVX1 INVX1_1874 ( .A(_abc_17692_n9668), .Y(_abc_17692_n9669) );
  INVX1 INVX1_1875 ( .A(_abc_17692_n9672), .Y(_abc_17692_n9673) );
  INVX1 INVX1_1876 ( .A(_abc_17692_n9438), .Y(_abc_17692_n9675) );
  INVX1 INVX1_1877 ( .A(_abc_17692_n9678), .Y(_abc_17692_n9679) );
  INVX1 INVX1_1878 ( .A(_abc_17692_n9680), .Y(_abc_17692_n9681) );
  INVX1 INVX1_1879 ( .A(_abc_17692_n9453), .Y(_abc_17692_n9687) );
  INVX1 INVX1_188 ( .A(_abc_17692_n1546), .Y(_abc_17692_n1547) );
  INVX1 INVX1_1880 ( .A(_abc_17692_n9692), .Y(_abc_17692_n9693) );
  INVX1 INVX1_1881 ( .A(_abc_17692_n9701), .Y(_abc_17692_n9702) );
  INVX1 INVX1_1882 ( .A(workunit2_16_bF_buf0), .Y(_abc_17692_n9717) );
  INVX1 INVX1_1883 ( .A(_abc_17692_n9740), .Y(_abc_17692_n9741) );
  INVX1 INVX1_1884 ( .A(_abc_17692_n9745), .Y(_abc_17692_n9746) );
  INVX1 INVX1_1885 ( .A(_abc_17692_n9747), .Y(_abc_17692_n9748) );
  INVX1 INVX1_1886 ( .A(_abc_17692_n9596), .Y(_abc_17692_n9749) );
  INVX1 INVX1_1887 ( .A(_abc_17692_n9750), .Y(_abc_17692_n9752) );
  INVX1 INVX1_1888 ( .A(_abc_17692_n9764), .Y(_abc_17692_n9765) );
  INVX1 INVX1_1889 ( .A(_abc_17692_n9766), .Y(_abc_17692_n9767) );
  INVX1 INVX1_189 ( .A(_abc_17692_n1555), .Y(_abc_17692_n1556) );
  INVX1 INVX1_1890 ( .A(_abc_17692_n9768), .Y(_abc_17692_n9769) );
  INVX1 INVX1_1891 ( .A(_abc_17692_n9783), .Y(_abc_17692_n9784) );
  INVX1 INVX1_1892 ( .A(_abc_17692_n9785), .Y(_abc_17692_n9786) );
  INVX1 INVX1_1893 ( .A(_abc_17692_n9777), .Y(_abc_17692_n9788) );
  INVX1 INVX1_1894 ( .A(_abc_17692_n9804), .Y(_abc_17692_n9805) );
  INVX1 INVX1_1895 ( .A(_abc_17692_n9806), .Y(_abc_17692_n9807) );
  INVX1 INVX1_1896 ( .A(_abc_17692_n9808), .Y(_abc_17692_n9810) );
  INVX1 INVX1_1897 ( .A(_abc_17692_n9816), .Y(_abc_17692_n9817) );
  INVX1 INVX1_1898 ( .A(_abc_17692_n9822), .Y(_abc_17692_n9823) );
  INVX1 INVX1_1899 ( .A(_abc_17692_n9824), .Y(_abc_17692_n9825) );
  INVX1 INVX1_19 ( .A(_abc_17692_n714_1), .Y(_abc_17692_n715_1) );
  INVX1 INVX1_190 ( .A(delta_23_), .Y(_abc_17692_n1557) );
  INVX1 INVX1_1900 ( .A(_abc_17692_n9830), .Y(_abc_17692_n9831) );
  INVX1 INVX1_1901 ( .A(_abc_17692_n9836), .Y(_abc_17692_n9837) );
  INVX1 INVX1_1902 ( .A(_abc_17692_n9854), .Y(_abc_17692_n9855) );
  INVX1 INVX1_1903 ( .A(_abc_17692_n9858), .Y(_abc_17692_n9859) );
  INVX1 INVX1_1904 ( .A(_abc_17692_n9865), .Y(_abc_17692_n9866) );
  INVX1 INVX1_1905 ( .A(_abc_17692_n9867), .Y(_abc_17692_n9874) );
  INVX1 INVX1_1906 ( .A(_abc_17692_n9881), .Y(_abc_17692_n9882) );
  INVX1 INVX1_1907 ( .A(_abc_17692_n9890), .Y(_abc_17692_n9891) );
  INVX1 INVX1_1908 ( .A(_abc_17692_n9894), .Y(_abc_17692_n9895) );
  INVX1 INVX1_1909 ( .A(_abc_17692_n1877_bF_buf1), .Y(_abc_17692_n9897) );
  INVX1 INVX1_191 ( .A(sum_23_), .Y(_abc_17692_n1558) );
  INVX1 INVX1_1910 ( .A(_abc_17692_n9885), .Y(_abc_17692_n9898) );
  INVX1 INVX1_1911 ( .A(_abc_17692_n9905), .Y(_abc_17692_n9906) );
  INVX1 INVX1_1912 ( .A(_abc_17692_n9912), .Y(_abc_17692_n9913) );
  INVX1 INVX1_1913 ( .A(_abc_17692_n9917), .Y(_abc_17692_n9918) );
  INVX1 INVX1_1914 ( .A(_abc_17692_n1846_bF_buf1), .Y(_abc_17692_n9920) );
  INVX1 INVX1_1915 ( .A(_abc_17692_n9908), .Y(_abc_17692_n9921) );
  INVX1 INVX1_1916 ( .A(_abc_17692_n9928), .Y(_abc_17692_n9929) );
  INVX1 INVX1_1917 ( .A(_abc_17692_n9931), .Y(_abc_17692_n9932) );
  INVX1 INVX1_1918 ( .A(_abc_17692_n9941), .Y(_abc_17692_n9942) );
  INVX1 INVX1_1919 ( .A(_abc_17692_n1830_bF_buf1), .Y(_abc_17692_n9944) );
  INVX1 INVX1_192 ( .A(_abc_17692_n1559), .Y(_abc_17692_n1560) );
  INVX1 INVX1_1920 ( .A(_abc_17692_n9953), .Y(_abc_17692_n9954) );
  INVX1 INVX1_1921 ( .A(_abc_17692_n9956), .Y(_abc_17692_n9957) );
  INVX1 INVX1_1922 ( .A(_abc_17692_n9965), .Y(_abc_17692_n9966) );
  INVX1 INVX1_1923 ( .A(_abc_17692_n9799), .Y(_abc_17692_n9976) );
  INVX1 INVX1_1924 ( .A(_abc_17692_n9575), .Y(_abc_17692_n9977) );
  INVX1 INVX1_1925 ( .A(_abc_17692_n9982), .Y(_abc_17692_n9984) );
  INVX1 INVX1_1926 ( .A(_abc_17692_n9988), .Y(_abc_17692_n9989) );
  INVX1 INVX1_1927 ( .A(_abc_17692_n9991), .Y(_abc_17692_n9992) );
  INVX1 INVX1_1928 ( .A(_abc_17692_n9994), .Y(_abc_17692_n9995) );
  INVX1 INVX1_1929 ( .A(_abc_17692_n9998), .Y(_abc_17692_n10001) );
  INVX1 INVX1_193 ( .A(_abc_17692_n1561), .Y(_abc_17692_n1562_1) );
  INVX1 INVX1_1930 ( .A(_abc_17692_n9390), .Y(_abc_17692_n10006) );
  INVX1 INVX1_1931 ( .A(_abc_17692_n9685), .Y(_abc_17692_n10007) );
  INVX1 INVX1_1932 ( .A(_abc_17692_n10008), .Y(_abc_17692_n10009) );
  INVX1 INVX1_1933 ( .A(_abc_17692_n9640), .Y(_abc_17692_n10012) );
  INVX1 INVX1_1934 ( .A(_abc_17692_n9759), .Y(_abc_17692_n10013) );
  INVX1 INVX1_1935 ( .A(_abc_17692_n10015), .Y(_abc_17692_n10016) );
  INVX1 INVX1_1936 ( .A(_abc_17692_n9689), .Y(_abc_17692_n10017) );
  INVX1 INVX1_1937 ( .A(_abc_17692_n10033), .Y(_abc_17692_n10034) );
  INVX1 INVX1_1938 ( .A(_abc_17692_n9397), .Y(_abc_17692_n10039) );
  INVX1 INVX1_1939 ( .A(_abc_17692_n9696), .Y(_abc_17692_n10044) );
  INVX1 INVX1_194 ( .A(_abc_17692_n1563), .Y(_abc_17692_n1564) );
  INVX1 INVX1_1940 ( .A(_abc_17692_n9699), .Y(_abc_17692_n10048) );
  INVX1 INVX1_1941 ( .A(_abc_17692_n8383_bF_buf2), .Y(_abc_17692_n10059) );
  INVX1 INVX1_1942 ( .A(_abc_17692_n10061), .Y(_abc_17692_n10062) );
  INVX1 INVX1_1943 ( .A(_abc_17692_n10065), .Y(workunit1_12__FF_INPUT) );
  INVX1 INVX1_1944 ( .A(_abc_17692_n10072), .Y(_abc_17692_n10073) );
  INVX1 INVX1_1945 ( .A(_abc_17692_n10075), .Y(_abc_17692_n10076) );
  INVX1 INVX1_1946 ( .A(_abc_17692_n10082), .Y(_abc_17692_n10084) );
  INVX1 INVX1_1947 ( .A(_abc_17692_n10086), .Y(_abc_17692_n10087) );
  INVX1 INVX1_1948 ( .A(_abc_17692_n10088), .Y(_abc_17692_n10090) );
  INVX1 INVX1_1949 ( .A(_abc_17692_n10096), .Y(_abc_17692_n10098) );
  INVX1 INVX1_195 ( .A(_abc_17692_n1569), .Y(_abc_17692_n1570) );
  INVX1 INVX1_1950 ( .A(_abc_17692_n10100), .Y(_abc_17692_n10101) );
  INVX1 INVX1_1951 ( .A(_abc_17692_n10102), .Y(_abc_17692_n10103) );
  INVX1 INVX1_1952 ( .A(_abc_17692_n10111), .Y(_abc_17692_n10112) );
  INVX1 INVX1_1953 ( .A(_abc_17692_n10114), .Y(_abc_17692_n10115) );
  INVX1 INVX1_1954 ( .A(_abc_17692_n10116), .Y(_abc_17692_n10118) );
  INVX1 INVX1_1955 ( .A(_abc_17692_n10130), .Y(_abc_17692_n10131) );
  INVX1 INVX1_1956 ( .A(_abc_17692_n9919), .Y(_abc_17692_n10132) );
  INVX1 INVX1_1957 ( .A(_abc_17692_n10133), .Y(_abc_17692_n10134) );
  INVX1 INVX1_1958 ( .A(_abc_17692_n9952), .Y(_abc_17692_n10144) );
  INVX1 INVX1_1959 ( .A(_abc_17692_n10146), .Y(_abc_17692_n10148) );
  INVX1 INVX1_196 ( .A(_abc_17692_n1571), .Y(_abc_17692_n1573) );
  INVX1 INVX1_1960 ( .A(_abc_17692_n10153), .Y(_abc_17692_n10155) );
  INVX1 INVX1_1961 ( .A(_abc_17692_n9927), .Y(_abc_17692_n10159) );
  INVX1 INVX1_1962 ( .A(_abc_17692_n10161), .Y(_abc_17692_n10162) );
  INVX1 INVX1_1963 ( .A(_abc_17692_n9904), .Y(_abc_17692_n10167) );
  INVX1 INVX1_1964 ( .A(_abc_17692_n10169), .Y(_abc_17692_n10171) );
  INVX1 INVX1_1965 ( .A(_abc_17692_n10071), .Y(_abc_17692_n10184) );
  INVX1 INVX1_1966 ( .A(_abc_17692_n10186), .Y(_abc_17692_n10187) );
  INVX1 INVX1_1967 ( .A(_abc_17692_n10190), .Y(_abc_17692_n10191) );
  INVX1 INVX1_1968 ( .A(_abc_17692_n10197), .Y(_abc_17692_n10198) );
  INVX1 INVX1_1969 ( .A(_abc_17692_n10196), .Y(_abc_17692_n10203) );
  INVX1 INVX1_197 ( .A(sum_24_), .Y(_abc_17692_n1581) );
  INVX1 INVX1_1970 ( .A(_abc_17692_n10206), .Y(_abc_17692_n10208) );
  INVX1 INVX1_1971 ( .A(_abc_17692_n10210), .Y(_abc_17692_n10211) );
  INVX1 INVX1_1972 ( .A(_abc_17692_n10085), .Y(_abc_17692_n10215) );
  INVX1 INVX1_1973 ( .A(_abc_17692_n10222), .Y(_abc_17692_n10223) );
  INVX1 INVX1_1974 ( .A(_abc_17692_n10229), .Y(_abc_17692_n10230) );
  INVX1 INVX1_1975 ( .A(_abc_17692_n10232), .Y(_abc_17692_n10233) );
  INVX1 INVX1_1976 ( .A(_abc_17692_n10099), .Y(_abc_17692_n10234) );
  INVX1 INVX1_1977 ( .A(_abc_17692_n10240), .Y(_abc_17692_n10241) );
  INVX1 INVX1_1978 ( .A(_abc_17692_n10247), .Y(_abc_17692_n10248) );
  INVX1 INVX1_1979 ( .A(_abc_17692_n10125), .Y(_abc_17692_n10252) );
  INVX1 INVX1_198 ( .A(_abc_17692_n1583), .Y(_abc_17692_n1584) );
  INVX1 INVX1_1980 ( .A(_abc_17692_n10258), .Y(_abc_17692_n10259) );
  INVX1 INVX1_1981 ( .A(_abc_17692_n10265), .Y(_abc_17692_n10266) );
  INVX1 INVX1_1982 ( .A(_abc_17692_n10275), .Y(_abc_17692_n10276) );
  INVX1 INVX1_1983 ( .A(_abc_17692_n10290), .Y(_abc_17692_n10291) );
  INVX1 INVX1_1984 ( .A(_abc_17692_n10251), .Y(_abc_17692_n10295) );
  INVX1 INVX1_1985 ( .A(_abc_17692_n10296), .Y(_abc_17692_n10297) );
  INVX1 INVX1_1986 ( .A(_abc_17692_n10299), .Y(_abc_17692_n10300) );
  INVX1 INVX1_1987 ( .A(_abc_17692_n10301), .Y(_abc_17692_n10302) );
  INVX1 INVX1_1988 ( .A(_abc_17692_n10305), .Y(_abc_17692_n10306) );
  INVX1 INVX1_1989 ( .A(_abc_17692_n10269), .Y(_abc_17692_n10310) );
  INVX1 INVX1_199 ( .A(_abc_17692_n1587), .Y(_abc_17692_n1588) );
  INVX1 INVX1_1990 ( .A(_abc_17692_n10110), .Y(_abc_17692_n10311) );
  INVX1 INVX1_1991 ( .A(_abc_17692_n10318), .Y(_abc_17692_n10319) );
  INVX1 INVX1_1992 ( .A(_abc_17692_n10214), .Y(_abc_17692_n10325) );
  INVX1 INVX1_1993 ( .A(_abc_17692_n10332), .Y(_abc_17692_n10333) );
  INVX1 INVX1_1994 ( .A(_abc_17692_n10348), .Y(_abc_17692_n10349) );
  INVX1 INVX1_1995 ( .A(_abc_17692_n10350), .Y(_abc_17692_n10355) );
  INVX1 INVX1_1996 ( .A(_abc_17692_n10364), .Y(_abc_17692_n10365) );
  INVX1 INVX1_1997 ( .A(_abc_17692_n10368), .Y(_abc_17692_n10369) );
  INVX1 INVX1_1998 ( .A(_abc_17692_n10228), .Y(_abc_17692_n10370) );
  INVX1 INVX1_1999 ( .A(_abc_17692_n10371), .Y(_abc_17692_n10372) );
  INVX1 INVX1_2 ( .A(state_7_bF_buf4), .Y(_abc_17692_n626) );
  INVX1 INVX1_20 ( .A(_abc_17692_n719), .Y(_abc_17692_n720) );
  INVX1 INVX1_200 ( .A(_abc_17692_n1593), .Y(_abc_17692_n1594) );
  INVX1 INVX1_2000 ( .A(_abc_17692_n10373), .Y(_abc_17692_n10375) );
  INVX1 INVX1_2001 ( .A(_abc_17692_n10388), .Y(_abc_17692_n10389) );
  INVX1 INVX1_2002 ( .A(_abc_17692_n10387), .Y(_abc_17692_n10391) );
  INVX1 INVX1_2003 ( .A(_abc_17692_n10404), .Y(_abc_17692_n10405) );
  INVX1 INVX1_2004 ( .A(_abc_17692_n10403), .Y(_abc_17692_n10407) );
  INVX1 INVX1_2005 ( .A(_abc_17692_n10414), .Y(_abc_17692_n10422) );
  INVX1 INVX1_2006 ( .A(_abc_17692_n10418), .Y(_abc_17692_n10423) );
  INVX1 INVX1_2007 ( .A(_abc_17692_n10420), .Y(_abc_17692_n10425) );
  INVX1 INVX1_2008 ( .A(_abc_17692_n10433), .Y(_abc_17692_n10435) );
  INVX1 INVX1_2009 ( .A(_abc_17692_n10439), .Y(_abc_17692_n10440) );
  INVX1 INVX1_201 ( .A(_abc_17692_n1597), .Y(_abc_17692_n1598_1) );
  INVX1 INVX1_2010 ( .A(_abc_17692_n10441), .Y(_abc_17692_n10442) );
  INVX1 INVX1_2011 ( .A(_abc_17692_n10447), .Y(_abc_17692_n10448) );
  INVX1 INVX1_2012 ( .A(_abc_17692_n10449), .Y(_abc_17692_n10450) );
  INVX1 INVX1_2013 ( .A(_abc_17692_n10457), .Y(_abc_17692_n10458) );
  INVX1 INVX1_2014 ( .A(_abc_17692_n10459), .Y(_abc_17692_n10460) );
  INVX1 INVX1_2015 ( .A(_abc_17692_n10473), .Y(_abc_17692_n10474) );
  INVX1 INVX1_2016 ( .A(_abc_17692_n10481), .Y(_abc_17692_n10482) );
  INVX1 INVX1_2017 ( .A(_abc_17692_n10487), .Y(_abc_17692_n10488) );
  INVX1 INVX1_2018 ( .A(_abc_17692_n10491), .Y(_abc_17692_n10498) );
  INVX1 INVX1_2019 ( .A(_abc_17692_n10505), .Y(_abc_17692_n10506) );
  INVX1 INVX1_202 ( .A(_abc_17692_n1600), .Y(_abc_17692_n1601) );
  INVX1 INVX1_2020 ( .A(_abc_17692_n10367), .Y(_abc_17692_n10511) );
  INVX1 INVX1_2021 ( .A(_abc_17692_n10518), .Y(_abc_17692_n10519) );
  INVX1 INVX1_2022 ( .A(_abc_17692_n10526), .Y(_abc_17692_n10527) );
  INVX1 INVX1_2023 ( .A(_abc_17692_n10532), .Y(_abc_17692_n10533) );
  INVX1 INVX1_2024 ( .A(_abc_17692_n10539), .Y(_abc_17692_n10540) );
  INVX1 INVX1_2025 ( .A(_abc_17692_n10542), .Y(_abc_17692_n10543) );
  INVX1 INVX1_2026 ( .A(_abc_17692_n10549), .Y(_abc_17692_n10550) );
  INVX1 INVX1_2027 ( .A(_abc_17692_n10563), .Y(_abc_17692_n10564) );
  INVX1 INVX1_2028 ( .A(_abc_17692_n10572), .Y(_abc_17692_n10573) );
  INVX1 INVX1_2029 ( .A(_abc_17692_n10586), .Y(_abc_17692_n10587) );
  INVX1 INVX1_203 ( .A(_abc_17692_n1585), .Y(_abc_17692_n1605) );
  INVX1 INVX1_2030 ( .A(_abc_17692_n10575), .Y(_abc_17692_n10592) );
  INVX1 INVX1_2031 ( .A(_abc_17692_n10212), .Y(_abc_17692_n10595) );
  INVX1 INVX1_2032 ( .A(_abc_17692_n10382), .Y(_abc_17692_n10596) );
  INVX1 INVX1_2033 ( .A(_abc_17692_n10604), .Y(_abc_17692_n10605) );
  INVX1 INVX1_2034 ( .A(_abc_17692_n10508), .Y(_abc_17692_n10608) );
  INVX1 INVX1_2035 ( .A(_abc_17692_n10236), .Y(_abc_17692_n10609) );
  INVX1 INVX1_2036 ( .A(_abc_17692_n10612), .Y(_abc_17692_n10613) );
  INVX1 INVX1_2037 ( .A(_abc_17692_n10616), .Y(_abc_17692_n10617) );
  INVX1 INVX1_2038 ( .A(_abc_17692_n10237), .Y(_abc_17692_n10618) );
  INVX1 INVX1_2039 ( .A(_abc_17692_n10619), .Y(_abc_17692_n10620) );
  INVX1 INVX1_204 ( .A(_abc_17692_n1615), .Y(_abc_17692_n1616) );
  INVX1 INVX1_2040 ( .A(_abc_17692_n10623), .Y(_abc_17692_n10624) );
  INVX1 INVX1_2041 ( .A(_abc_17692_n10552), .Y(_abc_17692_n10628) );
  INVX1 INVX1_2042 ( .A(_abc_17692_n10632), .Y(_abc_17692_n10633) );
  INVX1 INVX1_2043 ( .A(_abc_17692_n10638), .Y(_abc_17692_n10639) );
  INVX1 INVX1_2044 ( .A(_abc_17692_n10529), .Y(_abc_17692_n10643) );
  INVX1 INVX1_2045 ( .A(_abc_17692_n10249), .Y(_abc_17692_n10646) );
  INVX1 INVX1_2046 ( .A(_abc_17692_n10647), .Y(_abc_17692_n10648) );
  INVX1 INVX1_2047 ( .A(_abc_17692_n10649), .Y(_abc_17692_n10650) );
  INVX1 INVX1_2048 ( .A(_abc_17692_n10656), .Y(_abc_17692_n10657) );
  INVX1 INVX1_2049 ( .A(_abc_17692_n10672), .Y(_abc_17692_n10673) );
  INVX1 INVX1_205 ( .A(_abc_17692_n1622), .Y(_abc_17692_n1623) );
  INVX1 INVX1_2050 ( .A(_abc_17692_n10674), .Y(_abc_17692_n10675) );
  INVX1 INVX1_2051 ( .A(_abc_17692_n10676), .Y(_abc_17692_n10677) );
  INVX1 INVX1_2052 ( .A(_abc_17692_n10678), .Y(_abc_17692_n10679) );
  INVX1 INVX1_2053 ( .A(_abc_17692_n10681), .Y(_abc_17692_n10682) );
  INVX1 INVX1_2054 ( .A(_abc_17692_n10683), .Y(_abc_17692_n10685) );
  INVX1 INVX1_2055 ( .A(_abc_17692_n10688), .Y(_abc_17692_n10689) );
  INVX1 INVX1_2056 ( .A(_abc_17692_n10687), .Y(_abc_17692_n10690) );
  INVX1 INVX1_2057 ( .A(_abc_17692_n10691), .Y(_abc_17692_n10692) );
  INVX1 INVX1_2058 ( .A(_abc_17692_n10694), .Y(_abc_17692_n10695) );
  INVX1 INVX1_2059 ( .A(_abc_17692_n10693), .Y(_abc_17692_n10697) );
  INVX1 INVX1_206 ( .A(delta_25_), .Y(_abc_17692_n1624) );
  INVX1 INVX1_2060 ( .A(_abc_17692_n10704), .Y(_abc_17692_n10705) );
  INVX1 INVX1_2061 ( .A(_abc_17692_n10703), .Y(_abc_17692_n10706) );
  INVX1 INVX1_2062 ( .A(_abc_17692_n10707), .Y(_abc_17692_n10708) );
  INVX1 INVX1_2063 ( .A(_abc_17692_n10709), .Y(_abc_17692_n10712) );
  INVX1 INVX1_2064 ( .A(_abc_17692_n10710), .Y(_abc_17692_n10713) );
  INVX1 INVX1_2065 ( .A(_abc_17692_n10719), .Y(_abc_17692_n10720) );
  INVX1 INVX1_2066 ( .A(_abc_17692_n10724), .Y(_abc_17692_n10725) );
  INVX1 INVX1_2067 ( .A(_abc_17692_n10723), .Y(_abc_17692_n10727) );
  INVX1 INVX1_2068 ( .A(_abc_17692_n10733), .Y(_abc_17692_n10735) );
  INVX1 INVX1_2069 ( .A(_abc_17692_n10737), .Y(_abc_17692_n10740) );
  INVX1 INVX1_207 ( .A(sum_25_), .Y(_abc_17692_n1625) );
  INVX1 INVX1_2070 ( .A(_abc_17692_n10738), .Y(_abc_17692_n10741) );
  INVX1 INVX1_2071 ( .A(_abc_17692_n10571), .Y(_abc_17692_n10750) );
  INVX1 INVX1_2072 ( .A(_abc_17692_n10751), .Y(_abc_17692_n10752) );
  INVX1 INVX1_2073 ( .A(_abc_17692_n10753), .Y(_abc_17692_n10754) );
  INVX1 INVX1_2074 ( .A(_abc_17692_n10504), .Y(_abc_17692_n10759) );
  INVX1 INVX1_2075 ( .A(_abc_17692_n10760), .Y(_abc_17692_n10761) );
  INVX1 INVX1_2076 ( .A(_abc_17692_n10762), .Y(_abc_17692_n10764) );
  INVX1 INVX1_2077 ( .A(_abc_17692_n10525), .Y(_abc_17692_n10768) );
  INVX1 INVX1_2078 ( .A(_abc_17692_n10769), .Y(_abc_17692_n10770) );
  INVX1 INVX1_2079 ( .A(_abc_17692_n10771), .Y(_abc_17692_n10772) );
  INVX1 INVX1_208 ( .A(_abc_17692_n1626), .Y(_abc_17692_n1627) );
  INVX1 INVX1_2080 ( .A(_abc_17692_n10548), .Y(_abc_17692_n10777) );
  INVX1 INVX1_2081 ( .A(_abc_17692_n10778), .Y(_abc_17692_n10779) );
  INVX1 INVX1_2082 ( .A(_abc_17692_n10780), .Y(_abc_17692_n10782) );
  INVX1 INVX1_2083 ( .A(_abc_17692_n10802), .Y(_abc_17692_n10803) );
  INVX1 INVX1_2084 ( .A(_abc_17692_n10806), .Y(_abc_17692_n10807) );
  INVX1 INVX1_2085 ( .A(_abc_17692_n10799), .Y(_abc_17692_n10809) );
  INVX1 INVX1_2086 ( .A(_abc_17692_n10815), .Y(_abc_17692_n10816) );
  INVX1 INVX1_2087 ( .A(_abc_17692_n10826), .Y(_abc_17692_n10827) );
  INVX1 INVX1_2088 ( .A(_abc_17692_n10833), .Y(_abc_17692_n10834) );
  INVX1 INVX1_2089 ( .A(_abc_17692_n10836), .Y(_abc_17692_n10837) );
  INVX1 INVX1_209 ( .A(_abc_17692_n1628), .Y(_abc_17692_n1629) );
  INVX1 INVX1_2090 ( .A(_abc_17692_n10843), .Y(_abc_17692_n10844) );
  INVX1 INVX1_2091 ( .A(_abc_17692_n10850), .Y(_abc_17692_n10852) );
  INVX1 INVX1_2092 ( .A(_abc_17692_n10722), .Y(_abc_17692_n10855) );
  INVX1 INVX1_2093 ( .A(_abc_17692_n10861), .Y(_abc_17692_n10862) );
  INVX1 INVX1_2094 ( .A(_abc_17692_n10870), .Y(_abc_17692_n10871) );
  INVX1 INVX1_2095 ( .A(_abc_17692_n10872), .Y(_abc_17692_n10873) );
  INVX1 INVX1_2096 ( .A(_abc_17692_n10736), .Y(_abc_17692_n10874) );
  INVX1 INVX1_2097 ( .A(_abc_17692_n10651), .Y(_abc_17692_n10877) );
  INVX1 INVX1_2098 ( .A(_abc_17692_n10652), .Y(_abc_17692_n10878) );
  INVX1 INVX1_2099 ( .A(_abc_17692_n10881), .Y(_abc_17692_n10882) );
  INVX1 INVX1_21 ( .A(_abc_17692_n921), .Y(_abc_17692_n922) );
  INVX1 INVX1_210 ( .A(_abc_17692_n1631), .Y(_abc_17692_n1632) );
  INVX1 INVX1_2100 ( .A(_abc_17692_n10884), .Y(_abc_17692_n10885) );
  INVX1 INVX1_2101 ( .A(_abc_17692_n10886), .Y(_abc_17692_n10887) );
  INVX1 INVX1_2102 ( .A(_abc_17692_n10819), .Y(_abc_17692_n10895) );
  INVX1 INVX1_2103 ( .A(_abc_17692_n10896), .Y(_abc_17692_n10897) );
  INVX1 INVX1_2104 ( .A(_abc_17692_n10899), .Y(_abc_17692_n10900) );
  INVX1 INVX1_2105 ( .A(_abc_17692_n10905), .Y(_abc_17692_n10906) );
  INVX1 INVX1_2106 ( .A(_abc_17692_n10916), .Y(_abc_17692_n10917) );
  INVX1 INVX1_2107 ( .A(_abc_17692_n10854), .Y(_abc_17692_n10920) );
  INVX1 INVX1_2108 ( .A(_abc_17692_n10927), .Y(_abc_17692_n10928) );
  INVX1 INVX1_2109 ( .A(_abc_17692_n10932), .Y(_abc_17692_n10933) );
  INVX1 INVX1_211 ( .A(_abc_17692_n1640), .Y(_abc_17692_n1641) );
  INVX1 INVX1_2110 ( .A(_abc_17692_n10935), .Y(_abc_17692_n10936) );
  INVX1 INVX1_2111 ( .A(_abc_17692_n10941), .Y(_abc_17692_n10942) );
  INVX1 INVX1_2112 ( .A(_abc_17692_n10955), .Y(_abc_17692_n10956) );
  INVX1 INVX1_2113 ( .A(_abc_17692_n10959), .Y(_abc_17692_n10960) );
  INVX1 INVX1_2114 ( .A(_abc_17692_n10961), .Y(_abc_17692_n10962) );
  INVX1 INVX1_2115 ( .A(_abc_17692_n10963), .Y(_abc_17692_n10964) );
  INVX1 INVX1_2116 ( .A(_abc_17692_n10965), .Y(_abc_17692_n10966) );
  INVX1 INVX1_2117 ( .A(_abc_17692_n10967), .Y(_abc_17692_n10968) );
  INVX1 INVX1_2118 ( .A(_abc_17692_n10969), .Y(_abc_17692_n10970) );
  INVX1 INVX1_2119 ( .A(_abc_17692_n10982), .Y(_abc_17692_n10983) );
  INVX1 INVX1_212 ( .A(_abc_17692_n1642), .Y(_abc_17692_n1643) );
  INVX1 INVX1_2120 ( .A(_abc_17692_n10981), .Y(_abc_17692_n10986) );
  INVX1 INVX1_2121 ( .A(_abc_17692_n10984), .Y(_abc_17692_n10987) );
  INVX1 INVX1_2122 ( .A(_abc_17692_n10993), .Y(_abc_17692_n10994) );
  INVX1 INVX1_2123 ( .A(_abc_17692_n10998), .Y(_abc_17692_n10999) );
  INVX1 INVX1_2124 ( .A(_abc_17692_n10997), .Y(_abc_17692_n11001) );
  INVX1 INVX1_2125 ( .A(_abc_17692_n11014), .Y(_abc_17692_n11015) );
  INVX1 INVX1_2126 ( .A(_abc_17692_n10818), .Y(_abc_17692_n11034) );
  INVX1 INVX1_2127 ( .A(_abc_17692_n11035), .Y(_abc_17692_n11036) );
  INVX1 INVX1_2128 ( .A(_abc_17692_n11047), .Y(_abc_17692_n11048) );
  INVX1 INVX1_2129 ( .A(_abc_17692_n10832), .Y(_abc_17692_n11053) );
  INVX1 INVX1_213 ( .A(delta_26_), .Y(_abc_17692_n1652) );
  INVX1 INVX1_2130 ( .A(_abc_17692_n11054), .Y(_abc_17692_n11055) );
  INVX1 INVX1_2131 ( .A(_abc_17692_n11056), .Y(_abc_17692_n11058) );
  INVX1 INVX1_2132 ( .A(_abc_17692_n11062), .Y(_abc_17692_n11063) );
  INVX1 INVX1_2133 ( .A(_abc_17692_n11064), .Y(_abc_17692_n11065) );
  INVX1 INVX1_2134 ( .A(_abc_17692_n11070), .Y(_abc_17692_n11071) );
  INVX1 INVX1_2135 ( .A(_abc_17692_n11086), .Y(_abc_17692_n11087) );
  INVX1 INVX1_2136 ( .A(_abc_17692_n11089), .Y(_abc_17692_n11090) );
  INVX1 INVX1_2137 ( .A(_abc_17692_n10804), .Y(_abc_17692_n11091) );
  INVX1 INVX1_2138 ( .A(_abc_17692_n11098), .Y(_abc_17692_n11099) );
  INVX1 INVX1_2139 ( .A(_abc_17692_n11094), .Y(_abc_17692_n11105) );
  INVX1 INVX1_214 ( .A(sum_26_), .Y(_abc_17692_n1653) );
  INVX1 INVX1_2140 ( .A(_abc_17692_n11102), .Y(_abc_17692_n11107) );
  INVX1 INVX1_2141 ( .A(_abc_17692_n11113), .Y(_abc_17692_n11114) );
  INVX1 INVX1_2142 ( .A(_abc_17692_n11117), .Y(_abc_17692_n11118) );
  INVX1 INVX1_2143 ( .A(_abc_17692_n11119), .Y(_abc_17692_n11122) );
  INVX1 INVX1_2144 ( .A(_abc_17692_n11125), .Y(_abc_17692_n11126) );
  INVX1 INVX1_2145 ( .A(_abc_17692_n11127), .Y(_abc_17692_n11128) );
  INVX1 INVX1_2146 ( .A(_abc_17692_n11130), .Y(_abc_17692_n11131) );
  INVX1 INVX1_2147 ( .A(_abc_17692_n11138), .Y(_abc_17692_n11139) );
  INVX1 INVX1_2148 ( .A(_abc_17692_n10995), .Y(_abc_17692_n11144) );
  INVX1 INVX1_2149 ( .A(_abc_17692_n11146), .Y(_abc_17692_n11147) );
  INVX1 INVX1_215 ( .A(_abc_17692_n1655), .Y(_abc_17692_n1656) );
  INVX1 INVX1_2150 ( .A(_abc_17692_n11153), .Y(_abc_17692_n11154) );
  INVX1 INVX1_2151 ( .A(_abc_17692_n11159), .Y(_abc_17692_n11160) );
  INVX1 INVX1_2152 ( .A(_abc_17692_n11163), .Y(_abc_17692_n11164) );
  INVX1 INVX1_2153 ( .A(_abc_17692_n11173), .Y(_abc_17692_n11174) );
  INVX1 INVX1_2154 ( .A(_abc_17692_n11180), .Y(_abc_17692_n11181) );
  INVX1 INVX1_2155 ( .A(_abc_17692_n11184), .Y(_abc_17692_n11185) );
  INVX1 INVX1_2156 ( .A(_abc_17692_n11189), .Y(_abc_17692_n11190) );
  INVX1 INVX1_2157 ( .A(_abc_17692_n11186), .Y(_abc_17692_n11192) );
  INVX1 INVX1_2158 ( .A(_abc_17692_n11193), .Y(_abc_17692_n11194) );
  INVX1 INVX1_2159 ( .A(_abc_17692_n11196), .Y(_abc_17692_n11197) );
  INVX1 INVX1_216 ( .A(_abc_17692_n1657), .Y(_abc_17692_n1658) );
  INVX1 INVX1_2160 ( .A(_abc_17692_n11198), .Y(_abc_17692_n11199) );
  INVX1 INVX1_2161 ( .A(_abc_17692_n11218), .Y(_abc_17692_n11219) );
  INVX1 INVX1_2162 ( .A(_abc_17692_n11141), .Y(_abc_17692_n11222) );
  INVX1 INVX1_2163 ( .A(_abc_17692_n10839), .Y(_abc_17692_n11223) );
  INVX1 INVX1_2164 ( .A(_abc_17692_n11226), .Y(_abc_17692_n11227) );
  INVX1 INVX1_2165 ( .A(_abc_17692_n11230), .Y(_abc_17692_n11231) );
  INVX1 INVX1_2166 ( .A(_abc_17692_n11224), .Y(_abc_17692_n11232) );
  INVX1 INVX1_2167 ( .A(_abc_17692_n11236), .Y(_abc_17692_n11237) );
  INVX1 INVX1_2168 ( .A(_abc_17692_n11243), .Y(_abc_17692_n11244) );
  INVX1 INVX1_2169 ( .A(_abc_17692_n11247), .Y(_abc_17692_n11248) );
  INVX1 INVX1_217 ( .A(_abc_17692_n1661), .Y(_abc_17692_n1662) );
  INVX1 INVX1_2170 ( .A(_abc_17692_n11249), .Y(_abc_17692_n11250) );
  INVX1 INVX1_2171 ( .A(_abc_17692_n11254), .Y(_abc_17692_n11255) );
  INVX1 INVX1_2172 ( .A(_abc_17692_n10851), .Y(_abc_17692_n11261) );
  INVX1 INVX1_2173 ( .A(_abc_17692_n11264), .Y(_abc_17692_n11265) );
  INVX1 INVX1_2174 ( .A(_abc_17692_n10271), .Y(_abc_17692_n11266) );
  INVX1 INVX1_2175 ( .A(_abc_17692_n10272), .Y(_abc_17692_n11270) );
  INVX1 INVX1_2176 ( .A(_abc_17692_n11274), .Y(_abc_17692_n11275) );
  INVX1 INVX1_2177 ( .A(_abc_17692_n11277), .Y(_abc_17692_n11278) );
  INVX1 INVX1_2178 ( .A(_abc_17692_n11279), .Y(_abc_17692_n11280) );
  INVX1 INVX1_2179 ( .A(_abc_17692_n11296), .Y(_abc_17692_n11297) );
  INVX1 INVX1_218 ( .A(_abc_17692_n1663), .Y(_abc_17692_n1664) );
  INVX1 INVX1_2180 ( .A(_abc_17692_n11298), .Y(_abc_17692_n11299) );
  INVX1 INVX1_2181 ( .A(_abc_17692_n11300), .Y(_abc_17692_n11301) );
  INVX1 INVX1_2182 ( .A(_abc_17692_n11302), .Y(_abc_17692_n11303) );
  INVX1 INVX1_2183 ( .A(_abc_17692_n11304), .Y(_abc_17692_n11305) );
  INVX1 INVX1_2184 ( .A(_abc_17692_n11311), .Y(_abc_17692_n11313) );
  INVX1 INVX1_2185 ( .A(_abc_17692_n11316), .Y(_abc_17692_n11317) );
  INVX1 INVX1_2186 ( .A(_abc_17692_n11315), .Y(_abc_17692_n11319) );
  INVX1 INVX1_2187 ( .A(_abc_17692_n11325), .Y(_abc_17692_n11327) );
  INVX1 INVX1_2188 ( .A(_abc_17692_n11329), .Y(_abc_17692_n11330) );
  INVX1 INVX1_2189 ( .A(_abc_17692_n11332), .Y(_abc_17692_n11333) );
  INVX1 INVX1_219 ( .A(_abc_17692_n1666), .Y(_abc_17692_n1667) );
  INVX1 INVX1_2190 ( .A(_abc_17692_n11347), .Y(_abc_17692_n11348) );
  INVX1 INVX1_2191 ( .A(_abc_17692_n11183), .Y(_abc_17692_n11349) );
  INVX1 INVX1_2192 ( .A(_abc_17692_n11350), .Y(_abc_17692_n11351) );
  INVX1 INVX1_2193 ( .A(_abc_17692_n11360), .Y(_abc_17692_n11361) );
  INVX1 INVX1_2194 ( .A(_abc_17692_n11116), .Y(_abc_17692_n11365) );
  INVX1 INVX1_2195 ( .A(_abc_17692_n11364), .Y(_abc_17692_n11368) );
  INVX1 INVX1_2196 ( .A(_abc_17692_n11366), .Y(_abc_17692_n11369) );
  INVX1 INVX1_2197 ( .A(_abc_17692_n11376), .Y(_abc_17692_n11378) );
  INVX1 INVX1_2198 ( .A(_abc_17692_n11137), .Y(_abc_17692_n11382) );
  INVX1 INVX1_2199 ( .A(_abc_17692_n11383), .Y(_abc_17692_n11384) );
  INVX1 INVX1_22 ( .A(delta_1_), .Y(_abc_17692_n926_1) );
  INVX1 INVX1_220 ( .A(_abc_17692_n1673), .Y(_abc_17692_n1674) );
  INVX1 INVX1_2200 ( .A(_abc_17692_n11385), .Y(_abc_17692_n11386) );
  INVX1 INVX1_2201 ( .A(_abc_17692_n11391), .Y(_abc_17692_n11392) );
  INVX1 INVX1_2202 ( .A(_abc_17692_n11393), .Y(_abc_17692_n11394) );
  INVX1 INVX1_2203 ( .A(_abc_17692_n11399), .Y(_abc_17692_n11400) );
  INVX1 INVX1_2204 ( .A(_abc_17692_n11401), .Y(_abc_17692_n11403) );
  INVX1 INVX1_2205 ( .A(_abc_17692_n11416), .Y(_abc_17692_n11417) );
  INVX1 INVX1_2206 ( .A(_abc_17692_n11420), .Y(_abc_17692_n11421) );
  INVX1 INVX1_2207 ( .A(_abc_17692_n11425), .Y(_abc_17692_n11426) );
  INVX1 INVX1_2208 ( .A(_abc_17692_n11429), .Y(_abc_17692_n11433) );
  INVX1 INVX1_2209 ( .A(_abc_17692_n11435), .Y(_abc_17692_n11436) );
  INVX1 INVX1_221 ( .A(sum_27_), .Y(_abc_17692_n1682) );
  INVX1 INVX1_2210 ( .A(_abc_17692_n11440), .Y(_abc_17692_n11441) );
  INVX1 INVX1_2211 ( .A(_abc_17692_n11450), .Y(_abc_17692_n11451) );
  INVX1 INVX1_2212 ( .A(_abc_17692_n11457), .Y(_abc_17692_n11458) );
  INVX1 INVX1_2213 ( .A(_abc_17692_n11462), .Y(_abc_17692_n11463) );
  INVX1 INVX1_2214 ( .A(_abc_17692_n11465), .Y(_abc_17692_n11466) );
  INVX1 INVX1_2215 ( .A(_abc_17692_n11467), .Y(_abc_17692_n11468) );
  INVX1 INVX1_2216 ( .A(_abc_17692_n11471), .Y(_abc_17692_n11472) );
  INVX1 INVX1_2217 ( .A(_abc_17692_n11478), .Y(_abc_17692_n11479) );
  INVX1 INVX1_2218 ( .A(_abc_17692_n11482), .Y(_abc_17692_n11483) );
  INVX1 INVX1_2219 ( .A(_abc_17692_n11485), .Y(_abc_17692_n11486) );
  INVX1 INVX1_222 ( .A(_abc_17692_n1684), .Y(_abc_17692_n1685_1) );
  INVX1 INVX1_2220 ( .A(_abc_17692_n11487), .Y(_abc_17692_n11488) );
  INVX1 INVX1_2221 ( .A(_abc_17692_n11497), .Y(_abc_17692_n11498) );
  INVX1 INVX1_2222 ( .A(_abc_17692_n11501), .Y(_abc_17692_n11502) );
  INVX1 INVX1_2223 ( .A(_abc_17692_n11509), .Y(_abc_17692_n11510) );
  INVX1 INVX1_2224 ( .A(_abc_17692_n11363), .Y(_abc_17692_n11516) );
  INVX1 INVX1_2225 ( .A(_abc_17692_n11519), .Y(_abc_17692_n11520) );
  INVX1 INVX1_2226 ( .A(_abc_17692_n11523), .Y(_abc_17692_n11524) );
  INVX1 INVX1_2227 ( .A(_abc_17692_n11443), .Y(_abc_17692_n11528) );
  INVX1 INVX1_2228 ( .A(_abc_17692_n11529), .Y(_abc_17692_n11530) );
  INVX1 INVX1_2229 ( .A(_abc_17692_n11312), .Y(_abc_17692_n11532) );
  INVX1 INVX1_223 ( .A(_abc_17692_n1689), .Y(_abc_17692_n1690) );
  INVX1 INVX1_2230 ( .A(_abc_17692_n11534), .Y(_abc_17692_n11535) );
  INVX1 INVX1_2231 ( .A(_abc_17692_n11537), .Y(_abc_17692_n11538) );
  INVX1 INVX1_2232 ( .A(_abc_17692_n11461), .Y(_abc_17692_n11542) );
  INVX1 INVX1_2233 ( .A(_abc_17692_n11543), .Y(_abc_17692_n11544) );
  INVX1 INVX1_2234 ( .A(_abc_17692_n11346), .Y(_abc_17692_n11546) );
  INVX1 INVX1_2235 ( .A(_abc_17692_n11548), .Y(_abc_17692_n11549) );
  INVX1 INVX1_2236 ( .A(_abc_17692_n11552), .Y(_abc_17692_n11553) );
  INVX1 INVX1_2237 ( .A(_abc_17692_n11328), .Y(_abc_17692_n11556) );
  INVX1 INVX1_2238 ( .A(_abc_17692_n11562), .Y(_abc_17692_n11563) );
  INVX1 INVX1_2239 ( .A(_abc_17692_n11427), .Y(_abc_17692_n11576) );
  INVX1 INVX1_224 ( .A(_abc_17692_n1692), .Y(_abc_17692_n1693) );
  INVX1 INVX1_2240 ( .A(_abc_17692_n11581), .Y(_abc_17692_n11582) );
  INVX1 INVX1_2241 ( .A(_abc_17692_n11583), .Y(_abc_17692_n11584) );
  INVX1 INVX1_2242 ( .A(_abc_17692_n11585), .Y(_abc_17692_n11586) );
  INVX1 INVX1_2243 ( .A(_abc_17692_n11587), .Y(_abc_17692_n11588) );
  INVX1 INVX1_2244 ( .A(_abc_17692_n11605), .Y(_abc_17692_n11606) );
  INVX1 INVX1_2245 ( .A(_abc_17692_n11604), .Y(_abc_17692_n11608) );
  INVX1 INVX1_2246 ( .A(_abc_17692_n11620), .Y(_abc_17692_n11621) );
  INVX1 INVX1_2247 ( .A(_abc_17692_n11622), .Y(_abc_17692_n11623) );
  INVX1 INVX1_2248 ( .A(_abc_17692_n11624), .Y(_abc_17692_n11625) );
  INVX1 INVX1_2249 ( .A(_abc_17692_n11640), .Y(_abc_17692_n11641) );
  INVX1 INVX1_225 ( .A(_abc_17692_n1686), .Y(_abc_17692_n1698) );
  INVX1 INVX1_2250 ( .A(_abc_17692_n11661), .Y(_abc_17692_n11662) );
  INVX1 INVX1_2251 ( .A(_abc_17692_n11499), .Y(_abc_17692_n11672) );
  INVX1 INVX1_2252 ( .A(_abc_17692_n11673), .Y(_abc_17692_n11674) );
  INVX1 INVX1_2253 ( .A(_abc_17692_n11439), .Y(_abc_17692_n11679) );
  INVX1 INVX1_2254 ( .A(_abc_17692_n11680), .Y(_abc_17692_n11681) );
  INVX1 INVX1_2255 ( .A(_abc_17692_n11682), .Y(_abc_17692_n11683) );
  INVX1 INVX1_2256 ( .A(_abc_17692_n11688), .Y(_abc_17692_n11689) );
  INVX1 INVX1_2257 ( .A(_abc_17692_n11480), .Y(_abc_17692_n11694) );
  INVX1 INVX1_2258 ( .A(_abc_17692_n11695), .Y(_abc_17692_n11696) );
  INVX1 INVX1_2259 ( .A(_abc_17692_n11712), .Y(_abc_17692_n11713) );
  INVX1 INVX1_226 ( .A(_abc_17692_n1703), .Y(_abc_17692_n1704) );
  INVX1 INVX1_2260 ( .A(_abc_17692_n11716), .Y(_abc_17692_n11717) );
  INVX1 INVX1_2261 ( .A(_abc_17692_n11720), .Y(_abc_17692_n11721) );
  INVX1 INVX1_2262 ( .A(_abc_17692_n11729), .Y(_abc_17692_n11730) );
  INVX1 INVX1_2263 ( .A(_abc_17692_n11737), .Y(_abc_17692_n11739) );
  INVX1 INVX1_2264 ( .A(_abc_17692_n11743), .Y(_abc_17692_n11744) );
  INVX1 INVX1_2265 ( .A(_abc_17692_n11748), .Y(_abc_17692_n11749) );
  INVX1 INVX1_2266 ( .A(_abc_17692_n11753), .Y(_abc_17692_n11754) );
  INVX1 INVX1_2267 ( .A(_abc_17692_n11755), .Y(_abc_17692_n11756) );
  INVX1 INVX1_2268 ( .A(_abc_17692_n11757), .Y(_abc_17692_n11758) );
  INVX1 INVX1_2269 ( .A(_abc_17692_n11765), .Y(_abc_17692_n11766) );
  INVX1 INVX1_227 ( .A(_abc_17692_n1705), .Y(_abc_17692_n1706) );
  INVX1 INVX1_2270 ( .A(_abc_17692_n11768), .Y(_abc_17692_n11769) );
  INVX1 INVX1_2271 ( .A(_abc_17692_n11603), .Y(_abc_17692_n11774) );
  INVX1 INVX1_2272 ( .A(_abc_17692_n11782), .Y(_abc_17692_n11783) );
  INVX1 INVX1_2273 ( .A(_abc_17692_n11788), .Y(_abc_17692_n11790) );
  INVX1 INVX1_2274 ( .A(_abc_17692_n11805), .Y(_abc_17692_n11806) );
  INVX1 INVX1_2275 ( .A(_abc_17692_n11812), .Y(_abc_17692_n11814) );
  INVX1 INVX1_2276 ( .A(_abc_17692_n11826), .Y(_abc_17692_n11827) );
  INVX1 INVX1_2277 ( .A(_abc_17692_n11828), .Y(_abc_17692_n11829) );
  INVX1 INVX1_2278 ( .A(_abc_17692_n11741), .Y(_abc_17692_n11838) );
  INVX1 INVX1_2279 ( .A(_abc_17692_n11851), .Y(_abc_17692_n11852) );
  INVX1 INVX1_228 ( .A(sum_28_), .Y(_abc_17692_n1712) );
  INVX1 INVX1_2280 ( .A(_abc_17692_n11859), .Y(_abc_17692_n11860) );
  INVX1 INVX1_2281 ( .A(_abc_17692_n11233), .Y(_abc_17692_n11867) );
  INVX1 INVX1_2282 ( .A(_abc_17692_n11870), .Y(_abc_17692_n11871) );
  INVX1 INVX1_2283 ( .A(_abc_17692_n11872), .Y(_abc_17692_n11873) );
  INVX1 INVX1_2284 ( .A(_abc_17692_n11816), .Y(_abc_17692_n11877) );
  INVX1 INVX1_2285 ( .A(_abc_17692_n11882), .Y(_abc_17692_n11883) );
  INVX1 INVX1_2286 ( .A(_abc_17692_n11459), .Y(_abc_17692_n11884) );
  INVX1 INVX1_2287 ( .A(_abc_17692_n11891), .Y(_abc_17692_n11892) );
  INVX1 INVX1_2288 ( .A(_abc_17692_n11908), .Y(_abc_17692_n11909) );
  INVX1 INVX1_2289 ( .A(_abc_17692_n11792), .Y(_abc_17692_n11911) );
  INVX1 INVX1_229 ( .A(_abc_17692_n1714), .Y(_abc_17692_n1715) );
  INVX1 INVX1_2290 ( .A(_abc_17692_n11924), .Y(_abc_17692_n11925) );
  INVX1 INVX1_2291 ( .A(_abc_17692_n11928), .Y(_abc_17692_n11929) );
  INVX1 INVX1_2292 ( .A(_abc_17692_n11930), .Y(_abc_17692_n11931) );
  INVX1 INVX1_2293 ( .A(_abc_17692_n11932), .Y(_abc_17692_n11933) );
  INVX1 INVX1_2294 ( .A(_abc_17692_n11934), .Y(_abc_17692_n11935) );
  INVX1 INVX1_2295 ( .A(_abc_17692_n11948), .Y(_abc_17692_n11949) );
  INVX1 INVX1_2296 ( .A(_abc_17692_n11764), .Y(_abc_17692_n11950) );
  INVX1 INVX1_2297 ( .A(_abc_17692_n11951), .Y(_abc_17692_n11952) );
  INVX1 INVX1_2298 ( .A(_abc_17692_n11953), .Y(_abc_17692_n11955) );
  INVX1 INVX1_2299 ( .A(_abc_17692_n11968), .Y(_abc_17692_n11969) );
  INVX1 INVX1_23 ( .A(_abc_17692_n928), .Y(_abc_17692_n929) );
  INVX1 INVX1_230 ( .A(_abc_17692_n1718), .Y(_abc_17692_n1719) );
  INVX1 INVX1_2300 ( .A(_abc_17692_n11970), .Y(_abc_17692_n11971) );
  INVX1 INVX1_2301 ( .A(_abc_17692_n11967), .Y(_abc_17692_n11973) );
  INVX1 INVX1_2302 ( .A(_abc_17692_n11986), .Y(_abc_17692_n11987) );
  INVX1 INVX1_2303 ( .A(_abc_17692_n11985), .Y(_abc_17692_n11990) );
  INVX1 INVX1_2304 ( .A(_abc_17692_n11988), .Y(_abc_17692_n11991) );
  INVX1 INVX1_2305 ( .A(_abc_17692_n12000), .Y(_abc_17692_n12001) );
  INVX1 INVX1_2306 ( .A(_abc_17692_n12005), .Y(_abc_17692_n12006) );
  INVX1 INVX1_2307 ( .A(_abc_17692_n12008), .Y(_abc_17692_n12009) );
  INVX1 INVX1_2308 ( .A(_abc_17692_n12010), .Y(_abc_17692_n12013) );
  INVX1 INVX1_2309 ( .A(_abc_17692_n11738), .Y(_abc_17692_n12019) );
  INVX1 INVX1_231 ( .A(_abc_17692_n1720), .Y(_abc_17692_n1721) );
  INVX1 INVX1_2310 ( .A(_abc_17692_n12020), .Y(_abc_17692_n12021) );
  INVX1 INVX1_2311 ( .A(_abc_17692_n12026), .Y(_abc_17692_n12027) );
  INVX1 INVX1_2312 ( .A(_abc_17692_n11813), .Y(_abc_17692_n12032) );
  INVX1 INVX1_2313 ( .A(_abc_17692_n12033), .Y(_abc_17692_n12034) );
  INVX1 INVX1_2314 ( .A(_abc_17692_n11789), .Y(_abc_17692_n12039) );
  INVX1 INVX1_2315 ( .A(_abc_17692_n12040), .Y(_abc_17692_n12042) );
  INVX1 INVX1_2316 ( .A(_abc_17692_n12058), .Y(_abc_17692_n12059) );
  INVX1 INVX1_2317 ( .A(_abc_17692_n12065), .Y(_abc_17692_n12066) );
  INVX1 INVX1_2318 ( .A(_abc_17692_n12069), .Y(_abc_17692_n12070) );
  INVX1 INVX1_2319 ( .A(_abc_17692_n12073), .Y(_abc_17692_n12075) );
  INVX1 INVX1_232 ( .A(_abc_17692_n1716), .Y(_abc_17692_n1723) );
  INVX1 INVX1_2320 ( .A(_abc_17692_n12077), .Y(_abc_17692_n12078) );
  INVX1 INVX1_2321 ( .A(_abc_17692_n12082), .Y(_abc_17692_n12083) );
  INVX1 INVX1_2322 ( .A(_abc_17692_n12087), .Y(_abc_17692_n12088) );
  INVX1 INVX1_2323 ( .A(_abc_17692_n12093), .Y(_abc_17692_n12094) );
  INVX1 INVX1_2324 ( .A(_abc_17692_n12097), .Y(_abc_17692_n12098) );
  INVX1 INVX1_2325 ( .A(_abc_17692_n12099), .Y(_abc_17692_n12100) );
  INVX1 INVX1_2326 ( .A(_abc_17692_n12102), .Y(_abc_17692_n12103) );
  INVX1 INVX1_2327 ( .A(_abc_17692_n12110), .Y(_abc_17692_n12111) );
  INVX1 INVX1_2328 ( .A(_abc_17692_n12114), .Y(_abc_17692_n12115) );
  INVX1 INVX1_2329 ( .A(_abc_17692_n11962), .Y(_abc_17692_n12116) );
  INVX1 INVX1_233 ( .A(_abc_17692_n1728), .Y(_abc_17692_n1729) );
  INVX1 INVX1_2330 ( .A(_abc_17692_n12118), .Y(_abc_17692_n12119) );
  INVX1 INVX1_2331 ( .A(_abc_17692_n12123), .Y(_abc_17692_n12124) );
  INVX1 INVX1_2332 ( .A(_abc_17692_n12138), .Y(_abc_17692_n12140) );
  INVX1 INVX1_2333 ( .A(_abc_17692_n12142), .Y(_abc_17692_n12143) );
  INVX1 INVX1_2334 ( .A(_abc_17692_n12144), .Y(_abc_17692_n12145) );
  INVX1 INVX1_2335 ( .A(_abc_17692_n12157), .Y(_abc_17692_n12158) );
  INVX1 INVX1_2336 ( .A(_abc_17692_n12085), .Y(_abc_17692_n12162) );
  INVX1 INVX1_2337 ( .A(_abc_17692_n12163), .Y(_abc_17692_n12164) );
  INVX1 INVX1_2338 ( .A(_abc_17692_n12166), .Y(_abc_17692_n12167) );
  INVX1 INVX1_2339 ( .A(_abc_17692_n12171), .Y(_abc_17692_n12172) );
  INVX1 INVX1_234 ( .A(_abc_17692_n1731), .Y(_abc_17692_n1732) );
  INVX1 INVX1_2340 ( .A(_abc_17692_n12176), .Y(_abc_17692_n12177) );
  INVX1 INVX1_2341 ( .A(_abc_17692_n12179), .Y(_abc_17692_n12180) );
  INVX1 INVX1_2342 ( .A(_abc_17692_n12181), .Y(_abc_17692_n12182) );
  INVX1 INVX1_2343 ( .A(_abc_17692_n12186), .Y(_abc_17692_n12187) );
  INVX1 INVX1_2344 ( .A(_abc_17692_n12190), .Y(_abc_17692_n12191) );
  INVX1 INVX1_2345 ( .A(_abc_17692_n12195), .Y(_abc_17692_n12196) );
  INVX1 INVX1_2346 ( .A(_abc_17692_n12197), .Y(_abc_17692_n12199) );
  INVX1 INVX1_2347 ( .A(_abc_17692_n12213), .Y(_abc_17692_n12214) );
  INVX1 INVX1_2348 ( .A(_abc_17692_n12215), .Y(_abc_17692_n12216) );
  INVX1 INVX1_2349 ( .A(_abc_17692_n12217), .Y(_abc_17692_n12218) );
  INVX1 INVX1_235 ( .A(sum_29_), .Y(_abc_17692_n1738) );
  INVX1 INVX1_2350 ( .A(_abc_17692_n12219), .Y(_abc_17692_n12220) );
  INVX1 INVX1_2351 ( .A(_abc_17692_n12233), .Y(_abc_17692_n12234) );
  INVX1 INVX1_2352 ( .A(_abc_17692_n12235), .Y(_abc_17692_n12236) );
  INVX1 INVX1_2353 ( .A(_abc_17692_n12252), .Y(_abc_17692_n12253) );
  INVX1 INVX1_2354 ( .A(_abc_17692_n12254), .Y(_abc_17692_n12255) );
  INVX1 INVX1_2355 ( .A(_abc_17692_n12256), .Y(_abc_17692_n12257) );
  INVX1 INVX1_2356 ( .A(_abc_17692_n12271), .Y(_abc_17692_n12272) );
  INVX1 INVX1_2357 ( .A(_abc_17692_n12270), .Y(_abc_17692_n12274) );
  INVX1 INVX1_2358 ( .A(_abc_17692_n12287), .Y(_abc_17692_n12288) );
  INVX1 INVX1_2359 ( .A(_abc_17692_n12301), .Y(_abc_17692_n12302) );
  INVX1 INVX1_236 ( .A(_abc_17692_n1739), .Y(_abc_17692_n1740) );
  INVX1 INVX1_2360 ( .A(_abc_17692_n12081), .Y(_abc_17692_n12307) );
  INVX1 INVX1_2361 ( .A(_abc_17692_n12308), .Y(_abc_17692_n12309) );
  INVX1 INVX1_2362 ( .A(_abc_17692_n12310), .Y(_abc_17692_n12311) );
  INVX1 INVX1_2363 ( .A(_abc_17692_n12316), .Y(_abc_17692_n12317) );
  INVX1 INVX1_2364 ( .A(_abc_17692_n12318), .Y(_abc_17692_n12319) );
  INVX1 INVX1_2365 ( .A(_abc_17692_n12324), .Y(_abc_17692_n12325) );
  INVX1 INVX1_2366 ( .A(_abc_17692_n12344), .Y(_abc_17692_n12345) );
  INVX1 INVX1_2367 ( .A(_abc_17692_n12341), .Y(_abc_17692_n12347) );
  INVX1 INVX1_2368 ( .A(_abc_17692_n12353), .Y(_abc_17692_n12354) );
  INVX1 INVX1_2369 ( .A(_abc_17692_n12357), .Y(_abc_17692_n12358) );
  INVX1 INVX1_237 ( .A(delta_29_), .Y(_abc_17692_n1741) );
  INVX1 INVX1_2370 ( .A(_abc_17692_n12360), .Y(_abc_17692_n12361) );
  INVX1 INVX1_2371 ( .A(_abc_17692_n12366), .Y(_abc_17692_n12367) );
  INVX1 INVX1_2372 ( .A(_abc_17692_n12368), .Y(_abc_17692_n12369) );
  INVX1 INVX1_2373 ( .A(_abc_17692_n12371), .Y(_abc_17692_n12372) );
  INVX1 INVX1_2374 ( .A(_abc_17692_n12378), .Y(_abc_17692_n12379) );
  INVX1 INVX1_2375 ( .A(_abc_17692_n12381), .Y(_abc_17692_n12382) );
  INVX1 INVX1_2376 ( .A(_abc_17692_n12269), .Y(_abc_17692_n12387) );
  INVX1 INVX1_2377 ( .A(_abc_17692_n12392), .Y(_abc_17692_n12393) );
  INVX1 INVX1_2378 ( .A(_abc_17692_n12399), .Y(_abc_17692_n12400) );
  INVX1 INVX1_2379 ( .A(_abc_17692_n12403), .Y(_abc_17692_n12404) );
  INVX1 INVX1_238 ( .A(_abc_17692_n1742), .Y(_abc_17692_n1743) );
  INVX1 INVX1_2380 ( .A(_abc_17692_n12409), .Y(_abc_17692_n12410) );
  INVX1 INVX1_2381 ( .A(_abc_17692_n12417), .Y(_abc_17692_n12418) );
  INVX1 INVX1_2382 ( .A(_abc_17692_n12423), .Y(_abc_17692_n12424) );
  INVX1 INVX1_2383 ( .A(_abc_17692_n12427), .Y(_abc_17692_n12428) );
  INVX1 INVX1_2384 ( .A(_abc_17692_n12120), .Y(_abc_17692_n12429) );
  INVX1 INVX1_2385 ( .A(_abc_17692_n12435), .Y(_abc_17692_n12436) );
  INVX1 INVX1_2386 ( .A(_abc_17692_n12438), .Y(_abc_17692_n12439) );
  INVX1 INVX1_2387 ( .A(_abc_17692_n12440), .Y(_abc_17692_n12441) );
  INVX1 INVX1_2388 ( .A(_abc_17692_n12139), .Y(_abc_17692_n12455) );
  INVX1 INVX1_2389 ( .A(_abc_17692_n12460), .Y(_abc_17692_n12461) );
  INVX1 INVX1_239 ( .A(_abc_17692_n1744), .Y(_abc_17692_n1745) );
  INVX1 INVX1_2390 ( .A(_abc_17692_n12168), .Y(_abc_17692_n12465) );
  INVX1 INVX1_2391 ( .A(_abc_17692_n12470), .Y(_abc_17692_n12471) );
  INVX1 INVX1_2392 ( .A(_abc_17692_n12475), .Y(_abc_17692_n12476) );
  INVX1 INVX1_2393 ( .A(_abc_17692_n12477), .Y(_abc_17692_n12478) );
  INVX1 INVX1_2394 ( .A(_abc_17692_n12486), .Y(_abc_17692_n12487) );
  INVX1 INVX1_2395 ( .A(_abc_17692_n12491), .Y(_abc_17692_n12492) );
  INVX1 INVX1_2396 ( .A(_abc_17692_n12494), .Y(_abc_17692_n12495) );
  INVX1 INVX1_2397 ( .A(_abc_17692_n12095), .Y(_abc_17692_n12503) );
  INVX1 INVX1_2398 ( .A(_abc_17692_n12508), .Y(_abc_17692_n12509) );
  INVX1 INVX1_2399 ( .A(_abc_17692_n12523), .Y(_abc_17692_n12524) );
  INVX1 INVX1_24 ( .A(delta_0_), .Y(_abc_17692_n931) );
  INVX1 INVX1_240 ( .A(_abc_17692_n1746), .Y(_abc_17692_n1747) );
  INVX1 INVX1_2400 ( .A(_abc_17692_n12525), .Y(_abc_17692_n12526) );
  INVX1 INVX1_2401 ( .A(_abc_17692_n12527), .Y(_abc_17692_n12528) );
  INVX1 INVX1_2402 ( .A(_abc_17692_n12529), .Y(_abc_17692_n12530) );
  INVX1 INVX1_2403 ( .A(_abc_17692_n12544), .Y(_abc_17692_n12545) );
  INVX1 INVX1_2404 ( .A(_abc_17692_n12561), .Y(_abc_17692_n12562) );
  INVX1 INVX1_2405 ( .A(_abc_17692_n12377), .Y(_abc_17692_n12563) );
  INVX1 INVX1_2406 ( .A(_abc_17692_n12565), .Y(_abc_17692_n12566) );
  INVX1 INVX1_2407 ( .A(_abc_17692_n12580), .Y(_abc_17692_n12581) );
  INVX1 INVX1_2408 ( .A(_abc_17692_n12579), .Y(_abc_17692_n12584) );
  INVX1 INVX1_2409 ( .A(_abc_17692_n12582), .Y(_abc_17692_n12585) );
  INVX1 INVX1_241 ( .A(_abc_17692_n1748), .Y(_abc_17692_n1749) );
  INVX1 INVX1_2410 ( .A(_abc_17692_n12598), .Y(_abc_17692_n12599) );
  INVX1 INVX1_2411 ( .A(_abc_17692_n12600), .Y(_abc_17692_n12601) );
  INVX1 INVX1_2412 ( .A(_abc_17692_n12614), .Y(_abc_17692_n12615) );
  INVX1 INVX1_2413 ( .A(_abc_17692_n12620), .Y(_abc_17692_n12621) );
  INVX1 INVX1_2414 ( .A(_abc_17692_n12626), .Y(_abc_17692_n12628) );
  INVX1 INVX1_2415 ( .A(_abc_17692_n12632), .Y(_abc_17692_n12633) );
  INVX1 INVX1_2416 ( .A(_abc_17692_n7990), .Y(_abc_17692_n12647) );
  INVX1 INVX1_2417 ( .A(_abc_17692_n12650), .Y(_abc_17692_n12651) );
  INVX1 INVX1_2418 ( .A(_abc_17692_n12654), .Y(_abc_17692_n12655) );
  INVX1 INVX1_2419 ( .A(_abc_17692_n12667), .Y(_abc_17692_n12668) );
  INVX1 INVX1_242 ( .A(_abc_17692_n1755_1), .Y(_abc_17692_n1757) );
  INVX1 INVX1_2420 ( .A(_abc_17692_n12675), .Y(_abc_17692_n12676) );
  INVX1 INVX1_2421 ( .A(_abc_17692_n12681), .Y(_abc_17692_n12682) );
  INVX1 INVX1_2422 ( .A(_abc_17692_n12560), .Y(_abc_17692_n12688) );
  INVX1 INVX1_2423 ( .A(_abc_17692_n12692), .Y(_abc_17692_n12693) );
  INVX1 INVX1_2424 ( .A(_abc_17692_n12710), .Y(_abc_17692_n12711) );
  INVX1 INVX1_2425 ( .A(_abc_17692_n12724), .Y(_abc_17692_n12725) );
  INVX1 INVX1_2426 ( .A(_abc_17692_n12729), .Y(_abc_17692_n12730) );
  INVX1 INVX1_2427 ( .A(_abc_17692_n12734), .Y(_abc_17692_n12735) );
  INVX1 INVX1_2428 ( .A(_abc_17692_n11209), .Y(_abc_17692_n12745) );
  INVX1 INVX1_2429 ( .A(_abc_17692_n11046), .Y(_abc_17692_n12746) );
  INVX1 INVX1_243 ( .A(delta_30_), .Y(_abc_17692_n1764) );
  INVX1 INVX1_2430 ( .A(_abc_17692_n11211), .Y(_abc_17692_n12748) );
  INVX1 INVX1_2431 ( .A(_abc_17692_n11518), .Y(_abc_17692_n12754) );
  INVX1 INVX1_2432 ( .A(_abc_17692_n11843), .Y(_abc_17692_n12756) );
  INVX1 INVX1_2433 ( .A(_abc_17692_n10602), .Y(_abc_17692_n12761) );
  INVX1 INVX1_2434 ( .A(_abc_17692_n11214), .Y(_abc_17692_n12762) );
  INVX1 INVX1_2435 ( .A(_abc_17692_n12154), .Y(_abc_17692_n12766) );
  INVX1 INVX1_2436 ( .A(_abc_17692_n12151), .Y(_abc_17692_n12770) );
  INVX1 INVX1_2437 ( .A(_abc_17692_n12152), .Y(_abc_17692_n12771) );
  INVX1 INVX1_2438 ( .A(_abc_17692_n12454), .Y(_abc_17692_n12774) );
  INVX1 INVX1_2439 ( .A(_abc_17692_n12781), .Y(_abc_17692_n12782) );
  INVX1 INVX1_244 ( .A(sum_30_), .Y(_abc_17692_n1765) );
  INVX1 INVX1_2440 ( .A(_abc_17692_n12355), .Y(_abc_17692_n12789) );
  INVX1 INVX1_2441 ( .A(_abc_17692_n12685), .Y(_abc_17692_n12796) );
  INVX1 INVX1_2442 ( .A(_abc_17692_n12799), .Y(_abc_17692_n12800) );
  INVX1 INVX1_2443 ( .A(_abc_17692_n12803), .Y(_abc_17692_n12804) );
  INVX1 INVX1_2444 ( .A(_abc_17692_n12811), .Y(_abc_17692_n12812) );
  INVX1 INVX1_2445 ( .A(_abc_17692_n12815), .Y(_abc_17692_n12817) );
  INVX1 INVX1_2446 ( .A(_abc_17692_n12401), .Y(_abc_17692_n12824) );
  INVX1 INVX1_2447 ( .A(_abc_17692_n12828), .Y(_abc_17692_n12829) );
  INVX1 INVX1_2448 ( .A(_abc_17692_n12842), .Y(_abc_17692_n12843) );
  INVX1 INVX1_2449 ( .A(_abc_17692_n12844), .Y(_abc_17692_n12849) );
  INVX1 INVX1_245 ( .A(_abc_17692_n1767), .Y(_abc_17692_n1768) );
  INVX1 INVX1_2450 ( .A(_abc_17692_n12847), .Y(_abc_17692_n12850) );
  INVX1 INVX1_2451 ( .A(_abc_17692_n12853), .Y(_abc_17692_n12854) );
  INVX1 INVX1_2452 ( .A(_abc_17692_n12856), .Y(_abc_17692_n12857) );
  INVX1 INVX1_2453 ( .A(_abc_17692_n12860), .Y(_abc_17692_n12862) );
  INVX1 INVX1_2454 ( .A(_abc_17692_n12684), .Y(_abc_17692_n12866) );
  INVX1 INVX1_2455 ( .A(_abc_17692_n12867), .Y(_abc_17692_n12868) );
  INVX1 INVX1_2456 ( .A(_abc_17692_n12871), .Y(_abc_17692_n12872) );
  INVX1 INVX1_2457 ( .A(_abc_17692_n12878), .Y(_abc_17692_n12879) );
  INVX1 INVX1_2458 ( .A(_abc_17692_n12882), .Y(_abc_17692_n12884) );
  INVX1 INVX1_2459 ( .A(_abc_17692_n12888), .Y(_abc_17692_n12889) );
  INVX1 INVX1_246 ( .A(_abc_17692_n1769), .Y(_abc_17692_n1770) );
  INVX1 INVX1_2460 ( .A(_abc_17692_n12892), .Y(_abc_17692_n12894) );
  INVX1 INVX1_2461 ( .A(_abc_17692_n12737), .Y(_abc_17692_n12903) );
  INVX1 INVX1_2462 ( .A(_abc_17692_n12911), .Y(_abc_17692_n12912) );
  INVX1 INVX1_2463 ( .A(_abc_17692_n12913), .Y(_abc_17692_n12914) );
  INVX1 INVX1_2464 ( .A(_abc_17692_n12919), .Y(_abc_17692_n12920) );
  INVX1 INVX1_2465 ( .A(_abc_17692_n12662), .Y(_abc_17692_n12925) );
  INVX1 INVX1_2466 ( .A(_abc_17692_n12926), .Y(_abc_17692_n12927) );
  INVX1 INVX1_2467 ( .A(_abc_17692_n709), .Y(_abc_17692_n12941) );
  INVX1 INVX1_2468 ( .A(_abc_17692_n12942), .Y(_abc_17692_n12943) );
  INVX1 INVX1_2469 ( .A(modereg), .Y(_abc_17692_n12955) );
  INVX1 INVX1_247 ( .A(_abc_17692_n1773), .Y(_abc_17692_n1774) );
  INVX1 INVX1_248 ( .A(_abc_17692_n1782), .Y(_abc_17692_n1783) );
  INVX1 INVX1_249 ( .A(delta_31_), .Y(_abc_17692_n1790) );
  INVX1 INVX1_25 ( .A(_abc_17692_n933), .Y(_abc_17692_n934) );
  INVX1 INVX1_250 ( .A(_abc_17692_n1794), .Y(_abc_17692_n1795) );
  INVX1 INVX1_251 ( .A(_abc_17692_n1763), .Y(_abc_17692_n1796) );
  INVX1 INVX1_252 ( .A(_abc_17692_n1797), .Y(_abc_17692_n1798) );
  INVX1 INVX1_253 ( .A(_abc_17692_n1804_1), .Y(_abc_17692_n1805) );
  INVX1 INVX1_254 ( .A(_abc_17692_n1820), .Y(_abc_17692_n1821) );
  INVX1 INVX1_255 ( .A(_abc_17692_n1823), .Y(_abc_17692_n1824) );
  INVX1 INVX1_256 ( .A(_abc_17692_n1819), .Y(_abc_17692_n1826) );
  INVX1 INVX1_257 ( .A(_abc_17692_n1828), .Y(_abc_17692_n1831) );
  INVX1 INVX1_258 ( .A(_abc_17692_n1835), .Y(_abc_17692_n1836) );
  INVX1 INVX1_259 ( .A(_abc_17692_n1838), .Y(_abc_17692_n1839) );
  INVX1 INVX1_26 ( .A(_abc_17692_n930_1), .Y(_abc_17692_n940) );
  INVX1 INVX1_260 ( .A(_abc_17692_n1842), .Y(_abc_17692_n1843) );
  INVX1 INVX1_261 ( .A(selectslice_0_), .Y(_abc_17692_n1845) );
  INVX1 INVX1_262 ( .A(_abc_17692_n1851), .Y(_abc_17692_n1852_1) );
  INVX1 INVX1_263 ( .A(_abc_17692_n1854), .Y(_abc_17692_n1855_1) );
  INVX1 INVX1_264 ( .A(_abc_17692_n1858), .Y(_abc_17692_n1859) );
  INVX1 INVX1_265 ( .A(_abc_17692_n1860), .Y(_abc_17692_n1861) );
  INVX1 INVX1_266 ( .A(selectslice_1_), .Y(_abc_17692_n1862) );
  INVX1 INVX1_267 ( .A(_abc_17692_n1867_1), .Y(_abc_17692_n1868) );
  INVX1 INVX1_268 ( .A(_abc_17692_n1870), .Y(_abc_17692_n1871) );
  INVX1 INVX1_269 ( .A(_abc_17692_n1874), .Y(_abc_17692_n1875) );
  INVX1 INVX1_27 ( .A(sum_2_), .Y(_abc_17692_n946) );
  INVX1 INVX1_270 ( .A(_abc_17692_n1878), .Y(_abc_17692_n1879) );
  INVX1 INVX1_271 ( .A(_abc_17692_n1815_1), .Y(_abc_17692_n1890) );
  INVX1 INVX1_272 ( .A(_abc_17692_n1892), .Y(_abc_17692_n1893) );
  INVX1 INVX1_273 ( .A(_abc_17692_n1891), .Y(_abc_17692_n1896) );
  INVX1 INVX1_274 ( .A(_abc_17692_n1900), .Y(_abc_17692_n1901_1) );
  INVX1 INVX1_275 ( .A(_abc_17692_n1902), .Y(_abc_17692_n1905) );
  INVX1 INVX1_276 ( .A(_abc_17692_n1925), .Y(_abc_17692_n1926) );
  INVX1 INVX1_277 ( .A(_abc_17692_n1928), .Y(_abc_17692_n1929) );
  INVX1 INVX1_278 ( .A(_abc_17692_n1932), .Y(_abc_17692_n1933) );
  INVX1 INVX1_279 ( .A(_abc_17692_n1934), .Y(_abc_17692_n1935) );
  INVX1 INVX1_28 ( .A(_abc_17692_n947), .Y(_abc_17692_n948) );
  INVX1 INVX1_280 ( .A(_abc_17692_n1936), .Y(_abc_17692_n1939) );
  INVX1 INVX1_281 ( .A(_abc_17692_n1962), .Y(_abc_17692_n1963) );
  INVX1 INVX1_282 ( .A(_abc_17692_n1964), .Y(_abc_17692_n1965) );
  INVX1 INVX1_283 ( .A(sum_1_), .Y(_abc_17692_n1969) );
  INVX1 INVX1_284 ( .A(\key_in[33] ), .Y(_abc_17692_n1970) );
  INVX1 INVX1_285 ( .A(_abc_17692_n1987), .Y(_abc_17692_n1988) );
  INVX1 INVX1_286 ( .A(_abc_17692_n1995), .Y(_abc_17692_n1996) );
  INVX1 INVX1_287 ( .A(_abc_17692_n1999), .Y(_abc_17692_n2000) );
  INVX1 INVX1_288 ( .A(_abc_17692_n1997), .Y(_abc_17692_n2004_1) );
  INVX1 INVX1_289 ( .A(_abc_17692_n1994), .Y(_abc_17692_n2017) );
  INVX1 INVX1_29 ( .A(_abc_17692_n950), .Y(_abc_17692_n951) );
  INVX1 INVX1_290 ( .A(_abc_17692_n1829), .Y(_abc_17692_n2033) );
  INVX1 INVX1_291 ( .A(_abc_17692_n2034), .Y(_abc_17692_n2035) );
  INVX1 INVX1_292 ( .A(_abc_17692_n1847), .Y(_abc_17692_n2045) );
  INVX1 INVX1_293 ( .A(_abc_17692_n2065), .Y(_abc_17692_n2066) );
  INVX1 INVX1_294 ( .A(_abc_17692_n2072), .Y(_abc_17692_n2073) );
  INVX1 INVX1_295 ( .A(_abc_17692_n2075), .Y(_abc_17692_n2076) );
  INVX1 INVX1_296 ( .A(_abc_17692_n2099), .Y(_abc_17692_n2100) );
  INVX1 INVX1_297 ( .A(_abc_17692_n2105), .Y(_abc_17692_n2106) );
  INVX1 INVX1_298 ( .A(_abc_17692_n2108), .Y(_abc_17692_n2111) );
  INVX1 INVX1_299 ( .A(_abc_17692_n2128), .Y(_abc_17692_n2129) );
  INVX1 INVX1_3 ( .A(state_10_bF_buf4), .Y(_abc_17692_n627) );
  INVX1 INVX1_30 ( .A(_abc_17692_n952), .Y(_abc_17692_n953) );
  INVX1 INVX1_300 ( .A(_abc_17692_n2134), .Y(_abc_17692_n2135) );
  INVX1 INVX1_301 ( .A(_abc_17692_n2138), .Y(_abc_17692_n2139) );
  INVX1 INVX1_302 ( .A(_abc_17692_n2137_1), .Y(_abc_17692_n2144) );
  INVX1 INVX1_303 ( .A(_abc_17692_n2155), .Y(_abc_17692_n2156) );
  INVX1 INVX1_304 ( .A(_abc_17692_n2170), .Y(_abc_17692_n2171) );
  INVX1 INVX1_305 ( .A(_abc_17692_n2174), .Y(_abc_17692_n2175) );
  INVX1 INVX1_306 ( .A(_abc_17692_n2173), .Y(_abc_17692_n2180) );
  INVX1 INVX1_307 ( .A(_abc_17692_n2191), .Y(_abc_17692_n2192) );
  INVX1 INVX1_308 ( .A(_abc_17692_n2193), .Y(_abc_17692_n2198) );
  INVX1 INVX1_309 ( .A(_abc_17692_n2215), .Y(_abc_17692_n2216) );
  INVX1 INVX1_31 ( .A(_abc_17692_n954), .Y(_abc_17692_n955) );
  INVX1 INVX1_310 ( .A(_abc_17692_n2061), .Y(_abc_17692_n2254) );
  INVX1 INVX1_311 ( .A(_abc_17692_n2252), .Y(_abc_17692_n2256) );
  INVX1 INVX1_312 ( .A(_abc_17692_n2260), .Y(_abc_17692_n2261) );
  INVX1 INVX1_313 ( .A(_abc_17692_n2263), .Y(_abc_17692_n2264) );
  INVX1 INVX1_314 ( .A(_abc_17692_n2284), .Y(_abc_17692_n2285) );
  INVX1 INVX1_315 ( .A(_abc_17692_n2294), .Y(_abc_17692_n2295) );
  INVX1 INVX1_316 ( .A(_abc_17692_n2297), .Y(_abc_17692_n2298) );
  INVX1 INVX1_317 ( .A(_abc_17692_n2095), .Y(_abc_17692_n2315) );
  INVX1 INVX1_318 ( .A(_abc_17692_n2317), .Y(_abc_17692_n2318) );
  INVX1 INVX1_319 ( .A(_abc_17692_n2323), .Y(_abc_17692_n2324) );
  INVX1 INVX1_32 ( .A(_abc_17692_n962), .Y(_abc_17692_n963) );
  INVX1 INVX1_320 ( .A(_abc_17692_n2326_1), .Y(_abc_17692_n2329_1) );
  INVX1 INVX1_321 ( .A(_abc_17692_n2330), .Y(_abc_17692_n2334) );
  INVX1 INVX1_322 ( .A(_abc_17692_n2159), .Y(_abc_17692_n2349) );
  INVX1 INVX1_323 ( .A(_abc_17692_n2358), .Y(_abc_17692_n2359) );
  INVX1 INVX1_324 ( .A(_abc_17692_n2361_1), .Y(_abc_17692_n2364) );
  INVX1 INVX1_325 ( .A(_abc_17692_n2362), .Y(_abc_17692_n2368) );
  INVX1 INVX1_326 ( .A(_abc_17692_n2379), .Y(_abc_17692_n2380_1) );
  INVX1 INVX1_327 ( .A(_abc_17692_n2204), .Y(_abc_17692_n2393) );
  INVX1 INVX1_328 ( .A(_abc_17692_n2149), .Y(_abc_17692_n2401) );
  INVX1 INVX1_329 ( .A(_abc_17692_n2403), .Y(_abc_17692_n2404) );
  INVX1 INVX1_33 ( .A(sum_3_), .Y(_abc_17692_n969) );
  INVX1 INVX1_330 ( .A(_abc_17692_n2185), .Y(_abc_17692_n2411) );
  INVX1 INVX1_331 ( .A(_abc_17692_n2230), .Y(_abc_17692_n2419) );
  INVX1 INVX1_332 ( .A(_abc_17692_n2445), .Y(_abc_17692_n2453) );
  INVX1 INVX1_333 ( .A(_abc_17692_n2446), .Y(_abc_17692_n2454) );
  INVX1 INVX1_334 ( .A(_abc_17692_n2465), .Y(_abc_17692_n2466) );
  INVX1 INVX1_335 ( .A(_abc_17692_n2461), .Y(_abc_17692_n2470) );
  INVX1 INVX1_336 ( .A(_abc_17692_n2462_1), .Y(_abc_17692_n2471) );
  INVX1 INVX1_337 ( .A(_abc_17692_n2468), .Y(_abc_17692_n2474) );
  INVX1 INVX1_338 ( .A(_abc_17692_n2476), .Y(_abc_17692_n2478) );
  INVX1 INVX1_339 ( .A(_abc_17692_n2480), .Y(_abc_17692_n2483) );
  INVX1 INVX1_34 ( .A(_abc_17692_n970), .Y(_abc_17692_n971) );
  INVX1 INVX1_340 ( .A(_abc_17692_n2485), .Y(_abc_17692_n2486) );
  INVX1 INVX1_341 ( .A(_abc_17692_n2346), .Y(_abc_17692_n2489) );
  INVX1 INVX1_342 ( .A(_abc_17692_n2495), .Y(_abc_17692_n2496) );
  INVX1 INVX1_343 ( .A(_abc_17692_n2498), .Y(_abc_17692_n2505) );
  INVX1 INVX1_344 ( .A(_abc_17692_n2503), .Y(_abc_17692_n2506) );
  INVX1 INVX1_345 ( .A(_abc_17692_n2508), .Y(_abc_17692_n2510) );
  INVX1 INVX1_346 ( .A(_abc_17692_n2512), .Y(_abc_17692_n2514) );
  INVX1 INVX1_347 ( .A(_abc_17692_n2516), .Y(_abc_17692_n2517) );
  INVX1 INVX1_348 ( .A(_abc_17692_n2309), .Y(_abc_17692_n2518) );
  INVX1 INVX1_349 ( .A(_abc_17692_n2521), .Y(_abc_17692_n2522) );
  INVX1 INVX1_35 ( .A(delta_3_), .Y(_abc_17692_n972_1) );
  INVX1 INVX1_350 ( .A(_abc_17692_n2530), .Y(_abc_17692_n2531) );
  INVX1 INVX1_351 ( .A(_abc_17692_n2526), .Y(_abc_17692_n2535_1) );
  INVX1 INVX1_352 ( .A(_abc_17692_n2527), .Y(_abc_17692_n2536) );
  INVX1 INVX1_353 ( .A(_abc_17692_n2533), .Y(_abc_17692_n2539) );
  INVX1 INVX1_354 ( .A(_abc_17692_n2541), .Y(_abc_17692_n2543) );
  INVX1 INVX1_355 ( .A(_abc_17692_n2545), .Y(_abc_17692_n2547) );
  INVX1 INVX1_356 ( .A(_abc_17692_n2550), .Y(_abc_17692_n2551) );
  INVX1 INVX1_357 ( .A(_abc_17692_n2552_1), .Y(_abc_17692_n2553) );
  INVX1 INVX1_358 ( .A(_abc_17692_n2560), .Y(_abc_17692_n2561) );
  INVX1 INVX1_359 ( .A(_abc_17692_n2564), .Y(_abc_17692_n2565) );
  INVX1 INVX1_36 ( .A(_abc_17692_n973), .Y(_abc_17692_n974) );
  INVX1 INVX1_360 ( .A(_abc_17692_n2563), .Y(_abc_17692_n2570) );
  INVX1 INVX1_361 ( .A(_abc_17692_n2581_1), .Y(_abc_17692_n2586) );
  INVX1 INVX1_362 ( .A(_abc_17692_n2390), .Y(_abc_17692_n2592) );
  INVX1 INVX1_363 ( .A(_abc_17692_n2338), .Y(_abc_17692_n2600) );
  INVX1 INVX1_364 ( .A(_abc_17692_n2602), .Y(_abc_17692_n2603) );
  INVX1 INVX1_365 ( .A(_abc_17692_n2382), .Y(_abc_17692_n2610) );
  INVX1 INVX1_366 ( .A(_abc_17692_n2549), .Y(_abc_17692_n2618) );
  INVX1 INVX1_367 ( .A(_abc_17692_n2287), .Y(_abc_17692_n2619) );
  INVX1 INVX1_368 ( .A(workunit1_1_bF_buf3), .Y(_abc_17692_n2637) );
  INVX1 INVX1_369 ( .A(_abc_17692_n2636), .Y(_abc_17692_n2642) );
  INVX1 INVX1_37 ( .A(_abc_17692_n949_1), .Y(_abc_17692_n976) );
  INVX1 INVX1_370 ( .A(_abc_17692_n2655), .Y(_abc_17692_n2656) );
  INVX1 INVX1_371 ( .A(_abc_17692_n2658), .Y(_abc_17692_n2659) );
  INVX1 INVX1_372 ( .A(_abc_17692_n2661), .Y(_abc_17692_n2662) );
  INVX1 INVX1_373 ( .A(_abc_17692_n2663), .Y(_abc_17692_n2664) );
  INVX1 INVX1_374 ( .A(_abc_17692_n2670), .Y(_abc_17692_n2671) );
  INVX1 INVX1_375 ( .A(_abc_17692_n2675), .Y(_abc_17692_n2676) );
  INVX1 INVX1_376 ( .A(_abc_17692_n2678), .Y(_abc_17692_n2679) );
  INVX1 INVX1_377 ( .A(\key_in[5] ), .Y(_abc_17692_n2685) );
  INVX1 INVX1_378 ( .A(_abc_17692_n2689), .Y(_abc_17692_n2690) );
  INVX1 INVX1_379 ( .A(_abc_17692_n2691), .Y(_abc_17692_n2693) );
  INVX1 INVX1_38 ( .A(_abc_17692_n975), .Y(_abc_17692_n979) );
  INVX1 INVX1_380 ( .A(_abc_17692_n2695), .Y(_abc_17692_n2697) );
  INVX1 INVX1_381 ( .A(_abc_17692_n2699), .Y(_abc_17692_n2700) );
  INVX1 INVX1_382 ( .A(_abc_17692_n2701), .Y(_abc_17692_n2702) );
  INVX1 INVX1_383 ( .A(\key_in[37] ), .Y(_abc_17692_n2713_1) );
  INVX1 INVX1_384 ( .A(_abc_17692_n2715), .Y(_abc_17692_n2716_1) );
  INVX1 INVX1_385 ( .A(_abc_17692_n2732), .Y(_abc_17692_n2733) );
  INVX1 INVX1_386 ( .A(_abc_17692_n2737), .Y(_abc_17692_n2738) );
  INVX1 INVX1_387 ( .A(_abc_17692_n2744), .Y(_abc_17692_n2745_1) );
  INVX1 INVX1_388 ( .A(_abc_17692_n2747), .Y(_abc_17692_n2750) );
  INVX1 INVX1_389 ( .A(_abc_17692_n2751), .Y(_abc_17692_n2755) );
  INVX1 INVX1_39 ( .A(_abc_17692_n977), .Y(_abc_17692_n980_1) );
  INVX1 INVX1_390 ( .A(_abc_17692_n2765), .Y(_abc_17692_n2770) );
  INVX1 INVX1_391 ( .A(_abc_17692_n2674), .Y(_abc_17692_n2776) );
  INVX1 INVX1_392 ( .A(_abc_17692_n2513), .Y(_abc_17692_n2777) );
  INVX1 INVX1_393 ( .A(_abc_17692_n2786), .Y(_abc_17692_n2787) );
  INVX1 INVX1_394 ( .A(_abc_17692_n2575), .Y(_abc_17692_n2794) );
  INVX1 INVX1_395 ( .A(_abc_17692_n2546), .Y(_abc_17692_n2800_1) );
  INVX1 INVX1_396 ( .A(_abc_17692_n2822), .Y(_abc_17692_n2827) );
  INVX1 INVX1_397 ( .A(_abc_17692_n2817), .Y(_abc_17692_n2833) );
  INVX1 INVX1_398 ( .A(_abc_17692_n2841), .Y(_abc_17692_n2842) );
  INVX1 INVX1_399 ( .A(_abc_17692_n2846), .Y(_abc_17692_n2847) );
  INVX1 INVX1_4 ( .A(_abc_17692_n628), .Y(_abc_17692_n629) );
  INVX1 INVX1_40 ( .A(_abc_17692_n985), .Y(_abc_17692_n986) );
  INVX1 INVX1_400 ( .A(_abc_17692_n2849_1), .Y(_abc_17692_n2850) );
  INVX1 INVX1_401 ( .A(_abc_17692_n2853), .Y(_abc_17692_n2854) );
  INVX1 INVX1_402 ( .A(_abc_17692_n2856), .Y(_abc_17692_n2857) );
  INVX1 INVX1_403 ( .A(_abc_17692_n2860), .Y(_abc_17692_n2863) );
  INVX1 INVX1_404 ( .A(_abc_17692_n2672), .Y(_abc_17692_n2866) );
  INVX1 INVX1_405 ( .A(_abc_17692_n2869), .Y(_abc_17692_n2870) );
  INVX1 INVX1_406 ( .A(_abc_17692_n2873), .Y(_abc_17692_n2874) );
  INVX1 INVX1_407 ( .A(_abc_17692_n2686), .Y(_abc_17692_n2876) );
  INVX1 INVX1_408 ( .A(_abc_17692_n2880), .Y(_abc_17692_n2881) );
  INVX1 INVX1_409 ( .A(_abc_17692_n2879), .Y(_abc_17692_n2885) );
  INVX1 INVX1_41 ( .A(_abc_17692_n987), .Y(_abc_17692_n988_1) );
  INVX1 INVX1_410 ( .A(_abc_17692_n2883), .Y(_abc_17692_n2886) );
  INVX1 INVX1_411 ( .A(_abc_17692_n2888), .Y(_abc_17692_n2890) );
  INVX1 INVX1_412 ( .A(_abc_17692_n2893), .Y(_abc_17692_n2894) );
  INVX1 INVX1_413 ( .A(_abc_17692_n2896), .Y(_abc_17692_n2899) );
  INVX1 INVX1_414 ( .A(_abc_17692_n2696), .Y(_abc_17692_n2900) );
  INVX1 INVX1_415 ( .A(_abc_17692_n2714), .Y(_abc_17692_n2908) );
  INVX1 INVX1_416 ( .A(_abc_17692_n2912), .Y(_abc_17692_n2913) );
  INVX1 INVX1_417 ( .A(_abc_17692_n2906), .Y(_abc_17692_n2917) );
  INVX1 INVX1_418 ( .A(_abc_17692_n2910), .Y(_abc_17692_n2919_1) );
  INVX1 INVX1_419 ( .A(_abc_17692_n2915), .Y(_abc_17692_n2921) );
  INVX1 INVX1_42 ( .A(sum_4_), .Y(_abc_17692_n995) );
  INVX1 INVX1_420 ( .A(_abc_17692_n2923), .Y(_abc_17692_n2925) );
  INVX1 INVX1_421 ( .A(_abc_17692_n2927), .Y(_abc_17692_n2928) );
  INVX1 INVX1_422 ( .A(_abc_17692_n2931), .Y(_abc_17692_n2932) );
  INVX1 INVX1_423 ( .A(_abc_17692_n2935), .Y(_abc_17692_n2936) );
  INVX1 INVX1_424 ( .A(_abc_17692_n2734_1), .Y(_abc_17692_n2937) );
  INVX1 INVX1_425 ( .A(_abc_17692_n2940), .Y(_abc_17692_n2941) );
  INVX1 INVX1_426 ( .A(_abc_17692_n2943), .Y(_abc_17692_n2944) );
  INVX1 INVX1_427 ( .A(_abc_17692_n2952), .Y(_abc_17692_n2953) );
  INVX1 INVX1_428 ( .A(_abc_17692_n2955), .Y(_abc_17692_n2956) );
  INVX1 INVX1_429 ( .A(_abc_17692_n2959), .Y(_abc_17692_n2960_1) );
  INVX1 INVX1_43 ( .A(_abc_17692_n997), .Y(_abc_17692_n998) );
  INVX1 INVX1_430 ( .A(_abc_17692_n2962), .Y(_abc_17692_n2963) );
  INVX1 INVX1_431 ( .A(_abc_17692_n2966), .Y(_abc_17692_n2968) );
  INVX1 INVX1_432 ( .A(_abc_17692_n2971), .Y(_abc_17692_n2972) );
  INVX1 INVX1_433 ( .A(_abc_17692_n2970), .Y(_abc_17692_n2974) );
  INVX1 INVX1_434 ( .A(_abc_17692_n2980), .Y(_abc_17692_n2981) );
  INVX1 INVX1_435 ( .A(_abc_17692_n2983), .Y(_abc_17692_n2984) );
  INVX1 INVX1_436 ( .A(_abc_17692_n2727), .Y(_abc_17692_n2988) );
  INVX1 INVX1_437 ( .A(_abc_17692_n2992), .Y(_abc_17692_n2993) );
  INVX1 INVX1_438 ( .A(_abc_17692_n2759), .Y(_abc_17692_n2999) );
  INVX1 INVX1_439 ( .A(_abc_17692_n2865), .Y(_abc_17692_n3008) );
  INVX1 INVX1_44 ( .A(_abc_17692_n1000), .Y(_abc_17692_n1001) );
  INVX1 INVX1_440 ( .A(_abc_17692_n3005), .Y(_abc_17692_n3009_1) );
  INVX1 INVX1_441 ( .A(_abc_17692_n2832), .Y(_abc_17692_n3023) );
  INVX1 INVX1_442 ( .A(workunit1_12_bF_buf1), .Y(_abc_17692_n3026) );
  INVX1 INVX1_443 ( .A(_abc_17692_n3025), .Y(_abc_17692_n3030) );
  INVX1 INVX1_444 ( .A(_abc_17692_n3042), .Y(_abc_17692_n3043) );
  INVX1 INVX1_445 ( .A(_abc_17692_n3044), .Y(_abc_17692_n3045) );
  INVX1 INVX1_446 ( .A(_abc_17692_n3047), .Y(_abc_17692_n3049) );
  INVX1 INVX1_447 ( .A(_abc_17692_n3040), .Y(_abc_17692_n3054) );
  INVX1 INVX1_448 ( .A(_abc_17692_n3051), .Y(_abc_17692_n3056) );
  INVX1 INVX1_449 ( .A(_abc_17692_n3058_1), .Y(_abc_17692_n3061) );
  INVX1 INVX1_45 ( .A(_abc_17692_n1004), .Y(_abc_17692_n1005) );
  INVX1 INVX1_450 ( .A(_abc_17692_n3063), .Y(_abc_17692_n3064) );
  INVX1 INVX1_451 ( .A(_abc_17692_n3066), .Y(_abc_17692_n3067) );
  INVX1 INVX1_452 ( .A(_abc_17692_n3073), .Y(_abc_17692_n3074) );
  INVX1 INVX1_453 ( .A(_abc_17692_n3076), .Y(_abc_17692_n3077) );
  INVX1 INVX1_454 ( .A(_abc_17692_n3079), .Y(_abc_17692_n3080_1) );
  INVX1 INVX1_455 ( .A(_abc_17692_n3081), .Y(_abc_17692_n3082) );
  INVX1 INVX1_456 ( .A(_abc_17692_n3085), .Y(_abc_17692_n3086) );
  INVX1 INVX1_457 ( .A(_abc_17692_n3089), .Y(_abc_17692_n3090) );
  INVX1 INVX1_458 ( .A(_abc_17692_n3092), .Y(_abc_17692_n3093) );
  INVX1 INVX1_459 ( .A(_abc_17692_n3100), .Y(_abc_17692_n3101) );
  INVX1 INVX1_46 ( .A(_abc_17692_n999), .Y(_abc_17692_n1007) );
  INVX1 INVX1_460 ( .A(_abc_17692_n3103), .Y(_abc_17692_n3106) );
  INVX1 INVX1_461 ( .A(_abc_17692_n3120), .Y(_abc_17692_n3121) );
  INVX1 INVX1_462 ( .A(_abc_17692_n3122), .Y(_abc_17692_n3123) );
  INVX1 INVX1_463 ( .A(_abc_17692_n3124), .Y(_abc_17692_n3125) );
  INVX1 INVX1_464 ( .A(_abc_17692_n3133), .Y(_abc_17692_n3134) );
  INVX1 INVX1_465 ( .A(_abc_17692_n3136), .Y(_abc_17692_n3137) );
  INVX1 INVX1_466 ( .A(_abc_17692_n3139), .Y(_abc_17692_n3140) );
  INVX1 INVX1_467 ( .A(_abc_17692_n3141_1), .Y(_abc_17692_n3142) );
  INVX1 INVX1_468 ( .A(_abc_17692_n3145), .Y(_abc_17692_n3146) );
  INVX1 INVX1_469 ( .A(_abc_17692_n3150), .Y(_abc_17692_n3151) );
  INVX1 INVX1_47 ( .A(_abc_17692_n1014), .Y(_abc_17692_n1015) );
  INVX1 INVX1_470 ( .A(_abc_17692_n3149), .Y(_abc_17692_n3153_1) );
  INVX1 INVX1_471 ( .A(_abc_17692_n3159), .Y(_abc_17692_n3161) );
  INVX1 INVX1_472 ( .A(_abc_17692_n3165), .Y(_abc_17692_n3166_1) );
  INVX1 INVX1_473 ( .A(_abc_17692_n3172), .Y(_abc_17692_n3173) );
  INVX1 INVX1_474 ( .A(_abc_17692_n2861), .Y(_abc_17692_n3184) );
  INVX1 INVX1_475 ( .A(_abc_17692_n3204), .Y(_abc_17692_n3205) );
  INVX1 INVX1_476 ( .A(_abc_17692_n3217), .Y(_abc_17692_n3218) );
  INVX1 INVX1_477 ( .A(_abc_17692_n3237), .Y(_abc_17692_n3238) );
  INVX1 INVX1_478 ( .A(_abc_17692_n3236), .Y(_abc_17692_n3242) );
  INVX1 INVX1_479 ( .A(_abc_17692_n3240_1), .Y(_abc_17692_n3243) );
  INVX1 INVX1_48 ( .A(_abc_17692_n1021), .Y(_abc_17692_n1022) );
  INVX1 INVX1_480 ( .A(_abc_17692_n3245), .Y(_abc_17692_n3246) );
  INVX1 INVX1_481 ( .A(_abc_17692_n3228), .Y(_abc_17692_n3248) );
  INVX1 INVX1_482 ( .A(_abc_17692_n3250), .Y(_abc_17692_n3251) );
  INVX1 INVX1_483 ( .A(_abc_17692_n3254), .Y(_abc_17692_n3255) );
  INVX1 INVX1_484 ( .A(_abc_17692_n3087), .Y(_abc_17692_n3256) );
  INVX1 INVX1_485 ( .A(_abc_17692_n3260), .Y(_abc_17692_n3261) );
  INVX1 INVX1_486 ( .A(_abc_17692_n3115), .Y(_abc_17692_n3264) );
  INVX1 INVX1_487 ( .A(_abc_17692_n3269), .Y(_abc_17692_n3270) );
  INVX1 INVX1_488 ( .A(_abc_17692_n3279), .Y(_abc_17692_n3280) );
  INVX1 INVX1_489 ( .A(_abc_17692_n3272), .Y(_abc_17692_n3284) );
  INVX1 INVX1_49 ( .A(delta_5_), .Y(_abc_17692_n1023) );
  INVX1 INVX1_490 ( .A(_abc_17692_n3277), .Y(_abc_17692_n3286) );
  INVX1 INVX1_491 ( .A(_abc_17692_n3282), .Y(_abc_17692_n3288) );
  INVX1 INVX1_492 ( .A(_abc_17692_n3290), .Y(_abc_17692_n3291) );
  INVX1 INVX1_493 ( .A(_abc_17692_n3295_1), .Y(_abc_17692_n3296) );
  INVX1 INVX1_494 ( .A(_abc_17692_n3300), .Y(_abc_17692_n3301) );
  INVX1 INVX1_495 ( .A(_abc_17692_n3312), .Y(_abc_17692_n3313) );
  INVX1 INVX1_496 ( .A(_abc_17692_n3305), .Y(_abc_17692_n3317) );
  INVX1 INVX1_497 ( .A(_abc_17692_n3310), .Y(_abc_17692_n3319) );
  INVX1 INVX1_498 ( .A(_abc_17692_n3315), .Y(_abc_17692_n3321) );
  INVX1 INVX1_499 ( .A(_abc_17692_n3323), .Y(_abc_17692_n3324) );
  INVX1 INVX1_5 ( .A(_abc_17692_n667), .Y(_abc_17692_n668) );
  INVX1 INVX1_50 ( .A(sum_5_), .Y(_abc_17692_n1024) );
  INVX1 INVX1_500 ( .A(_abc_17692_n3328), .Y(_abc_17692_n3329) );
  INVX1 INVX1_501 ( .A(_abc_17692_n3062), .Y(_abc_17692_n3332) );
  INVX1 INVX1_502 ( .A(_abc_17692_n3059), .Y(_abc_17692_n3334) );
  INVX1 INVX1_503 ( .A(_abc_17692_n3335), .Y(_abc_17692_n3336) );
  INVX1 INVX1_504 ( .A(_abc_17692_n3340), .Y(_abc_17692_n3341) );
  INVX1 INVX1_505 ( .A(_abc_17692_n3346_1), .Y(_abc_17692_n3347) );
  INVX1 INVX1_506 ( .A(_abc_17692_n3348), .Y(_abc_17692_n3349_1) );
  INVX1 INVX1_507 ( .A(_abc_17692_n3351), .Y(_abc_17692_n3361) );
  INVX1 INVX1_508 ( .A(_abc_17692_n3356), .Y(_abc_17692_n3362) );
  INVX1 INVX1_509 ( .A(_abc_17692_n3358), .Y(_abc_17692_n3363) );
  INVX1 INVX1_51 ( .A(_abc_17692_n1025_1), .Y(_abc_17692_n1026) );
  INVX1 INVX1_510 ( .A(_abc_17692_n3366_1), .Y(_abc_17692_n3368) );
  INVX1 INVX1_511 ( .A(_abc_17692_n3371), .Y(_abc_17692_n3372) );
  INVX1 INVX1_512 ( .A(_abc_17692_n3376_1), .Y(_abc_17692_n3377) );
  INVX1 INVX1_513 ( .A(_abc_17692_n3374), .Y(_abc_17692_n3382) );
  INVX1 INVX1_514 ( .A(_abc_17692_n3383), .Y(_abc_17692_n3384) );
  INVX1 INVX1_515 ( .A(_abc_17692_n3388_1), .Y(_abc_17692_n3389) );
  INVX1 INVX1_516 ( .A(_abc_17692_n3393), .Y(_abc_17692_n3394) );
  INVX1 INVX1_517 ( .A(_abc_17692_n3395), .Y(_abc_17692_n3396) );
  INVX1 INVX1_518 ( .A(_abc_17692_n3398), .Y(_abc_17692_n3399) );
  INVX1 INVX1_519 ( .A(_abc_17692_n3298), .Y(_abc_17692_n3403) );
  INVX1 INVX1_52 ( .A(_abc_17692_n1027), .Y(_abc_17692_n1028_1) );
  INVX1 INVX1_520 ( .A(_abc_17692_n2929), .Y(_abc_17692_n3405) );
  INVX1 INVX1_521 ( .A(_abc_17692_n3412), .Y(_abc_17692_n3413) );
  INVX1 INVX1_522 ( .A(_abc_17692_n3331), .Y(_abc_17692_n3416) );
  INVX1 INVX1_523 ( .A(_abc_17692_n3423), .Y(_abc_17692_n3424_1) );
  INVX1 INVX1_524 ( .A(_abc_17692_n3253), .Y(_abc_17692_n3437) );
  INVX1 INVX1_525 ( .A(_abc_17692_n3439), .Y(_abc_17692_n3440) );
  INVX1 INVX1_526 ( .A(_abc_17692_n3441), .Y(_abc_17692_n3442) );
  INVX1 INVX1_527 ( .A(_abc_17692_n3443), .Y(_abc_17692_n3446) );
  INVX1 INVX1_528 ( .A(_abc_17692_n3449), .Y(_abc_17692_n3450) );
  INVX1 INVX1_529 ( .A(_abc_17692_n3454), .Y(_abc_17692_n3455) );
  INVX1 INVX1_53 ( .A(_abc_17692_n1029), .Y(_abc_17692_n1030) );
  INVX1 INVX1_530 ( .A(_abc_17692_n3456), .Y(_abc_17692_n3457) );
  INVX1 INVX1_531 ( .A(_abc_17692_n3459), .Y(_abc_17692_n3461) );
  INVX1 INVX1_532 ( .A(_abc_17692_n3463), .Y(_abc_17692_n3466) );
  INVX1 INVX1_533 ( .A(_abc_17692_n3468), .Y(_abc_17692_n3469) );
  INVX1 INVX1_534 ( .A(_abc_17692_n3438), .Y(_abc_17692_n3475) );
  INVX1 INVX1_535 ( .A(_abc_17692_n3473), .Y(_abc_17692_n3476) );
  INVX1 INVX1_536 ( .A(_abc_17692_n3480), .Y(_abc_17692_n3481) );
  INVX1 INVX1_537 ( .A(_abc_17692_n3482), .Y(_abc_17692_n3483) );
  INVX1 INVX1_538 ( .A(_abc_17692_n3484), .Y(_abc_17692_n3485) );
  INVX1 INVX1_539 ( .A(_abc_17692_n3489), .Y(_abc_17692_n3490) );
  INVX1 INVX1_54 ( .A(_abc_17692_n1031), .Y(_abc_17692_n1033) );
  INVX1 INVX1_540 ( .A(_abc_17692_n3488), .Y(_abc_17692_n3493) );
  INVX1 INVX1_541 ( .A(_abc_17692_n3502), .Y(_abc_17692_n3503_1) );
  INVX1 INVX1_542 ( .A(_abc_17692_n3508), .Y(_abc_17692_n3509) );
  INVX1 INVX1_543 ( .A(_abc_17692_n3511), .Y(_abc_17692_n3512) );
  INVX1 INVX1_544 ( .A(_abc_17692_n3514), .Y(_abc_17692_n3515) );
  INVX1 INVX1_545 ( .A(_abc_17692_n3517), .Y(_abc_17692_n3518) );
  INVX1 INVX1_546 ( .A(_abc_17692_n3519), .Y(_abc_17692_n3521) );
  INVX1 INVX1_547 ( .A(_abc_17692_n3523), .Y(_abc_17692_n3524) );
  INVX1 INVX1_548 ( .A(_abc_17692_n3527), .Y(_abc_17692_n3528) );
  INVX1 INVX1_549 ( .A(_abc_17692_n3537), .Y(_abc_17692_n3538) );
  INVX1 INVX1_55 ( .A(_abc_17692_n1039), .Y(_abc_17692_n1040) );
  INVX1 INVX1_550 ( .A(_abc_17692_n3540), .Y(_abc_17692_n3541) );
  INVX1 INVX1_551 ( .A(_abc_17692_n3543), .Y(_abc_17692_n3544) );
  INVX1 INVX1_552 ( .A(_abc_17692_n3545), .Y(_abc_17692_n3547) );
  INVX1 INVX1_553 ( .A(_abc_17692_n3549), .Y(_abc_17692_n3550) );
  INVX1 INVX1_554 ( .A(_abc_17692_n3553), .Y(_abc_17692_n3554) );
  INVX1 INVX1_555 ( .A(_abc_17692_n3535), .Y(_abc_17692_n3556) );
  INVX1 INVX1_556 ( .A(_abc_17692_n3370), .Y(_abc_17692_n3562) );
  INVX1 INVX1_557 ( .A(_abc_17692_n3563), .Y(_abc_17692_n3564) );
  INVX1 INVX1_558 ( .A(_abc_17692_n3565), .Y(_abc_17692_n3566) );
  INVX1 INVX1_559 ( .A(_abc_17692_n3571), .Y(_abc_17692_n3572) );
  INVX1 INVX1_56 ( .A(sum_6_), .Y(_abc_17692_n1047) );
  INVX1 INVX1_560 ( .A(_abc_17692_n3573), .Y(_abc_17692_n3574) );
  INVX1 INVX1_561 ( .A(_abc_17692_n3327), .Y(_abc_17692_n3579) );
  INVX1 INVX1_562 ( .A(_abc_17692_n3580), .Y(_abc_17692_n3581) );
  INVX1 INVX1_563 ( .A(_abc_17692_n3582), .Y(_abc_17692_n3584) );
  INVX1 INVX1_564 ( .A(_abc_17692_n3294), .Y(_abc_17692_n3588) );
  INVX1 INVX1_565 ( .A(_abc_17692_n3589), .Y(_abc_17692_n3590) );
  INVX1 INVX1_566 ( .A(_abc_17692_n3591), .Y(_abc_17692_n3592) );
  INVX1 INVX1_567 ( .A(_abc_17692_n3606), .Y(_abc_17692_n3607) );
  INVX1 INVX1_568 ( .A(_abc_17692_n3448), .Y(_abc_17692_n3609) );
  INVX1 INVX1_569 ( .A(_abc_17692_n3445), .Y(_abc_17692_n3625) );
  INVX1 INVX1_57 ( .A(_abc_17692_n1049), .Y(_abc_17692_n1050) );
  INVX1 INVX1_570 ( .A(_abc_17692_n3458), .Y(_abc_17692_n3637) );
  INVX1 INVX1_571 ( .A(_abc_17692_n3639), .Y(_abc_17692_n3640_1) );
  INVX1 INVX1_572 ( .A(_abc_17692_n3642), .Y(_abc_17692_n3643) );
  INVX1 INVX1_573 ( .A(_abc_17692_n3641), .Y(_abc_17692_n3647) );
  INVX1 INVX1_574 ( .A(_abc_17692_n3645), .Y(_abc_17692_n3648) );
  INVX1 INVX1_575 ( .A(_abc_17692_n3650_1), .Y(_abc_17692_n3651) );
  INVX1 INVX1_576 ( .A(_abc_17692_n3634), .Y(_abc_17692_n3653) );
  INVX1 INVX1_577 ( .A(_abc_17692_n3656), .Y(_abc_17692_n3657) );
  INVX1 INVX1_578 ( .A(_abc_17692_n3258_1), .Y(_abc_17692_n3660) );
  INVX1 INVX1_579 ( .A(_abc_17692_n3661_1), .Y(_abc_17692_n3662) );
  INVX1 INVX1_58 ( .A(_abc_17692_n1051), .Y(_abc_17692_n1052) );
  INVX1 INVX1_580 ( .A(_abc_17692_n3666), .Y(_abc_17692_n3667) );
  INVX1 INVX1_581 ( .A(_abc_17692_n3668), .Y(_abc_17692_n3669) );
  INVX1 INVX1_582 ( .A(_abc_17692_n3671), .Y(_abc_17692_n3672) );
  INVX1 INVX1_583 ( .A(_abc_17692_n3680), .Y(_abc_17692_n3681) );
  INVX1 INVX1_584 ( .A(_abc_17692_n3676), .Y(_abc_17692_n3685) );
  INVX1 INVX1_585 ( .A(_abc_17692_n3678), .Y(_abc_17692_n3686) );
  INVX1 INVX1_586 ( .A(_abc_17692_n3683), .Y(_abc_17692_n3688) );
  INVX1 INVX1_587 ( .A(_abc_17692_n3690), .Y(_abc_17692_n3692) );
  INVX1 INVX1_588 ( .A(_abc_17692_n3695), .Y(_abc_17692_n3696_1) );
  INVX1 INVX1_589 ( .A(_abc_17692_n3698), .Y(_abc_17692_n3699_1) );
  INVX1 INVX1_59 ( .A(_abc_17692_n1056), .Y(_abc_17692_n1057_1) );
  INVX1 INVX1_590 ( .A(_abc_17692_n3702), .Y(_abc_17692_n3703) );
  INVX1 INVX1_591 ( .A(_abc_17692_n3706), .Y(_abc_17692_n3707) );
  INVX1 INVX1_592 ( .A(_abc_17692_n3708), .Y(_abc_17692_n3709) );
  INVX1 INVX1_593 ( .A(_abc_17692_n3718), .Y(_abc_17692_n3719) );
  INVX1 INVX1_594 ( .A(_abc_17692_n3717), .Y(_abc_17692_n3723) );
  INVX1 INVX1_595 ( .A(_abc_17692_n3721), .Y(_abc_17692_n3724) );
  INVX1 INVX1_596 ( .A(_abc_17692_n3726), .Y(_abc_17692_n3727) );
  INVX1 INVX1_597 ( .A(_abc_17692_n3732), .Y(_abc_17692_n3733_1) );
  INVX1 INVX1_598 ( .A(_abc_17692_n3735), .Y(_abc_17692_n3736) );
  INVX1 INVX1_599 ( .A(_abc_17692_n3738), .Y(_abc_17692_n3739) );
  INVX1 INVX1_6 ( .A(_abc_17692_n671), .Y(_abc_17692_n672) );
  INVX1 INVX1_60 ( .A(_abc_17692_n1062), .Y(_abc_17692_n1064) );
  INVX1 INVX1_600 ( .A(_abc_17692_n3741), .Y(_abc_17692_n3742) );
  INVX1 INVX1_601 ( .A(_abc_17692_n3744), .Y(_abc_17692_n3745) );
  INVX1 INVX1_602 ( .A(_abc_17692_n3539), .Y(_abc_17692_n3754_1) );
  INVX1 INVX1_603 ( .A(_abc_17692_n3756), .Y(_abc_17692_n3757) );
  INVX1 INVX1_604 ( .A(_abc_17692_n3759), .Y(_abc_17692_n3760) );
  INVX1 INVX1_605 ( .A(_abc_17692_n3758), .Y(_abc_17692_n3764) );
  INVX1 INVX1_606 ( .A(_abc_17692_n3762), .Y(_abc_17692_n3765) );
  INVX1 INVX1_607 ( .A(_abc_17692_n3767), .Y(_abc_17692_n3768) );
  INVX1 INVX1_608 ( .A(_abc_17692_n3771), .Y(_abc_17692_n3773) );
  INVX1 INVX1_609 ( .A(_abc_17692_n3775), .Y(_abc_17692_n3776_1) );
  INVX1 INVX1_61 ( .A(sum_7_), .Y(_abc_17692_n1070) );
  INVX1 INVX1_610 ( .A(_abc_17692_n3777), .Y(_abc_17692_n3778) );
  INVX1 INVX1_611 ( .A(_abc_17692_n3780), .Y(_abc_17692_n3781) );
  INVX1 INVX1_612 ( .A(_abc_17692_n3786), .Y(_abc_17692_n3787) );
  INVX1 INVX1_613 ( .A(_abc_17692_n3793), .Y(_abc_17692_n3794) );
  INVX1 INVX1_614 ( .A(_abc_17692_n3551), .Y(_abc_17692_n3796) );
  INVX1 INVX1_615 ( .A(_abc_17692_n3798), .Y(_abc_17692_n3799) );
  INVX1 INVX1_616 ( .A(_abc_17692_n3800), .Y(_abc_17692_n3801) );
  INVX1 INVX1_617 ( .A(_abc_17692_n3803), .Y(_abc_17692_n3804) );
  INVX1 INVX1_618 ( .A(_abc_17692_n3659), .Y(_abc_17692_n3807) );
  INVX1 INVX1_619 ( .A(_abc_17692_n3808), .Y(_abc_17692_n3809) );
  INVX1 INVX1_62 ( .A(_abc_17692_n1072), .Y(_abc_17692_n1073) );
  INVX1 INVX1_620 ( .A(_abc_17692_n3470), .Y(_abc_17692_n3811) );
  INVX1 INVX1_621 ( .A(_abc_17692_n3813), .Y(_abc_17692_n3814) );
  INVX1 INVX1_622 ( .A(_abc_17692_n3816), .Y(_abc_17692_n3817) );
  INVX1 INVX1_623 ( .A(_abc_17692_n3407), .Y(_abc_17692_n3821) );
  INVX1 INVX1_624 ( .A(_abc_17692_n3408), .Y(_abc_17692_n3823) );
  INVX1 INVX1_625 ( .A(_abc_17692_n3826), .Y(_abc_17692_n3827) );
  INVX1 INVX1_626 ( .A(_abc_17692_n3497), .Y(_abc_17692_n3829) );
  INVX1 INVX1_627 ( .A(_abc_17692_n3831), .Y(_abc_17692_n3832) );
  INVX1 INVX1_628 ( .A(_abc_17692_n3833), .Y(_abc_17692_n3834_1) );
  INVX1 INVX1_629 ( .A(_abc_17692_n3836), .Y(_abc_17692_n3837_1) );
  INVX1 INVX1_63 ( .A(_abc_17692_n1074), .Y(_abc_17692_n1075) );
  INVX1 INVX1_630 ( .A(_abc_17692_n3734), .Y(_abc_17692_n3840) );
  INVX1 INVX1_631 ( .A(_abc_17692_n3422), .Y(_abc_17692_n3841) );
  INVX1 INVX1_632 ( .A(_abc_17692_n3842), .Y(_abc_17692_n3843_1) );
  INVX1 INVX1_633 ( .A(_abc_17692_n3525), .Y(_abc_17692_n3845) );
  INVX1 INVX1_634 ( .A(_abc_17692_n3847), .Y(_abc_17692_n3848) );
  INVX1 INVX1_635 ( .A(_abc_17692_n3849), .Y(_abc_17692_n3850) );
  INVX1 INVX1_636 ( .A(_abc_17692_n3851), .Y(_abc_17692_n3852) );
  INVX1 INVX1_637 ( .A(workunit1_16_bF_buf2), .Y(_abc_17692_n3867) );
  INVX1 INVX1_638 ( .A(_abc_17692_n3885), .Y(_abc_17692_n3886) );
  INVX1 INVX1_639 ( .A(_abc_17692_n3887), .Y(_abc_17692_n3888) );
  INVX1 INVX1_64 ( .A(_abc_17692_n1076), .Y(_abc_17692_n1077) );
  INVX1 INVX1_640 ( .A(_abc_17692_n3891), .Y(_abc_17692_n3892) );
  INVX1 INVX1_641 ( .A(_abc_17692_n3890), .Y(_abc_17692_n3893) );
  INVX1 INVX1_642 ( .A(_abc_17692_n3894), .Y(_abc_17692_n3895) );
  INVX1 INVX1_643 ( .A(_abc_17692_n3910), .Y(_abc_17692_n3911) );
  INVX1 INVX1_644 ( .A(_abc_17692_n3865), .Y(_abc_17692_n3913) );
  INVX1 INVX1_645 ( .A(_abc_17692_n3918), .Y(_abc_17692_n3919) );
  INVX1 INVX1_646 ( .A(_abc_17692_n3684), .Y(_abc_17692_n3920) );
  INVX1 INVX1_647 ( .A(_abc_17692_n3922), .Y(_abc_17692_n3923) );
  INVX1 INVX1_648 ( .A(_abc_17692_n3925), .Y(_abc_17692_n3928) );
  INVX1 INVX1_649 ( .A(_abc_17692_n3929), .Y(_abc_17692_n3933) );
  INVX1 INVX1_65 ( .A(_abc_17692_n1078), .Y(_abc_17692_n1080) );
  INVX1 INVX1_650 ( .A(_abc_17692_n3942), .Y(_abc_17692_n3943) );
  INVX1 INVX1_651 ( .A(_abc_17692_n3948), .Y(_abc_17692_n3949) );
  INVX1 INVX1_652 ( .A(_abc_17692_n3950), .Y(_abc_17692_n3951) );
  INVX1 INVX1_653 ( .A(_abc_17692_n3952), .Y(_abc_17692_n3953) );
  INVX1 INVX1_654 ( .A(_abc_17692_n3955), .Y(_abc_17692_n3957) );
  INVX1 INVX1_655 ( .A(_abc_17692_n3959), .Y(_abc_17692_n3961) );
  INVX1 INVX1_656 ( .A(_abc_17692_n3969), .Y(_abc_17692_n3970) );
  INVX1 INVX1_657 ( .A(_abc_17692_n3977), .Y(_abc_17692_n3978_1) );
  INVX1 INVX1_658 ( .A(_abc_17692_n3980), .Y(_abc_17692_n3981) );
  INVX1 INVX1_659 ( .A(_abc_17692_n3982), .Y(_abc_17692_n3983) );
  INVX1 INVX1_66 ( .A(_abc_17692_n1087), .Y(_abc_17692_n1088) );
  INVX1 INVX1_660 ( .A(_abc_17692_n3985), .Y(_abc_17692_n3987) );
  INVX1 INVX1_661 ( .A(_abc_17692_n3988), .Y(_abc_17692_n3992) );
  INVX1 INVX1_662 ( .A(_abc_17692_n4001), .Y(_abc_17692_n4002_1) );
  INVX1 INVX1_663 ( .A(_abc_17692_n3979), .Y(_abc_17692_n4004) );
  INVX1 INVX1_664 ( .A(_abc_17692_n4010), .Y(_abc_17692_n4011) );
  INVX1 INVX1_665 ( .A(_abc_17692_n3655), .Y(_abc_17692_n4016) );
  INVX1 INVX1_666 ( .A(_abc_17692_n4017), .Y(_abc_17692_n4018) );
  INVX1 INVX1_667 ( .A(_abc_17692_n4019), .Y(_abc_17692_n4020) );
  INVX1 INVX1_668 ( .A(_abc_17692_n4025), .Y(_abc_17692_n4026) );
  INVX1 INVX1_669 ( .A(_abc_17692_n4032), .Y(_abc_17692_n4033) );
  INVX1 INVX1_67 ( .A(_abc_17692_n1089), .Y(_abc_17692_n1090) );
  INVX1 INVX1_670 ( .A(_abc_17692_n4051), .Y(_abc_17692_n4052) );
  INVX1 INVX1_671 ( .A(_abc_17692_n4055), .Y(_abc_17692_n4056) );
  INVX1 INVX1_672 ( .A(_abc_17692_n4063), .Y(_abc_17692_n4064_1) );
  INVX1 INVX1_673 ( .A(_abc_17692_n4066), .Y(_abc_17692_n4072) );
  INVX1 INVX1_674 ( .A(_abc_17692_n4083), .Y(_abc_17692_n4084_1) );
  INVX1 INVX1_675 ( .A(_abc_17692_n4079), .Y(_abc_17692_n4088) );
  INVX1 INVX1_676 ( .A(_abc_17692_n4081), .Y(_abc_17692_n4089) );
  INVX1 INVX1_677 ( .A(_abc_17692_n4086), .Y(_abc_17692_n4091) );
  INVX1 INVX1_678 ( .A(_abc_17692_n4093), .Y(_abc_17692_n4094) );
  INVX1 INVX1_679 ( .A(_abc_17692_n4099), .Y(_abc_17692_n4100) );
  INVX1 INVX1_68 ( .A(delta_8_), .Y(_abc_17692_n1097) );
  INVX1 INVX1_680 ( .A(_abc_17692_n3782), .Y(_abc_17692_n4103) );
  INVX1 INVX1_681 ( .A(_abc_17692_n4104), .Y(_abc_17692_n4105) );
  INVX1 INVX1_682 ( .A(_abc_17692_n3996), .Y(_abc_17692_n4108) );
  INVX1 INVX1_683 ( .A(_abc_17692_n4113), .Y(_abc_17692_n4114) );
  INVX1 INVX1_684 ( .A(_abc_17692_n4115), .Y(_abc_17692_n4116) );
  INVX1 INVX1_685 ( .A(workunit2_12_bF_buf0), .Y(_abc_17692_n4120) );
  INVX1 INVX1_686 ( .A(_abc_17692_n4129), .Y(_abc_17692_n4130) );
  INVX1 INVX1_687 ( .A(_abc_17692_n4128), .Y(_abc_17692_n4134) );
  INVX1 INVX1_688 ( .A(_abc_17692_n4132), .Y(_abc_17692_n4135) );
  INVX1 INVX1_689 ( .A(_abc_17692_n4137), .Y(_abc_17692_n4138) );
  INVX1 INVX1_69 ( .A(sum_8_), .Y(_abc_17692_n1098) );
  INVX1 INVX1_690 ( .A(_abc_17692_n4141), .Y(_abc_17692_n4142) );
  INVX1 INVX1_691 ( .A(_abc_17692_n4145), .Y(_abc_17692_n4146) );
  INVX1 INVX1_692 ( .A(_abc_17692_n4157), .Y(_abc_17692_n4158) );
  INVX1 INVX1_693 ( .A(_abc_17692_n4169_1), .Y(_abc_17692_n4170) );
  INVX1 INVX1_694 ( .A(_abc_17692_n4168), .Y(_abc_17692_n4174) );
  INVX1 INVX1_695 ( .A(_abc_17692_n4172), .Y(_abc_17692_n4175) );
  INVX1 INVX1_696 ( .A(_abc_17692_n4177), .Y(_abc_17692_n4178) );
  INVX1 INVX1_697 ( .A(_abc_17692_n4182), .Y(_abc_17692_n4183) );
  INVX1 INVX1_698 ( .A(_abc_17692_n3964), .Y(_abc_17692_n4191) );
  INVX1 INVX1_699 ( .A(_abc_17692_n4196), .Y(_abc_17692_n4197) );
  INVX1 INVX1_7 ( .A(_abc_17692_n675), .Y(_abc_17692_n676_1) );
  INVX1 INVX1_70 ( .A(_abc_17692_n1100), .Y(_abc_17692_n1101) );
  INVX1 INVX1_700 ( .A(_abc_17692_n4199), .Y(_abc_17692_n4200) );
  INVX1 INVX1_701 ( .A(_abc_17692_n4211), .Y(_abc_17692_n4212) );
  INVX1 INVX1_702 ( .A(_abc_17692_n4207), .Y(_abc_17692_n4216) );
  INVX1 INVX1_703 ( .A(_abc_17692_n4209), .Y(_abc_17692_n4217) );
  INVX1 INVX1_704 ( .A(_abc_17692_n4214), .Y(_abc_17692_n4219) );
  INVX1 INVX1_705 ( .A(_abc_17692_n4221), .Y(_abc_17692_n4222) );
  INVX1 INVX1_706 ( .A(_abc_17692_n4226), .Y(_abc_17692_n4227) );
  INVX1 INVX1_707 ( .A(_abc_17692_n3937), .Y(_abc_17692_n4231) );
  INVX1 INVX1_708 ( .A(_abc_17692_n4237), .Y(_abc_17692_n4238) );
  INVX1 INVX1_709 ( .A(_abc_17692_n4240), .Y(_abc_17692_n4241) );
  INVX1 INVX1_71 ( .A(_abc_17692_n1102), .Y(_abc_17692_n1103) );
  INVX1 INVX1_710 ( .A(_abc_17692_n4102), .Y(_abc_17692_n4249) );
  INVX1 INVX1_711 ( .A(_abc_17692_n3772), .Y(_abc_17692_n4255) );
  INVX1 INVX1_712 ( .A(_abc_17692_n4261), .Y(_abc_17692_n4262) );
  INVX1 INVX1_713 ( .A(_abc_17692_n3904), .Y(_abc_17692_n4269_1) );
  INVX1 INVX1_714 ( .A(_abc_17692_n4274), .Y(_abc_17692_n4275) );
  INVX1 INVX1_715 ( .A(_abc_17692_n4277), .Y(_abc_17692_n4278) );
  INVX1 INVX1_716 ( .A(_abc_17692_n4229), .Y(_abc_17692_n4281) );
  INVX1 INVX1_717 ( .A(_abc_17692_n4292), .Y(_abc_17692_n4293) );
  INVX1 INVX1_718 ( .A(_abc_17692_n4185), .Y(_abc_17692_n4296) );
  INVX1 INVX1_719 ( .A(_abc_17692_n4031), .Y(_abc_17692_n4302) );
  INVX1 INVX1_72 ( .A(_abc_17692_n1104_1), .Y(_abc_17692_n1105) );
  INVX1 INVX1_720 ( .A(_abc_17692_n4307), .Y(_abc_17692_n4308) );
  INVX1 INVX1_721 ( .A(_abc_17692_n4327), .Y(_abc_17692_n4328) );
  INVX1 INVX1_722 ( .A(_abc_17692_n4330), .Y(_abc_17692_n4331) );
  INVX1 INVX1_723 ( .A(_abc_17692_n4335), .Y(_abc_17692_n4336) );
  INVX1 INVX1_724 ( .A(_abc_17692_n4337), .Y(_abc_17692_n4338) );
  INVX1 INVX1_725 ( .A(_abc_17692_n4340), .Y(_abc_17692_n4342) );
  INVX1 INVX1_726 ( .A(_abc_17692_n4344_1), .Y(_abc_17692_n4346) );
  INVX1 INVX1_727 ( .A(_abc_17692_n4348), .Y(_abc_17692_n4349) );
  INVX1 INVX1_728 ( .A(_abc_17692_n4353), .Y(_abc_17692_n4354) );
  INVX1 INVX1_729 ( .A(_abc_17692_n4144), .Y(_abc_17692_n4355) );
  INVX1 INVX1_73 ( .A(_abc_17692_n1113), .Y(_abc_17692_n1114) );
  INVX1 INVX1_730 ( .A(_abc_17692_n4356), .Y(_abc_17692_n4358) );
  INVX1 INVX1_731 ( .A(_abc_17692_n4362), .Y(_abc_17692_n4363) );
  INVX1 INVX1_732 ( .A(_abc_17692_n4364), .Y(_abc_17692_n4365) );
  INVX1 INVX1_733 ( .A(_abc_17692_n4369), .Y(_abc_17692_n4370) );
  INVX1 INVX1_734 ( .A(_abc_17692_n4368), .Y(_abc_17692_n4373) );
  INVX1 INVX1_735 ( .A(_abc_17692_n4382), .Y(_abc_17692_n4383) );
  INVX1 INVX1_736 ( .A(_abc_17692_n4384), .Y(_abc_17692_n4385) );
  INVX1 INVX1_737 ( .A(_abc_17692_n4391), .Y(_abc_17692_n4392_1) );
  INVX1 INVX1_738 ( .A(_abc_17692_n4394), .Y(_abc_17692_n4395) );
  INVX1 INVX1_739 ( .A(_abc_17692_n4397), .Y(_abc_17692_n4398) );
  INVX1 INVX1_74 ( .A(_abc_17692_n1121), .Y(_abc_17692_n1122) );
  INVX1 INVX1_740 ( .A(_abc_17692_n4399), .Y(_abc_17692_n4401) );
  INVX1 INVX1_741 ( .A(_abc_17692_n4403), .Y(_abc_17692_n4404) );
  INVX1 INVX1_742 ( .A(_abc_17692_n4407), .Y(_abc_17692_n4408) );
  INVX1 INVX1_743 ( .A(_abc_17692_n4409), .Y(_abc_17692_n4410) );
  INVX1 INVX1_744 ( .A(_abc_17692_n4418), .Y(_abc_17692_n4419) );
  INVX1 INVX1_745 ( .A(_abc_17692_n4421), .Y(_abc_17692_n4422) );
  INVX1 INVX1_746 ( .A(_abc_17692_n4424), .Y(_abc_17692_n4425) );
  INVX1 INVX1_747 ( .A(_abc_17692_n4426), .Y(_abc_17692_n4428) );
  INVX1 INVX1_748 ( .A(_abc_17692_n4430), .Y(_abc_17692_n4431) );
  INVX1 INVX1_749 ( .A(_abc_17692_n4434), .Y(_abc_17692_n4435) );
  INVX1 INVX1_75 ( .A(delta_9_), .Y(_abc_17692_n1123) );
  INVX1 INVX1_750 ( .A(_abc_17692_n4436), .Y(_abc_17692_n4437) );
  INVX1 INVX1_751 ( .A(_abc_17692_n4098), .Y(_abc_17692_n4444_1) );
  INVX1 INVX1_752 ( .A(_abc_17692_n4445), .Y(_abc_17692_n4446) );
  INVX1 INVX1_753 ( .A(_abc_17692_n4447_1), .Y(_abc_17692_n4449) );
  INVX1 INVX1_754 ( .A(_abc_17692_n4453), .Y(_abc_17692_n4454) );
  INVX1 INVX1_755 ( .A(_abc_17692_n4455), .Y(_abc_17692_n4456) );
  INVX1 INVX1_756 ( .A(_abc_17692_n4225), .Y(_abc_17692_n4461) );
  INVX1 INVX1_757 ( .A(_abc_17692_n4462), .Y(_abc_17692_n4463) );
  INVX1 INVX1_758 ( .A(_abc_17692_n4464), .Y(_abc_17692_n4465) );
  INVX1 INVX1_759 ( .A(_abc_17692_n4181), .Y(_abc_17692_n4470) );
  INVX1 INVX1_76 ( .A(sum_9_), .Y(_abc_17692_n1124) );
  INVX1 INVX1_760 ( .A(_abc_17692_n4471), .Y(_abc_17692_n4472) );
  INVX1 INVX1_761 ( .A(_abc_17692_n4473), .Y(_abc_17692_n4475) );
  INVX1 INVX1_762 ( .A(_abc_17692_n4329), .Y(_abc_17692_n4488) );
  INVX1 INVX1_763 ( .A(_abc_17692_n4498), .Y(_abc_17692_n4499) );
  INVX1 INVX1_764 ( .A(_abc_17692_n4492), .Y(_abc_17692_n4505) );
  INVX1 INVX1_765 ( .A(_abc_17692_n4500), .Y(_abc_17692_n4507_1) );
  INVX1 INVX1_766 ( .A(_abc_17692_n4420), .Y(_abc_17692_n4513) );
  INVX1 INVX1_767 ( .A(_abc_17692_n4515), .Y(_abc_17692_n4516) );
  INVX1 INVX1_768 ( .A(_abc_17692_n4518), .Y(_abc_17692_n4519) );
  INVX1 INVX1_769 ( .A(_abc_17692_n4512), .Y(_abc_17692_n4523) );
  INVX1 INVX1_77 ( .A(_abc_17692_n1125), .Y(_abc_17692_n1126) );
  INVX1 INVX1_770 ( .A(_abc_17692_n4521), .Y(_abc_17692_n4525) );
  INVX1 INVX1_771 ( .A(_abc_17692_n4527), .Y(_abc_17692_n4528) );
  INVX1 INVX1_772 ( .A(_abc_17692_n4510_1), .Y(_abc_17692_n4530) );
  INVX1 INVX1_773 ( .A(_abc_17692_n4534), .Y(_abc_17692_n4535) );
  INVX1 INVX1_774 ( .A(_abc_17692_n4537), .Y(_abc_17692_n4538) );
  INVX1 INVX1_775 ( .A(_abc_17692_n4540), .Y(_abc_17692_n4541) );
  INVX1 INVX1_776 ( .A(_abc_17692_n4546), .Y(_abc_17692_n4547) );
  INVX1 INVX1_777 ( .A(_abc_17692_n4339), .Y(_abc_17692_n4552) );
  INVX1 INVX1_778 ( .A(_abc_17692_n4554), .Y(_abc_17692_n4555) );
  INVX1 INVX1_779 ( .A(_abc_17692_n4557), .Y(_abc_17692_n4558) );
  INVX1 INVX1_78 ( .A(_abc_17692_n1096), .Y(_abc_17692_n1128) );
  INVX1 INVX1_780 ( .A(_abc_17692_n4556), .Y(_abc_17692_n4562) );
  INVX1 INVX1_781 ( .A(_abc_17692_n4560), .Y(_abc_17692_n4563) );
  INVX1 INVX1_782 ( .A(_abc_17692_n4565), .Y(_abc_17692_n4566) );
  INVX1 INVX1_783 ( .A(_abc_17692_n4570), .Y(_abc_17692_n4571) );
  INVX1 INVX1_784 ( .A(_abc_17692_n4580), .Y(_abc_17692_n4581) );
  INVX1 INVX1_785 ( .A(_abc_17692_n4393), .Y(_abc_17692_n4587_1) );
  INVX1 INVX1_786 ( .A(_abc_17692_n4589), .Y(_abc_17692_n4590) );
  INVX1 INVX1_787 ( .A(_abc_17692_n4592), .Y(_abc_17692_n4593) );
  INVX1 INVX1_788 ( .A(_abc_17692_n4591), .Y(_abc_17692_n4597) );
  INVX1 INVX1_789 ( .A(_abc_17692_n4595), .Y(_abc_17692_n4598) );
  INVX1 INVX1_79 ( .A(_abc_17692_n1129), .Y(_abc_17692_n1130) );
  INVX1 INVX1_790 ( .A(_abc_17692_n4600), .Y(_abc_17692_n4601) );
  INVX1 INVX1_791 ( .A(_abc_17692_n4606), .Y(_abc_17692_n4607) );
  INVX1 INVX1_792 ( .A(_abc_17692_n4609), .Y(_abc_17692_n4610) );
  INVX1 INVX1_793 ( .A(_abc_17692_n4612), .Y(_abc_17692_n4613) );
  INVX1 INVX1_794 ( .A(_abc_17692_n4614), .Y(_abc_17692_n4615) );
  INVX1 INVX1_795 ( .A(_abc_17692_n4618), .Y(_abc_17692_n4619) );
  INVX1 INVX1_796 ( .A(workunit2_14_bF_buf0), .Y(_abc_17692_n4623) );
  INVX1 INVX1_797 ( .A(_abc_17692_n4366), .Y(_abc_17692_n4626) );
  INVX1 INVX1_798 ( .A(_abc_17692_n4628), .Y(_abc_17692_n4629) );
  INVX1 INVX1_799 ( .A(_abc_17692_n4631), .Y(_abc_17692_n4632) );
  INVX1 INVX1_8 ( .A(_abc_17692_n679), .Y(_abc_17692_n680) );
  INVX1 INVX1_80 ( .A(_abc_17692_n1136), .Y(_abc_17692_n1137) );
  INVX1 INVX1_800 ( .A(_abc_17692_n4625), .Y(_abc_17692_n4636) );
  INVX1 INVX1_801 ( .A(_abc_17692_n4634), .Y(_abc_17692_n4638) );
  INVX1 INVX1_802 ( .A(_abc_17692_n4640), .Y(_abc_17692_n4642) );
  INVX1 INVX1_803 ( .A(_abc_17692_n4644), .Y(_abc_17692_n4645) );
  INVX1 INVX1_804 ( .A(_abc_17692_n4648), .Y(_abc_17692_n4649) );
  INVX1 INVX1_805 ( .A(_abc_17692_n4650), .Y(_abc_17692_n4651) );
  INVX1 INVX1_806 ( .A(_abc_17692_n4653), .Y(_abc_17692_n4654) );
  INVX1 INVX1_807 ( .A(_abc_17692_n4655), .Y(_abc_17692_n4656) );
  INVX1 INVX1_808 ( .A(_abc_17692_n4659), .Y(_abc_17692_n4660) );
  INVX1 INVX1_809 ( .A(_abc_17692_n4536), .Y(_abc_17692_n4669) );
  INVX1 INVX1_81 ( .A(_abc_17692_n1141), .Y(_abc_17692_n1142) );
  INVX1 INVX1_810 ( .A(_abc_17692_n4432), .Y(_abc_17692_n4670) );
  INVX1 INVX1_811 ( .A(_abc_17692_n4676), .Y(_abc_17692_n4677) );
  INVX1 INVX1_812 ( .A(_abc_17692_n4573), .Y(_abc_17692_n4681) );
  INVX1 INVX1_813 ( .A(_abc_17692_n4350), .Y(_abc_17692_n4682) );
  INVX1 INVX1_814 ( .A(_abc_17692_n4684), .Y(_abc_17692_n4685) );
  INVX1 INVX1_815 ( .A(_abc_17692_n4686), .Y(_abc_17692_n4687) );
  INVX1 INVX1_816 ( .A(_abc_17692_n4690), .Y(_abc_17692_n4691) );
  INVX1 INVX1_817 ( .A(_abc_17692_n4381), .Y(_abc_17692_n4695) );
  INVX1 INVX1_818 ( .A(_abc_17692_n4697), .Y(_abc_17692_n4698) );
  INVX1 INVX1_819 ( .A(_abc_17692_n4702), .Y(_abc_17692_n4703) );
  INVX1 INVX1_82 ( .A(delta_10_), .Y(_abc_17692_n1151) );
  INVX1 INVX1_820 ( .A(_abc_17692_n4608), .Y(_abc_17692_n4707) );
  INVX1 INVX1_821 ( .A(_abc_17692_n4406), .Y(_abc_17692_n4708) );
  INVX1 INVX1_822 ( .A(_abc_17692_n4710), .Y(_abc_17692_n4711) );
  INVX1 INVX1_823 ( .A(_abc_17692_n4715), .Y(_abc_17692_n4716) );
  INVX1 INVX1_824 ( .A(_abc_17692_n4735_1), .Y(_abc_17692_n4736) );
  INVX1 INVX1_825 ( .A(_abc_17692_n4734), .Y(_abc_17692_n4741) );
  INVX1 INVX1_826 ( .A(_abc_17692_n4745), .Y(_abc_17692_n4746) );
  INVX1 INVX1_827 ( .A(_abc_17692_n4747), .Y(_abc_17692_n4748) );
  INVX1 INVX1_828 ( .A(_abc_17692_n4751), .Y(_abc_17692_n4752) );
  INVX1 INVX1_829 ( .A(_abc_17692_n4750), .Y(_abc_17692_n4753) );
  INVX1 INVX1_83 ( .A(sum_10_), .Y(_abc_17692_n1152_1) );
  INVX1 INVX1_830 ( .A(_abc_17692_n4754), .Y(_abc_17692_n4755) );
  INVX1 INVX1_831 ( .A(_abc_17692_n4771), .Y(_abc_17692_n4772) );
  INVX1 INVX1_832 ( .A(_abc_17692_n4770), .Y(_abc_17692_n4774) );
  INVX1 INVX1_833 ( .A(_abc_17692_n4778), .Y(_abc_17692_n4779) );
  INVX1 INVX1_834 ( .A(_abc_17692_n4780), .Y(_abc_17692_n4781) );
  INVX1 INVX1_835 ( .A(_abc_17692_n4783), .Y(_abc_17692_n4785) );
  INVX1 INVX1_836 ( .A(_abc_17692_n4787), .Y(_abc_17692_n4789_1) );
  INVX1 INVX1_837 ( .A(_abc_17692_n4797), .Y(_abc_17692_n4800) );
  INVX1 INVX1_838 ( .A(_abc_17692_n4798), .Y(_abc_17692_n4801) );
  INVX1 INVX1_839 ( .A(_abc_17692_n4635), .Y(_abc_17692_n4805) );
  INVX1 INVX1_84 ( .A(_abc_17692_n1154), .Y(_abc_17692_n1155) );
  INVX1 INVX1_840 ( .A(_abc_17692_n4807), .Y(_abc_17692_n4808) );
  INVX1 INVX1_841 ( .A(_abc_17692_n4810), .Y(_abc_17692_n4813) );
  INVX1 INVX1_842 ( .A(_abc_17692_n4814), .Y(_abc_17692_n4818) );
  INVX1 INVX1_843 ( .A(_abc_17692_n4827), .Y(_abc_17692_n4828) );
  INVX1 INVX1_844 ( .A(_abc_17692_n4829), .Y(_abc_17692_n4830) );
  INVX1 INVX1_845 ( .A(_abc_17692_n4831), .Y(_abc_17692_n4832) );
  INVX1 INVX1_846 ( .A(_abc_17692_n4522), .Y(_abc_17692_n4840) );
  INVX1 INVX1_847 ( .A(_abc_17692_n4842), .Y(_abc_17692_n4843) );
  INVX1 INVX1_848 ( .A(_abc_17692_n4845), .Y(_abc_17692_n4848) );
  INVX1 INVX1_849 ( .A(_abc_17692_n4849), .Y(_abc_17692_n4853) );
  INVX1 INVX1_85 ( .A(_abc_17692_n1159), .Y(_abc_17692_n1160) );
  INVX1 INVX1_850 ( .A(_abc_17692_n4863), .Y(_abc_17692_n4864) );
  INVX1 INVX1_851 ( .A(_abc_17692_n4862), .Y(_abc_17692_n4866) );
  INVX1 INVX1_852 ( .A(_abc_17692_n4532), .Y(_abc_17692_n4872) );
  INVX1 INVX1_853 ( .A(_abc_17692_n4873), .Y(_abc_17692_n4874) );
  INVX1 INVX1_854 ( .A(_abc_17692_n4875), .Y(_abc_17692_n4876) );
  INVX1 INVX1_855 ( .A(_abc_17692_n4569), .Y(_abc_17692_n4881) );
  INVX1 INVX1_856 ( .A(_abc_17692_n4882), .Y(_abc_17692_n4883) );
  INVX1 INVX1_857 ( .A(_abc_17692_n4884), .Y(_abc_17692_n4885) );
  INVX1 INVX1_858 ( .A(_abc_17692_n4890), .Y(_abc_17692_n4891) );
  INVX1 INVX1_859 ( .A(_abc_17692_n4604), .Y(_abc_17692_n4896_1) );
  INVX1 INVX1_86 ( .A(_abc_17692_n1161), .Y(_abc_17692_n1162) );
  INVX1 INVX1_860 ( .A(_abc_17692_n4897), .Y(_abc_17692_n4898) );
  INVX1 INVX1_861 ( .A(_abc_17692_n4899), .Y(_abc_17692_n4901) );
  INVX1 INVX1_862 ( .A(_abc_17692_n4928), .Y(_abc_17692_n4929) );
  INVX1 INVX1_863 ( .A(_abc_17692_n4932), .Y(_abc_17692_n4933) );
  INVX1 INVX1_864 ( .A(_abc_17692_n4914), .Y(_abc_17692_n4935) );
  INVX1 INVX1_865 ( .A(_abc_17692_n4922), .Y(_abc_17692_n4940) );
  INVX1 INVX1_866 ( .A(_abc_17692_n4956), .Y(_abc_17692_n4957) );
  INVX1 INVX1_867 ( .A(_abc_17692_n4955), .Y(_abc_17692_n4961) );
  INVX1 INVX1_868 ( .A(_abc_17692_n4959), .Y(_abc_17692_n4962) );
  INVX1 INVX1_869 ( .A(_abc_17692_n4964), .Y(_abc_17692_n4965) );
  INVX1 INVX1_87 ( .A(_abc_17692_n1167), .Y(_abc_17692_n1168) );
  INVX1 INVX1_870 ( .A(_abc_17692_n4970), .Y(_abc_17692_n4971) );
  INVX1 INVX1_871 ( .A(_abc_17692_n4983), .Y(_abc_17692_n4984) );
  INVX1 INVX1_872 ( .A(_abc_17692_n4999), .Y(_abc_17692_n5000) );
  INVX1 INVX1_873 ( .A(_abc_17692_n4990), .Y(_abc_17692_n5004) );
  INVX1 INVX1_874 ( .A(_abc_17692_n4997), .Y(_abc_17692_n5006) );
  INVX1 INVX1_875 ( .A(_abc_17692_n5002), .Y(_abc_17692_n5008) );
  INVX1 INVX1_876 ( .A(_abc_17692_n5010), .Y(_abc_17692_n5011) );
  INVX1 INVX1_877 ( .A(_abc_17692_n5015), .Y(_abc_17692_n5016) );
  INVX1 INVX1_878 ( .A(_abc_17692_n4822), .Y(_abc_17692_n5021) );
  INVX1 INVX1_879 ( .A(_abc_17692_n5027), .Y(_abc_17692_n5028) );
  INVX1 INVX1_88 ( .A(_abc_17692_n1169), .Y(_abc_17692_n1170) );
  INVX1 INVX1_880 ( .A(_abc_17692_n5029), .Y(_abc_17692_n5030) );
  INVX1 INVX1_881 ( .A(_abc_17692_n5045), .Y(_abc_17692_n5046) );
  INVX1 INVX1_882 ( .A(_abc_17692_n5036), .Y(_abc_17692_n5050) );
  INVX1 INVX1_883 ( .A(_abc_17692_n5043), .Y(_abc_17692_n5052) );
  INVX1 INVX1_884 ( .A(_abc_17692_n5048), .Y(_abc_17692_n5054) );
  INVX1 INVX1_885 ( .A(_abc_17692_n5056), .Y(_abc_17692_n5057) );
  INVX1 INVX1_886 ( .A(_abc_17692_n5061), .Y(_abc_17692_n5062) );
  INVX1 INVX1_887 ( .A(_abc_17692_n4792_1), .Y(_abc_17692_n5067) );
  INVX1 INVX1_888 ( .A(_abc_17692_n5073), .Y(_abc_17692_n5074) );
  INVX1 INVX1_889 ( .A(_abc_17692_n5075), .Y(_abc_17692_n5076) );
  INVX1 INVX1_89 ( .A(_abc_17692_n1171), .Y(_abc_17692_n1172) );
  INVX1 INVX1_890 ( .A(_abc_17692_n5093), .Y(_abc_17692_n5094) );
  INVX1 INVX1_891 ( .A(_abc_17692_n5085), .Y(_abc_17692_n5098) );
  INVX1 INVX1_892 ( .A(_abc_17692_n5091), .Y(_abc_17692_n5099) );
  INVX1 INVX1_893 ( .A(_abc_17692_n5096), .Y(_abc_17692_n5101) );
  INVX1 INVX1_894 ( .A(_abc_17692_n5103), .Y(_abc_17692_n5104) );
  INVX1 INVX1_895 ( .A(_abc_17692_n5108), .Y(_abc_17692_n5109) );
  INVX1 INVX1_896 ( .A(_abc_17692_n4857), .Y(_abc_17692_n5114) );
  INVX1 INVX1_897 ( .A(_abc_17692_n4542), .Y(_abc_17692_n5118) );
  INVX1 INVX1_898 ( .A(_abc_17692_n5121), .Y(_abc_17692_n5122) );
  INVX1 INVX1_899 ( .A(_abc_17692_n5124), .Y(_abc_17692_n5125) );
  INVX1 INVX1_9 ( .A(_abc_17692_n683), .Y(_abc_17692_n684) );
  INVX1 INVX1_90 ( .A(sum_11_), .Y(_abc_17692_n1180) );
  INVX1 INVX1_900 ( .A(_abc_17692_n5111), .Y(_abc_17692_n5130) );
  INVX1 INVX1_901 ( .A(_abc_17692_n5141), .Y(_abc_17692_n5142) );
  INVX1 INVX1_902 ( .A(_abc_17692_n4973), .Y(_abc_17692_n5145) );
  INVX1 INVX1_903 ( .A(_abc_17692_n4769), .Y(_abc_17692_n5148) );
  INVX1 INVX1_904 ( .A(_abc_17692_n5150), .Y(_abc_17692_n5151) );
  INVX1 INVX1_905 ( .A(_abc_17692_n5155), .Y(_abc_17692_n5156) );
  INVX1 INVX1_906 ( .A(_abc_17692_n5157), .Y(_abc_17692_n5158) );
  INVX1 INVX1_907 ( .A(_abc_17692_n5018), .Y(_abc_17692_n5162) );
  INVX1 INVX1_908 ( .A(_abc_17692_n4646_1), .Y(_abc_17692_n5166) );
  INVX1 INVX1_909 ( .A(_abc_17692_n5174), .Y(_abc_17692_n5175) );
  INVX1 INVX1_91 ( .A(_abc_17692_n1181), .Y(_abc_17692_n1182) );
  INVX1 INVX1_910 ( .A(_abc_17692_n5064), .Y(_abc_17692_n5178) );
  INVX1 INVX1_911 ( .A(_abc_17692_n5188), .Y(_abc_17692_n5189) );
  INVX1 INVX1_912 ( .A(_abc_17692_n5207), .Y(_abc_17692_n5208) );
  INVX1 INVX1_913 ( .A(_abc_17692_n5209), .Y(_abc_17692_n5210) );
  INVX1 INVX1_914 ( .A(_abc_17692_n5211), .Y(_abc_17692_n5212_1) );
  INVX1 INVX1_915 ( .A(_abc_17692_n5213), .Y(_abc_17692_n5214) );
  INVX1 INVX1_916 ( .A(_abc_17692_n5216), .Y(_abc_17692_n5217) );
  INVX1 INVX1_917 ( .A(_abc_17692_n5049), .Y(_abc_17692_n5219) );
  INVX1 INVX1_918 ( .A(_abc_17692_n5221), .Y(_abc_17692_n5222) );
  INVX1 INVX1_919 ( .A(_abc_17692_n5225), .Y(_abc_17692_n5226) );
  INVX1 INVX1_92 ( .A(_abc_17692_n1150), .Y(_abc_17692_n1186) );
  INVX1 INVX1_920 ( .A(_abc_17692_n5218), .Y(_abc_17692_n5230) );
  INVX1 INVX1_921 ( .A(_abc_17692_n5228), .Y(_abc_17692_n5231) );
  INVX1 INVX1_922 ( .A(_abc_17692_n5234), .Y(_abc_17692_n5235) );
  INVX1 INVX1_923 ( .A(_abc_17692_n5237), .Y(_abc_17692_n5238) );
  INVX1 INVX1_924 ( .A(_abc_17692_n5202), .Y(_abc_17692_n5240) );
  INVX1 INVX1_925 ( .A(_abc_17692_n4960), .Y(_abc_17692_n5244) );
  INVX1 INVX1_926 ( .A(_abc_17692_n5246), .Y(_abc_17692_n5247) );
  INVX1 INVX1_927 ( .A(_abc_17692_n5250), .Y(_abc_17692_n5251) );
  INVX1 INVX1_928 ( .A(_abc_17692_n5253), .Y(_abc_17692_n5255) );
  INVX1 INVX1_929 ( .A(_abc_17692_n5258), .Y(_abc_17692_n5259) );
  INVX1 INVX1_93 ( .A(_abc_17692_n1187), .Y(_abc_17692_n1188) );
  INVX1 INVX1_930 ( .A(_abc_17692_n5257), .Y(_abc_17692_n5261) );
  INVX1 INVX1_931 ( .A(_abc_17692_n5262), .Y(_abc_17692_n5263) );
  INVX1 INVX1_932 ( .A(_abc_17692_n5264), .Y(_abc_17692_n5265) );
  INVX1 INVX1_933 ( .A(_abc_17692_n5269), .Y(_abc_17692_n5270) );
  INVX1 INVX1_934 ( .A(_abc_17692_n5275_1), .Y(_abc_17692_n5276) );
  INVX1 INVX1_935 ( .A(_abc_17692_n5003), .Y(_abc_17692_n5277) );
  INVX1 INVX1_936 ( .A(_abc_17692_n5279), .Y(_abc_17692_n5280) );
  INVX1 INVX1_937 ( .A(_abc_17692_n5283), .Y(_abc_17692_n5284) );
  INVX1 INVX1_938 ( .A(_abc_17692_n5286), .Y(_abc_17692_n5287) );
  INVX1 INVX1_939 ( .A(_abc_17692_n5290), .Y(_abc_17692_n5292) );
  INVX1 INVX1_94 ( .A(_abc_17692_n1194), .Y(_abc_17692_n1195_1) );
  INVX1 INVX1_940 ( .A(_abc_17692_n5294), .Y(_abc_17692_n5295) );
  INVX1 INVX1_941 ( .A(_abc_17692_n5097_1), .Y(_abc_17692_n5303) );
  INVX1 INVX1_942 ( .A(_abc_17692_n5305), .Y(_abc_17692_n5306) );
  INVX1 INVX1_943 ( .A(_abc_17692_n5309), .Y(_abc_17692_n5310) );
  INVX1 INVX1_944 ( .A(_abc_17692_n5312), .Y(_abc_17692_n5314) );
  INVX1 INVX1_945 ( .A(_abc_17692_n5317), .Y(_abc_17692_n5318) );
  INVX1 INVX1_946 ( .A(_abc_17692_n5316), .Y(_abc_17692_n5319) );
  INVX1 INVX1_947 ( .A(_abc_17692_n5320), .Y(_abc_17692_n5321) );
  INVX1 INVX1_948 ( .A(_abc_17692_n5322), .Y(_abc_17692_n5323) );
  INVX1 INVX1_949 ( .A(_abc_17692_n5302), .Y(_abc_17692_n5325) );
  INVX1 INVX1_95 ( .A(_abc_17692_n1196), .Y(_abc_17692_n1198) );
  INVX1 INVX1_950 ( .A(_abc_17692_n5107), .Y(_abc_17692_n5331) );
  INVX1 INVX1_951 ( .A(_abc_17692_n5332), .Y(_abc_17692_n5333) );
  INVX1 INVX1_952 ( .A(_abc_17692_n5334), .Y(_abc_17692_n5335) );
  INVX1 INVX1_953 ( .A(_abc_17692_n4969), .Y(_abc_17692_n5340) );
  INVX1 INVX1_954 ( .A(_abc_17692_n5341), .Y(_abc_17692_n5342) );
  INVX1 INVX1_955 ( .A(_abc_17692_n5343), .Y(_abc_17692_n5344) );
  INVX1 INVX1_956 ( .A(_abc_17692_n5014), .Y(_abc_17692_n5349) );
  INVX1 INVX1_957 ( .A(_abc_17692_n5350), .Y(_abc_17692_n5351) );
  INVX1 INVX1_958 ( .A(_abc_17692_n5352), .Y(_abc_17692_n5353) );
  INVX1 INVX1_959 ( .A(_abc_17692_n5060), .Y(_abc_17692_n5358) );
  INVX1 INVX1_96 ( .A(delta_12_), .Y(_abc_17692_n1205) );
  INVX1 INVX1_960 ( .A(_abc_17692_n5359), .Y(_abc_17692_n5360) );
  INVX1 INVX1_961 ( .A(_abc_17692_n5361), .Y(_abc_17692_n5362) );
  INVX1 INVX1_962 ( .A(_abc_17692_n5380), .Y(_abc_17692_n5381) );
  INVX1 INVX1_963 ( .A(_abc_17692_n5384), .Y(_abc_17692_n5385) );
  INVX1 INVX1_964 ( .A(_abc_17692_n5390), .Y(_abc_17692_n5392) );
  INVX1 INVX1_965 ( .A(_abc_17692_n5395), .Y(_abc_17692_n5396) );
  INVX1 INVX1_966 ( .A(_abc_17692_n5398), .Y(_abc_17692_n5399) );
  INVX1 INVX1_967 ( .A(_abc_17692_n5401), .Y(_abc_17692_n5402) );
  INVX1 INVX1_968 ( .A(_abc_17692_n5403), .Y(_abc_17692_n5404) );
  INVX1 INVX1_969 ( .A(_abc_17692_n5407), .Y(_abc_17692_n5408) );
  INVX1 INVX1_97 ( .A(sum_12_), .Y(_abc_17692_n1206_1) );
  INVX1 INVX1_970 ( .A(_abc_17692_n5394), .Y(_abc_17692_n5412) );
  INVX1 INVX1_971 ( .A(_abc_17692_n5410), .Y(_abc_17692_n5413) );
  INVX1 INVX1_972 ( .A(_abc_17692_n5416), .Y(_abc_17692_n5417) );
  INVX1 INVX1_973 ( .A(_abc_17692_n5420_1), .Y(_abc_17692_n5421) );
  INVX1 INVX1_974 ( .A(_abc_17692_n5423_1), .Y(_abc_17692_n5424) );
  INVX1 INVX1_975 ( .A(_abc_17692_n5425), .Y(_abc_17692_n5426) );
  INVX1 INVX1_976 ( .A(_abc_17692_n5431), .Y(_abc_17692_n5432) );
  INVX1 INVX1_977 ( .A(_abc_17692_n5434), .Y(_abc_17692_n5441) );
  INVX1 INVX1_978 ( .A(_abc_17692_n5439), .Y(_abc_17692_n5442) );
  INVX1 INVX1_979 ( .A(_abc_17692_n5444), .Y(_abc_17692_n5446) );
  INVX1 INVX1_98 ( .A(_abc_17692_n1208), .Y(_abc_17692_n1209) );
  INVX1 INVX1_980 ( .A(_abc_17692_n5448), .Y(_abc_17692_n5450) );
  INVX1 INVX1_981 ( .A(_abc_17692_n5452), .Y(_abc_17692_n5453) );
  INVX1 INVX1_982 ( .A(_abc_17692_n5454), .Y(_abc_17692_n5455) );
  INVX1 INVX1_983 ( .A(_abc_17692_n5457), .Y(_abc_17692_n5458) );
  INVX1 INVX1_984 ( .A(_abc_17692_n5462), .Y(_abc_17692_n5463) );
  INVX1 INVX1_985 ( .A(_abc_17692_n5223), .Y(_abc_17692_n5469) );
  INVX1 INVX1_986 ( .A(_abc_17692_n5471), .Y(_abc_17692_n5472) );
  INVX1 INVX1_987 ( .A(_abc_17692_n5474), .Y(_abc_17692_n5475) );
  INVX1 INVX1_988 ( .A(_abc_17692_n5473), .Y(_abc_17692_n5479) );
  INVX1 INVX1_989 ( .A(_abc_17692_n5477), .Y(_abc_17692_n5480) );
  INVX1 INVX1_99 ( .A(_abc_17692_n1210), .Y(_abc_17692_n1211) );
  INVX1 INVX1_990 ( .A(_abc_17692_n5482), .Y(_abc_17692_n5483) );
  INVX1 INVX1_991 ( .A(_abc_17692_n5486), .Y(_abc_17692_n5488) );
  INVX1 INVX1_992 ( .A(_abc_17692_n5490), .Y(_abc_17692_n5491) );
  INVX1 INVX1_993 ( .A(_abc_17692_n5494), .Y(_abc_17692_n5495) );
  INVX1 INVX1_994 ( .A(_abc_17692_n5500), .Y(_abc_17692_n5501) );
  INVX1 INVX1_995 ( .A(_abc_17692_n5307), .Y(_abc_17692_n5508) );
  INVX1 INVX1_996 ( .A(_abc_17692_n5510), .Y(_abc_17692_n5511) );
  INVX1 INVX1_997 ( .A(_abc_17692_n5513), .Y(_abc_17692_n5514) );
  INVX1 INVX1_998 ( .A(_abc_17692_n5512), .Y(_abc_17692_n5518) );
  INVX1 INVX1_999 ( .A(_abc_17692_n5516), .Y(_abc_17692_n5519) );
  INVX2 INVX2_1 ( .A(_abc_17692_n1127_1), .Y(_abc_17692_n1132) );
  INVX2 INVX2_10 ( .A(workunit1_7_), .Y(_abc_17692_n2063) );
  INVX2 INVX2_11 ( .A(workunit1_8_bF_buf1), .Y(_abc_17692_n2250) );
  INVX2 INVX2_12 ( .A(workunit1_9_), .Y(_abc_17692_n2435) );
  INVX2 INVX2_13 ( .A(_abc_17692_n2458), .Y(_abc_17692_n2459_1) );
  INVX2 INVX2_14 ( .A(workunit1_10_), .Y(_abc_17692_n2638) );
  INVX2 INVX2_15 ( .A(workunit1_6_), .Y(_abc_17692_n2821) );
  INVX2 INVX2_16 ( .A(workunit1_11_bF_buf1), .Y(_abc_17692_n2823) );
  INVX2 INVX2_17 ( .A(workunit2_8_bF_buf2), .Y(_abc_17692_n3198) );
  INVX2 INVX2_18 ( .A(workunit1_13_bF_buf2), .Y(_abc_17692_n3208) );
  INVX2 INVX2_19 ( .A(_abc_17692_n3453), .Y(_abc_17692_n3465) );
  INVX2 INVX2_2 ( .A(_abc_17692_n1184), .Y(_abc_17692_n1185) );
  INVX2 INVX2_20 ( .A(workunit2_9_), .Y(_abc_17692_n3471) );
  INVX2 INVX2_21 ( .A(workunit1_15_), .Y(_abc_17692_n3614) );
  INVX2 INVX2_22 ( .A(workunit2_10_bF_buf0), .Y(_abc_17692_n3751) );
  INVX2 INVX2_23 ( .A(workunit2_11_), .Y(_abc_17692_n3905) );
  INVX2 INVX2_24 ( .A(workunit1_17_), .Y(_abc_17692_n4059) );
  INVX2 INVX2_25 ( .A(_abc_17692_n4074), .Y(_abc_17692_n4096_1) );
  INVX2 INVX2_26 ( .A(workunit1_18_), .Y(_abc_17692_n4322) );
  INVX2 INVX2_27 ( .A(_abc_17692_n4333), .Y(_abc_17692_n4334) );
  INVX2 INVX2_28 ( .A(workunit2_13_), .Y(_abc_17692_n4351) );
  INVX2 INVX2_29 ( .A(workunit1_19_), .Y(_abc_17692_n4494) );
  INVX2 INVX2_3 ( .A(_abc_17692_n1250), .Y(_abc_17692_n1251) );
  INVX2 INVX2_30 ( .A(workunit1_20_), .Y(_abc_17692_n4730) );
  INVX2 INVX2_31 ( .A(workunit2_15_), .Y(_abc_17692_n4765) );
  INVX2 INVX2_32 ( .A(workunit1_21_), .Y(_abc_17692_n4926) );
  INVX2 INVX2_33 ( .A(_abc_17692_n4944), .Y(_abc_17692_n4967) );
  INVX2 INVX2_34 ( .A(workunit1_22_), .Y(_abc_17692_n5205) );
  INVX2 INVX2_35 ( .A(workunit2_17_), .Y(_abc_17692_n5260) );
  INVX2 INVX2_36 ( .A(workunit1_14_bF_buf2), .Y(_abc_17692_n5376) );
  INVX2 INVX2_37 ( .A(workunit1_23_), .Y(_abc_17692_n5378) );
  INVX2 INVX2_38 ( .A(workunit2_18_), .Y(_abc_17692_n5430) );
  INVX2 INVX2_39 ( .A(workunit1_24_), .Y(_abc_17692_n5598) );
  INVX2 INVX2_4 ( .A(_abc_17692_n1307), .Y(_abc_17692_n1312) );
  INVX2 INVX2_40 ( .A(_abc_17692_n5610), .Y(_abc_17692_n5611_1) );
  INVX2 INVX2_41 ( .A(workunit2_19_), .Y(_abc_17692_n5626) );
  INVX2 INVX2_42 ( .A(workunit2_20_), .Y(_abc_17692_n5769) );
  INVX2 INVX2_43 ( .A(workunit1_25_), .Y(_abc_17692_n5782) );
  INVX2 INVX2_44 ( .A(_abc_17692_n5795), .Y(_abc_17692_n5817) );
  INVX2 INVX2_45 ( .A(workunit1_26_), .Y(_abc_17692_n6065) );
  INVX2 INVX2_46 ( .A(workunit2_21_), .Y(_abc_17692_n6095) );
  INVX2 INVX2_47 ( .A(workunit1_27_), .Y(_abc_17692_n6242) );
  INVX2 INVX2_48 ( .A(workunit2_22_), .Y(_abc_17692_n6293) );
  INVX2 INVX2_49 ( .A(_abc_17692_n6397), .Y(_abc_17692_n6398) );
  INVX2 INVX2_5 ( .A(sum_31_), .Y(_abc_17692_n1792) );
  INVX2 INVX2_50 ( .A(workunit1_28_), .Y(_abc_17692_n6468_1) );
  INVX2 INVX2_51 ( .A(workunit2_23_), .Y(_abc_17692_n6505) );
  INVX2 INVX2_52 ( .A(workunit2_24_), .Y(_abc_17692_n6657_1) );
  INVX2 INVX2_53 ( .A(workunit1_29_), .Y(_abc_17692_n6659_1) );
  INVX2 INVX2_54 ( .A(_abc_17692_n6681), .Y(_abc_17692_n6702) );
  INVX2 INVX2_55 ( .A(workunit2_25_), .Y(_abc_17692_n6952) );
  INVX2 INVX2_56 ( .A(workunit1_30_), .Y(_abc_17692_n6956) );
  INVX2 INVX2_57 ( .A(workunit2_26_), .Y(_abc_17692_n7128) );
  INVX2 INVX2_58 ( .A(workunit2_27_), .Y(_abc_17692_n7385) );
  INVX2 INVX2_59 ( .A(workunit2_28_), .Y(_abc_17692_n7535) );
  INVX2 INVX2_6 ( .A(workunit2_0_), .Y(_abc_17692_n1814) );
  INVX2 INVX2_60 ( .A(_abc_17692_n7792), .Y(_abc_17692_n7805) );
  INVX2 INVX2_61 ( .A(workunit2_29_), .Y(_abc_17692_n7812) );
  INVX2 INVX2_62 ( .A(workunit2_30_), .Y(_abc_17692_n7968) );
  INVX2 INVX2_63 ( .A(_abc_17692_n8056), .Y(_abc_17692_n8058) );
  INVX2 INVX2_64 ( .A(_abc_17692_n8215), .Y(_abc_17692_n8218) );
  INVX2 INVX2_65 ( .A(_abc_17692_n8765), .Y(_abc_17692_n8767) );
  INVX2 INVX2_66 ( .A(_abc_17692_n9297), .Y(_abc_17692_n9298) );
  INVX2 INVX2_67 ( .A(_abc_17692_n9433), .Y(_abc_17692_n9434) );
  INVX2 INVX2_68 ( .A(_abc_17692_n9877), .Y(_abc_17692_n9878) );
  INVX2 INVX2_69 ( .A(_abc_17692_n10078), .Y(_abc_17692_n10080) );
  INVX2 INVX2_7 ( .A(workunit1_0_), .Y(_abc_17692_n1816) );
  INVX2 INVX2_70 ( .A(_abc_17692_n10500), .Y(_abc_17692_n10501) );
  INVX2 INVX2_71 ( .A(_abc_17692_n10811), .Y(_abc_17692_n10812) );
  INVX2 INVX2_72 ( .A(_abc_17692_n11109), .Y(_abc_17692_n11110) );
  INVX2 INVX2_73 ( .A(_abc_17692_n11307), .Y(_abc_17692_n11309) );
  INVX2 INVX2_74 ( .A(_abc_17692_n11733), .Y(_abc_17692_n11734) );
  INVX2 INVX2_75 ( .A(_abc_17692_n11938), .Y(_abc_17692_n11940) );
  INVX2 INVX2_76 ( .A(_abc_17692_n12222), .Y(_abc_17692_n12224) );
  INVX2 INVX2_77 ( .A(_abc_17692_n12349), .Y(_abc_17692_n12350) );
  INVX2 INVX2_78 ( .A(_abc_17692_n12532), .Y(_abc_17692_n12534) );
  INVX2 INVX2_79 ( .A(_abc_17692_n12657), .Y(_abc_17692_n12659) );
  INVX2 INVX2_8 ( .A(workunit1_5_), .Y(_abc_17692_n1817) );
  INVX2 INVX2_9 ( .A(workunit1_2_), .Y(_abc_17692_n2062_1) );
  INVX4 INVX4_1 ( .A(state_8_bF_buf7), .Y(_abc_17692_n632) );
  INVX4 INVX4_10 ( .A(workunit2_6_), .Y(_abc_17692_n2862) );
  INVX4 INVX4_11 ( .A(workunit2_7_), .Y(_abc_17692_n3060) );
  INVX4 INVX4_2 ( .A(_abc_17692_n721), .Y(_abc_17692_n722) );
  INVX4 INVX4_3 ( .A(workunit2_1_bF_buf1), .Y(_abc_17692_n1919_1) );
  INVX4 INVX4_4 ( .A(workunit2_2_), .Y(_abc_17692_n2091) );
  INVX4 INVX4_5 ( .A(workunit2_3_), .Y(_abc_17692_n2246) );
  INVX4 INVX4_6 ( .A(workunit1_3_), .Y(_abc_17692_n2249) );
  INVX4 INVX4_7 ( .A(workunit1_4_), .Y(_abc_17692_n2433) );
  INVX4 INVX4_8 ( .A(workunit2_4_), .Y(_abc_17692_n2482) );
  INVX4 INVX4_9 ( .A(workunit2_5_), .Y(_abc_17692_n2633) );
  INVX8 INVX8_1 ( .A(_abc_17692_n725_bF_buf6), .Y(_abc_17692_n727) );
  INVX8 INVX8_2 ( .A(_abc_17692_n1863_bF_buf9), .Y(_abc_17692_n4047) );
  INVX8 INVX8_3 ( .A(reset), .Y(_abc_17692_n6660) );
  OR2X2 OR2X2_1 ( .A(_abc_17692_n624), .B(state_12_), .Y(_abc_10892_n1037) );
  OR2X2 OR2X2_10 ( .A(state_8_bF_buf1), .B(delta_8_), .Y(delta_8__FF_INPUT) );
  OR2X2 OR2X2_100 ( .A(_abc_17692_n725_bF_buf1), .B(_auto_iopadmap_cc_313_execute_30065_29_), .Y(_abc_17692_n814_1) );
  OR2X2 OR2X2_1000 ( .A(_abc_17692_n3092), .B(_abc_17692_n3256), .Y(_abc_17692_n3257) );
  OR2X2 OR2X2_1001 ( .A(_abc_17692_n3258_1), .B(_abc_17692_n3255), .Y(_abc_17692_n3259) );
  OR2X2 OR2X2_1002 ( .A(_abc_17692_n3119), .B(_abc_17692_n3123), .Y(_abc_17692_n3265) );
  OR2X2 OR2X2_1003 ( .A(_abc_17692_n3120), .B(_abc_17692_n2931), .Y(_abc_17692_n3267) );
  OR2X2 OR2X2_1004 ( .A(_abc_17692_n3267), .B(_abc_17692_n2940), .Y(_abc_17692_n3268) );
  OR2X2 OR2X2_1005 ( .A(_abc_17692_n3275), .B(_abc_17692_n3100), .Y(_abc_17692_n3276) );
  OR2X2 OR2X2_1006 ( .A(_abc_17692_n3274), .B(_abc_17692_n3276), .Y(_abc_17692_n3277) );
  OR2X2 OR2X2_1007 ( .A(_abc_17692_n3273), .B(_abc_17692_n3277), .Y(_abc_17692_n3278_1) );
  OR2X2 OR2X2_1008 ( .A(sum_8_), .B(\key_in[40] ), .Y(_abc_17692_n3281) );
  OR2X2 OR2X2_1009 ( .A(_abc_17692_n2538_1), .B(_abc_17692_n3284), .Y(_abc_17692_n3285) );
  OR2X2 OR2X2_101 ( .A(_abc_17692_n727_bF_buf2), .B(workunit2_29_), .Y(_abc_17692_n815_1) );
  OR2X2 OR2X2_1010 ( .A(_abc_17692_n3289), .B(_abc_17692_n3283), .Y(_abc_17692_n3290) );
  OR2X2 OR2X2_1011 ( .A(_abc_17692_n3291), .B(_abc_17692_n3228), .Y(_abc_17692_n3292) );
  OR2X2 OR2X2_1012 ( .A(_abc_17692_n3248), .B(_abc_17692_n3290), .Y(_abc_17692_n3293) );
  OR2X2 OR2X2_1013 ( .A(_abc_17692_n3294), .B(workunit2_8_bF_buf3), .Y(_abc_17692_n3297) );
  OR2X2 OR2X2_1014 ( .A(_abc_17692_n3270), .B(_abc_17692_n3298), .Y(_abc_17692_n3299) );
  OR2X2 OR2X2_1015 ( .A(_abc_17692_n3308), .B(_abc_17692_n3044), .Y(_abc_17692_n3309) );
  OR2X2 OR2X2_1016 ( .A(_abc_17692_n3307), .B(_abc_17692_n3309), .Y(_abc_17692_n3310) );
  OR2X2 OR2X2_1017 ( .A(_abc_17692_n3306), .B(_abc_17692_n3310), .Y(_abc_17692_n3311) );
  OR2X2 OR2X2_1018 ( .A(sum_8_), .B(\key_in[8] ), .Y(_abc_17692_n3314) );
  OR2X2 OR2X2_1019 ( .A(_abc_17692_n2473), .B(_abc_17692_n3317), .Y(_abc_17692_n3318) );
  OR2X2 OR2X2_102 ( .A(_abc_17692_n725_bF_buf0), .B(_auto_iopadmap_cc_313_execute_30065_30_), .Y(_abc_17692_n817) );
  OR2X2 OR2X2_1020 ( .A(_abc_17692_n3322), .B(_abc_17692_n3316), .Y(_abc_17692_n3323) );
  OR2X2 OR2X2_1021 ( .A(_abc_17692_n3324), .B(_abc_17692_n3228), .Y(_abc_17692_n3325) );
  OR2X2 OR2X2_1022 ( .A(_abc_17692_n3248), .B(_abc_17692_n3323), .Y(_abc_17692_n3326) );
  OR2X2 OR2X2_1023 ( .A(_abc_17692_n3327), .B(workunit2_8_bF_buf1), .Y(_abc_17692_n3330) );
  OR2X2 OR2X2_1024 ( .A(_abc_17692_n3333), .B(_abc_17692_n3336), .Y(_abc_17692_n3337) );
  OR2X2 OR2X2_1025 ( .A(_abc_17692_n3338), .B(_abc_17692_n3331), .Y(_abc_17692_n3339) );
  OR2X2 OR2X2_1026 ( .A(_abc_17692_n3343), .B(_abc_17692_n3303), .Y(_abc_17692_n3344) );
  OR2X2 OR2X2_1027 ( .A(_abc_17692_n3344), .B(_abc_17692_n3263), .Y(_abc_17692_n3345) );
  OR2X2 OR2X2_1028 ( .A(sum_8_), .B(\key_in[104] ), .Y(_abc_17692_n3350) );
  OR2X2 OR2X2_1029 ( .A(_abc_17692_n3352), .B(_abc_17692_n3133), .Y(_abc_17692_n3353) );
  OR2X2 OR2X2_103 ( .A(_abc_17692_n727_bF_buf1), .B(workunit2_30_), .Y(_abc_17692_n818) );
  OR2X2 OR2X2_1030 ( .A(_abc_17692_n3355_1), .B(_abc_17692_n3353), .Y(_abc_17692_n3356) );
  OR2X2 OR2X2_1031 ( .A(_abc_17692_n3358), .B(_abc_17692_n3356), .Y(_abc_17692_n3359) );
  OR2X2 OR2X2_1032 ( .A(_abc_17692_n3365), .B(_abc_17692_n3360), .Y(_abc_17692_n3366_1) );
  OR2X2 OR2X2_1033 ( .A(_abc_17692_n3369), .B(_abc_17692_n3367), .Y(_abc_17692_n3370) );
  OR2X2 OR2X2_1034 ( .A(_abc_17692_n3370), .B(workunit2_8_bF_buf3), .Y(_abc_17692_n3373) );
  OR2X2 OR2X2_1035 ( .A(_abc_17692_n3347), .B(_abc_17692_n3374), .Y(_abc_17692_n3375) );
  OR2X2 OR2X2_1036 ( .A(_abc_17692_n3345), .B(_abc_17692_n3379), .Y(_abc_17692_n3380) );
  OR2X2 OR2X2_1037 ( .A(_abc_17692_n3145), .B(_abc_17692_n3060), .Y(_abc_17692_n3383) );
  OR2X2 OR2X2_1038 ( .A(_abc_17692_n3385), .B(_abc_17692_n3384), .Y(_abc_17692_n3386) );
  OR2X2 OR2X2_1039 ( .A(_abc_17692_n3386), .B(_abc_17692_n3382), .Y(_abc_17692_n3387) );
  OR2X2 OR2X2_104 ( .A(_abc_17692_n725_bF_buf7), .B(_auto_iopadmap_cc_313_execute_30065_31_), .Y(_abc_17692_n820) );
  OR2X2 OR2X2_1040 ( .A(_abc_17692_n3392), .B(_abc_17692_n3396), .Y(_abc_17692_n3397) );
  OR2X2 OR2X2_1041 ( .A(_abc_17692_n3397), .B(_abc_17692_n3254), .Y(_abc_17692_n3400) );
  OR2X2 OR2X2_1042 ( .A(_abc_17692_n3406), .B(_abc_17692_n3404), .Y(_abc_17692_n3407) );
  OR2X2 OR2X2_1043 ( .A(_abc_17692_n3409), .B(_abc_17692_n3407), .Y(_abc_17692_n3410) );
  OR2X2 OR2X2_1044 ( .A(_abc_17692_n3410), .B(_abc_17692_n3403), .Y(_abc_17692_n3411) );
  OR2X2 OR2X2_1045 ( .A(_abc_17692_n3418), .B(_abc_17692_n3417), .Y(_abc_17692_n3419) );
  OR2X2 OR2X2_1046 ( .A(_abc_17692_n3419), .B(_abc_17692_n3421), .Y(_abc_17692_n3422) );
  OR2X2 OR2X2_1047 ( .A(_abc_17692_n3422), .B(_abc_17692_n3416), .Y(_abc_17692_n3425) );
  OR2X2 OR2X2_1048 ( .A(_abc_17692_n3415), .B(_abc_17692_n3427_1), .Y(_abc_17692_n3428) );
  OR2X2 OR2X2_1049 ( .A(_abc_17692_n3428), .B(_abc_17692_n3402), .Y(_abc_17692_n3429) );
  OR2X2 OR2X2_105 ( .A(_abc_17692_n727_bF_buf0), .B(workunit2_31_), .Y(_abc_17692_n821) );
  OR2X2 OR2X2_1050 ( .A(_abc_17692_n3429), .B(_abc_17692_n3391), .Y(_abc_17692_n3430) );
  OR2X2 OR2X2_1051 ( .A(_abc_17692_n3432), .B(_abc_17692_n3433), .Y(_abc_17692_n3434) );
  OR2X2 OR2X2_1052 ( .A(_abc_17692_n3431), .B(_abc_17692_n3434), .Y(_abc_17692_n3435) );
  OR2X2 OR2X2_1053 ( .A(_abc_17692_n3435), .B(_abc_17692_n3381), .Y(workunit2_8__FF_INPUT) );
  OR2X2 OR2X2_1054 ( .A(_abc_17692_n3219), .B(_abc_17692_n3212), .Y(_abc_17692_n3439) );
  OR2X2 OR2X2_1055 ( .A(workunit1_5_), .B(workunit1_14_bF_buf1), .Y(_abc_17692_n3443) );
  OR2X2 OR2X2_1056 ( .A(_abc_17692_n3446), .B(_abc_17692_n3441), .Y(_abc_17692_n3447) );
  OR2X2 OR2X2_1057 ( .A(_abc_17692_n3448), .B(_abc_17692_n3445), .Y(_abc_17692_n3449) );
  OR2X2 OR2X2_1058 ( .A(_abc_17692_n3451), .B(_abc_17692_n3452), .Y(_abc_17692_n3453) );
  OR2X2 OR2X2_1059 ( .A(_abc_17692_n3241), .B(_abc_17692_n3237), .Y(_abc_17692_n3454) );
  OR2X2 OR2X2_106 ( .A(_abc_17692_n725_bF_buf6), .B(_auto_iopadmap_cc_313_execute_30032_0_), .Y(_abc_17692_n823) );
  OR2X2 OR2X2_1060 ( .A(sum_9_), .B(\key_in[73] ), .Y(_abc_17692_n3458) );
  OR2X2 OR2X2_1061 ( .A(_abc_17692_n3460), .B(_abc_17692_n3462), .Y(_abc_17692_n3463) );
  OR2X2 OR2X2_1062 ( .A(_abc_17692_n3467), .B(_abc_17692_n3464), .Y(_abc_17692_n3468) );
  OR2X2 OR2X2_1063 ( .A(_abc_17692_n3470), .B(_abc_17692_n3472_1), .Y(_abc_17692_n3473) );
  OR2X2 OR2X2_1064 ( .A(_abc_17692_n3477), .B(_abc_17692_n3474), .Y(_abc_17692_n3478) );
  OR2X2 OR2X2_1065 ( .A(_abc_17692_n3283), .B(_abc_17692_n3279), .Y(_abc_17692_n3482) );
  OR2X2 OR2X2_1066 ( .A(sum_9_), .B(\key_in[41] ), .Y(_abc_17692_n3486) );
  OR2X2 OR2X2_1067 ( .A(_abc_17692_n3483), .B(_abc_17692_n3487), .Y(_abc_17692_n3489) );
  OR2X2 OR2X2_1068 ( .A(_abc_17692_n3490), .B(_abc_17692_n3488), .Y(_abc_17692_n3491) );
  OR2X2 OR2X2_1069 ( .A(_abc_17692_n3465), .B(_abc_17692_n3491), .Y(_abc_17692_n3492) );
  OR2X2 OR2X2_107 ( .A(_abc_17692_n727_bF_buf7), .B(workunit1_0_), .Y(_abc_17692_n824) );
  OR2X2 OR2X2_1070 ( .A(_abc_17692_n3494), .B(_abc_17692_n3453), .Y(_abc_17692_n3495) );
  OR2X2 OR2X2_1071 ( .A(_abc_17692_n3496), .B(_abc_17692_n3471), .Y(_abc_17692_n3497) );
  OR2X2 OR2X2_1072 ( .A(_abc_17692_n3465), .B(_abc_17692_n3494), .Y(_abc_17692_n3498) );
  OR2X2 OR2X2_1073 ( .A(_abc_17692_n3491), .B(_abc_17692_n3453), .Y(_abc_17692_n3499) );
  OR2X2 OR2X2_1074 ( .A(_abc_17692_n3500), .B(workunit2_9_), .Y(_abc_17692_n3501) );
  OR2X2 OR2X2_1075 ( .A(_abc_17692_n3481), .B(_abc_17692_n3503_1), .Y(_abc_17692_n3504) );
  OR2X2 OR2X2_1076 ( .A(_abc_17692_n3480), .B(_abc_17692_n3502), .Y(_abc_17692_n3505) );
  OR2X2 OR2X2_1077 ( .A(_abc_17692_n3316), .B(_abc_17692_n3312), .Y(_abc_17692_n3510) );
  OR2X2 OR2X2_1078 ( .A(sum_9_), .B(\key_in[9] ), .Y(_abc_17692_n3513) );
  OR2X2 OR2X2_1079 ( .A(_abc_17692_n3510), .B(_abc_17692_n3515), .Y(_abc_17692_n3516) );
  OR2X2 OR2X2_108 ( .A(_abc_17692_n725_bF_buf5), .B(_auto_iopadmap_cc_313_execute_30032_1_), .Y(_abc_17692_n826) );
  OR2X2 OR2X2_1080 ( .A(_abc_17692_n3465), .B(_abc_17692_n3519), .Y(_abc_17692_n3520) );
  OR2X2 OR2X2_1081 ( .A(_abc_17692_n3521), .B(_abc_17692_n3453), .Y(_abc_17692_n3522) );
  OR2X2 OR2X2_1082 ( .A(_abc_17692_n3524), .B(_abc_17692_n3471), .Y(_abc_17692_n3525) );
  OR2X2 OR2X2_1083 ( .A(_abc_17692_n3523), .B(workunit2_9_), .Y(_abc_17692_n3526) );
  OR2X2 OR2X2_1084 ( .A(_abc_17692_n3509), .B(_abc_17692_n3528), .Y(_abc_17692_n3529) );
  OR2X2 OR2X2_1085 ( .A(_abc_17692_n3508), .B(_abc_17692_n3527), .Y(_abc_17692_n3530) );
  OR2X2 OR2X2_1086 ( .A(_abc_17692_n3532), .B(_abc_17692_n3507), .Y(_abc_17692_n3533_1) );
  OR2X2 OR2X2_1087 ( .A(_abc_17692_n3479), .B(_abc_17692_n3533_1), .Y(_abc_17692_n3534) );
  OR2X2 OR2X2_1088 ( .A(_abc_17692_n3360), .B(_abc_17692_n3348), .Y(_abc_17692_n3536) );
  OR2X2 OR2X2_1089 ( .A(sum_9_), .B(\key_in[105] ), .Y(_abc_17692_n3539) );
  OR2X2 OR2X2_109 ( .A(_abc_17692_n727_bF_buf6), .B(workunit1_1_bF_buf3), .Y(_abc_17692_n827) );
  OR2X2 OR2X2_1090 ( .A(_abc_17692_n3536), .B(_abc_17692_n3541), .Y(_abc_17692_n3542) );
  OR2X2 OR2X2_1091 ( .A(_abc_17692_n3545), .B(_abc_17692_n3465), .Y(_abc_17692_n3546) );
  OR2X2 OR2X2_1092 ( .A(_abc_17692_n3547), .B(_abc_17692_n3453), .Y(_abc_17692_n3548) );
  OR2X2 OR2X2_1093 ( .A(_abc_17692_n3550), .B(_abc_17692_n3471), .Y(_abc_17692_n3551) );
  OR2X2 OR2X2_1094 ( .A(_abc_17692_n3549), .B(workunit2_9_), .Y(_abc_17692_n3552) );
  OR2X2 OR2X2_1095 ( .A(_abc_17692_n3557), .B(_abc_17692_n3555), .Y(_abc_17692_n3558) );
  OR2X2 OR2X2_1096 ( .A(_abc_17692_n3534), .B(_abc_17692_n3559), .Y(_abc_17692_n3560) );
  OR2X2 OR2X2_1097 ( .A(_abc_17692_n3567), .B(_abc_17692_n3568), .Y(_abc_17692_n3569) );
  OR2X2 OR2X2_1098 ( .A(_abc_17692_n3574), .B(_abc_17692_n3476), .Y(_abc_17692_n3575) );
  OR2X2 OR2X2_1099 ( .A(_abc_17692_n3573), .B(_abc_17692_n3473), .Y(_abc_17692_n3576) );
  OR2X2 OR2X2_11 ( .A(state_8_bF_buf0), .B(delta_11_), .Y(delta_11__FF_INPUT) );
  OR2X2 OR2X2_110 ( .A(_abc_17692_n725_bF_buf4), .B(_auto_iopadmap_cc_313_execute_30032_2_), .Y(_abc_17692_n829) );
  OR2X2 OR2X2_1100 ( .A(_abc_17692_n3582), .B(_abc_17692_n3528), .Y(_abc_17692_n3583) );
  OR2X2 OR2X2_1101 ( .A(_abc_17692_n3584), .B(_abc_17692_n3527), .Y(_abc_17692_n3585) );
  OR2X2 OR2X2_1102 ( .A(_abc_17692_n3592), .B(_abc_17692_n3502), .Y(_abc_17692_n3593) );
  OR2X2 OR2X2_1103 ( .A(_abc_17692_n3591), .B(_abc_17692_n3503_1), .Y(_abc_17692_n3594) );
  OR2X2 OR2X2_1104 ( .A(_abc_17692_n3587), .B(_abc_17692_n3596), .Y(_abc_17692_n3597) );
  OR2X2 OR2X2_1105 ( .A(_abc_17692_n3597), .B(_abc_17692_n3578), .Y(_abc_17692_n3598) );
  OR2X2 OR2X2_1106 ( .A(_abc_17692_n3598), .B(_abc_17692_n3570), .Y(_abc_17692_n3599) );
  OR2X2 OR2X2_1107 ( .A(_abc_17692_n3601), .B(_abc_17692_n3602), .Y(_abc_17692_n3603) );
  OR2X2 OR2X2_1108 ( .A(_abc_17692_n3600), .B(_abc_17692_n3603), .Y(_abc_17692_n3604) );
  OR2X2 OR2X2_1109 ( .A(_abc_17692_n3604), .B(_abc_17692_n3561), .Y(workunit2_9__FF_INPUT) );
  OR2X2 OR2X2_111 ( .A(_abc_17692_n727_bF_buf5), .B(workunit1_2_), .Y(_abc_17692_n830) );
  OR2X2 OR2X2_1110 ( .A(_abc_17692_n3449), .B(_abc_17692_n3217), .Y(_abc_17692_n3606) );
  OR2X2 OR2X2_1111 ( .A(_abc_17692_n3212), .B(_abc_17692_n3445), .Y(_abc_17692_n3610) );
  OR2X2 OR2X2_1112 ( .A(_abc_17692_n3608), .B(_abc_17692_n3611), .Y(_abc_17692_n3612) );
  OR2X2 OR2X2_1113 ( .A(_abc_17692_n2821), .B(workunit1_15_), .Y(_abc_17692_n3613) );
  OR2X2 OR2X2_1114 ( .A(_abc_17692_n3614), .B(workunit1_6_), .Y(_abc_17692_n3615) );
  OR2X2 OR2X2_1115 ( .A(_abc_17692_n3616), .B(_abc_17692_n2638), .Y(_abc_17692_n3617) );
  OR2X2 OR2X2_1116 ( .A(_abc_17692_n3618_1), .B(_abc_17692_n3619), .Y(_abc_17692_n3620) );
  OR2X2 OR2X2_1117 ( .A(_abc_17692_n3620), .B(workunit1_10_), .Y(_abc_17692_n3621_1) );
  OR2X2 OR2X2_1118 ( .A(_abc_17692_n3226), .B(_abc_17692_n3606), .Y(_abc_17692_n3624) );
  OR2X2 OR2X2_1119 ( .A(_abc_17692_n3215), .B(_abc_17692_n2250), .Y(_abc_17692_n3626) );
  OR2X2 OR2X2_112 ( .A(_abc_17692_n725_bF_buf3), .B(_auto_iopadmap_cc_313_execute_30032_3_), .Y(_abc_17692_n832) );
  OR2X2 OR2X2_1120 ( .A(_abc_17692_n3448), .B(_abc_17692_n3626), .Y(_abc_17692_n3627) );
  OR2X2 OR2X2_1121 ( .A(_abc_17692_n3630_1), .B(_abc_17692_n3631), .Y(_abc_17692_n3632) );
  OR2X2 OR2X2_1122 ( .A(_abc_17692_n3633), .B(_abc_17692_n3623), .Y(_abc_17692_n3634) );
  OR2X2 OR2X2_1123 ( .A(_abc_17692_n3638), .B(_abc_17692_n3637), .Y(_abc_17692_n3639) );
  OR2X2 OR2X2_1124 ( .A(_abc_17692_n3636), .B(_abc_17692_n3640_1), .Y(_abc_17692_n3641) );
  OR2X2 OR2X2_1125 ( .A(sum_10_), .B(\key_in[74] ), .Y(_abc_17692_n3644) );
  OR2X2 OR2X2_1126 ( .A(_abc_17692_n3649), .B(_abc_17692_n3646), .Y(_abc_17692_n3650_1) );
  OR2X2 OR2X2_1127 ( .A(_abc_17692_n3651), .B(_abc_17692_n3634), .Y(_abc_17692_n3652) );
  OR2X2 OR2X2_1128 ( .A(_abc_17692_n3653), .B(_abc_17692_n3650_1), .Y(_abc_17692_n3654) );
  OR2X2 OR2X2_1129 ( .A(_abc_17692_n3655), .B(workunit2_10_bF_buf1), .Y(_abc_17692_n3658) );
  OR2X2 OR2X2_113 ( .A(_abc_17692_n727_bF_buf4), .B(workunit1_3_), .Y(_abc_17692_n833) );
  OR2X2 OR2X2_1130 ( .A(_abc_17692_n3660), .B(_abc_17692_n3662), .Y(_abc_17692_n3663) );
  OR2X2 OR2X2_1131 ( .A(_abc_17692_n3665), .B(_abc_17692_n3664), .Y(_abc_17692_n3666) );
  OR2X2 OR2X2_1132 ( .A(_abc_17692_n3669), .B(_abc_17692_n3659), .Y(_abc_17692_n3670) );
  OR2X2 OR2X2_1133 ( .A(_abc_17692_n3279), .B(_abc_17692_n3484), .Y(_abc_17692_n3677) );
  OR2X2 OR2X2_1134 ( .A(_abc_17692_n3676), .B(_abc_17692_n3678), .Y(_abc_17692_n3679) );
  OR2X2 OR2X2_1135 ( .A(sum_10_), .B(\key_in[42] ), .Y(_abc_17692_n3682) );
  OR2X2 OR2X2_1136 ( .A(_abc_17692_n3689), .B(_abc_17692_n3684), .Y(_abc_17692_n3690) );
  OR2X2 OR2X2_1137 ( .A(_abc_17692_n3691), .B(_abc_17692_n3693), .Y(_abc_17692_n3694) );
  OR2X2 OR2X2_1138 ( .A(_abc_17692_n3694), .B(workunit2_10_bF_buf3), .Y(_abc_17692_n3697) );
  OR2X2 OR2X2_1139 ( .A(_abc_17692_n3502), .B(_abc_17692_n3403), .Y(_abc_17692_n3700) );
  OR2X2 OR2X2_114 ( .A(_abc_17692_n725_bF_buf2), .B(_auto_iopadmap_cc_313_execute_30032_4_), .Y(_abc_17692_n835) );
  OR2X2 OR2X2_1140 ( .A(_abc_17692_n3269), .B(_abc_17692_n3700), .Y(_abc_17692_n3701) );
  OR2X2 OR2X2_1141 ( .A(_abc_17692_n3502), .B(_abc_17692_n3296), .Y(_abc_17692_n3704) );
  OR2X2 OR2X2_1142 ( .A(_abc_17692_n3707), .B(_abc_17692_n3699_1), .Y(_abc_17692_n3710) );
  OR2X2 OR2X2_1143 ( .A(_abc_17692_n3312), .B(_abc_17692_n3511), .Y(_abc_17692_n3715) );
  OR2X2 OR2X2_1144 ( .A(_abc_17692_n3714), .B(_abc_17692_n3716), .Y(_abc_17692_n3717) );
  OR2X2 OR2X2_1145 ( .A(sum_10_), .B(\key_in[10] ), .Y(_abc_17692_n3720) );
  OR2X2 OR2X2_1146 ( .A(_abc_17692_n3725), .B(_abc_17692_n3722), .Y(_abc_17692_n3726) );
  OR2X2 OR2X2_1147 ( .A(_abc_17692_n3727), .B(_abc_17692_n3634), .Y(_abc_17692_n3728) );
  OR2X2 OR2X2_1148 ( .A(_abc_17692_n3653), .B(_abc_17692_n3726), .Y(_abc_17692_n3729) );
  OR2X2 OR2X2_1149 ( .A(_abc_17692_n3730), .B(workunit2_10_bF_buf2), .Y(_abc_17692_n3731) );
  OR2X2 OR2X2_115 ( .A(_abc_17692_n727_bF_buf3), .B(workunit1_4_), .Y(_abc_17692_n836_1) );
  OR2X2 OR2X2_1150 ( .A(_abc_17692_n3527), .B(_abc_17692_n3416), .Y(_abc_17692_n3735) );
  OR2X2 OR2X2_1151 ( .A(_abc_17692_n3527), .B(_abc_17692_n3329), .Y(_abc_17692_n3740) );
  OR2X2 OR2X2_1152 ( .A(_abc_17692_n3737), .B(_abc_17692_n3742), .Y(_abc_17692_n3743) );
  OR2X2 OR2X2_1153 ( .A(_abc_17692_n3743), .B(_abc_17692_n3734), .Y(_abc_17692_n3746) );
  OR2X2 OR2X2_1154 ( .A(_abc_17692_n3748), .B(_abc_17692_n3712_1), .Y(_abc_17692_n3749) );
  OR2X2 OR2X2_1155 ( .A(_abc_17692_n3674), .B(_abc_17692_n3749), .Y(_abc_17692_n3750) );
  OR2X2 OR2X2_1156 ( .A(_abc_17692_n3755), .B(_abc_17692_n3754_1), .Y(_abc_17692_n3756) );
  OR2X2 OR2X2_1157 ( .A(_abc_17692_n3753), .B(_abc_17692_n3757), .Y(_abc_17692_n3758) );
  OR2X2 OR2X2_1158 ( .A(sum_10_), .B(\key_in[106] ), .Y(_abc_17692_n3761) );
  OR2X2 OR2X2_1159 ( .A(_abc_17692_n3766), .B(_abc_17692_n3763), .Y(_abc_17692_n3767) );
  OR2X2 OR2X2_116 ( .A(_abc_17692_n725_bF_buf1), .B(_auto_iopadmap_cc_313_execute_30032_5_), .Y(_abc_17692_n838) );
  OR2X2 OR2X2_1160 ( .A(_abc_17692_n3768), .B(_abc_17692_n3634), .Y(_abc_17692_n3769) );
  OR2X2 OR2X2_1161 ( .A(_abc_17692_n3767), .B(_abc_17692_n3653), .Y(_abc_17692_n3770) );
  OR2X2 OR2X2_1162 ( .A(_abc_17692_n3771), .B(_abc_17692_n3751), .Y(_abc_17692_n3772) );
  OR2X2 OR2X2_1163 ( .A(_abc_17692_n3773), .B(workunit2_10_bF_buf3), .Y(_abc_17692_n3774) );
  OR2X2 OR2X2_1164 ( .A(_abc_17692_n3553), .B(_abc_17692_n3372), .Y(_abc_17692_n3779) );
  OR2X2 OR2X2_1165 ( .A(_abc_17692_n3783), .B(_abc_17692_n3781), .Y(_abc_17692_n3784) );
  OR2X2 OR2X2_1166 ( .A(_abc_17692_n3784), .B(_abc_17692_n3776_1), .Y(_abc_17692_n3785) );
  OR2X2 OR2X2_1167 ( .A(_abc_17692_n3750), .B(_abc_17692_n3789), .Y(_abc_17692_n3790) );
  OR2X2 OR2X2_1168 ( .A(_abc_17692_n3792), .B(_abc_17692_n3794), .Y(_abc_17692_n3795) );
  OR2X2 OR2X2_1169 ( .A(_abc_17692_n3796), .B(_abc_17692_n3797), .Y(_abc_17692_n3798) );
  OR2X2 OR2X2_117 ( .A(_abc_17692_n727_bF_buf2), .B(workunit1_5_), .Y(_abc_17692_n839) );
  OR2X2 OR2X2_1170 ( .A(_abc_17692_n3801), .B(_abc_17692_n3775), .Y(_abc_17692_n3802) );
  OR2X2 OR2X2_1171 ( .A(_abc_17692_n3473), .B(_abc_17692_n3255), .Y(_abc_17692_n3808) );
  OR2X2 OR2X2_1172 ( .A(_abc_17692_n3472_1), .B(_abc_17692_n3572), .Y(_abc_17692_n3812) );
  OR2X2 OR2X2_1173 ( .A(_abc_17692_n3810), .B(_abc_17692_n3814), .Y(_abc_17692_n3815) );
  OR2X2 OR2X2_1174 ( .A(_abc_17692_n3815), .B(_abc_17692_n3807), .Y(_abc_17692_n3818) );
  OR2X2 OR2X2_1175 ( .A(_abc_17692_n3822), .B(_abc_17692_n3823), .Y(_abc_17692_n3824) );
  OR2X2 OR2X2_1176 ( .A(_abc_17692_n3825), .B(_abc_17692_n3827), .Y(_abc_17692_n3828) );
  OR2X2 OR2X2_1177 ( .A(_abc_17692_n3829), .B(_abc_17692_n3589), .Y(_abc_17692_n3830) );
  OR2X2 OR2X2_1178 ( .A(_abc_17692_n3834_1), .B(_abc_17692_n3698), .Y(_abc_17692_n3835) );
  OR2X2 OR2X2_1179 ( .A(_abc_17692_n3841), .B(_abc_17692_n3843_1), .Y(_abc_17692_n3844) );
  OR2X2 OR2X2_118 ( .A(_abc_17692_n725_bF_buf0), .B(_auto_iopadmap_cc_313_execute_30032_6_), .Y(_abc_17692_n841) );
  OR2X2 OR2X2_1180 ( .A(_abc_17692_n3845), .B(_abc_17692_n3846), .Y(_abc_17692_n3847) );
  OR2X2 OR2X2_1181 ( .A(_abc_17692_n3850), .B(_abc_17692_n3840), .Y(_abc_17692_n3853) );
  OR2X2 OR2X2_1182 ( .A(_abc_17692_n3855_1), .B(_abc_17692_n3839), .Y(_abc_17692_n3856) );
  OR2X2 OR2X2_1183 ( .A(_abc_17692_n3856), .B(_abc_17692_n3820), .Y(_abc_17692_n3857) );
  OR2X2 OR2X2_1184 ( .A(_abc_17692_n3857), .B(_abc_17692_n3806), .Y(_abc_17692_n3858) );
  OR2X2 OR2X2_1185 ( .A(_abc_17692_n3860), .B(_abc_17692_n3861), .Y(_abc_17692_n3862) );
  OR2X2 OR2X2_1186 ( .A(_abc_17692_n3859), .B(_abc_17692_n3862), .Y(_abc_17692_n3863) );
  OR2X2 OR2X2_1187 ( .A(_abc_17692_n3791), .B(_abc_17692_n3863), .Y(workunit2_10__FF_INPUT) );
  OR2X2 OR2X2_1188 ( .A(_abc_17692_n3623), .B(_abc_17692_n3630_1), .Y(_abc_17692_n3866_1) );
  OR2X2 OR2X2_1189 ( .A(_abc_17692_n3868), .B(_abc_17692_n3869), .Y(_abc_17692_n3870) );
  OR2X2 OR2X2_119 ( .A(_abc_17692_n727_bF_buf1), .B(workunit1_6_), .Y(_abc_17692_n842) );
  OR2X2 OR2X2_1190 ( .A(_abc_17692_n2063), .B(workunit1_16_bF_buf0), .Y(_abc_17692_n3872) );
  OR2X2 OR2X2_1191 ( .A(_abc_17692_n3867), .B(workunit1_7_), .Y(_abc_17692_n3873) );
  OR2X2 OR2X2_1192 ( .A(_abc_17692_n3871), .B(_abc_17692_n3875), .Y(_abc_17692_n3876) );
  OR2X2 OR2X2_1193 ( .A(_abc_17692_n3866_1), .B(_abc_17692_n3876), .Y(_abc_17692_n3877_1) );
  OR2X2 OR2X2_1194 ( .A(_abc_17692_n3629), .B(_abc_17692_n3632), .Y(_abc_17692_n3878) );
  OR2X2 OR2X2_1195 ( .A(_abc_17692_n3874), .B(_abc_17692_n2823), .Y(_abc_17692_n3880) );
  OR2X2 OR2X2_1196 ( .A(_abc_17692_n3870), .B(workunit1_11_bF_buf2), .Y(_abc_17692_n3881) );
  OR2X2 OR2X2_1197 ( .A(_abc_17692_n3879), .B(_abc_17692_n3882), .Y(_abc_17692_n3883) );
  OR2X2 OR2X2_1198 ( .A(_abc_17692_n3646), .B(_abc_17692_n3642), .Y(_abc_17692_n3885) );
  OR2X2 OR2X2_1199 ( .A(sum_11_), .B(\key_in[75] ), .Y(_abc_17692_n3889) );
  OR2X2 OR2X2_12 ( .A(state_8_bF_buf9), .B(delta_12_), .Y(delta_12__FF_INPUT) );
  OR2X2 OR2X2_120 ( .A(_abc_17692_n725_bF_buf7), .B(_auto_iopadmap_cc_313_execute_30032_7_), .Y(_abc_17692_n844) );
  OR2X2 OR2X2_1200 ( .A(_abc_17692_n3896), .B(_abc_17692_n3884), .Y(_abc_17692_n3897) );
  OR2X2 OR2X2_1201 ( .A(_abc_17692_n3898), .B(_abc_17692_n3899), .Y(_abc_17692_n3900) );
  OR2X2 OR2X2_1202 ( .A(_abc_17692_n3891), .B(_abc_17692_n3894), .Y(_abc_17692_n3901) );
  OR2X2 OR2X2_1203 ( .A(_abc_17692_n3901), .B(_abc_17692_n3900), .Y(_abc_17692_n3902) );
  OR2X2 OR2X2_1204 ( .A(_abc_17692_n3901), .B(_abc_17692_n3884), .Y(_abc_17692_n3906) );
  OR2X2 OR2X2_1205 ( .A(_abc_17692_n3896), .B(_abc_17692_n3900), .Y(_abc_17692_n3907) );
  OR2X2 OR2X2_1206 ( .A(_abc_17692_n3904), .B(_abc_17692_n3909), .Y(_abc_17692_n3910) );
  OR2X2 OR2X2_1207 ( .A(_abc_17692_n3865), .B(_abc_17692_n3911), .Y(_abc_17692_n3912_1) );
  OR2X2 OR2X2_1208 ( .A(_abc_17692_n3913), .B(_abc_17692_n3910), .Y(_abc_17692_n3914) );
  OR2X2 OR2X2_1209 ( .A(_abc_17692_n3694), .B(_abc_17692_n3751), .Y(_abc_17692_n3917) );
  OR2X2 OR2X2_121 ( .A(_abc_17692_n727_bF_buf0), .B(workunit1_7_), .Y(_abc_17692_n845) );
  OR2X2 OR2X2_1210 ( .A(sum_11_), .B(\key_in[43] ), .Y(_abc_17692_n3924) );
  OR2X2 OR2X2_1211 ( .A(_abc_17692_n3684), .B(_abc_17692_n3680), .Y(_abc_17692_n3927) );
  OR2X2 OR2X2_1212 ( .A(_abc_17692_n3926), .B(_abc_17692_n3929), .Y(_abc_17692_n3930_1) );
  OR2X2 OR2X2_1213 ( .A(_abc_17692_n3884), .B(_abc_17692_n3930_1), .Y(_abc_17692_n3931) );
  OR2X2 OR2X2_1214 ( .A(_abc_17692_n3927), .B(_abc_17692_n3928), .Y(_abc_17692_n3932) );
  OR2X2 OR2X2_1215 ( .A(_abc_17692_n3900), .B(_abc_17692_n3934), .Y(_abc_17692_n3935) );
  OR2X2 OR2X2_1216 ( .A(_abc_17692_n3884), .B(_abc_17692_n3934), .Y(_abc_17692_n3938) );
  OR2X2 OR2X2_1217 ( .A(_abc_17692_n3900), .B(_abc_17692_n3930_1), .Y(_abc_17692_n3939) );
  OR2X2 OR2X2_1218 ( .A(_abc_17692_n3937), .B(_abc_17692_n3941), .Y(_abc_17692_n3942) );
  OR2X2 OR2X2_1219 ( .A(_abc_17692_n3919), .B(_abc_17692_n3943), .Y(_abc_17692_n3944) );
  OR2X2 OR2X2_122 ( .A(_abc_17692_n725_bF_buf6), .B(_auto_iopadmap_cc_313_execute_30032_8_), .Y(_abc_17692_n847) );
  OR2X2 OR2X2_1220 ( .A(_abc_17692_n3918), .B(_abc_17692_n3942), .Y(_abc_17692_n3945) );
  OR2X2 OR2X2_1221 ( .A(_abc_17692_n3722), .B(_abc_17692_n3718), .Y(_abc_17692_n3950) );
  OR2X2 OR2X2_1222 ( .A(sum_11_), .B(\key_in[11] ), .Y(_abc_17692_n3954_1) );
  OR2X2 OR2X2_1223 ( .A(_abc_17692_n3956), .B(_abc_17692_n3958), .Y(_abc_17692_n3959) );
  OR2X2 OR2X2_1224 ( .A(_abc_17692_n3959), .B(_abc_17692_n3884), .Y(_abc_17692_n3960) );
  OR2X2 OR2X2_1225 ( .A(_abc_17692_n3961), .B(_abc_17692_n3900), .Y(_abc_17692_n3962) );
  OR2X2 OR2X2_1226 ( .A(_abc_17692_n3961), .B(_abc_17692_n3884), .Y(_abc_17692_n3965) );
  OR2X2 OR2X2_1227 ( .A(_abc_17692_n3959), .B(_abc_17692_n3900), .Y(_abc_17692_n3966) );
  OR2X2 OR2X2_1228 ( .A(_abc_17692_n3964), .B(_abc_17692_n3968), .Y(_abc_17692_n3969) );
  OR2X2 OR2X2_1229 ( .A(_abc_17692_n3949), .B(_abc_17692_n3970), .Y(_abc_17692_n3971) );
  OR2X2 OR2X2_123 ( .A(_abc_17692_n727_bF_buf7), .B(workunit1_8_bF_buf3), .Y(_abc_17692_n848) );
  OR2X2 OR2X2_1230 ( .A(_abc_17692_n3948), .B(_abc_17692_n3969), .Y(_abc_17692_n3972) );
  OR2X2 OR2X2_1231 ( .A(_abc_17692_n3974), .B(_abc_17692_n3947), .Y(_abc_17692_n3975) );
  OR2X2 OR2X2_1232 ( .A(_abc_17692_n3916), .B(_abc_17692_n3975), .Y(_abc_17692_n3976) );
  OR2X2 OR2X2_1233 ( .A(_abc_17692_n3763), .B(_abc_17692_n3759), .Y(_abc_17692_n3980) );
  OR2X2 OR2X2_1234 ( .A(sum_11_), .B(\key_in[107] ), .Y(_abc_17692_n3984) );
  OR2X2 OR2X2_1235 ( .A(_abc_17692_n3986), .B(_abc_17692_n3988), .Y(_abc_17692_n3989) );
  OR2X2 OR2X2_1236 ( .A(_abc_17692_n3989), .B(_abc_17692_n3884), .Y(_abc_17692_n3990) );
  OR2X2 OR2X2_1237 ( .A(_abc_17692_n3980), .B(_abc_17692_n3987), .Y(_abc_17692_n3991) );
  OR2X2 OR2X2_1238 ( .A(_abc_17692_n3993), .B(_abc_17692_n3900), .Y(_abc_17692_n3994) );
  OR2X2 OR2X2_1239 ( .A(_abc_17692_n3993), .B(_abc_17692_n3884), .Y(_abc_17692_n3997) );
  OR2X2 OR2X2_124 ( .A(_abc_17692_n725_bF_buf5), .B(_auto_iopadmap_cc_313_execute_30032_9_), .Y(_abc_17692_n850_1) );
  OR2X2 OR2X2_1240 ( .A(_abc_17692_n3989), .B(_abc_17692_n3900), .Y(_abc_17692_n3998) );
  OR2X2 OR2X2_1241 ( .A(_abc_17692_n3996), .B(_abc_17692_n4000), .Y(_abc_17692_n4001) );
  OR2X2 OR2X2_1242 ( .A(_abc_17692_n4005), .B(_abc_17692_n4003), .Y(_abc_17692_n4006) );
  OR2X2 OR2X2_1243 ( .A(_abc_17692_n3976), .B(_abc_17692_n4007), .Y(_abc_17692_n4008) );
  OR2X2 OR2X2_1244 ( .A(_abc_17692_n4012), .B(_abc_17692_n4013), .Y(_abc_17692_n4014) );
  OR2X2 OR2X2_1245 ( .A(_abc_17692_n4020), .B(_abc_17692_n3911), .Y(_abc_17692_n4021) );
  OR2X2 OR2X2_1246 ( .A(_abc_17692_n4019), .B(_abc_17692_n3910), .Y(_abc_17692_n4022) );
  OR2X2 OR2X2_1247 ( .A(_abc_17692_n4026), .B(_abc_17692_n3942), .Y(_abc_17692_n4027) );
  OR2X2 OR2X2_1248 ( .A(_abc_17692_n4025), .B(_abc_17692_n3943), .Y(_abc_17692_n4028) );
  OR2X2 OR2X2_1249 ( .A(_abc_17692_n3730), .B(_abc_17692_n3751), .Y(_abc_17692_n4031) );
  OR2X2 OR2X2_125 ( .A(_abc_17692_n727_bF_buf6), .B(workunit1_9_), .Y(_abc_17692_n851_1) );
  OR2X2 OR2X2_1250 ( .A(_abc_17692_n4033), .B(_abc_17692_n3969), .Y(_abc_17692_n4034) );
  OR2X2 OR2X2_1251 ( .A(_abc_17692_n4032), .B(_abc_17692_n3970), .Y(_abc_17692_n4035) );
  OR2X2 OR2X2_1252 ( .A(_abc_17692_n4037), .B(_abc_17692_n4030), .Y(_abc_17692_n4038) );
  OR2X2 OR2X2_1253 ( .A(_abc_17692_n4038), .B(_abc_17692_n4024), .Y(_abc_17692_n4039) );
  OR2X2 OR2X2_1254 ( .A(_abc_17692_n4039), .B(_abc_17692_n4015), .Y(_abc_17692_n4040) );
  OR2X2 OR2X2_1255 ( .A(_abc_17692_n4042), .B(_abc_17692_n4043), .Y(_abc_17692_n4044) );
  OR2X2 OR2X2_1256 ( .A(_abc_17692_n4041), .B(_abc_17692_n4044), .Y(_abc_17692_n4045) );
  OR2X2 OR2X2_1257 ( .A(_abc_17692_n4009), .B(_abc_17692_n4045), .Y(workunit2_11__FF_INPUT) );
  OR2X2 OR2X2_1258 ( .A(_abc_17692_n4050), .B(_abc_17692_n3875), .Y(_abc_17692_n4051) );
  OR2X2 OR2X2_1259 ( .A(_abc_17692_n4049), .B(_abc_17692_n4052), .Y(_abc_17692_n4053) );
  OR2X2 OR2X2_126 ( .A(_abc_17692_n725_bF_buf4), .B(_auto_iopadmap_cc_313_execute_30032_10_), .Y(_abc_17692_n853) );
  OR2X2 OR2X2_1260 ( .A(_abc_17692_n3632), .B(_abc_17692_n3876), .Y(_abc_17692_n4054) );
  OR2X2 OR2X2_1261 ( .A(_abc_17692_n3606), .B(_abc_17692_n4054), .Y(_abc_17692_n4055) );
  OR2X2 OR2X2_1262 ( .A(_abc_17692_n4057), .B(_abc_17692_n4053), .Y(_abc_17692_n4058) );
  OR2X2 OR2X2_1263 ( .A(_abc_17692_n4060), .B(_abc_17692_n4061), .Y(_abc_17692_n4062) );
  OR2X2 OR2X2_1264 ( .A(_abc_17692_n4062), .B(workunit1_12_bF_buf2), .Y(_abc_17692_n4065) );
  OR2X2 OR2X2_1265 ( .A(_abc_17692_n4054), .B(_abc_17692_n3628), .Y(_abc_17692_n4068) );
  OR2X2 OR2X2_1266 ( .A(_abc_17692_n3226), .B(_abc_17692_n4055), .Y(_abc_17692_n4070) );
  OR2X2 OR2X2_1267 ( .A(_abc_17692_n4073_1), .B(_abc_17692_n4067_1), .Y(_abc_17692_n4074) );
  OR2X2 OR2X2_1268 ( .A(_abc_17692_n4077), .B(_abc_17692_n3982), .Y(_abc_17692_n4078) );
  OR2X2 OR2X2_1269 ( .A(_abc_17692_n4076), .B(_abc_17692_n4078), .Y(_abc_17692_n4079) );
  OR2X2 OR2X2_127 ( .A(_abc_17692_n727_bF_buf5), .B(workunit1_10_), .Y(_abc_17692_n854) );
  OR2X2 OR2X2_1270 ( .A(_abc_17692_n4081), .B(_abc_17692_n4079), .Y(_abc_17692_n4082) );
  OR2X2 OR2X2_1271 ( .A(sum_12_), .B(\key_in[108] ), .Y(_abc_17692_n4085) );
  OR2X2 OR2X2_1272 ( .A(_abc_17692_n4092), .B(_abc_17692_n4087), .Y(_abc_17692_n4093) );
  OR2X2 OR2X2_1273 ( .A(_abc_17692_n4094), .B(_abc_17692_n4074), .Y(_abc_17692_n4095) );
  OR2X2 OR2X2_1274 ( .A(_abc_17692_n4093), .B(_abc_17692_n4096_1), .Y(_abc_17692_n4097) );
  OR2X2 OR2X2_1275 ( .A(_abc_17692_n4098), .B(workunit2_12_bF_buf1), .Y(_abc_17692_n4101) );
  OR2X2 OR2X2_1276 ( .A(_abc_17692_n4105), .B(_abc_17692_n4103), .Y(_abc_17692_n4106) );
  OR2X2 OR2X2_1277 ( .A(_abc_17692_n4106), .B(_abc_17692_n3346_1), .Y(_abc_17692_n4107_1) );
  OR2X2 OR2X2_1278 ( .A(_abc_17692_n4109), .B(_abc_17692_n4000), .Y(_abc_17692_n4110) );
  OR2X2 OR2X2_1279 ( .A(_abc_17692_n4105), .B(_abc_17692_n3780), .Y(_abc_17692_n4111) );
  OR2X2 OR2X2_128 ( .A(_abc_17692_n725_bF_buf3), .B(_auto_iopadmap_cc_313_execute_30032_11_), .Y(_abc_17692_n856) );
  OR2X2 OR2X2_1280 ( .A(_abc_17692_n4114), .B(_abc_17692_n4102), .Y(_abc_17692_n4117) );
  OR2X2 OR2X2_1281 ( .A(_abc_17692_n4118), .B(_abc_17692_n4047_bF_buf4), .Y(_abc_17692_n4119) );
  OR2X2 OR2X2_1282 ( .A(_abc_17692_n4123), .B(_abc_17692_n3887), .Y(_abc_17692_n4124) );
  OR2X2 OR2X2_1283 ( .A(_abc_17692_n4122), .B(_abc_17692_n4124), .Y(_abc_17692_n4125) );
  OR2X2 OR2X2_1284 ( .A(_abc_17692_n4127), .B(_abc_17692_n4125), .Y(_abc_17692_n4128) );
  OR2X2 OR2X2_1285 ( .A(sum_12_), .B(\key_in[76] ), .Y(_abc_17692_n4131) );
  OR2X2 OR2X2_1286 ( .A(_abc_17692_n4136), .B(_abc_17692_n4133), .Y(_abc_17692_n4137) );
  OR2X2 OR2X2_1287 ( .A(_abc_17692_n4138), .B(_abc_17692_n4074), .Y(_abc_17692_n4139) );
  OR2X2 OR2X2_1288 ( .A(_abc_17692_n4096_1), .B(_abc_17692_n4137), .Y(_abc_17692_n4140_1) );
  OR2X2 OR2X2_1289 ( .A(_abc_17692_n4143_1), .B(_abc_17692_n4144), .Y(_abc_17692_n4145) );
  OR2X2 OR2X2_129 ( .A(_abc_17692_n727_bF_buf4), .B(workunit1_11_bF_buf3), .Y(_abc_17692_n857) );
  OR2X2 OR2X2_1290 ( .A(_abc_17692_n4152_1), .B(_abc_17692_n4151), .Y(_abc_17692_n4153) );
  OR2X2 OR2X2_1291 ( .A(_abc_17692_n4153), .B(_abc_17692_n4150), .Y(_abc_17692_n4154) );
  OR2X2 OR2X2_1292 ( .A(_abc_17692_n4149), .B(_abc_17692_n4154), .Y(_abc_17692_n4155) );
  OR2X2 OR2X2_1293 ( .A(_abc_17692_n4155), .B(_abc_17692_n4146), .Y(_abc_17692_n4156) );
  OR2X2 OR2X2_1294 ( .A(_abc_17692_n4163), .B(_abc_17692_n3952), .Y(_abc_17692_n4164) );
  OR2X2 OR2X2_1295 ( .A(_abc_17692_n4162), .B(_abc_17692_n4164), .Y(_abc_17692_n4165) );
  OR2X2 OR2X2_1296 ( .A(_abc_17692_n4167), .B(_abc_17692_n4165), .Y(_abc_17692_n4168) );
  OR2X2 OR2X2_1297 ( .A(sum_12_), .B(\key_in[12] ), .Y(_abc_17692_n4171) );
  OR2X2 OR2X2_1298 ( .A(_abc_17692_n4176), .B(_abc_17692_n4173), .Y(_abc_17692_n4177) );
  OR2X2 OR2X2_1299 ( .A(_abc_17692_n4178), .B(_abc_17692_n4074), .Y(_abc_17692_n4179) );
  OR2X2 OR2X2_13 ( .A(state_8_bF_buf8), .B(delta_13_), .Y(delta_13__FF_INPUT) );
  OR2X2 OR2X2_130 ( .A(_abc_17692_n725_bF_buf2), .B(_auto_iopadmap_cc_313_execute_30032_12_), .Y(_abc_17692_n859) );
  OR2X2 OR2X2_1300 ( .A(_abc_17692_n4096_1), .B(_abc_17692_n4177), .Y(_abc_17692_n4180) );
  OR2X2 OR2X2_1301 ( .A(_abc_17692_n4181), .B(workunit2_12_bF_buf1), .Y(_abc_17692_n4184) );
  OR2X2 OR2X2_1302 ( .A(_abc_17692_n4186_1), .B(_abc_17692_n3062), .Y(_abc_17692_n4187) );
  OR2X2 OR2X2_1303 ( .A(_abc_17692_n3969), .B(_abc_17692_n3840), .Y(_abc_17692_n4188) );
  OR2X2 OR2X2_1304 ( .A(_abc_17692_n4188), .B(_abc_17692_n3735), .Y(_abc_17692_n4189) );
  OR2X2 OR2X2_1305 ( .A(_abc_17692_n4187), .B(_abc_17692_n4189), .Y(_abc_17692_n4190) );
  OR2X2 OR2X2_1306 ( .A(_abc_17692_n3968), .B(_abc_17692_n3733_1), .Y(_abc_17692_n4192) );
  OR2X2 OR2X2_1307 ( .A(_abc_17692_n4188), .B(_abc_17692_n3741), .Y(_abc_17692_n4194) );
  OR2X2 OR2X2_1308 ( .A(_abc_17692_n4197), .B(_abc_17692_n4185), .Y(_abc_17692_n4198) );
  OR2X2 OR2X2_1309 ( .A(_abc_17692_n4205), .B(_abc_17692_n3922), .Y(_abc_17692_n4206) );
  OR2X2 OR2X2_131 ( .A(_abc_17692_n727_bF_buf3), .B(workunit1_12_bF_buf3), .Y(_abc_17692_n860) );
  OR2X2 OR2X2_1310 ( .A(_abc_17692_n4204), .B(_abc_17692_n4206), .Y(_abc_17692_n4207) );
  OR2X2 OR2X2_1311 ( .A(_abc_17692_n4209), .B(_abc_17692_n4207), .Y(_abc_17692_n4210) );
  OR2X2 OR2X2_1312 ( .A(sum_12_), .B(\key_in[44] ), .Y(_abc_17692_n4213) );
  OR2X2 OR2X2_1313 ( .A(_abc_17692_n4220), .B(_abc_17692_n4215), .Y(_abc_17692_n4221) );
  OR2X2 OR2X2_1314 ( .A(_abc_17692_n4222), .B(_abc_17692_n4074), .Y(_abc_17692_n4223) );
  OR2X2 OR2X2_1315 ( .A(_abc_17692_n4096_1), .B(_abc_17692_n4221), .Y(_abc_17692_n4224) );
  OR2X2 OR2X2_1316 ( .A(_abc_17692_n4225), .B(workunit2_12_bF_buf3), .Y(_abc_17692_n4228) );
  OR2X2 OR2X2_1317 ( .A(_abc_17692_n3942), .B(_abc_17692_n3698), .Y(_abc_17692_n4230) );
  OR2X2 OR2X2_1318 ( .A(_abc_17692_n3941), .B(_abc_17692_n3917), .Y(_abc_17692_n4232) );
  OR2X2 OR2X2_1319 ( .A(_abc_17692_n4236), .B(_abc_17692_n4234), .Y(_abc_17692_n4237) );
  OR2X2 OR2X2_132 ( .A(_abc_17692_n725_bF_buf1), .B(_auto_iopadmap_cc_313_execute_30032_13_), .Y(_abc_17692_n862) );
  OR2X2 OR2X2_1320 ( .A(_abc_17692_n4238), .B(_abc_17692_n4229), .Y(_abc_17692_n4239) );
  OR2X2 OR2X2_1321 ( .A(_abc_17692_n4243), .B(_abc_17692_n1863_bF_buf8), .Y(_abc_17692_n4244) );
  OR2X2 OR2X2_1322 ( .A(_abc_17692_n4244), .B(_abc_17692_n4202_1), .Y(_abc_17692_n4245) );
  OR2X2 OR2X2_1323 ( .A(_abc_17692_n4245), .B(_abc_17692_n4160), .Y(_abc_17692_n4246) );
  OR2X2 OR2X2_1324 ( .A(_abc_17692_n4256), .B(_abc_17692_n4254), .Y(_abc_17692_n4257) );
  OR2X2 OR2X2_1325 ( .A(_abc_17692_n4257), .B(_abc_17692_n4253_1), .Y(_abc_17692_n4258_1) );
  OR2X2 OR2X2_1326 ( .A(_abc_17692_n4258_1), .B(_abc_17692_n4252), .Y(_abc_17692_n4259) );
  OR2X2 OR2X2_1327 ( .A(_abc_17692_n4259), .B(_abc_17692_n4249), .Y(_abc_17692_n4260) );
  OR2X2 OR2X2_1328 ( .A(_abc_17692_n3910), .B(_abc_17692_n3659), .Y(_abc_17692_n4266) );
  OR2X2 OR2X2_1329 ( .A(_abc_17692_n4266), .B(_abc_17692_n3808), .Y(_abc_17692_n4267) );
  OR2X2 OR2X2_133 ( .A(_abc_17692_n727_bF_buf2), .B(workunit1_13_bF_buf3), .Y(_abc_17692_n863) );
  OR2X2 OR2X2_1330 ( .A(_abc_17692_n4265), .B(_abc_17692_n4267), .Y(_abc_17692_n4268) );
  OR2X2 OR2X2_1331 ( .A(_abc_17692_n3909), .B(_abc_17692_n4018), .Y(_abc_17692_n4270) );
  OR2X2 OR2X2_1332 ( .A(_abc_17692_n4266), .B(_abc_17692_n3813), .Y(_abc_17692_n4272) );
  OR2X2 OR2X2_1333 ( .A(_abc_17692_n4275), .B(_abc_17692_n4145), .Y(_abc_17692_n4276) );
  OR2X2 OR2X2_1334 ( .A(_abc_17692_n4287), .B(_abc_17692_n4286), .Y(_abc_17692_n4288) );
  OR2X2 OR2X2_1335 ( .A(_abc_17692_n4288), .B(_abc_17692_n4285), .Y(_abc_17692_n4289_1) );
  OR2X2 OR2X2_1336 ( .A(_abc_17692_n4289_1), .B(_abc_17692_n4284), .Y(_abc_17692_n4290) );
  OR2X2 OR2X2_1337 ( .A(_abc_17692_n4290), .B(_abc_17692_n4281), .Y(_abc_17692_n4291) );
  OR2X2 OR2X2_1338 ( .A(_abc_17692_n4303), .B(_abc_17692_n4301), .Y(_abc_17692_n4304) );
  OR2X2 OR2X2_1339 ( .A(_abc_17692_n4304), .B(_abc_17692_n4300), .Y(_abc_17692_n4305) );
  OR2X2 OR2X2_134 ( .A(_abc_17692_n725_bF_buf0), .B(_auto_iopadmap_cc_313_execute_30032_14_), .Y(_abc_17692_n865) );
  OR2X2 OR2X2_1340 ( .A(_abc_17692_n4305), .B(_abc_17692_n4299), .Y(_abc_17692_n4306) );
  OR2X2 OR2X2_1341 ( .A(_abc_17692_n4306), .B(_abc_17692_n4296), .Y(_abc_17692_n4309) );
  OR2X2 OR2X2_1342 ( .A(_abc_17692_n4311), .B(_abc_17692_n4295), .Y(_abc_17692_n4312) );
  OR2X2 OR2X2_1343 ( .A(_abc_17692_n4280), .B(_abc_17692_n4312), .Y(_abc_17692_n4313) );
  OR2X2 OR2X2_1344 ( .A(_abc_17692_n4313), .B(_abc_17692_n4264), .Y(_abc_17692_n4314) );
  OR2X2 OR2X2_1345 ( .A(_abc_17692_n4316), .B(_abc_17692_n4317_1), .Y(_abc_17692_n4318) );
  OR2X2 OR2X2_1346 ( .A(_abc_17692_n4315), .B(_abc_17692_n4318), .Y(_abc_17692_n4319) );
  OR2X2 OR2X2_1347 ( .A(_abc_17692_n4319), .B(_abc_17692_n4248), .Y(workunit2_12__FF_INPUT) );
  OR2X2 OR2X2_1348 ( .A(_abc_17692_n4067_1), .B(_abc_17692_n4063), .Y(_abc_17692_n4321) );
  OR2X2 OR2X2_1349 ( .A(_abc_17692_n4323), .B(_abc_17692_n4324), .Y(_abc_17692_n4325) );
  OR2X2 OR2X2_135 ( .A(_abc_17692_n727_bF_buf1), .B(workunit1_14_bF_buf3), .Y(_abc_17692_n866) );
  OR2X2 OR2X2_1350 ( .A(_abc_17692_n4325), .B(workunit1_13_bF_buf2), .Y(_abc_17692_n4327) );
  OR2X2 OR2X2_1351 ( .A(_abc_17692_n4328), .B(_abc_17692_n4326), .Y(_abc_17692_n4329) );
  OR2X2 OR2X2_1352 ( .A(_abc_17692_n4321), .B(_abc_17692_n4329), .Y(_abc_17692_n4332) );
  OR2X2 OR2X2_1353 ( .A(_abc_17692_n4133), .B(_abc_17692_n4129), .Y(_abc_17692_n4335) );
  OR2X2 OR2X2_1354 ( .A(sum_13_), .B(\key_in[77] ), .Y(_abc_17692_n4339) );
  OR2X2 OR2X2_1355 ( .A(_abc_17692_n4341), .B(_abc_17692_n4343), .Y(_abc_17692_n4344_1) );
  OR2X2 OR2X2_1356 ( .A(_abc_17692_n4347_1), .B(_abc_17692_n4345), .Y(_abc_17692_n4348) );
  OR2X2 OR2X2_1357 ( .A(_abc_17692_n4350), .B(_abc_17692_n4352), .Y(_abc_17692_n4353) );
  OR2X2 OR2X2_1358 ( .A(_abc_17692_n4356), .B(_abc_17692_n4354), .Y(_abc_17692_n4357) );
  OR2X2 OR2X2_1359 ( .A(_abc_17692_n4358), .B(_abc_17692_n4353), .Y(_abc_17692_n4359) );
  OR2X2 OR2X2_136 ( .A(_abc_17692_n725_bF_buf7), .B(_auto_iopadmap_cc_313_execute_30032_15_), .Y(_abc_17692_n868) );
  OR2X2 OR2X2_1360 ( .A(_abc_17692_n4215), .B(_abc_17692_n4211), .Y(_abc_17692_n4362) );
  OR2X2 OR2X2_1361 ( .A(sum_13_), .B(\key_in[45] ), .Y(_abc_17692_n4366) );
  OR2X2 OR2X2_1362 ( .A(_abc_17692_n4363), .B(_abc_17692_n4367), .Y(_abc_17692_n4369) );
  OR2X2 OR2X2_1363 ( .A(_abc_17692_n4370), .B(_abc_17692_n4368), .Y(_abc_17692_n4371) );
  OR2X2 OR2X2_1364 ( .A(_abc_17692_n4371), .B(_abc_17692_n4333), .Y(_abc_17692_n4372) );
  OR2X2 OR2X2_1365 ( .A(_abc_17692_n4334), .B(_abc_17692_n4374), .Y(_abc_17692_n4375) );
  OR2X2 OR2X2_1366 ( .A(_abc_17692_n4376), .B(_abc_17692_n4351), .Y(_abc_17692_n4377) );
  OR2X2 OR2X2_1367 ( .A(_abc_17692_n4374), .B(_abc_17692_n4333), .Y(_abc_17692_n4378) );
  OR2X2 OR2X2_1368 ( .A(_abc_17692_n4371), .B(_abc_17692_n4334), .Y(_abc_17692_n4379) );
  OR2X2 OR2X2_1369 ( .A(_abc_17692_n4380), .B(workunit2_13_), .Y(_abc_17692_n4381) );
  OR2X2 OR2X2_137 ( .A(_abc_17692_n727_bF_buf0), .B(workunit1_15_), .Y(_abc_17692_n869) );
  OR2X2 OR2X2_1370 ( .A(_abc_17692_n4385), .B(_abc_17692_n4383), .Y(_abc_17692_n4386) );
  OR2X2 OR2X2_1371 ( .A(_abc_17692_n4384), .B(_abc_17692_n4382), .Y(_abc_17692_n4387) );
  OR2X2 OR2X2_1372 ( .A(_abc_17692_n4173), .B(_abc_17692_n4169_1), .Y(_abc_17692_n4390) );
  OR2X2 OR2X2_1373 ( .A(sum_13_), .B(\key_in[13] ), .Y(_abc_17692_n4393) );
  OR2X2 OR2X2_1374 ( .A(_abc_17692_n4390), .B(_abc_17692_n4395), .Y(_abc_17692_n4396) );
  OR2X2 OR2X2_1375 ( .A(_abc_17692_n4333), .B(_abc_17692_n4399), .Y(_abc_17692_n4400) );
  OR2X2 OR2X2_1376 ( .A(_abc_17692_n4334), .B(_abc_17692_n4401), .Y(_abc_17692_n4402) );
  OR2X2 OR2X2_1377 ( .A(_abc_17692_n4404), .B(_abc_17692_n4351), .Y(_abc_17692_n4405) );
  OR2X2 OR2X2_1378 ( .A(_abc_17692_n4403), .B(workunit2_13_), .Y(_abc_17692_n4406) );
  OR2X2 OR2X2_1379 ( .A(_abc_17692_n4410), .B(_abc_17692_n4408), .Y(_abc_17692_n4411) );
  OR2X2 OR2X2_138 ( .A(_abc_17692_n725_bF_buf6), .B(_auto_iopadmap_cc_313_execute_30032_16_), .Y(_abc_17692_n871) );
  OR2X2 OR2X2_1380 ( .A(_abc_17692_n4409), .B(_abc_17692_n4407), .Y(_abc_17692_n4412) );
  OR2X2 OR2X2_1381 ( .A(_abc_17692_n4414), .B(_abc_17692_n4389_1), .Y(_abc_17692_n4415) );
  OR2X2 OR2X2_1382 ( .A(_abc_17692_n4415), .B(_abc_17692_n4361), .Y(_abc_17692_n4416) );
  OR2X2 OR2X2_1383 ( .A(_abc_17692_n4087), .B(_abc_17692_n4083), .Y(_abc_17692_n4417) );
  OR2X2 OR2X2_1384 ( .A(sum_13_), .B(\key_in[109] ), .Y(_abc_17692_n4420) );
  OR2X2 OR2X2_1385 ( .A(_abc_17692_n4417), .B(_abc_17692_n4422), .Y(_abc_17692_n4423) );
  OR2X2 OR2X2_1386 ( .A(_abc_17692_n4426), .B(_abc_17692_n4333), .Y(_abc_17692_n4427) );
  OR2X2 OR2X2_1387 ( .A(_abc_17692_n4428), .B(_abc_17692_n4334), .Y(_abc_17692_n4429) );
  OR2X2 OR2X2_1388 ( .A(_abc_17692_n4431), .B(_abc_17692_n4351), .Y(_abc_17692_n4432) );
  OR2X2 OR2X2_1389 ( .A(_abc_17692_n4430), .B(workunit2_13_), .Y(_abc_17692_n4433) );
  OR2X2 OR2X2_139 ( .A(_abc_17692_n727_bF_buf7), .B(workunit1_16_bF_buf3), .Y(_abc_17692_n872) );
  OR2X2 OR2X2_1390 ( .A(_abc_17692_n4437), .B(_abc_17692_n4435), .Y(_abc_17692_n4438) );
  OR2X2 OR2X2_1391 ( .A(_abc_17692_n4436), .B(_abc_17692_n4434), .Y(_abc_17692_n4439) );
  OR2X2 OR2X2_1392 ( .A(_abc_17692_n4416), .B(_abc_17692_n4441), .Y(_abc_17692_n4442) );
  OR2X2 OR2X2_1393 ( .A(_abc_17692_n4447_1), .B(_abc_17692_n4435), .Y(_abc_17692_n4448) );
  OR2X2 OR2X2_1394 ( .A(_abc_17692_n4449), .B(_abc_17692_n4434), .Y(_abc_17692_n4450) );
  OR2X2 OR2X2_1395 ( .A(_abc_17692_n4457), .B(_abc_17692_n4458), .Y(_abc_17692_n4459) );
  OR2X2 OR2X2_1396 ( .A(_abc_17692_n4465), .B(_abc_17692_n4382), .Y(_abc_17692_n4466) );
  OR2X2 OR2X2_1397 ( .A(_abc_17692_n4464), .B(_abc_17692_n4383), .Y(_abc_17692_n4467) );
  OR2X2 OR2X2_1398 ( .A(_abc_17692_n4473), .B(_abc_17692_n4408), .Y(_abc_17692_n4474) );
  OR2X2 OR2X2_1399 ( .A(_abc_17692_n4475), .B(_abc_17692_n4407), .Y(_abc_17692_n4476) );
  OR2X2 OR2X2_14 ( .A(state_8_bF_buf7), .B(delta_14_), .Y(delta_14__FF_INPUT) );
  OR2X2 OR2X2_140 ( .A(_abc_17692_n725_bF_buf5), .B(_auto_iopadmap_cc_313_execute_30032_17_), .Y(_abc_17692_n874) );
  OR2X2 OR2X2_1400 ( .A(_abc_17692_n4478), .B(_abc_17692_n4469), .Y(_abc_17692_n4479) );
  OR2X2 OR2X2_1401 ( .A(_abc_17692_n4479), .B(_abc_17692_n4460), .Y(_abc_17692_n4480) );
  OR2X2 OR2X2_1402 ( .A(_abc_17692_n4480), .B(_abc_17692_n4452), .Y(_abc_17692_n4481) );
  OR2X2 OR2X2_1403 ( .A(_abc_17692_n4483), .B(_abc_17692_n4484), .Y(_abc_17692_n4485) );
  OR2X2 OR2X2_1404 ( .A(_abc_17692_n4482), .B(_abc_17692_n4485), .Y(_abc_17692_n4486) );
  OR2X2 OR2X2_1405 ( .A(_abc_17692_n4486), .B(_abc_17692_n4443), .Y(workunit2_13__FF_INPUT) );
  OR2X2 OR2X2_1406 ( .A(_abc_17692_n4063), .B(_abc_17692_n4326), .Y(_abc_17692_n4491) );
  OR2X2 OR2X2_1407 ( .A(_abc_17692_n4490), .B(_abc_17692_n4492), .Y(_abc_17692_n4493) );
  OR2X2 OR2X2_1408 ( .A(_abc_17692_n4495), .B(_abc_17692_n4496), .Y(_abc_17692_n4497) );
  OR2X2 OR2X2_1409 ( .A(_abc_17692_n4497), .B(workunit1_14_bF_buf3), .Y(_abc_17692_n4500) );
  OR2X2 OR2X2_141 ( .A(_abc_17692_n727_bF_buf6), .B(workunit1_17_), .Y(_abc_17692_n875_1) );
  OR2X2 OR2X2_1410 ( .A(_abc_17692_n4072), .B(_abc_17692_n4329), .Y(_abc_17692_n4503) );
  OR2X2 OR2X2_1411 ( .A(_abc_17692_n4071), .B(_abc_17692_n4503), .Y(_abc_17692_n4504) );
  OR2X2 OR2X2_1412 ( .A(_abc_17692_n4507_1), .B(_abc_17692_n4498), .Y(_abc_17692_n4508) );
  OR2X2 OR2X2_1413 ( .A(_abc_17692_n4509), .B(_abc_17692_n4502), .Y(_abc_17692_n4510_1) );
  OR2X2 OR2X2_1414 ( .A(_abc_17692_n4514), .B(_abc_17692_n4513), .Y(_abc_17692_n4515) );
  OR2X2 OR2X2_1415 ( .A(_abc_17692_n4512), .B(_abc_17692_n4516), .Y(_abc_17692_n4517) );
  OR2X2 OR2X2_1416 ( .A(sum_14_), .B(\key_in[110] ), .Y(_abc_17692_n4520) );
  OR2X2 OR2X2_1417 ( .A(_abc_17692_n4526), .B(_abc_17692_n4522), .Y(_abc_17692_n4527) );
  OR2X2 OR2X2_1418 ( .A(_abc_17692_n4528), .B(_abc_17692_n4510_1), .Y(_abc_17692_n4529) );
  OR2X2 OR2X2_1419 ( .A(_abc_17692_n4527), .B(_abc_17692_n4530), .Y(_abc_17692_n4531) );
  OR2X2 OR2X2_142 ( .A(_abc_17692_n725_bF_buf4), .B(_auto_iopadmap_cc_313_execute_30032_18_), .Y(_abc_17692_n877) );
  OR2X2 OR2X2_1420 ( .A(_abc_17692_n4532), .B(workunit2_14_bF_buf2), .Y(_abc_17692_n4533) );
  OR2X2 OR2X2_1421 ( .A(_abc_17692_n4434), .B(_abc_17692_n4100), .Y(_abc_17692_n4539) );
  OR2X2 OR2X2_1422 ( .A(_abc_17692_n4543), .B(_abc_17692_n4541), .Y(_abc_17692_n4544) );
  OR2X2 OR2X2_1423 ( .A(_abc_17692_n4544), .B(_abc_17692_n4536), .Y(_abc_17692_n4545) );
  OR2X2 OR2X2_1424 ( .A(_abc_17692_n4548), .B(_abc_17692_n4047_bF_buf3), .Y(_abc_17692_n4549) );
  OR2X2 OR2X2_1425 ( .A(_abc_17692_n4553), .B(_abc_17692_n4552), .Y(_abc_17692_n4554) );
  OR2X2 OR2X2_1426 ( .A(_abc_17692_n4551), .B(_abc_17692_n4555), .Y(_abc_17692_n4556) );
  OR2X2 OR2X2_1427 ( .A(sum_14_), .B(\key_in[78] ), .Y(_abc_17692_n4559) );
  OR2X2 OR2X2_1428 ( .A(_abc_17692_n4564), .B(_abc_17692_n4561), .Y(_abc_17692_n4565) );
  OR2X2 OR2X2_1429 ( .A(_abc_17692_n4566), .B(_abc_17692_n4510_1), .Y(_abc_17692_n4567) );
  OR2X2 OR2X2_143 ( .A(_abc_17692_n727_bF_buf5), .B(workunit1_18_), .Y(_abc_17692_n878) );
  OR2X2 OR2X2_1430 ( .A(_abc_17692_n4530), .B(_abc_17692_n4565), .Y(_abc_17692_n4568) );
  OR2X2 OR2X2_1431 ( .A(_abc_17692_n4569), .B(workunit2_14_bF_buf3), .Y(_abc_17692_n4572) );
  OR2X2 OR2X2_1432 ( .A(_abc_17692_n4575), .B(_abc_17692_n4574), .Y(_abc_17692_n4576) );
  OR2X2 OR2X2_1433 ( .A(_abc_17692_n4578), .B(_abc_17692_n4576), .Y(_abc_17692_n4579) );
  OR2X2 OR2X2_1434 ( .A(_abc_17692_n4579), .B(_abc_17692_n4573), .Y(_abc_17692_n4582) );
  OR2X2 OR2X2_1435 ( .A(_abc_17692_n4588), .B(_abc_17692_n4587_1), .Y(_abc_17692_n4589) );
  OR2X2 OR2X2_1436 ( .A(_abc_17692_n4586), .B(_abc_17692_n4590), .Y(_abc_17692_n4591) );
  OR2X2 OR2X2_1437 ( .A(sum_14_), .B(\key_in[14] ), .Y(_abc_17692_n4594) );
  OR2X2 OR2X2_1438 ( .A(_abc_17692_n4599), .B(_abc_17692_n4596), .Y(_abc_17692_n4600) );
  OR2X2 OR2X2_1439 ( .A(_abc_17692_n4601), .B(_abc_17692_n4510_1), .Y(_abc_17692_n4602) );
  OR2X2 OR2X2_144 ( .A(_abc_17692_n725_bF_buf3), .B(_auto_iopadmap_cc_313_execute_30032_19_), .Y(_abc_17692_n880) );
  OR2X2 OR2X2_1440 ( .A(_abc_17692_n4530), .B(_abc_17692_n4600), .Y(_abc_17692_n4603) );
  OR2X2 OR2X2_1441 ( .A(_abc_17692_n4604), .B(workunit2_14_bF_buf2), .Y(_abc_17692_n4605) );
  OR2X2 OR2X2_1442 ( .A(_abc_17692_n4407), .B(_abc_17692_n4183), .Y(_abc_17692_n4611) );
  OR2X2 OR2X2_1443 ( .A(_abc_17692_n4407), .B(_abc_17692_n4296), .Y(_abc_17692_n4614) );
  OR2X2 OR2X2_1444 ( .A(_abc_17692_n4616), .B(_abc_17692_n4613), .Y(_abc_17692_n4617) );
  OR2X2 OR2X2_1445 ( .A(_abc_17692_n4617), .B(_abc_17692_n4608), .Y(_abc_17692_n4620) );
  OR2X2 OR2X2_1446 ( .A(_abc_17692_n4627), .B(_abc_17692_n4626), .Y(_abc_17692_n4628) );
  OR2X2 OR2X2_1447 ( .A(_abc_17692_n4625), .B(_abc_17692_n4629), .Y(_abc_17692_n4630) );
  OR2X2 OR2X2_1448 ( .A(sum_14_), .B(\key_in[46] ), .Y(_abc_17692_n4633) );
  OR2X2 OR2X2_1449 ( .A(_abc_17692_n4639), .B(_abc_17692_n4635), .Y(_abc_17692_n4640) );
  OR2X2 OR2X2_145 ( .A(_abc_17692_n727_bF_buf4), .B(workunit1_19_), .Y(_abc_17692_n881) );
  OR2X2 OR2X2_1450 ( .A(_abc_17692_n4641), .B(_abc_17692_n4643_1), .Y(_abc_17692_n4644) );
  OR2X2 OR2X2_1451 ( .A(_abc_17692_n4645), .B(_abc_17692_n4623), .Y(_abc_17692_n4646_1) );
  OR2X2 OR2X2_1452 ( .A(_abc_17692_n4644), .B(workunit2_14_bF_buf3), .Y(_abc_17692_n4647) );
  OR2X2 OR2X2_1453 ( .A(_abc_17692_n4382), .B(_abc_17692_n4227), .Y(_abc_17692_n4652) );
  OR2X2 OR2X2_1454 ( .A(_abc_17692_n4382), .B(_abc_17692_n4281), .Y(_abc_17692_n4655) );
  OR2X2 OR2X2_1455 ( .A(_abc_17692_n4657), .B(_abc_17692_n4654), .Y(_abc_17692_n4658) );
  OR2X2 OR2X2_1456 ( .A(_abc_17692_n4658), .B(_abc_17692_n4649), .Y(_abc_17692_n4661) );
  OR2X2 OR2X2_1457 ( .A(_abc_17692_n4663), .B(_abc_17692_n1863_bF_buf4), .Y(_abc_17692_n4664) );
  OR2X2 OR2X2_1458 ( .A(_abc_17692_n4664), .B(_abc_17692_n4622), .Y(_abc_17692_n4665) );
  OR2X2 OR2X2_1459 ( .A(_abc_17692_n4665), .B(_abc_17692_n4584_1), .Y(_abc_17692_n4666) );
  OR2X2 OR2X2_146 ( .A(_abc_17692_n725_bF_buf2), .B(_auto_iopadmap_cc_313_execute_30032_20_), .Y(_abc_17692_n883) );
  OR2X2 OR2X2_1460 ( .A(_abc_17692_n4670), .B(_abc_17692_n4671), .Y(_abc_17692_n4672) );
  OR2X2 OR2X2_1461 ( .A(_abc_17692_n4674), .B(_abc_17692_n4672), .Y(_abc_17692_n4675) );
  OR2X2 OR2X2_1462 ( .A(_abc_17692_n4675), .B(_abc_17692_n4669), .Y(_abc_17692_n4678) );
  OR2X2 OR2X2_1463 ( .A(_abc_17692_n4352), .B(_abc_17692_n4454), .Y(_abc_17692_n4683) );
  OR2X2 OR2X2_1464 ( .A(_abc_17692_n4353), .B(_abc_17692_n4146), .Y(_abc_17692_n4686) );
  OR2X2 OR2X2_1465 ( .A(_abc_17692_n4688), .B(_abc_17692_n4685), .Y(_abc_17692_n4689) );
  OR2X2 OR2X2_1466 ( .A(_abc_17692_n4689), .B(_abc_17692_n4681), .Y(_abc_17692_n4692) );
  OR2X2 OR2X2_1467 ( .A(_abc_17692_n4696), .B(_abc_17692_n4695), .Y(_abc_17692_n4697) );
  OR2X2 OR2X2_1468 ( .A(_abc_17692_n4700), .B(_abc_17692_n4698), .Y(_abc_17692_n4701) );
  OR2X2 OR2X2_1469 ( .A(_abc_17692_n4701), .B(_abc_17692_n4648), .Y(_abc_17692_n4704) );
  OR2X2 OR2X2_147 ( .A(_abc_17692_n727_bF_buf3), .B(workunit1_20_), .Y(_abc_17692_n884) );
  OR2X2 OR2X2_1470 ( .A(_abc_17692_n4709), .B(_abc_17692_n4708), .Y(_abc_17692_n4710) );
  OR2X2 OR2X2_1471 ( .A(_abc_17692_n4713), .B(_abc_17692_n4711), .Y(_abc_17692_n4714) );
  OR2X2 OR2X2_1472 ( .A(_abc_17692_n4714), .B(_abc_17692_n4707), .Y(_abc_17692_n4717) );
  OR2X2 OR2X2_1473 ( .A(_abc_17692_n4719), .B(_abc_17692_n4706), .Y(_abc_17692_n4720) );
  OR2X2 OR2X2_1474 ( .A(_abc_17692_n4720), .B(_abc_17692_n4694), .Y(_abc_17692_n4721) );
  OR2X2 OR2X2_1475 ( .A(_abc_17692_n4721), .B(_abc_17692_n4680), .Y(_abc_17692_n4722) );
  OR2X2 OR2X2_1476 ( .A(_abc_17692_n4724), .B(_abc_17692_n4725), .Y(_abc_17692_n4726) );
  OR2X2 OR2X2_1477 ( .A(_abc_17692_n4723), .B(_abc_17692_n4726), .Y(_abc_17692_n4727) );
  OR2X2 OR2X2_1478 ( .A(_abc_17692_n4727), .B(_abc_17692_n4668), .Y(workunit2_14__FF_INPUT) );
  OR2X2 OR2X2_1479 ( .A(_abc_17692_n4502), .B(_abc_17692_n4498), .Y(_abc_17692_n4729) );
  OR2X2 OR2X2_148 ( .A(_abc_17692_n725_bF_buf1), .B(_auto_iopadmap_cc_313_execute_30032_21_), .Y(_abc_17692_n886) );
  OR2X2 OR2X2_1480 ( .A(_abc_17692_n4731), .B(_abc_17692_n4732), .Y(_abc_17692_n4733) );
  OR2X2 OR2X2_1481 ( .A(_abc_17692_n4733), .B(workunit1_15_), .Y(_abc_17692_n4735_1) );
  OR2X2 OR2X2_1482 ( .A(_abc_17692_n4736), .B(_abc_17692_n4734), .Y(_abc_17692_n4737) );
  OR2X2 OR2X2_1483 ( .A(_abc_17692_n4729), .B(_abc_17692_n4737), .Y(_abc_17692_n4738_1) );
  OR2X2 OR2X2_1484 ( .A(_abc_17692_n4506), .B(_abc_17692_n4508), .Y(_abc_17692_n4739) );
  OR2X2 OR2X2_1485 ( .A(_abc_17692_n4740), .B(_abc_17692_n4742), .Y(_abc_17692_n4743) );
  OR2X2 OR2X2_1486 ( .A(_abc_17692_n4561), .B(_abc_17692_n4557), .Y(_abc_17692_n4745) );
  OR2X2 OR2X2_1487 ( .A(sum_15_), .B(\key_in[79] ), .Y(_abc_17692_n4749) );
  OR2X2 OR2X2_1488 ( .A(_abc_17692_n4756), .B(_abc_17692_n4744), .Y(_abc_17692_n4757) );
  OR2X2 OR2X2_1489 ( .A(_abc_17692_n4758), .B(_abc_17692_n4759), .Y(_abc_17692_n4760) );
  OR2X2 OR2X2_149 ( .A(_abc_17692_n727_bF_buf2), .B(workunit1_21_), .Y(_abc_17692_n887) );
  OR2X2 OR2X2_1490 ( .A(_abc_17692_n4751), .B(_abc_17692_n4754), .Y(_abc_17692_n4761) );
  OR2X2 OR2X2_1491 ( .A(_abc_17692_n4761), .B(_abc_17692_n4760), .Y(_abc_17692_n4762) );
  OR2X2 OR2X2_1492 ( .A(_abc_17692_n4761), .B(_abc_17692_n4744), .Y(_abc_17692_n4766) );
  OR2X2 OR2X2_1493 ( .A(_abc_17692_n4756), .B(_abc_17692_n4760), .Y(_abc_17692_n4767) );
  OR2X2 OR2X2_1494 ( .A(_abc_17692_n4764), .B(_abc_17692_n4769), .Y(_abc_17692_n4770) );
  OR2X2 OR2X2_1495 ( .A(_abc_17692_n4772), .B(_abc_17692_n4770), .Y(_abc_17692_n4773) );
  OR2X2 OR2X2_1496 ( .A(_abc_17692_n4771), .B(_abc_17692_n4774), .Y(_abc_17692_n4775) );
  OR2X2 OR2X2_1497 ( .A(_abc_17692_n4596), .B(_abc_17692_n4592), .Y(_abc_17692_n4778) );
  OR2X2 OR2X2_1498 ( .A(sum_15_), .B(\key_in[15] ), .Y(_abc_17692_n4782) );
  OR2X2 OR2X2_1499 ( .A(_abc_17692_n4784), .B(_abc_17692_n4786), .Y(_abc_17692_n4787) );
  OR2X2 OR2X2_15 ( .A(state_8_bF_buf6), .B(delta_16_), .Y(delta_16__FF_INPUT) );
  OR2X2 OR2X2_150 ( .A(_abc_17692_n725_bF_buf0), .B(_auto_iopadmap_cc_313_execute_30032_22_), .Y(_abc_17692_n889_1) );
  OR2X2 OR2X2_1500 ( .A(_abc_17692_n4787), .B(_abc_17692_n4744), .Y(_abc_17692_n4788) );
  OR2X2 OR2X2_1501 ( .A(_abc_17692_n4789_1), .B(_abc_17692_n4760), .Y(_abc_17692_n4790) );
  OR2X2 OR2X2_1502 ( .A(_abc_17692_n4789_1), .B(_abc_17692_n4744), .Y(_abc_17692_n4793) );
  OR2X2 OR2X2_1503 ( .A(_abc_17692_n4787), .B(_abc_17692_n4760), .Y(_abc_17692_n4794) );
  OR2X2 OR2X2_1504 ( .A(_abc_17692_n4792_1), .B(_abc_17692_n4796), .Y(_abc_17692_n4797) );
  OR2X2 OR2X2_1505 ( .A(_abc_17692_n4798), .B(_abc_17692_n4797), .Y(_abc_17692_n4799) );
  OR2X2 OR2X2_1506 ( .A(_abc_17692_n4801), .B(_abc_17692_n4800), .Y(_abc_17692_n4802) );
  OR2X2 OR2X2_1507 ( .A(sum_15_), .B(\key_in[47] ), .Y(_abc_17692_n4809) );
  OR2X2 OR2X2_1508 ( .A(_abc_17692_n4635), .B(_abc_17692_n4631), .Y(_abc_17692_n4812) );
  OR2X2 OR2X2_1509 ( .A(_abc_17692_n4811), .B(_abc_17692_n4814), .Y(_abc_17692_n4815) );
  OR2X2 OR2X2_151 ( .A(_abc_17692_n727_bF_buf1), .B(workunit1_22_), .Y(_abc_17692_n890_1) );
  OR2X2 OR2X2_1510 ( .A(_abc_17692_n4744), .B(_abc_17692_n4815), .Y(_abc_17692_n4816) );
  OR2X2 OR2X2_1511 ( .A(_abc_17692_n4812), .B(_abc_17692_n4813), .Y(_abc_17692_n4817) );
  OR2X2 OR2X2_1512 ( .A(_abc_17692_n4760), .B(_abc_17692_n4819), .Y(_abc_17692_n4820) );
  OR2X2 OR2X2_1513 ( .A(_abc_17692_n4744), .B(_abc_17692_n4819), .Y(_abc_17692_n4823) );
  OR2X2 OR2X2_1514 ( .A(_abc_17692_n4760), .B(_abc_17692_n4815), .Y(_abc_17692_n4824) );
  OR2X2 OR2X2_1515 ( .A(_abc_17692_n4822), .B(_abc_17692_n4826), .Y(_abc_17692_n4827) );
  OR2X2 OR2X2_1516 ( .A(_abc_17692_n4832), .B(_abc_17692_n4828), .Y(_abc_17692_n4833) );
  OR2X2 OR2X2_1517 ( .A(_abc_17692_n4831), .B(_abc_17692_n4827), .Y(_abc_17692_n4834) );
  OR2X2 OR2X2_1518 ( .A(_abc_17692_n4836), .B(_abc_17692_n1863_bF_buf2), .Y(_abc_17692_n4837) );
  OR2X2 OR2X2_1519 ( .A(_abc_17692_n4804), .B(_abc_17692_n4837), .Y(_abc_17692_n4838) );
  OR2X2 OR2X2_152 ( .A(_abc_17692_n725_bF_buf7), .B(_auto_iopadmap_cc_313_execute_30032_23_), .Y(_abc_17692_n892) );
  OR2X2 OR2X2_1520 ( .A(_abc_17692_n4838), .B(_abc_17692_n4777), .Y(_abc_17692_n4839) );
  OR2X2 OR2X2_1521 ( .A(sum_15_), .B(\key_in[111] ), .Y(_abc_17692_n4844) );
  OR2X2 OR2X2_1522 ( .A(_abc_17692_n4522), .B(_abc_17692_n4518), .Y(_abc_17692_n4847) );
  OR2X2 OR2X2_1523 ( .A(_abc_17692_n4846), .B(_abc_17692_n4849), .Y(_abc_17692_n4850) );
  OR2X2 OR2X2_1524 ( .A(_abc_17692_n4850), .B(_abc_17692_n4744), .Y(_abc_17692_n4851) );
  OR2X2 OR2X2_1525 ( .A(_abc_17692_n4847), .B(_abc_17692_n4848), .Y(_abc_17692_n4852) );
  OR2X2 OR2X2_1526 ( .A(_abc_17692_n4854), .B(_abc_17692_n4760), .Y(_abc_17692_n4855) );
  OR2X2 OR2X2_1527 ( .A(_abc_17692_n4854), .B(_abc_17692_n4744), .Y(_abc_17692_n4858) );
  OR2X2 OR2X2_1528 ( .A(_abc_17692_n4850), .B(_abc_17692_n4760), .Y(_abc_17692_n4859) );
  OR2X2 OR2X2_1529 ( .A(_abc_17692_n4857), .B(_abc_17692_n4861), .Y(_abc_17692_n4862) );
  OR2X2 OR2X2_153 ( .A(_abc_17692_n727_bF_buf0), .B(workunit1_23_), .Y(_abc_17692_n893) );
  OR2X2 OR2X2_1530 ( .A(_abc_17692_n4867), .B(_abc_17692_n4047_bF_buf2), .Y(_abc_17692_n4868) );
  OR2X2 OR2X2_1531 ( .A(_abc_17692_n4868), .B(_abc_17692_n4865), .Y(_abc_17692_n4869) );
  OR2X2 OR2X2_1532 ( .A(_abc_17692_n4876), .B(_abc_17692_n4862), .Y(_abc_17692_n4877) );
  OR2X2 OR2X2_1533 ( .A(_abc_17692_n4875), .B(_abc_17692_n4866), .Y(_abc_17692_n4878) );
  OR2X2 OR2X2_1534 ( .A(_abc_17692_n4885), .B(_abc_17692_n4774), .Y(_abc_17692_n4886) );
  OR2X2 OR2X2_1535 ( .A(_abc_17692_n4884), .B(_abc_17692_n4770), .Y(_abc_17692_n4887) );
  OR2X2 OR2X2_1536 ( .A(_abc_17692_n4891), .B(_abc_17692_n4827), .Y(_abc_17692_n4892) );
  OR2X2 OR2X2_1537 ( .A(_abc_17692_n4890), .B(_abc_17692_n4828), .Y(_abc_17692_n4893_1) );
  OR2X2 OR2X2_1538 ( .A(_abc_17692_n4899), .B(_abc_17692_n4800), .Y(_abc_17692_n4900) );
  OR2X2 OR2X2_1539 ( .A(_abc_17692_n4901), .B(_abc_17692_n4797), .Y(_abc_17692_n4902) );
  OR2X2 OR2X2_154 ( .A(_abc_17692_n725_bF_buf6), .B(_auto_iopadmap_cc_313_execute_30032_24_), .Y(_abc_17692_n895) );
  OR2X2 OR2X2_1540 ( .A(_abc_17692_n4904), .B(_abc_17692_n4895), .Y(_abc_17692_n4905) );
  OR2X2 OR2X2_1541 ( .A(_abc_17692_n4905), .B(_abc_17692_n4889), .Y(_abc_17692_n4906) );
  OR2X2 OR2X2_1542 ( .A(_abc_17692_n4906), .B(_abc_17692_n4880), .Y(_abc_17692_n4907) );
  OR2X2 OR2X2_1543 ( .A(_abc_17692_n4909), .B(_abc_17692_n4910), .Y(_abc_17692_n4911) );
  OR2X2 OR2X2_1544 ( .A(_abc_17692_n4908), .B(_abc_17692_n4911), .Y(_abc_17692_n4912) );
  OR2X2 OR2X2_1545 ( .A(_abc_17692_n4912), .B(_abc_17692_n4871), .Y(workunit2_15__FF_INPUT) );
  OR2X2 OR2X2_1546 ( .A(_abc_17692_n4920), .B(_abc_17692_n4734), .Y(_abc_17692_n4921) );
  OR2X2 OR2X2_1547 ( .A(_abc_17692_n4919), .B(_abc_17692_n4921), .Y(_abc_17692_n4922) );
  OR2X2 OR2X2_1548 ( .A(_abc_17692_n4918), .B(_abc_17692_n4922), .Y(_abc_17692_n4923) );
  OR2X2 OR2X2_1549 ( .A(_abc_17692_n4923), .B(_abc_17692_n4917), .Y(_abc_17692_n4924) );
  OR2X2 OR2X2_155 ( .A(_abc_17692_n727_bF_buf7), .B(workunit1_24_), .Y(_abc_17692_n896) );
  OR2X2 OR2X2_1550 ( .A(_abc_17692_n3026), .B(workunit1_21_), .Y(_abc_17692_n4925) );
  OR2X2 OR2X2_1551 ( .A(_abc_17692_n4926), .B(workunit1_12_bF_buf1), .Y(_abc_17692_n4927) );
  OR2X2 OR2X2_1552 ( .A(_abc_17692_n4930), .B(_abc_17692_n4931), .Y(_abc_17692_n4932) );
  OR2X2 OR2X2_1553 ( .A(_abc_17692_n4503), .B(_abc_17692_n4935), .Y(_abc_17692_n4936) );
  OR2X2 OR2X2_1554 ( .A(_abc_17692_n4936), .B(_abc_17692_n4055), .Y(_abc_17692_n4937) );
  OR2X2 OR2X2_1555 ( .A(_abc_17692_n3226), .B(_abc_17692_n4937), .Y(_abc_17692_n4938) );
  OR2X2 OR2X2_1556 ( .A(_abc_17692_n4069), .B(_abc_17692_n4936), .Y(_abc_17692_n4939) );
  OR2X2 OR2X2_1557 ( .A(_abc_17692_n4943), .B(_abc_17692_n4934), .Y(_abc_17692_n4944) );
  OR2X2 OR2X2_1558 ( .A(_abc_17692_n4951), .B(_abc_17692_n4747), .Y(_abc_17692_n4952) );
  OR2X2 OR2X2_1559 ( .A(_abc_17692_n4950), .B(_abc_17692_n4952), .Y(_abc_17692_n4953) );
  OR2X2 OR2X2_156 ( .A(_abc_17692_n725_bF_buf5), .B(_auto_iopadmap_cc_313_execute_30032_25_), .Y(_abc_17692_n898) );
  OR2X2 OR2X2_1560 ( .A(_abc_17692_n4949), .B(_abc_17692_n4953), .Y(_abc_17692_n4954) );
  OR2X2 OR2X2_1561 ( .A(_abc_17692_n4948), .B(_abc_17692_n4954), .Y(_abc_17692_n4955) );
  OR2X2 OR2X2_1562 ( .A(sum_16_), .B(\key_in[80] ), .Y(_abc_17692_n4958) );
  OR2X2 OR2X2_1563 ( .A(_abc_17692_n4963_1), .B(_abc_17692_n4960), .Y(_abc_17692_n4964) );
  OR2X2 OR2X2_1564 ( .A(_abc_17692_n4965), .B(_abc_17692_n4944), .Y(_abc_17692_n4966_1) );
  OR2X2 OR2X2_1565 ( .A(_abc_17692_n4967), .B(_abc_17692_n4964), .Y(_abc_17692_n4968) );
  OR2X2 OR2X2_1566 ( .A(_abc_17692_n4969), .B(workunit2_16_bF_buf1), .Y(_abc_17692_n4972) );
  OR2X2 OR2X2_1567 ( .A(_abc_17692_n4977), .B(_abc_17692_n4976), .Y(_abc_17692_n4978) );
  OR2X2 OR2X2_1568 ( .A(_abc_17692_n4978), .B(_abc_17692_n4975), .Y(_abc_17692_n4979) );
  OR2X2 OR2X2_1569 ( .A(_abc_17692_n4981), .B(_abc_17692_n4979), .Y(_abc_17692_n4982) );
  OR2X2 OR2X2_157 ( .A(_abc_17692_n727_bF_buf6), .B(workunit1_25_), .Y(_abc_17692_n899) );
  OR2X2 OR2X2_1570 ( .A(_abc_17692_n4982), .B(_abc_17692_n4973), .Y(_abc_17692_n4985) );
  OR2X2 OR2X2_1571 ( .A(_abc_17692_n4994), .B(_abc_17692_n4807), .Y(_abc_17692_n4995) );
  OR2X2 OR2X2_1572 ( .A(_abc_17692_n4993), .B(_abc_17692_n4995), .Y(_abc_17692_n4996) );
  OR2X2 OR2X2_1573 ( .A(_abc_17692_n4992), .B(_abc_17692_n4996), .Y(_abc_17692_n4997) );
  OR2X2 OR2X2_1574 ( .A(_abc_17692_n4991), .B(_abc_17692_n4997), .Y(_abc_17692_n4998) );
  OR2X2 OR2X2_1575 ( .A(sum_16_), .B(\key_in[48] ), .Y(_abc_17692_n5001) );
  OR2X2 OR2X2_1576 ( .A(_abc_17692_n3287), .B(_abc_17692_n5004), .Y(_abc_17692_n5005) );
  OR2X2 OR2X2_1577 ( .A(_abc_17692_n5009), .B(_abc_17692_n5003), .Y(_abc_17692_n5010) );
  OR2X2 OR2X2_1578 ( .A(_abc_17692_n5011), .B(_abc_17692_n4944), .Y(_abc_17692_n5012) );
  OR2X2 OR2X2_1579 ( .A(_abc_17692_n4967), .B(_abc_17692_n5010), .Y(_abc_17692_n5013) );
  OR2X2 OR2X2_158 ( .A(_abc_17692_n725_bF_buf4), .B(_auto_iopadmap_cc_313_execute_30032_26_), .Y(_abc_17692_n901) );
  OR2X2 OR2X2_1580 ( .A(_abc_17692_n5014), .B(workunit2_16_bF_buf3), .Y(_abc_17692_n5017) );
  OR2X2 OR2X2_1581 ( .A(_abc_17692_n4827), .B(_abc_17692_n4648), .Y(_abc_17692_n5019) );
  OR2X2 OR2X2_1582 ( .A(_abc_17692_n5019), .B(_abc_17692_n4653), .Y(_abc_17692_n5020) );
  OR2X2 OR2X2_1583 ( .A(_abc_17692_n4826), .B(_abc_17692_n4830), .Y(_abc_17692_n5022) );
  OR2X2 OR2X2_1584 ( .A(_abc_17692_n5019), .B(_abc_17692_n4655), .Y(_abc_17692_n5025) );
  OR2X2 OR2X2_1585 ( .A(_abc_17692_n5025), .B(_abc_17692_n4237), .Y(_abc_17692_n5026) );
  OR2X2 OR2X2_1586 ( .A(_abc_17692_n5028), .B(_abc_17692_n5018), .Y(_abc_17692_n5031) );
  OR2X2 OR2X2_1587 ( .A(_abc_17692_n5040), .B(_abc_17692_n4780), .Y(_abc_17692_n5041) );
  OR2X2 OR2X2_1588 ( .A(_abc_17692_n5039), .B(_abc_17692_n5041), .Y(_abc_17692_n5042) );
  OR2X2 OR2X2_1589 ( .A(_abc_17692_n5038), .B(_abc_17692_n5042), .Y(_abc_17692_n5043) );
  OR2X2 OR2X2_159 ( .A(_abc_17692_n727_bF_buf5), .B(workunit1_26_), .Y(_abc_17692_n902) );
  OR2X2 OR2X2_1590 ( .A(_abc_17692_n5037), .B(_abc_17692_n5043), .Y(_abc_17692_n5044_1) );
  OR2X2 OR2X2_1591 ( .A(sum_16_), .B(\key_in[16] ), .Y(_abc_17692_n5047_1) );
  OR2X2 OR2X2_1592 ( .A(_abc_17692_n3320), .B(_abc_17692_n5050), .Y(_abc_17692_n5051) );
  OR2X2 OR2X2_1593 ( .A(_abc_17692_n5055), .B(_abc_17692_n5049), .Y(_abc_17692_n5056) );
  OR2X2 OR2X2_1594 ( .A(_abc_17692_n5057), .B(_abc_17692_n4944), .Y(_abc_17692_n5058) );
  OR2X2 OR2X2_1595 ( .A(_abc_17692_n4967), .B(_abc_17692_n5056), .Y(_abc_17692_n5059) );
  OR2X2 OR2X2_1596 ( .A(_abc_17692_n5060), .B(workunit2_16_bF_buf1), .Y(_abc_17692_n5063) );
  OR2X2 OR2X2_1597 ( .A(_abc_17692_n4797), .B(_abc_17692_n4707), .Y(_abc_17692_n5065) );
  OR2X2 OR2X2_1598 ( .A(_abc_17692_n5065), .B(_abc_17692_n4612), .Y(_abc_17692_n5066) );
  OR2X2 OR2X2_1599 ( .A(_abc_17692_n4796), .B(_abc_17692_n4607), .Y(_abc_17692_n5068) );
  OR2X2 OR2X2_16 ( .A(state_8_bF_buf5), .B(delta_17_), .Y(delta_17__FF_INPUT) );
  OR2X2 OR2X2_160 ( .A(_abc_17692_n725_bF_buf3), .B(_auto_iopadmap_cc_313_execute_30032_27_), .Y(_abc_17692_n904) );
  OR2X2 OR2X2_1600 ( .A(_abc_17692_n5065), .B(_abc_17692_n4614), .Y(_abc_17692_n5071) );
  OR2X2 OR2X2_1601 ( .A(_abc_17692_n4196), .B(_abc_17692_n5071), .Y(_abc_17692_n5072) );
  OR2X2 OR2X2_1602 ( .A(_abc_17692_n5074), .B(_abc_17692_n5064), .Y(_abc_17692_n5077) );
  OR2X2 OR2X2_1603 ( .A(_abc_17692_n5079), .B(_abc_17692_n5033), .Y(_abc_17692_n5080) );
  OR2X2 OR2X2_1604 ( .A(_abc_17692_n5080), .B(_abc_17692_n4987), .Y(_abc_17692_n5081) );
  OR2X2 OR2X2_1605 ( .A(_abc_17692_n5088), .B(_abc_17692_n4842), .Y(_abc_17692_n5089) );
  OR2X2 OR2X2_1606 ( .A(_abc_17692_n5087), .B(_abc_17692_n5089), .Y(_abc_17692_n5090) );
  OR2X2 OR2X2_1607 ( .A(_abc_17692_n5086), .B(_abc_17692_n5090), .Y(_abc_17692_n5091) );
  OR2X2 OR2X2_1608 ( .A(_abc_17692_n5085), .B(_abc_17692_n5091), .Y(_abc_17692_n5092) );
  OR2X2 OR2X2_1609 ( .A(sum_16_), .B(\key_in[112] ), .Y(_abc_17692_n5095) );
  OR2X2 OR2X2_161 ( .A(_abc_17692_n727_bF_buf4), .B(workunit1_27_), .Y(_abc_17692_n905) );
  OR2X2 OR2X2_1610 ( .A(_abc_17692_n5102), .B(_abc_17692_n5097_1), .Y(_abc_17692_n5103) );
  OR2X2 OR2X2_1611 ( .A(_abc_17692_n5104), .B(_abc_17692_n4944), .Y(_abc_17692_n5105) );
  OR2X2 OR2X2_1612 ( .A(_abc_17692_n5103), .B(_abc_17692_n4967), .Y(_abc_17692_n5106) );
  OR2X2 OR2X2_1613 ( .A(_abc_17692_n5107), .B(workunit2_16_bF_buf3), .Y(_abc_17692_n5110) );
  OR2X2 OR2X2_1614 ( .A(_abc_17692_n4862), .B(_abc_17692_n4669), .Y(_abc_17692_n5112) );
  OR2X2 OR2X2_1615 ( .A(_abc_17692_n5112), .B(_abc_17692_n4540), .Y(_abc_17692_n5113) );
  OR2X2 OR2X2_1616 ( .A(_abc_17692_n5115), .B(_abc_17692_n4861), .Y(_abc_17692_n5116) );
  OR2X2 OR2X2_1617 ( .A(_abc_17692_n5112), .B(_abc_17692_n5118), .Y(_abc_17692_n5119) );
  OR2X2 OR2X2_1618 ( .A(_abc_17692_n4113), .B(_abc_17692_n5119), .Y(_abc_17692_n5120) );
  OR2X2 OR2X2_1619 ( .A(_abc_17692_n5122), .B(_abc_17692_n5111), .Y(_abc_17692_n5123) );
  OR2X2 OR2X2_162 ( .A(_abc_17692_n725_bF_buf2), .B(_auto_iopadmap_cc_313_execute_30032_28_), .Y(_abc_17692_n907) );
  OR2X2 OR2X2_1620 ( .A(_abc_17692_n5127), .B(_abc_17692_n5081), .Y(_abc_17692_n5128) );
  OR2X2 OR2X2_1621 ( .A(_abc_17692_n5134), .B(_abc_17692_n5133), .Y(_abc_17692_n5135) );
  OR2X2 OR2X2_1622 ( .A(_abc_17692_n5135), .B(_abc_17692_n5132), .Y(_abc_17692_n5136) );
  OR2X2 OR2X2_1623 ( .A(_abc_17692_n5138), .B(_abc_17692_n5136), .Y(_abc_17692_n5139) );
  OR2X2 OR2X2_1624 ( .A(_abc_17692_n5139), .B(_abc_17692_n5130), .Y(_abc_17692_n5140) );
  OR2X2 OR2X2_1625 ( .A(_abc_17692_n4770), .B(_abc_17692_n4573), .Y(_abc_17692_n5146) );
  OR2X2 OR2X2_1626 ( .A(_abc_17692_n5146), .B(_abc_17692_n4684), .Y(_abc_17692_n5147) );
  OR2X2 OR2X2_1627 ( .A(_abc_17692_n4764), .B(_abc_17692_n4882), .Y(_abc_17692_n5149) );
  OR2X2 OR2X2_1628 ( .A(_abc_17692_n5146), .B(_abc_17692_n4686), .Y(_abc_17692_n5153) );
  OR2X2 OR2X2_1629 ( .A(_abc_17692_n4274), .B(_abc_17692_n5153), .Y(_abc_17692_n5154) );
  OR2X2 OR2X2_163 ( .A(_abc_17692_n727_bF_buf3), .B(workunit1_28_), .Y(_abc_17692_n908) );
  OR2X2 OR2X2_1630 ( .A(_abc_17692_n5156), .B(_abc_17692_n5145), .Y(_abc_17692_n5159) );
  OR2X2 OR2X2_1631 ( .A(_abc_17692_n5167), .B(_abc_17692_n5165), .Y(_abc_17692_n5168) );
  OR2X2 OR2X2_1632 ( .A(_abc_17692_n5168), .B(_abc_17692_n5164), .Y(_abc_17692_n5169) );
  OR2X2 OR2X2_1633 ( .A(_abc_17692_n5169), .B(_abc_17692_n5171), .Y(_abc_17692_n5172) );
  OR2X2 OR2X2_1634 ( .A(_abc_17692_n5172), .B(_abc_17692_n5162), .Y(_abc_17692_n5173) );
  OR2X2 OR2X2_1635 ( .A(_abc_17692_n5182), .B(_abc_17692_n5181), .Y(_abc_17692_n5183) );
  OR2X2 OR2X2_1636 ( .A(_abc_17692_n5183), .B(_abc_17692_n5180), .Y(_abc_17692_n5184) );
  OR2X2 OR2X2_1637 ( .A(_abc_17692_n5184), .B(_abc_17692_n5186), .Y(_abc_17692_n5187) );
  OR2X2 OR2X2_1638 ( .A(_abc_17692_n5187), .B(_abc_17692_n5178), .Y(_abc_17692_n5190) );
  OR2X2 OR2X2_1639 ( .A(_abc_17692_n5192), .B(_abc_17692_n5177), .Y(_abc_17692_n5193) );
  OR2X2 OR2X2_164 ( .A(_abc_17692_n725_bF_buf1), .B(_auto_iopadmap_cc_313_execute_30032_29_), .Y(_abc_17692_n910_1) );
  OR2X2 OR2X2_1640 ( .A(_abc_17692_n5193), .B(_abc_17692_n5161), .Y(_abc_17692_n5194) );
  OR2X2 OR2X2_1641 ( .A(_abc_17692_n5194), .B(_abc_17692_n5144), .Y(_abc_17692_n5195) );
  OR2X2 OR2X2_1642 ( .A(_abc_17692_n5197), .B(_abc_17692_n5198), .Y(_abc_17692_n5199) );
  OR2X2 OR2X2_1643 ( .A(_abc_17692_n5196), .B(_abc_17692_n5199), .Y(_abc_17692_n5200) );
  OR2X2 OR2X2_1644 ( .A(_abc_17692_n5129), .B(_abc_17692_n5200), .Y(workunit2_16__FF_INPUT) );
  OR2X2 OR2X2_1645 ( .A(_abc_17692_n4934), .B(_abc_17692_n4930), .Y(_abc_17692_n5203) );
  OR2X2 OR2X2_1646 ( .A(_abc_17692_n3208), .B(workunit1_22_), .Y(_abc_17692_n5204) );
  OR2X2 OR2X2_1647 ( .A(_abc_17692_n5205), .B(workunit1_13_bF_buf1), .Y(_abc_17692_n5206) );
  OR2X2 OR2X2_1648 ( .A(_abc_17692_n5203), .B(_abc_17692_n5214), .Y(_abc_17692_n5215_1) );
  OR2X2 OR2X2_1649 ( .A(sum_17_), .B(\key_in[17] ), .Y(_abc_17692_n5223) );
  OR2X2 OR2X2_165 ( .A(_abc_17692_n727_bF_buf2), .B(workunit1_29_), .Y(_abc_17692_n911_1) );
  OR2X2 OR2X2_1650 ( .A(_abc_17692_n5220), .B(_abc_17692_n5224), .Y(_abc_17692_n5227) );
  OR2X2 OR2X2_1651 ( .A(_abc_17692_n5228), .B(_abc_17692_n5218), .Y(_abc_17692_n5229) );
  OR2X2 OR2X2_1652 ( .A(_abc_17692_n5231), .B(_abc_17692_n5230), .Y(_abc_17692_n5232) );
  OR2X2 OR2X2_1653 ( .A(_abc_17692_n5233), .B(workunit2_17_), .Y(_abc_17692_n5236) );
  OR2X2 OR2X2_1654 ( .A(_abc_17692_n5241), .B(_abc_17692_n5239), .Y(_abc_17692_n5242) );
  OR2X2 OR2X2_1655 ( .A(sum_17_), .B(\key_in[81] ), .Y(_abc_17692_n5248) );
  OR2X2 OR2X2_1656 ( .A(_abc_17692_n5245), .B(_abc_17692_n5249), .Y(_abc_17692_n5252) );
  OR2X2 OR2X2_1657 ( .A(_abc_17692_n5253), .B(_abc_17692_n5218), .Y(_abc_17692_n5254) );
  OR2X2 OR2X2_1658 ( .A(_abc_17692_n5255), .B(_abc_17692_n5230), .Y(_abc_17692_n5256) );
  OR2X2 OR2X2_1659 ( .A(_abc_17692_n5265), .B(_abc_17692_n4970), .Y(_abc_17692_n5266) );
  OR2X2 OR2X2_166 ( .A(_abc_17692_n725_bF_buf0), .B(_auto_iopadmap_cc_313_execute_30032_30_), .Y(_abc_17692_n913) );
  OR2X2 OR2X2_1660 ( .A(_abc_17692_n4983), .B(_abc_17692_n5266), .Y(_abc_17692_n5267) );
  OR2X2 OR2X2_1661 ( .A(_abc_17692_n5264), .B(_abc_17692_n4971), .Y(_abc_17692_n5271) );
  OR2X2 OR2X2_1662 ( .A(sum_17_), .B(\key_in[49] ), .Y(_abc_17692_n5281) );
  OR2X2 OR2X2_1663 ( .A(_abc_17692_n5278_1), .B(_abc_17692_n5282), .Y(_abc_17692_n5285) );
  OR2X2 OR2X2_1664 ( .A(_abc_17692_n5288), .B(_abc_17692_n5289), .Y(_abc_17692_n5290) );
  OR2X2 OR2X2_1665 ( .A(_abc_17692_n5290), .B(_abc_17692_n5260), .Y(_abc_17692_n5291) );
  OR2X2 OR2X2_1666 ( .A(_abc_17692_n5292), .B(workunit2_17_), .Y(_abc_17692_n5293) );
  OR2X2 OR2X2_1667 ( .A(_abc_17692_n5276), .B(_abc_17692_n5295), .Y(_abc_17692_n5296) );
  OR2X2 OR2X2_1668 ( .A(_abc_17692_n5275_1), .B(_abc_17692_n5294), .Y(_abc_17692_n5297) );
  OR2X2 OR2X2_1669 ( .A(_abc_17692_n5299), .B(_abc_17692_n5274), .Y(_abc_17692_n5300) );
  OR2X2 OR2X2_167 ( .A(_abc_17692_n727_bF_buf1), .B(workunit1_30_), .Y(_abc_17692_n914) );
  OR2X2 OR2X2_1670 ( .A(_abc_17692_n5243), .B(_abc_17692_n5300), .Y(_abc_17692_n5301) );
  OR2X2 OR2X2_1671 ( .A(sum_17_), .B(\key_in[113] ), .Y(_abc_17692_n5307) );
  OR2X2 OR2X2_1672 ( .A(_abc_17692_n5304), .B(_abc_17692_n5308), .Y(_abc_17692_n5311) );
  OR2X2 OR2X2_1673 ( .A(_abc_17692_n5312), .B(_abc_17692_n5218), .Y(_abc_17692_n5313) );
  OR2X2 OR2X2_1674 ( .A(_abc_17692_n5314), .B(_abc_17692_n5230), .Y(_abc_17692_n5315) );
  OR2X2 OR2X2_1675 ( .A(_abc_17692_n5326), .B(_abc_17692_n5324), .Y(_abc_17692_n5327) );
  OR2X2 OR2X2_1676 ( .A(_abc_17692_n5328), .B(_abc_17692_n5301), .Y(_abc_17692_n5329) );
  OR2X2 OR2X2_1677 ( .A(_abc_17692_n5336), .B(_abc_17692_n5337), .Y(_abc_17692_n5338) );
  OR2X2 OR2X2_1678 ( .A(_abc_17692_n5344), .B(_abc_17692_n5264), .Y(_abc_17692_n5345) );
  OR2X2 OR2X2_1679 ( .A(_abc_17692_n5343), .B(_abc_17692_n5265), .Y(_abc_17692_n5346) );
  OR2X2 OR2X2_168 ( .A(_abc_17692_n725_bF_buf7), .B(_auto_iopadmap_cc_313_execute_30032_31_), .Y(_abc_17692_n916) );
  OR2X2 OR2X2_1680 ( .A(_abc_17692_n5353), .B(_abc_17692_n5294), .Y(_abc_17692_n5354) );
  OR2X2 OR2X2_1681 ( .A(_abc_17692_n5352), .B(_abc_17692_n5295), .Y(_abc_17692_n5355) );
  OR2X2 OR2X2_1682 ( .A(_abc_17692_n5362), .B(_abc_17692_n5237), .Y(_abc_17692_n5363) );
  OR2X2 OR2X2_1683 ( .A(_abc_17692_n5361), .B(_abc_17692_n5238), .Y(_abc_17692_n5364) );
  OR2X2 OR2X2_1684 ( .A(_abc_17692_n5366_1), .B(_abc_17692_n5357), .Y(_abc_17692_n5367) );
  OR2X2 OR2X2_1685 ( .A(_abc_17692_n5367), .B(_abc_17692_n5348), .Y(_abc_17692_n5368) );
  OR2X2 OR2X2_1686 ( .A(_abc_17692_n5368), .B(_abc_17692_n5339), .Y(_abc_17692_n5369_1) );
  OR2X2 OR2X2_1687 ( .A(_abc_17692_n5371), .B(_abc_17692_n5372), .Y(_abc_17692_n5373) );
  OR2X2 OR2X2_1688 ( .A(_abc_17692_n5370), .B(_abc_17692_n5373), .Y(_abc_17692_n5374) );
  OR2X2 OR2X2_1689 ( .A(_abc_17692_n5330), .B(_abc_17692_n5374), .Y(workunit2_17__FF_INPUT) );
  OR2X2 OR2X2_169 ( .A(_abc_17692_n727_bF_buf0), .B(workunit1_31_), .Y(_abc_17692_n917) );
  OR2X2 OR2X2_1690 ( .A(_abc_17692_n5376), .B(workunit1_23_), .Y(_abc_17692_n5377) );
  OR2X2 OR2X2_1691 ( .A(_abc_17692_n5378), .B(workunit1_14_bF_buf1), .Y(_abc_17692_n5379) );
  OR2X2 OR2X2_1692 ( .A(_abc_17692_n5382), .B(_abc_17692_n5383), .Y(_abc_17692_n5384) );
  OR2X2 OR2X2_1693 ( .A(_abc_17692_n5386), .B(_abc_17692_n5209), .Y(_abc_17692_n5387) );
  OR2X2 OR2X2_1694 ( .A(_abc_17692_n5389), .B(_abc_17692_n5387), .Y(_abc_17692_n5390) );
  OR2X2 OR2X2_1695 ( .A(_abc_17692_n5393), .B(_abc_17692_n5391), .Y(_abc_17692_n5394) );
  OR2X2 OR2X2_1696 ( .A(sum_18_), .B(\key_in[82] ), .Y(_abc_17692_n5397) );
  OR2X2 OR2X2_1697 ( .A(_abc_17692_n5400), .B(_abc_17692_n5246), .Y(_abc_17692_n5401) );
  OR2X2 OR2X2_1698 ( .A(_abc_17692_n4961), .B(_abc_17692_n5404), .Y(_abc_17692_n5405) );
  OR2X2 OR2X2_1699 ( .A(_abc_17692_n5406), .B(_abc_17692_n5399), .Y(_abc_17692_n5407) );
  OR2X2 OR2X2_17 ( .A(state_8_bF_buf4), .B(delta_18_), .Y(delta_18__FF_INPUT) );
  OR2X2 OR2X2_170 ( .A(delta_0_), .B(sum_0_), .Y(_abc_17692_n920) );
  OR2X2 OR2X2_1700 ( .A(_abc_17692_n5408), .B(_abc_17692_n5409), .Y(_abc_17692_n5410) );
  OR2X2 OR2X2_1701 ( .A(_abc_17692_n5414), .B(_abc_17692_n5411), .Y(_abc_17692_n5415) );
  OR2X2 OR2X2_1702 ( .A(_abc_17692_n5415), .B(workunit2_18_), .Y(_abc_17692_n5418) );
  OR2X2 OR2X2_1703 ( .A(_abc_17692_n5424), .B(_abc_17692_n5419), .Y(_abc_17692_n5427) );
  OR2X2 OR2X2_1704 ( .A(sum_18_), .B(\key_in[50] ), .Y(_abc_17692_n5433) );
  OR2X2 OR2X2_1705 ( .A(_abc_17692_n5435), .B(_abc_17692_n5279), .Y(_abc_17692_n5436) );
  OR2X2 OR2X2_1706 ( .A(_abc_17692_n5438), .B(_abc_17692_n5436), .Y(_abc_17692_n5439) );
  OR2X2 OR2X2_1707 ( .A(_abc_17692_n5443), .B(_abc_17692_n5440), .Y(_abc_17692_n5444) );
  OR2X2 OR2X2_1708 ( .A(_abc_17692_n5447), .B(_abc_17692_n5445), .Y(_abc_17692_n5448) );
  OR2X2 OR2X2_1709 ( .A(_abc_17692_n5448), .B(_abc_17692_n5430), .Y(_abc_17692_n5449) );
  OR2X2 OR2X2_171 ( .A(_abc_17692_n919), .B(_abc_17692_n924), .Y(sum_0__FF_INPUT) );
  OR2X2 OR2X2_1710 ( .A(_abc_17692_n5450), .B(workunit2_18_), .Y(_abc_17692_n5451) );
  OR2X2 OR2X2_1711 ( .A(_abc_17692_n5294), .B(_abc_17692_n5016), .Y(_abc_17692_n5456) );
  OR2X2 OR2X2_1712 ( .A(_abc_17692_n5460), .B(_abc_17692_n5458), .Y(_abc_17692_n5461) );
  OR2X2 OR2X2_1713 ( .A(_abc_17692_n5461), .B(_abc_17692_n5453), .Y(_abc_17692_n5464) );
  OR2X2 OR2X2_1714 ( .A(_abc_17692_n5470), .B(_abc_17692_n5469), .Y(_abc_17692_n5471) );
  OR2X2 OR2X2_1715 ( .A(_abc_17692_n5468), .B(_abc_17692_n5472), .Y(_abc_17692_n5473) );
  OR2X2 OR2X2_1716 ( .A(sum_18_), .B(\key_in[18] ), .Y(_abc_17692_n5476) );
  OR2X2 OR2X2_1717 ( .A(_abc_17692_n5481), .B(_abc_17692_n5478), .Y(_abc_17692_n5482) );
  OR2X2 OR2X2_1718 ( .A(_abc_17692_n5483), .B(_abc_17692_n5394), .Y(_abc_17692_n5484) );
  OR2X2 OR2X2_1719 ( .A(_abc_17692_n5412), .B(_abc_17692_n5482), .Y(_abc_17692_n5485) );
  OR2X2 OR2X2_172 ( .A(_abc_17692_n926_1), .B(sum_1_), .Y(_abc_17692_n927_1) );
  OR2X2 OR2X2_1720 ( .A(_abc_17692_n5486), .B(_abc_17692_n5430), .Y(_abc_17692_n5487) );
  OR2X2 OR2X2_1721 ( .A(_abc_17692_n5488), .B(workunit2_18_), .Y(_abc_17692_n5489) );
  OR2X2 OR2X2_1722 ( .A(_abc_17692_n5233), .B(_abc_17692_n5260), .Y(_abc_17692_n5492) );
  OR2X2 OR2X2_1723 ( .A(_abc_17692_n5237), .B(_abc_17692_n5062), .Y(_abc_17692_n5493) );
  OR2X2 OR2X2_1724 ( .A(_abc_17692_n5497), .B(_abc_17692_n5495), .Y(_abc_17692_n5498) );
  OR2X2 OR2X2_1725 ( .A(_abc_17692_n5498), .B(_abc_17692_n5491), .Y(_abc_17692_n5499) );
  OR2X2 OR2X2_1726 ( .A(_abc_17692_n5503), .B(_abc_17692_n5466), .Y(_abc_17692_n5504) );
  OR2X2 OR2X2_1727 ( .A(_abc_17692_n5504), .B(_abc_17692_n5429), .Y(_abc_17692_n5505) );
  OR2X2 OR2X2_1728 ( .A(_abc_17692_n5509), .B(_abc_17692_n5508), .Y(_abc_17692_n5510) );
  OR2X2 OR2X2_1729 ( .A(_abc_17692_n5507), .B(_abc_17692_n5511), .Y(_abc_17692_n5512) );
  OR2X2 OR2X2_173 ( .A(_abc_17692_n931), .B(sum_0_), .Y(_abc_17692_n932) );
  OR2X2 OR2X2_1730 ( .A(sum_18_), .B(\key_in[114] ), .Y(_abc_17692_n5515) );
  OR2X2 OR2X2_1731 ( .A(_abc_17692_n5520), .B(_abc_17692_n5517), .Y(_abc_17692_n5521) );
  OR2X2 OR2X2_1732 ( .A(_abc_17692_n5522), .B(_abc_17692_n5394), .Y(_abc_17692_n5523) );
  OR2X2 OR2X2_1733 ( .A(_abc_17692_n5521), .B(_abc_17692_n5412), .Y(_abc_17692_n5524) );
  OR2X2 OR2X2_1734 ( .A(_abc_17692_n5527), .B(_abc_17692_n5528), .Y(_abc_17692_n5529) );
  OR2X2 OR2X2_1735 ( .A(_abc_17692_n5322), .B(_abc_17692_n5109), .Y(_abc_17692_n5533) );
  OR2X2 OR2X2_1736 ( .A(_abc_17692_n5537), .B(_abc_17692_n5535), .Y(_abc_17692_n5538) );
  OR2X2 OR2X2_1737 ( .A(_abc_17692_n5538), .B(_abc_17692_n5530), .Y(_abc_17692_n5541) );
  OR2X2 OR2X2_1738 ( .A(_abc_17692_n5505), .B(_abc_17692_n5543), .Y(_abc_17692_n5544) );
  OR2X2 OR2X2_1739 ( .A(_abc_17692_n5317), .B(_abc_17692_n5332), .Y(_abc_17692_n5546) );
  OR2X2 OR2X2_174 ( .A(_abc_17692_n930_1), .B(_abc_17692_n932), .Y(_abc_17692_n935) );
  OR2X2 OR2X2_1740 ( .A(_abc_17692_n5549), .B(_abc_17692_n5547), .Y(_abc_17692_n5550) );
  OR2X2 OR2X2_1741 ( .A(_abc_17692_n5550), .B(_abc_17692_n5529), .Y(_abc_17692_n5553) );
  OR2X2 OR2X2_1742 ( .A(_abc_17692_n5557), .B(_abc_17692_n5258), .Y(_abc_17692_n5558) );
  OR2X2 OR2X2_1743 ( .A(_abc_17692_n5558), .B(_abc_17692_n5556), .Y(_abc_17692_n5561) );
  OR2X2 OR2X2_1744 ( .A(_abc_17692_n5234), .B(_abc_17692_n5359), .Y(_abc_17692_n5564) );
  OR2X2 OR2X2_1745 ( .A(_abc_17692_n5567), .B(_abc_17692_n5565), .Y(_abc_17692_n5568) );
  OR2X2 OR2X2_1746 ( .A(_abc_17692_n5568), .B(_abc_17692_n5490), .Y(_abc_17692_n5571) );
  OR2X2 OR2X2_1747 ( .A(_abc_17692_n5574), .B(_abc_17692_n5575), .Y(_abc_17692_n5576) );
  OR2X2 OR2X2_1748 ( .A(_abc_17692_n5579), .B(_abc_17692_n5577), .Y(_abc_17692_n5580) );
  OR2X2 OR2X2_1749 ( .A(_abc_17692_n5580), .B(_abc_17692_n5452), .Y(_abc_17692_n5583) );
  OR2X2 OR2X2_175 ( .A(_abc_17692_n930_1), .B(_abc_17692_n922), .Y(_abc_17692_n939) );
  OR2X2 OR2X2_1750 ( .A(_abc_17692_n5573), .B(_abc_17692_n5585), .Y(_abc_17692_n5586) );
  OR2X2 OR2X2_1751 ( .A(_abc_17692_n5563), .B(_abc_17692_n5586), .Y(_abc_17692_n5587) );
  OR2X2 OR2X2_1752 ( .A(_abc_17692_n5587), .B(_abc_17692_n5555), .Y(_abc_17692_n5588) );
  OR2X2 OR2X2_1753 ( .A(_abc_17692_n5590), .B(_abc_17692_n5591), .Y(_abc_17692_n5592) );
  OR2X2 OR2X2_1754 ( .A(_abc_17692_n5589), .B(_abc_17692_n5592), .Y(_abc_17692_n5593) );
  OR2X2 OR2X2_1755 ( .A(_abc_17692_n5593), .B(_abc_17692_n5545_1), .Y(workunit2_18__FF_INPUT) );
  OR2X2 OR2X2_1756 ( .A(_abc_17692_n5391), .B(_abc_17692_n5382), .Y(_abc_17692_n5595) );
  OR2X2 OR2X2_1757 ( .A(_abc_17692_n3614), .B(workunit1_24_), .Y(_abc_17692_n5597) );
  OR2X2 OR2X2_1758 ( .A(_abc_17692_n5598), .B(workunit1_15_), .Y(_abc_17692_n5599) );
  OR2X2 OR2X2_1759 ( .A(_abc_17692_n5607), .B(_abc_17692_n5609), .Y(_abc_17692_n5610) );
  OR2X2 OR2X2_176 ( .A(_abc_17692_n940), .B(_abc_17692_n921), .Y(_abc_17692_n941) );
  OR2X2 OR2X2_1760 ( .A(sum_19_), .B(\key_in[83] ), .Y(_abc_17692_n5615) );
  OR2X2 OR2X2_1761 ( .A(_abc_17692_n5612), .B(_abc_17692_n5616), .Y(_abc_17692_n5619) );
  OR2X2 OR2X2_1762 ( .A(_abc_17692_n5611_1), .B(_abc_17692_n5620), .Y(_abc_17692_n5621) );
  OR2X2 OR2X2_1763 ( .A(_abc_17692_n5622), .B(_abc_17692_n5610), .Y(_abc_17692_n5623) );
  OR2X2 OR2X2_1764 ( .A(_abc_17692_n5628), .B(_abc_17692_n5625), .Y(_abc_17692_n5629) );
  OR2X2 OR2X2_1765 ( .A(_abc_17692_n5559), .B(_abc_17692_n5631), .Y(_abc_17692_n5632) );
  OR2X2 OR2X2_1766 ( .A(_abc_17692_n5636), .B(_abc_17692_n5633), .Y(_abc_17692_n5637) );
  OR2X2 OR2X2_1767 ( .A(_abc_17692_n5517), .B(_abc_17692_n5513), .Y(_abc_17692_n5639) );
  OR2X2 OR2X2_1768 ( .A(sum_19_), .B(\key_in[115] ), .Y(_abc_17692_n5643) );
  OR2X2 OR2X2_1769 ( .A(_abc_17692_n5640), .B(_abc_17692_n5644), .Y(_abc_17692_n5647) );
  OR2X2 OR2X2_177 ( .A(_abc_17692_n943), .B(_abc_17692_n938), .Y(_abc_17692_n944) );
  OR2X2 OR2X2_1770 ( .A(_abc_17692_n5648), .B(_abc_17692_n5611_1), .Y(_abc_17692_n5649) );
  OR2X2 OR2X2_1771 ( .A(_abc_17692_n5650), .B(_abc_17692_n5645), .Y(_abc_17692_n5651) );
  OR2X2 OR2X2_1772 ( .A(_abc_17692_n5651), .B(_abc_17692_n5610), .Y(_abc_17692_n5652) );
  OR2X2 OR2X2_1773 ( .A(_abc_17692_n5651), .B(_abc_17692_n5611_1), .Y(_abc_17692_n5655) );
  OR2X2 OR2X2_1774 ( .A(_abc_17692_n5648), .B(_abc_17692_n5610), .Y(_abc_17692_n5656) );
  OR2X2 OR2X2_1775 ( .A(_abc_17692_n5654), .B(_abc_17692_n5658), .Y(_abc_17692_n5659) );
  OR2X2 OR2X2_1776 ( .A(_abc_17692_n5662), .B(_abc_17692_n5659), .Y(_abc_17692_n5663) );
  OR2X2 OR2X2_1777 ( .A(_abc_17692_n5657), .B(_abc_17692_n5626), .Y(_abc_17692_n5664) );
  OR2X2 OR2X2_1778 ( .A(_abc_17692_n5653), .B(workunit2_19_), .Y(_abc_17692_n5665) );
  OR2X2 OR2X2_1779 ( .A(_abc_17692_n5667), .B(_abc_17692_n5666), .Y(_abc_17692_n5668) );
  OR2X2 OR2X2_178 ( .A(_abc_17692_n944), .B(_abc_17692_n937_1), .Y(sum_1__FF_INPUT) );
  OR2X2 OR2X2_1780 ( .A(_abc_17692_n5440), .B(_abc_17692_n5431), .Y(_abc_17692_n5671) );
  OR2X2 OR2X2_1781 ( .A(sum_19_), .B(\key_in[51] ), .Y(_abc_17692_n5675) );
  OR2X2 OR2X2_1782 ( .A(_abc_17692_n5672), .B(_abc_17692_n5676), .Y(_abc_17692_n5678) );
  OR2X2 OR2X2_1783 ( .A(_abc_17692_n5679), .B(_abc_17692_n5677), .Y(_abc_17692_n5680) );
  OR2X2 OR2X2_1784 ( .A(_abc_17692_n5611_1), .B(_abc_17692_n5680), .Y(_abc_17692_n5681) );
  OR2X2 OR2X2_1785 ( .A(_abc_17692_n5683), .B(_abc_17692_n5610), .Y(_abc_17692_n5684) );
  OR2X2 OR2X2_1786 ( .A(_abc_17692_n5685), .B(_abc_17692_n5626), .Y(_abc_17692_n5686) );
  OR2X2 OR2X2_1787 ( .A(_abc_17692_n5611_1), .B(_abc_17692_n5683), .Y(_abc_17692_n5687) );
  OR2X2 OR2X2_1788 ( .A(_abc_17692_n5680), .B(_abc_17692_n5610), .Y(_abc_17692_n5688) );
  OR2X2 OR2X2_1789 ( .A(_abc_17692_n5689), .B(workunit2_19_), .Y(_abc_17692_n5690) );
  OR2X2 OR2X2_179 ( .A(_abc_17692_n946), .B(delta_2_), .Y(_abc_17692_n949_1) );
  OR2X2 OR2X2_1790 ( .A(_abc_17692_n5693), .B(_abc_17692_n5691), .Y(_abc_17692_n5694) );
  OR2X2 OR2X2_1791 ( .A(_abc_17692_n5692_1), .B(_abc_17692_n5695_1), .Y(_abc_17692_n5696) );
  OR2X2 OR2X2_1792 ( .A(_abc_17692_n5478), .B(_abc_17692_n5474), .Y(_abc_17692_n5699) );
  OR2X2 OR2X2_1793 ( .A(sum_19_), .B(\key_in[19] ), .Y(_abc_17692_n5703) );
  OR2X2 OR2X2_1794 ( .A(_abc_17692_n5700), .B(_abc_17692_n5704), .Y(_abc_17692_n5706) );
  OR2X2 OR2X2_1795 ( .A(_abc_17692_n5707), .B(_abc_17692_n5705), .Y(_abc_17692_n5708) );
  OR2X2 OR2X2_1796 ( .A(_abc_17692_n5611_1), .B(_abc_17692_n5708), .Y(_abc_17692_n5709) );
  OR2X2 OR2X2_1797 ( .A(_abc_17692_n5711), .B(_abc_17692_n5610), .Y(_abc_17692_n5712) );
  OR2X2 OR2X2_1798 ( .A(_abc_17692_n5713), .B(_abc_17692_n5626), .Y(_abc_17692_n5714) );
  OR2X2 OR2X2_1799 ( .A(_abc_17692_n5611_1), .B(_abc_17692_n5711), .Y(_abc_17692_n5715) );
  OR2X2 OR2X2_18 ( .A(state_8_bF_buf3), .B(delta_20_), .Y(delta_20__FF_INPUT) );
  OR2X2 OR2X2_180 ( .A(_abc_17692_n955), .B(_abc_17692_n951), .Y(_abc_17692_n956) );
  OR2X2 OR2X2_1800 ( .A(_abc_17692_n5708), .B(_abc_17692_n5610), .Y(_abc_17692_n5716) );
  OR2X2 OR2X2_1801 ( .A(_abc_17692_n5717), .B(workunit2_19_), .Y(_abc_17692_n5718) );
  OR2X2 OR2X2_1802 ( .A(_abc_17692_n5721), .B(_abc_17692_n5720), .Y(_abc_17692_n5722) );
  OR2X2 OR2X2_1803 ( .A(_abc_17692_n5723), .B(_abc_17692_n5719), .Y(_abc_17692_n5724) );
  OR2X2 OR2X2_1804 ( .A(_abc_17692_n5726), .B(_abc_17692_n5698), .Y(_abc_17692_n5727) );
  OR2X2 OR2X2_1805 ( .A(_abc_17692_n5670), .B(_abc_17692_n5727), .Y(_abc_17692_n5728) );
  OR2X2 OR2X2_1806 ( .A(_abc_17692_n5638), .B(_abc_17692_n5728), .Y(_abc_17692_n5729) );
  OR2X2 OR2X2_1807 ( .A(_abc_17692_n5735), .B(_abc_17692_n4047_bF_buf1), .Y(_abc_17692_n5736) );
  OR2X2 OR2X2_1808 ( .A(_abc_17692_n5736), .B(_abc_17692_n5734), .Y(_abc_17692_n5737) );
  OR2X2 OR2X2_1809 ( .A(_abc_17692_n5739), .B(_abc_17692_n5629), .Y(_abc_17692_n5740) );
  OR2X2 OR2X2_181 ( .A(_abc_17692_n954), .B(_abc_17692_n950), .Y(_abc_17692_n957) );
  OR2X2 OR2X2_1810 ( .A(_abc_17692_n5738), .B(_abc_17692_n5634), .Y(_abc_17692_n5741) );
  OR2X2 OR2X2_1811 ( .A(_abc_17692_n5500), .B(_abc_17692_n5744), .Y(_abc_17692_n5745_1) );
  OR2X2 OR2X2_1812 ( .A(_abc_17692_n5746), .B(_abc_17692_n5719), .Y(_abc_17692_n5747) );
  OR2X2 OR2X2_1813 ( .A(_abc_17692_n5745_1), .B(_abc_17692_n5720), .Y(_abc_17692_n5748_1) );
  OR2X2 OR2X2_1814 ( .A(_abc_17692_n5754), .B(_abc_17692_n5695_1), .Y(_abc_17692_n5755) );
  OR2X2 OR2X2_1815 ( .A(_abc_17692_n5753), .B(_abc_17692_n5691), .Y(_abc_17692_n5756) );
  OR2X2 OR2X2_1816 ( .A(_abc_17692_n5758), .B(_abc_17692_n1863_bF_buf4), .Y(_abc_17692_n5759) );
  OR2X2 OR2X2_1817 ( .A(_abc_17692_n5759), .B(_abc_17692_n5750), .Y(_abc_17692_n5760) );
  OR2X2 OR2X2_1818 ( .A(_abc_17692_n5743), .B(_abc_17692_n5760), .Y(_abc_17692_n5761) );
  OR2X2 OR2X2_1819 ( .A(_abc_17692_n5764), .B(_abc_17692_n5765), .Y(_abc_17692_n5766) );
  OR2X2 OR2X2_182 ( .A(_abc_17692_n933), .B(_abc_17692_n928), .Y(_abc_17692_n961) );
  OR2X2 OR2X2_1820 ( .A(_abc_17692_n5763), .B(_abc_17692_n5766), .Y(_abc_17692_n5767) );
  OR2X2 OR2X2_1821 ( .A(_abc_17692_n5767), .B(_abc_17692_n5730), .Y(workunit2_19__FF_INPUT) );
  OR2X2 OR2X2_1822 ( .A(_abc_17692_n5776), .B(_abc_17692_n5604), .Y(_abc_17692_n5777) );
  OR2X2 OR2X2_1823 ( .A(_abc_17692_n5772), .B(_abc_17692_n5779), .Y(_abc_17692_n5780) );
  OR2X2 OR2X2_1824 ( .A(_abc_17692_n3867), .B(workunit1_25_), .Y(_abc_17692_n5781) );
  OR2X2 OR2X2_1825 ( .A(_abc_17692_n5782), .B(workunit1_16_bF_buf2), .Y(_abc_17692_n5783) );
  OR2X2 OR2X2_1826 ( .A(_abc_17692_n5786), .B(_abc_17692_n5787), .Y(_abc_17692_n5788) );
  OR2X2 OR2X2_1827 ( .A(_abc_17692_n4942), .B(_abc_17692_n5791), .Y(_abc_17692_n5792) );
  OR2X2 OR2X2_1828 ( .A(_abc_17692_n5794), .B(_abc_17692_n5790), .Y(_abc_17692_n5795) );
  OR2X2 OR2X2_1829 ( .A(_abc_17692_n5800), .B(_abc_17692_n5641), .Y(_abc_17692_n5801) );
  OR2X2 OR2X2_183 ( .A(_abc_17692_n961), .B(_abc_17692_n950), .Y(_abc_17692_n964_1) );
  OR2X2 OR2X2_1830 ( .A(_abc_17692_n5799), .B(_abc_17692_n5801), .Y(_abc_17692_n5802) );
  OR2X2 OR2X2_1831 ( .A(_abc_17692_n5798), .B(_abc_17692_n5802), .Y(_abc_17692_n5803) );
  OR2X2 OR2X2_1832 ( .A(sum_20_), .B(\key_in[116] ), .Y(_abc_17692_n5806) );
  OR2X2 OR2X2_1833 ( .A(_abc_17692_n5813), .B(_abc_17692_n5808), .Y(_abc_17692_n5814) );
  OR2X2 OR2X2_1834 ( .A(_abc_17692_n5815), .B(_abc_17692_n5795), .Y(_abc_17692_n5816) );
  OR2X2 OR2X2_1835 ( .A(_abc_17692_n5814), .B(_abc_17692_n5817), .Y(_abc_17692_n5818) );
  OR2X2 OR2X2_1836 ( .A(_abc_17692_n5821), .B(_abc_17692_n5822), .Y(_abc_17692_n5823) );
  OR2X2 OR2X2_1837 ( .A(_abc_17692_n5121), .B(_abc_17692_n5827), .Y(_abc_17692_n5828) );
  OR2X2 OR2X2_1838 ( .A(_abc_17692_n5832), .B(_abc_17692_n5831), .Y(_abc_17692_n5833) );
  OR2X2 OR2X2_1839 ( .A(_abc_17692_n5837), .B(_abc_17692_n5824), .Y(_abc_17692_n5840) );
  OR2X2 OR2X2_184 ( .A(_abc_17692_n966), .B(_abc_17692_n960), .Y(_abc_17692_n967_1) );
  OR2X2 OR2X2_1840 ( .A(_abc_17692_n5841), .B(_abc_17692_n4047_bF_buf0), .Y(_abc_17692_n5842) );
  OR2X2 OR2X2_1841 ( .A(_abc_17692_n5847), .B(_abc_17692_n5613), .Y(_abc_17692_n5848) );
  OR2X2 OR2X2_1842 ( .A(_abc_17692_n5846_1), .B(_abc_17692_n5848), .Y(_abc_17692_n5849) );
  OR2X2 OR2X2_1843 ( .A(_abc_17692_n5845), .B(_abc_17692_n5849), .Y(_abc_17692_n5850) );
  OR2X2 OR2X2_1844 ( .A(sum_20_), .B(\key_in[84] ), .Y(_abc_17692_n5853) );
  OR2X2 OR2X2_1845 ( .A(_abc_17692_n5858), .B(_abc_17692_n5855), .Y(_abc_17692_n5859) );
  OR2X2 OR2X2_1846 ( .A(_abc_17692_n5860), .B(_abc_17692_n5795), .Y(_abc_17692_n5861) );
  OR2X2 OR2X2_1847 ( .A(_abc_17692_n5817), .B(_abc_17692_n5859), .Y(_abc_17692_n5862) );
  OR2X2 OR2X2_1848 ( .A(_abc_17692_n5863), .B(workunit2_20_), .Y(_abc_17692_n5866) );
  OR2X2 OR2X2_1849 ( .A(_abc_17692_n5869), .B(_abc_17692_n5422), .Y(_abc_17692_n5870) );
  OR2X2 OR2X2_185 ( .A(_abc_17692_n967_1), .B(_abc_17692_n959), .Y(sum_2__FF_INPUT) );
  OR2X2 OR2X2_1850 ( .A(_abc_17692_n5872), .B(_abc_17692_n5871), .Y(_abc_17692_n5873) );
  OR2X2 OR2X2_1851 ( .A(_abc_17692_n5880), .B(_abc_17692_n5867), .Y(_abc_17692_n5883) );
  OR2X2 OR2X2_1852 ( .A(_abc_17692_n5890), .B(_abc_17692_n5701), .Y(_abc_17692_n5891) );
  OR2X2 OR2X2_1853 ( .A(_abc_17692_n5889), .B(_abc_17692_n5891), .Y(_abc_17692_n5892) );
  OR2X2 OR2X2_1854 ( .A(_abc_17692_n5888), .B(_abc_17692_n5892), .Y(_abc_17692_n5893) );
  OR2X2 OR2X2_1855 ( .A(sum_20_), .B(\key_in[20] ), .Y(_abc_17692_n5896) );
  OR2X2 OR2X2_1856 ( .A(_abc_17692_n5053), .B(_abc_17692_n5899), .Y(_abc_17692_n5900_1) );
  OR2X2 OR2X2_1857 ( .A(_abc_17692_n5904), .B(_abc_17692_n5898), .Y(_abc_17692_n5905) );
  OR2X2 OR2X2_1858 ( .A(_abc_17692_n5906), .B(_abc_17692_n5795), .Y(_abc_17692_n5907) );
  OR2X2 OR2X2_1859 ( .A(_abc_17692_n5817), .B(_abc_17692_n5905), .Y(_abc_17692_n5908) );
  OR2X2 OR2X2_186 ( .A(_abc_17692_n962), .B(_abc_17692_n976), .Y(_abc_17692_n977) );
  OR2X2 OR2X2_1860 ( .A(_abc_17692_n5911), .B(_abc_17692_n5912), .Y(_abc_17692_n5913) );
  OR2X2 OR2X2_1861 ( .A(_abc_17692_n5915), .B(_abc_17692_n5494), .Y(_abc_17692_n5916) );
  OR2X2 OR2X2_1862 ( .A(_abc_17692_n5073), .B(_abc_17692_n5924), .Y(_abc_17692_n5925) );
  OR2X2 OR2X2_1863 ( .A(_abc_17692_n5926), .B(_abc_17692_n5913), .Y(_abc_17692_n5927) );
  OR2X2 OR2X2_1864 ( .A(_abc_17692_n5929), .B(_abc_17692_n5928), .Y(_abc_17692_n5930) );
  OR2X2 OR2X2_1865 ( .A(_abc_17692_n5937), .B(_abc_17692_n5673), .Y(_abc_17692_n5938) );
  OR2X2 OR2X2_1866 ( .A(_abc_17692_n5936), .B(_abc_17692_n5938), .Y(_abc_17692_n5939) );
  OR2X2 OR2X2_1867 ( .A(_abc_17692_n5935), .B(_abc_17692_n5939), .Y(_abc_17692_n5940) );
  OR2X2 OR2X2_1868 ( .A(sum_20_), .B(\key_in[52] ), .Y(_abc_17692_n5943) );
  OR2X2 OR2X2_1869 ( .A(_abc_17692_n5007), .B(_abc_17692_n5946), .Y(_abc_17692_n5947) );
  OR2X2 OR2X2_187 ( .A(_abc_17692_n977), .B(_abc_17692_n975), .Y(_abc_17692_n978) );
  OR2X2 OR2X2_1870 ( .A(_abc_17692_n5951), .B(_abc_17692_n5945), .Y(_abc_17692_n5952) );
  OR2X2 OR2X2_1871 ( .A(_abc_17692_n5953), .B(_abc_17692_n5795), .Y(_abc_17692_n5954) );
  OR2X2 OR2X2_1872 ( .A(_abc_17692_n5817), .B(_abc_17692_n5952), .Y(_abc_17692_n5955) );
  OR2X2 OR2X2_1873 ( .A(_abc_17692_n5958), .B(_abc_17692_n5959), .Y(_abc_17692_n5960) );
  OR2X2 OR2X2_1874 ( .A(_abc_17692_n5691), .B(_abc_17692_n5452), .Y(_abc_17692_n5961) );
  OR2X2 OR2X2_1875 ( .A(_abc_17692_n5961), .B(_abc_17692_n5457), .Y(_abc_17692_n5962) );
  OR2X2 OR2X2_1876 ( .A(_abc_17692_n5691), .B(_abc_17692_n5752), .Y(_abc_17692_n5965) );
  OR2X2 OR2X2_1877 ( .A(_abc_17692_n5027), .B(_abc_17692_n5970), .Y(_abc_17692_n5971) );
  OR2X2 OR2X2_1878 ( .A(_abc_17692_n5972), .B(_abc_17692_n5960), .Y(_abc_17692_n5973) );
  OR2X2 OR2X2_1879 ( .A(_abc_17692_n5975), .B(_abc_17692_n5974), .Y(_abc_17692_n5976) );
  OR2X2 OR2X2_188 ( .A(_abc_17692_n980_1), .B(_abc_17692_n979), .Y(_abc_17692_n981) );
  OR2X2 OR2X2_1880 ( .A(_abc_17692_n5978), .B(_abc_17692_n1863_bF_buf3), .Y(_abc_17692_n5979) );
  OR2X2 OR2X2_1881 ( .A(_abc_17692_n5979), .B(_abc_17692_n5932), .Y(_abc_17692_n5980) );
  OR2X2 OR2X2_1882 ( .A(_abc_17692_n5885), .B(_abc_17692_n5980), .Y(_abc_17692_n5981_1) );
  OR2X2 OR2X2_1883 ( .A(_abc_17692_n5658), .B(_abc_17692_n5661), .Y(_abc_17692_n5986) );
  OR2X2 OR2X2_1884 ( .A(_abc_17692_n5985), .B(_abc_17692_n5988), .Y(_abc_17692_n5989) );
  OR2X2 OR2X2_1885 ( .A(_abc_17692_n5991), .B(_abc_17692_n5989), .Y(_abc_17692_n5992) );
  OR2X2 OR2X2_1886 ( .A(_abc_17692_n5992), .B(_abc_17692_n5823), .Y(_abc_17692_n5993) );
  OR2X2 OR2X2_1887 ( .A(_abc_17692_n5999), .B(_abc_17692_n5262), .Y(_abc_17692_n6000) );
  OR2X2 OR2X2_1888 ( .A(_abc_17692_n5629), .B(_abc_17692_n5419), .Y(_abc_17692_n6001) );
  OR2X2 OR2X2_1889 ( .A(_abc_17692_n6001), .B(_abc_17692_n6000), .Y(_abc_17692_n6002) );
  OR2X2 OR2X2_189 ( .A(_abc_17692_n988_1), .B(_abc_17692_n979), .Y(_abc_17692_n989) );
  OR2X2 OR2X2_1890 ( .A(_abc_17692_n5628), .B(_abc_17692_n6004), .Y(_abc_17692_n6005) );
  OR2X2 OR2X2_1891 ( .A(_abc_17692_n5155), .B(_abc_17692_n6011), .Y(_abc_17692_n6012) );
  OR2X2 OR2X2_1892 ( .A(_abc_17692_n6014), .B(_abc_17692_n5998), .Y(_abc_17692_n6017) );
  OR2X2 OR2X2_1893 ( .A(_abc_17692_n6024), .B(_abc_17692_n6022), .Y(_abc_17692_n6025) );
  OR2X2 OR2X2_1894 ( .A(_abc_17692_n6021), .B(_abc_17692_n6025), .Y(_abc_17692_n6026) );
  OR2X2 OR2X2_1895 ( .A(_abc_17692_n6032), .B(_abc_17692_n5960), .Y(_abc_17692_n6033) );
  OR2X2 OR2X2_1896 ( .A(_abc_17692_n6042), .B(_abc_17692_n6040), .Y(_abc_17692_n6043) );
  OR2X2 OR2X2_1897 ( .A(_abc_17692_n6039), .B(_abc_17692_n6043), .Y(_abc_17692_n6044) );
  OR2X2 OR2X2_1898 ( .A(_abc_17692_n6046), .B(_abc_17692_n6044), .Y(_abc_17692_n6047) );
  OR2X2 OR2X2_1899 ( .A(_abc_17692_n6047), .B(_abc_17692_n5913), .Y(_abc_17692_n6050) );
  OR2X2 OR2X2_19 ( .A(state_8_bF_buf2), .B(delta_21_), .Y(delta_21__FF_INPUT) );
  OR2X2 OR2X2_190 ( .A(_abc_17692_n987), .B(_abc_17692_n975), .Y(_abc_17692_n990) );
  OR2X2 OR2X2_1900 ( .A(_abc_17692_n6037), .B(_abc_17692_n6052), .Y(_abc_17692_n6053) );
  OR2X2 OR2X2_1901 ( .A(_abc_17692_n6053), .B(_abc_17692_n6019), .Y(_abc_17692_n6054) );
  OR2X2 OR2X2_1902 ( .A(_abc_17692_n6054), .B(_abc_17692_n5997), .Y(_abc_17692_n6055) );
  OR2X2 OR2X2_1903 ( .A(_abc_17692_n6057), .B(_abc_17692_n6058), .Y(_abc_17692_n6059) );
  OR2X2 OR2X2_1904 ( .A(_abc_17692_n6056), .B(_abc_17692_n6059), .Y(_abc_17692_n6060) );
  OR2X2 OR2X2_1905 ( .A(_abc_17692_n6060), .B(_abc_17692_n5983), .Y(workunit2_20__FF_INPUT) );
  OR2X2 OR2X2_1906 ( .A(_abc_17692_n5790), .B(_abc_17692_n5786), .Y(_abc_17692_n6062) );
  OR2X2 OR2X2_1907 ( .A(_abc_17692_n4059), .B(workunit1_26_), .Y(_abc_17692_n6064) );
  OR2X2 OR2X2_1908 ( .A(_abc_17692_n6065), .B(workunit1_17_), .Y(_abc_17692_n6066) );
  OR2X2 OR2X2_1909 ( .A(_abc_17692_n6063), .B(_abc_17692_n6073), .Y(_abc_17692_n6076) );
  OR2X2 OR2X2_191 ( .A(_abc_17692_n992), .B(_abc_17692_n984), .Y(_abc_17692_n993) );
  OR2X2 OR2X2_1910 ( .A(_abc_17692_n5855), .B(_abc_17692_n5851), .Y(_abc_17692_n6078) );
  OR2X2 OR2X2_1911 ( .A(sum_21_), .B(\key_in[85] ), .Y(_abc_17692_n6082) );
  OR2X2 OR2X2_1912 ( .A(_abc_17692_n6084), .B(_abc_17692_n6086), .Y(_abc_17692_n6087) );
  OR2X2 OR2X2_1913 ( .A(_abc_17692_n6077), .B(_abc_17692_n6088), .Y(_abc_17692_n6089) );
  OR2X2 OR2X2_1914 ( .A(_abc_17692_n6090), .B(_abc_17692_n6074), .Y(_abc_17692_n6091) );
  OR2X2 OR2X2_1915 ( .A(_abc_17692_n6091), .B(_abc_17692_n6087), .Y(_abc_17692_n6092) );
  OR2X2 OR2X2_1916 ( .A(_abc_17692_n6097), .B(_abc_17692_n6094), .Y(_abc_17692_n6098) );
  OR2X2 OR2X2_1917 ( .A(_abc_17692_n6100), .B(_abc_17692_n6098), .Y(_abc_17692_n6101) );
  OR2X2 OR2X2_1918 ( .A(_abc_17692_n6099), .B(_abc_17692_n6102), .Y(_abc_17692_n6103) );
  OR2X2 OR2X2_1919 ( .A(_abc_17692_n5898), .B(_abc_17692_n5894), .Y(_abc_17692_n6106) );
  OR2X2 OR2X2_192 ( .A(_abc_17692_n993), .B(_abc_17692_n983), .Y(sum_3__FF_INPUT) );
  OR2X2 OR2X2_1920 ( .A(sum_21_), .B(\key_in[21] ), .Y(_abc_17692_n6109) );
  OR2X2 OR2X2_1921 ( .A(_abc_17692_n6106), .B(_abc_17692_n6111), .Y(_abc_17692_n6112) );
  OR2X2 OR2X2_1922 ( .A(_abc_17692_n6117), .B(_abc_17692_n6118), .Y(_abc_17692_n6119) );
  OR2X2 OR2X2_1923 ( .A(_abc_17692_n6121), .B(_abc_17692_n6122), .Y(_abc_17692_n6123) );
  OR2X2 OR2X2_1924 ( .A(_abc_17692_n6126), .B(_abc_17692_n6123), .Y(_abc_17692_n6127) );
  OR2X2 OR2X2_1925 ( .A(_abc_17692_n6125), .B(_abc_17692_n6130), .Y(_abc_17692_n6131) );
  OR2X2 OR2X2_1926 ( .A(_abc_17692_n5945), .B(_abc_17692_n5941), .Y(_abc_17692_n6134) );
  OR2X2 OR2X2_1927 ( .A(sum_21_), .B(\key_in[53] ), .Y(_abc_17692_n6138) );
  OR2X2 OR2X2_1928 ( .A(_abc_17692_n6135), .B(_abc_17692_n6139), .Y(_abc_17692_n6142) );
  OR2X2 OR2X2_1929 ( .A(_abc_17692_n6145), .B(_abc_17692_n6146), .Y(_abc_17692_n6147) );
  OR2X2 OR2X2_193 ( .A(_abc_17692_n995), .B(delta_4_), .Y(_abc_17692_n997) );
  OR2X2 OR2X2_1930 ( .A(_abc_17692_n6147), .B(_abc_17692_n6095), .Y(_abc_17692_n6148) );
  OR2X2 OR2X2_1931 ( .A(_abc_17692_n6077), .B(_abc_17692_n6143), .Y(_abc_17692_n6149) );
  OR2X2 OR2X2_1932 ( .A(_abc_17692_n6091), .B(_abc_17692_n6144), .Y(_abc_17692_n6150) );
  OR2X2 OR2X2_1933 ( .A(_abc_17692_n6151), .B(workunit2_21_), .Y(_abc_17692_n6152) );
  OR2X2 OR2X2_1934 ( .A(_abc_17692_n6157), .B(_abc_17692_n6154), .Y(_abc_17692_n6158) );
  OR2X2 OR2X2_1935 ( .A(_abc_17692_n6156), .B(_abc_17692_n6153), .Y(_abc_17692_n6159) );
  OR2X2 OR2X2_1936 ( .A(_abc_17692_n6161), .B(_abc_17692_n1863_bF_buf1), .Y(_abc_17692_n6162) );
  OR2X2 OR2X2_1937 ( .A(_abc_17692_n6162), .B(_abc_17692_n6133), .Y(_abc_17692_n6163) );
  OR2X2 OR2X2_1938 ( .A(_abc_17692_n6105), .B(_abc_17692_n6163), .Y(_abc_17692_n6164) );
  OR2X2 OR2X2_1939 ( .A(_abc_17692_n5808), .B(_abc_17692_n5804), .Y(_abc_17692_n6165) );
  OR2X2 OR2X2_194 ( .A(_abc_17692_n998), .B(_abc_17692_n996_1), .Y(_abc_17692_n999) );
  OR2X2 OR2X2_1940 ( .A(sum_21_), .B(\key_in[117] ), .Y(_abc_17692_n6168) );
  OR2X2 OR2X2_1941 ( .A(_abc_17692_n6165), .B(_abc_17692_n6170), .Y(_abc_17692_n6171) );
  OR2X2 OR2X2_1942 ( .A(_abc_17692_n6174), .B(_abc_17692_n6077), .Y(_abc_17692_n6175) );
  OR2X2 OR2X2_1943 ( .A(_abc_17692_n6176), .B(_abc_17692_n6091), .Y(_abc_17692_n6177) );
  OR2X2 OR2X2_1944 ( .A(_abc_17692_n6190), .B(_abc_17692_n4047_bF_buf4), .Y(_abc_17692_n6191) );
  OR2X2 OR2X2_1945 ( .A(_abc_17692_n6191), .B(_abc_17692_n6188), .Y(_abc_17692_n6192) );
  OR2X2 OR2X2_1946 ( .A(_abc_17692_n6197), .B(_abc_17692_n6189), .Y(_abc_17692_n6198) );
  OR2X2 OR2X2_1947 ( .A(_abc_17692_n6199), .B(_abc_17692_n6184), .Y(_abc_17692_n6200) );
  OR2X2 OR2X2_1948 ( .A(_abc_17692_n6206), .B(_abc_17692_n6098), .Y(_abc_17692_n6207) );
  OR2X2 OR2X2_1949 ( .A(_abc_17692_n6208), .B(_abc_17692_n6102), .Y(_abc_17692_n6209) );
  OR2X2 OR2X2_195 ( .A(_abc_17692_n987), .B(_abc_17692_n1002), .Y(_abc_17692_n1003) );
  OR2X2 OR2X2_1950 ( .A(_abc_17692_n6214), .B(_abc_17692_n6123), .Y(_abc_17692_n6215) );
  OR2X2 OR2X2_1951 ( .A(_abc_17692_n6216), .B(_abc_17692_n6130), .Y(_abc_17692_n6217) );
  OR2X2 OR2X2_1952 ( .A(_abc_17692_n6034), .B(_abc_17692_n6220), .Y(_abc_17692_n6221) );
  OR2X2 OR2X2_1953 ( .A(_abc_17692_n6221), .B(_abc_17692_n6153), .Y(_abc_17692_n6222_1) );
  OR2X2 OR2X2_1954 ( .A(_abc_17692_n6223), .B(_abc_17692_n6154), .Y(_abc_17692_n6224) );
  OR2X2 OR2X2_1955 ( .A(_abc_17692_n6219), .B(_abc_17692_n6226), .Y(_abc_17692_n6227) );
  OR2X2 OR2X2_1956 ( .A(_abc_17692_n6227), .B(_abc_17692_n6211), .Y(_abc_17692_n6228) );
  OR2X2 OR2X2_1957 ( .A(_abc_17692_n6228), .B(_abc_17692_n6202), .Y(_abc_17692_n6229) );
  OR2X2 OR2X2_1958 ( .A(_abc_17692_n6231), .B(_abc_17692_n6232), .Y(_abc_17692_n6233) );
  OR2X2 OR2X2_1959 ( .A(_abc_17692_n6230), .B(_abc_17692_n6233), .Y(_abc_17692_n6234) );
  OR2X2 OR2X2_196 ( .A(_abc_17692_n1005), .B(_abc_17692_n999), .Y(_abc_17692_n1006) );
  OR2X2 OR2X2_1960 ( .A(_abc_17692_n6234), .B(_abc_17692_n6194), .Y(workunit2_21__FF_INPUT) );
  OR2X2 OR2X2_1961 ( .A(_abc_17692_n6238), .B(_abc_17692_n6069), .Y(_abc_17692_n6239) );
  OR2X2 OR2X2_1962 ( .A(_abc_17692_n6237), .B(_abc_17692_n6239), .Y(_abc_17692_n6240) );
  OR2X2 OR2X2_1963 ( .A(_abc_17692_n4322), .B(workunit1_27_), .Y(_abc_17692_n6241) );
  OR2X2 OR2X2_1964 ( .A(_abc_17692_n6242), .B(workunit1_18_), .Y(_abc_17692_n6243) );
  OR2X2 OR2X2_1965 ( .A(_abc_17692_n6246), .B(_abc_17692_n6247), .Y(_abc_17692_n6248) );
  OR2X2 OR2X2_1966 ( .A(_abc_17692_n5793), .B(_abc_17692_n6251), .Y(_abc_17692_n6252) );
  OR2X2 OR2X2_1967 ( .A(_abc_17692_n6255), .B(_abc_17692_n6250), .Y(_abc_17692_n6256) );
  OR2X2 OR2X2_1968 ( .A(_abc_17692_n6261), .B(_abc_17692_n6260), .Y(_abc_17692_n6262) );
  OR2X2 OR2X2_1969 ( .A(sum_22_), .B(\key_in[86] ), .Y(_abc_17692_n6267) );
  OR2X2 OR2X2_197 ( .A(_abc_17692_n1004), .B(_abc_17692_n1007), .Y(_abc_17692_n1008) );
  OR2X2 OR2X2_1970 ( .A(_abc_17692_n6269), .B(_abc_17692_n6271), .Y(_abc_17692_n6272) );
  OR2X2 OR2X2_1971 ( .A(_abc_17692_n6273), .B(_abc_17692_n6256), .Y(_abc_17692_n6274) );
  OR2X2 OR2X2_1972 ( .A(_abc_17692_n6272), .B(_abc_17692_n6275), .Y(_abc_17692_n6276) );
  OR2X2 OR2X2_1973 ( .A(_abc_17692_n6277), .B(workunit2_22_), .Y(_abc_17692_n6280) );
  OR2X2 OR2X2_1974 ( .A(_abc_17692_n6283), .B(_abc_17692_n6282), .Y(_abc_17692_n6284) );
  OR2X2 OR2X2_1975 ( .A(_abc_17692_n6286), .B(_abc_17692_n6284), .Y(_abc_17692_n6287) );
  OR2X2 OR2X2_1976 ( .A(_abc_17692_n6287), .B(_abc_17692_n6281), .Y(_abc_17692_n6290) );
  OR2X2 OR2X2_1977 ( .A(_abc_17692_n6297), .B(_abc_17692_n6296), .Y(_abc_17692_n6298) );
  OR2X2 OR2X2_1978 ( .A(_abc_17692_n6295), .B(_abc_17692_n6299), .Y(_abc_17692_n6300) );
  OR2X2 OR2X2_1979 ( .A(sum_22_), .B(\key_in[22] ), .Y(_abc_17692_n6303) );
  OR2X2 OR2X2_198 ( .A(_abc_17692_n1012), .B(_abc_17692_n973), .Y(_abc_17692_n1013) );
  OR2X2 OR2X2_1980 ( .A(_abc_17692_n5902), .B(_abc_17692_n6306), .Y(_abc_17692_n6307) );
  OR2X2 OR2X2_1981 ( .A(_abc_17692_n6310), .B(_abc_17692_n6305), .Y(_abc_17692_n6311) );
  OR2X2 OR2X2_1982 ( .A(_abc_17692_n6312), .B(_abc_17692_n6314), .Y(_abc_17692_n6315) );
  OR2X2 OR2X2_1983 ( .A(_abc_17692_n6316_1), .B(_abc_17692_n6293), .Y(_abc_17692_n6317) );
  OR2X2 OR2X2_1984 ( .A(_abc_17692_n6315), .B(workunit2_22_), .Y(_abc_17692_n6318) );
  OR2X2 OR2X2_1985 ( .A(_abc_17692_n6322), .B(_abc_17692_n6321), .Y(_abc_17692_n6323) );
  OR2X2 OR2X2_1986 ( .A(_abc_17692_n6325), .B(_abc_17692_n6323), .Y(_abc_17692_n6326) );
  OR2X2 OR2X2_1987 ( .A(_abc_17692_n6326), .B(_abc_17692_n6320), .Y(_abc_17692_n6329) );
  OR2X2 OR2X2_1988 ( .A(_abc_17692_n6335), .B(_abc_17692_n6334), .Y(_abc_17692_n6336) );
  OR2X2 OR2X2_1989 ( .A(_abc_17692_n6333), .B(_abc_17692_n6337), .Y(_abc_17692_n6338) );
  OR2X2 OR2X2_199 ( .A(_abc_17692_n1013), .B(_abc_17692_n1007), .Y(_abc_17692_n1016) );
  OR2X2 OR2X2_1990 ( .A(sum_22_), .B(\key_in[54] ), .Y(_abc_17692_n6341) );
  OR2X2 OR2X2_1991 ( .A(_abc_17692_n5949), .B(_abc_17692_n6344), .Y(_abc_17692_n6345) );
  OR2X2 OR2X2_1992 ( .A(_abc_17692_n6348), .B(_abc_17692_n6343), .Y(_abc_17692_n6349) );
  OR2X2 OR2X2_1993 ( .A(_abc_17692_n6350), .B(_abc_17692_n6256), .Y(_abc_17692_n6351) );
  OR2X2 OR2X2_1994 ( .A(_abc_17692_n6275), .B(_abc_17692_n6349), .Y(_abc_17692_n6352) );
  OR2X2 OR2X2_1995 ( .A(_abc_17692_n6355), .B(_abc_17692_n6356), .Y(_abc_17692_n6357) );
  OR2X2 OR2X2_1996 ( .A(_abc_17692_n6153), .B(_abc_17692_n6155), .Y(_abc_17692_n6361) );
  OR2X2 OR2X2_1997 ( .A(_abc_17692_n6153), .B(_abc_17692_n5960), .Y(_abc_17692_n6363) );
  OR2X2 OR2X2_1998 ( .A(_abc_17692_n5972), .B(_abc_17692_n6363), .Y(_abc_17692_n6364) );
  OR2X2 OR2X2_1999 ( .A(_abc_17692_n6366), .B(_abc_17692_n6358), .Y(_abc_17692_n6367) );
  OR2X2 OR2X2_2 ( .A(_abc_17692_n629), .B(state_8_bF_buf9), .Y(_abc_10892_n1125) );
  OR2X2 OR2X2_20 ( .A(state_8_bF_buf1), .B(delta_25_), .Y(delta_25__FF_INPUT) );
  OR2X2 OR2X2_200 ( .A(_abc_17692_n1018), .B(_abc_17692_n1011), .Y(_abc_17692_n1019) );
  OR2X2 OR2X2_2000 ( .A(_abc_17692_n6365), .B(_abc_17692_n6357), .Y(_abc_17692_n6368) );
  OR2X2 OR2X2_2001 ( .A(_abc_17692_n6331), .B(_abc_17692_n6370), .Y(_abc_17692_n6371_1) );
  OR2X2 OR2X2_2002 ( .A(_abc_17692_n6292), .B(_abc_17692_n6371_1), .Y(_abc_17692_n6372) );
  OR2X2 OR2X2_2003 ( .A(_abc_17692_n6376), .B(_abc_17692_n6375), .Y(_abc_17692_n6377) );
  OR2X2 OR2X2_2004 ( .A(_abc_17692_n6374_1), .B(_abc_17692_n6378), .Y(_abc_17692_n6379) );
  OR2X2 OR2X2_2005 ( .A(sum_22_), .B(\key_in[118] ), .Y(_abc_17692_n6382) );
  OR2X2 OR2X2_2006 ( .A(_abc_17692_n6388), .B(_abc_17692_n6384), .Y(_abc_17692_n6389) );
  OR2X2 OR2X2_2007 ( .A(_abc_17692_n6392), .B(_abc_17692_n6390), .Y(_abc_17692_n6393) );
  OR2X2 OR2X2_2008 ( .A(_abc_17692_n6394), .B(_abc_17692_n6293), .Y(_abc_17692_n6395) );
  OR2X2 OR2X2_2009 ( .A(_abc_17692_n6393), .B(workunit2_22_), .Y(_abc_17692_n6396) );
  OR2X2 OR2X2_201 ( .A(_abc_17692_n1019), .B(_abc_17692_n1010), .Y(sum_4__FF_INPUT) );
  OR2X2 OR2X2_2010 ( .A(_abc_17692_n6400), .B(_abc_17692_n6399), .Y(_abc_17692_n6401) );
  OR2X2 OR2X2_2011 ( .A(_abc_17692_n6403), .B(_abc_17692_n6401), .Y(_abc_17692_n6404) );
  OR2X2 OR2X2_2012 ( .A(_abc_17692_n6404), .B(_abc_17692_n6398), .Y(_abc_17692_n6407) );
  OR2X2 OR2X2_2013 ( .A(_abc_17692_n6372), .B(_abc_17692_n6409), .Y(_abc_17692_n6410) );
  OR2X2 OR2X2_2014 ( .A(_abc_17692_n6413), .B(_abc_17692_n6182), .Y(_abc_17692_n6414) );
  OR2X2 OR2X2_2015 ( .A(_abc_17692_n6414), .B(_abc_17692_n6398), .Y(_abc_17692_n6415) );
  OR2X2 OR2X2_2016 ( .A(_abc_17692_n6416), .B(_abc_17692_n6397), .Y(_abc_17692_n6417) );
  OR2X2 OR2X2_2017 ( .A(_abc_17692_n6098), .B(_abc_17692_n5867), .Y(_abc_17692_n6421) );
  OR2X2 OR2X2_2018 ( .A(_abc_17692_n6425), .B(_abc_17692_n6097), .Y(_abc_17692_n6426) );
  OR2X2 OR2X2_2019 ( .A(_abc_17692_n6423), .B(_abc_17692_n6427), .Y(_abc_17692_n6428) );
  OR2X2 OR2X2_202 ( .A(_abc_17692_n1031), .B(_abc_17692_n1028_1), .Y(_abc_17692_n1032) );
  OR2X2 OR2X2_2020 ( .A(_abc_17692_n6428), .B(_abc_17692_n6420), .Y(_abc_17692_n6431) );
  OR2X2 OR2X2_2021 ( .A(_abc_17692_n6434), .B(_abc_17692_n6220), .Y(_abc_17692_n6435) );
  OR2X2 OR2X2_2022 ( .A(_abc_17692_n6031), .B(_abc_17692_n6439), .Y(_abc_17692_n6440) );
  OR2X2 OR2X2_2023 ( .A(_abc_17692_n6441), .B(_abc_17692_n6358), .Y(_abc_17692_n6442) );
  OR2X2 OR2X2_2024 ( .A(_abc_17692_n6443), .B(_abc_17692_n6357), .Y(_abc_17692_n6444) );
  OR2X2 OR2X2_2025 ( .A(_abc_17692_n6121), .B(_abc_17692_n6212), .Y(_abc_17692_n6447) );
  OR2X2 OR2X2_2026 ( .A(_abc_17692_n6450), .B(_abc_17692_n6448), .Y(_abc_17692_n6451) );
  OR2X2 OR2X2_2027 ( .A(_abc_17692_n6451), .B(_abc_17692_n6319_1), .Y(_abc_17692_n6454) );
  OR2X2 OR2X2_2028 ( .A(_abc_17692_n6446), .B(_abc_17692_n6456), .Y(_abc_17692_n6457) );
  OR2X2 OR2X2_2029 ( .A(_abc_17692_n6457), .B(_abc_17692_n6433), .Y(_abc_17692_n6458) );
  OR2X2 OR2X2_203 ( .A(_abc_17692_n1033), .B(_abc_17692_n1027), .Y(_abc_17692_n1034) );
  OR2X2 OR2X2_2030 ( .A(_abc_17692_n6419), .B(_abc_17692_n6458), .Y(_abc_17692_n6459) );
  OR2X2 OR2X2_2031 ( .A(_abc_17692_n6461), .B(_abc_17692_n6462), .Y(_abc_17692_n6463) );
  OR2X2 OR2X2_2032 ( .A(_abc_17692_n6460), .B(_abc_17692_n6463), .Y(_abc_17692_n6464) );
  OR2X2 OR2X2_2033 ( .A(_abc_17692_n6464), .B(_abc_17692_n6411), .Y(workunit2_22__FF_INPUT) );
  OR2X2 OR2X2_2034 ( .A(_abc_17692_n6250), .B(_abc_17692_n6246), .Y(_abc_17692_n6466) );
  OR2X2 OR2X2_2035 ( .A(_abc_17692_n4494), .B(workunit1_28_), .Y(_abc_17692_n6467) );
  OR2X2 OR2X2_2036 ( .A(_abc_17692_n6468_1), .B(workunit1_19_), .Y(_abc_17692_n6469) );
  OR2X2 OR2X2_2037 ( .A(_abc_17692_n6466), .B(_abc_17692_n6477), .Y(_abc_17692_n6478) );
  OR2X2 OR2X2_2038 ( .A(_abc_17692_n6254), .B(_abc_17692_n6248), .Y(_abc_17692_n6480) );
  OR2X2 OR2X2_2039 ( .A(_abc_17692_n6481), .B(_abc_17692_n6476), .Y(_abc_17692_n6482) );
  OR2X2 OR2X2_204 ( .A(_abc_17692_n1014), .B(_abc_17692_n998), .Y(_abc_17692_n1037) );
  OR2X2 OR2X2_2040 ( .A(_abc_17692_n6263), .B(_abc_17692_n6270), .Y(_abc_17692_n6484) );
  OR2X2 OR2X2_2041 ( .A(sum_23_), .B(\key_in[87] ), .Y(_abc_17692_n6488) );
  OR2X2 OR2X2_2042 ( .A(_abc_17692_n6485), .B(_abc_17692_n6489), .Y(_abc_17692_n6492) );
  OR2X2 OR2X2_2043 ( .A(_abc_17692_n6493), .B(_abc_17692_n6483), .Y(_abc_17692_n6494) );
  OR2X2 OR2X2_2044 ( .A(_abc_17692_n6495), .B(_abc_17692_n6496), .Y(_abc_17692_n6497) );
  OR2X2 OR2X2_2045 ( .A(_abc_17692_n6500), .B(_abc_17692_n6490), .Y(_abc_17692_n6501) );
  OR2X2 OR2X2_2046 ( .A(_abc_17692_n6501), .B(_abc_17692_n6497), .Y(_abc_17692_n6502) );
  OR2X2 OR2X2_2047 ( .A(_abc_17692_n6501), .B(_abc_17692_n6483), .Y(_abc_17692_n6506) );
  OR2X2 OR2X2_2048 ( .A(_abc_17692_n6493), .B(_abc_17692_n6497), .Y(_abc_17692_n6507) );
  OR2X2 OR2X2_2049 ( .A(_abc_17692_n6504), .B(_abc_17692_n6509), .Y(_abc_17692_n6510) );
  OR2X2 OR2X2_205 ( .A(_abc_17692_n1037), .B(_abc_17692_n1028_1), .Y(_abc_17692_n1038) );
  OR2X2 OR2X2_2050 ( .A(_abc_17692_n6512), .B(_abc_17692_n6510), .Y(_abc_17692_n6513) );
  OR2X2 OR2X2_2051 ( .A(_abc_17692_n6511), .B(_abc_17692_n6514), .Y(_abc_17692_n6515) );
  OR2X2 OR2X2_2052 ( .A(_abc_17692_n6346), .B(_abc_17692_n6347), .Y(_abc_17692_n6518) );
  OR2X2 OR2X2_2053 ( .A(sum_23_), .B(\key_in[55] ), .Y(_abc_17692_n6522) );
  OR2X2 OR2X2_2054 ( .A(_abc_17692_n6343), .B(_abc_17692_n6339), .Y(_abc_17692_n6525) );
  OR2X2 OR2X2_2055 ( .A(_abc_17692_n6524), .B(_abc_17692_n6527), .Y(_abc_17692_n6528) );
  OR2X2 OR2X2_2056 ( .A(_abc_17692_n6483), .B(_abc_17692_n6528), .Y(_abc_17692_n6529) );
  OR2X2 OR2X2_2057 ( .A(_abc_17692_n6525), .B(_abc_17692_n6526_1), .Y(_abc_17692_n6530) );
  OR2X2 OR2X2_2058 ( .A(_abc_17692_n6519), .B(_abc_17692_n6523_1), .Y(_abc_17692_n6531) );
  OR2X2 OR2X2_2059 ( .A(_abc_17692_n6497), .B(_abc_17692_n6532), .Y(_abc_17692_n6533) );
  OR2X2 OR2X2_206 ( .A(_abc_17692_n1043), .B(state_8_bF_buf6), .Y(_abc_17692_n1044) );
  OR2X2 OR2X2_2060 ( .A(_abc_17692_n6534), .B(_abc_17692_n6505), .Y(_abc_17692_n6535) );
  OR2X2 OR2X2_2061 ( .A(_abc_17692_n6483), .B(_abc_17692_n6532), .Y(_abc_17692_n6536) );
  OR2X2 OR2X2_2062 ( .A(_abc_17692_n6497), .B(_abc_17692_n6528), .Y(_abc_17692_n6537) );
  OR2X2 OR2X2_2063 ( .A(_abc_17692_n6538), .B(workunit2_23_), .Y(_abc_17692_n6539) );
  OR2X2 OR2X2_2064 ( .A(_abc_17692_n6544), .B(_abc_17692_n6541), .Y(_abc_17692_n6545) );
  OR2X2 OR2X2_2065 ( .A(_abc_17692_n6543), .B(_abc_17692_n6540), .Y(_abc_17692_n6546) );
  OR2X2 OR2X2_2066 ( .A(_abc_17692_n6308), .B(_abc_17692_n6309), .Y(_abc_17692_n6549) );
  OR2X2 OR2X2_2067 ( .A(sum_23_), .B(\key_in[23] ), .Y(_abc_17692_n6553) );
  OR2X2 OR2X2_2068 ( .A(_abc_17692_n6305), .B(_abc_17692_n6301), .Y(_abc_17692_n6556) );
  OR2X2 OR2X2_2069 ( .A(_abc_17692_n6555), .B(_abc_17692_n6558), .Y(_abc_17692_n6559) );
  OR2X2 OR2X2_207 ( .A(_abc_17692_n1042), .B(_abc_17692_n1044), .Y(_abc_17692_n1045) );
  OR2X2 OR2X2_2070 ( .A(_abc_17692_n6483), .B(_abc_17692_n6559), .Y(_abc_17692_n6560) );
  OR2X2 OR2X2_2071 ( .A(_abc_17692_n6556), .B(_abc_17692_n6557), .Y(_abc_17692_n6561) );
  OR2X2 OR2X2_2072 ( .A(_abc_17692_n6550), .B(_abc_17692_n6554), .Y(_abc_17692_n6562) );
  OR2X2 OR2X2_2073 ( .A(_abc_17692_n6497), .B(_abc_17692_n6563), .Y(_abc_17692_n6564) );
  OR2X2 OR2X2_2074 ( .A(_abc_17692_n6565), .B(_abc_17692_n6505), .Y(_abc_17692_n6566) );
  OR2X2 OR2X2_2075 ( .A(_abc_17692_n6483), .B(_abc_17692_n6563), .Y(_abc_17692_n6567) );
  OR2X2 OR2X2_2076 ( .A(_abc_17692_n6497), .B(_abc_17692_n6559), .Y(_abc_17692_n6568) );
  OR2X2 OR2X2_2077 ( .A(_abc_17692_n6569), .B(workunit2_23_), .Y(_abc_17692_n6570) );
  OR2X2 OR2X2_2078 ( .A(_abc_17692_n6576), .B(_abc_17692_n6572), .Y(_abc_17692_n6577) );
  OR2X2 OR2X2_2079 ( .A(_abc_17692_n6575), .B(_abc_17692_n6571), .Y(_abc_17692_n6578) );
  OR2X2 OR2X2_208 ( .A(_abc_17692_n1045), .B(_abc_17692_n1036), .Y(sum_5__FF_INPUT) );
  OR2X2 OR2X2_2080 ( .A(_abc_17692_n6580), .B(_abc_17692_n6548), .Y(_abc_17692_n6581) );
  OR2X2 OR2X2_2081 ( .A(_abc_17692_n6517), .B(_abc_17692_n6581), .Y(_abc_17692_n6582) );
  OR2X2 OR2X2_2082 ( .A(_abc_17692_n6384), .B(_abc_17692_n6380), .Y(_abc_17692_n6583) );
  OR2X2 OR2X2_2083 ( .A(sum_23_), .B(\key_in[119] ), .Y(_abc_17692_n6586) );
  OR2X2 OR2X2_2084 ( .A(_abc_17692_n6583), .B(_abc_17692_n6588), .Y(_abc_17692_n6589) );
  OR2X2 OR2X2_2085 ( .A(_abc_17692_n6592), .B(_abc_17692_n6483), .Y(_abc_17692_n6593) );
  OR2X2 OR2X2_2086 ( .A(_abc_17692_n6596), .B(_abc_17692_n6590), .Y(_abc_17692_n6597_1) );
  OR2X2 OR2X2_2087 ( .A(_abc_17692_n6597_1), .B(_abc_17692_n6497), .Y(_abc_17692_n6598) );
  OR2X2 OR2X2_2088 ( .A(_abc_17692_n6597_1), .B(_abc_17692_n6483), .Y(_abc_17692_n6601) );
  OR2X2 OR2X2_2089 ( .A(_abc_17692_n6592), .B(_abc_17692_n6497), .Y(_abc_17692_n6602) );
  OR2X2 OR2X2_209 ( .A(_abc_17692_n1047), .B(delta_6_), .Y(_abc_17692_n1049) );
  OR2X2 OR2X2_2090 ( .A(_abc_17692_n6600_1), .B(_abc_17692_n6604), .Y(_abc_17692_n6605) );
  OR2X2 OR2X2_2091 ( .A(_abc_17692_n6393), .B(_abc_17692_n6293), .Y(_abc_17692_n6606) );
  OR2X2 OR2X2_2092 ( .A(_abc_17692_n6405), .B(_abc_17692_n6607), .Y(_abc_17692_n6608) );
  OR2X2 OR2X2_2093 ( .A(_abc_17692_n6603), .B(_abc_17692_n6505), .Y(_abc_17692_n6611) );
  OR2X2 OR2X2_2094 ( .A(_abc_17692_n6599), .B(workunit2_23_), .Y(_abc_17692_n6612) );
  OR2X2 OR2X2_2095 ( .A(_abc_17692_n6610), .B(_abc_17692_n6614), .Y(_abc_17692_n6615) );
  OR2X2 OR2X2_2096 ( .A(_abc_17692_n6582), .B(_abc_17692_n6616), .Y(_abc_17692_n6617) );
  OR2X2 OR2X2_2097 ( .A(_abc_17692_n6620), .B(_abc_17692_n6613), .Y(_abc_17692_n6621) );
  OR2X2 OR2X2_2098 ( .A(_abc_17692_n6619), .B(_abc_17692_n6605), .Y(_abc_17692_n6622) );
  OR2X2 OR2X2_2099 ( .A(_abc_17692_n6429), .B(_abc_17692_n6626), .Y(_abc_17692_n6627) );
  OR2X2 OR2X2_21 ( .A(state_8_bF_buf0), .B(delta_26_), .Y(delta_26__FF_INPUT) );
  OR2X2 OR2X2_210 ( .A(_abc_17692_n1050), .B(_abc_17692_n1048), .Y(_abc_17692_n1051) );
  OR2X2 OR2X2_2100 ( .A(_abc_17692_n6630), .B(_abc_17692_n6628), .Y(_abc_17692_n6631) );
  OR2X2 OR2X2_2101 ( .A(_abc_17692_n6636), .B(_abc_17692_n6540), .Y(_abc_17692_n6637) );
  OR2X2 OR2X2_2102 ( .A(_abc_17692_n6635), .B(_abc_17692_n6541), .Y(_abc_17692_n6638) );
  OR2X2 OR2X2_2103 ( .A(_abc_17692_n6452), .B(_abc_17692_n6641), .Y(_abc_17692_n6642) );
  OR2X2 OR2X2_2104 ( .A(_abc_17692_n6643), .B(_abc_17692_n6572), .Y(_abc_17692_n6644_1) );
  OR2X2 OR2X2_2105 ( .A(_abc_17692_n6642), .B(_abc_17692_n6571), .Y(_abc_17692_n6645) );
  OR2X2 OR2X2_2106 ( .A(_abc_17692_n6647_1), .B(_abc_17692_n6640), .Y(_abc_17692_n6648) );
  OR2X2 OR2X2_2107 ( .A(_abc_17692_n6632), .B(_abc_17692_n6648), .Y(_abc_17692_n6649) );
  OR2X2 OR2X2_2108 ( .A(_abc_17692_n6624), .B(_abc_17692_n6649), .Y(_abc_17692_n6650) );
  OR2X2 OR2X2_2109 ( .A(_abc_17692_n6652_1), .B(_abc_17692_n6653), .Y(_abc_17692_n6654_1) );
  OR2X2 OR2X2_211 ( .A(_abc_17692_n1039), .B(_abc_17692_n1053), .Y(_abc_17692_n1054) );
  OR2X2 OR2X2_2110 ( .A(_abc_17692_n6651), .B(_abc_17692_n6654_1), .Y(_abc_17692_n6655) );
  OR2X2 OR2X2_2111 ( .A(_abc_17692_n6655), .B(_abc_17692_n6618), .Y(workunit2_23__FF_INPUT) );
  OR2X2 OR2X2_2112 ( .A(_abc_17692_n4730), .B(workunit1_29_), .Y(_abc_17692_n6658_1) );
  OR2X2 OR2X2_2113 ( .A(_abc_17692_n6659_1), .B(workunit1_20_), .Y(_abc_17692_n6660_1) );
  OR2X2 OR2X2_2114 ( .A(_abc_17692_n6663), .B(_abc_17692_n6664), .Y(_abc_17692_n6665) );
  OR2X2 OR2X2_2115 ( .A(_abc_17692_n6667), .B(_abc_17692_n6474), .Y(_abc_17692_n6668) );
  OR2X2 OR2X2_2116 ( .A(_abc_17692_n6669), .B(_abc_17692_n6670), .Y(_abc_17692_n6671) );
  OR2X2 OR2X2_2117 ( .A(_abc_17692_n6237), .B(_abc_17692_n6673), .Y(_abc_17692_n6674) );
  OR2X2 OR2X2_2118 ( .A(_abc_17692_n6678), .B(_abc_17692_n6677), .Y(_abc_17692_n6679) );
  OR2X2 OR2X2_2119 ( .A(_abc_17692_n6680), .B(_abc_17692_n6676), .Y(_abc_17692_n6681) );
  OR2X2 OR2X2_212 ( .A(_abc_17692_n1054), .B(_abc_17692_n1052), .Y(_abc_17692_n1055) );
  OR2X2 OR2X2_2120 ( .A(sum_24_), .B(\key_in[120] ), .Y(_abc_17692_n6684) );
  OR2X2 OR2X2_2121 ( .A(_abc_17692_n6686), .B(_abc_17692_n6584), .Y(_abc_17692_n6687) );
  OR2X2 OR2X2_2122 ( .A(_abc_17692_n6374_1), .B(_abc_17692_n6690), .Y(_abc_17692_n6691) );
  OR2X2 OR2X2_2123 ( .A(_abc_17692_n6692), .B(_abc_17692_n6687), .Y(_abc_17692_n6693) );
  OR2X2 OR2X2_2124 ( .A(_abc_17692_n6698), .B(_abc_17692_n6695), .Y(_abc_17692_n6699) );
  OR2X2 OR2X2_2125 ( .A(_abc_17692_n6700), .B(_abc_17692_n6681), .Y(_abc_17692_n6701) );
  OR2X2 OR2X2_2126 ( .A(_abc_17692_n6699), .B(_abc_17692_n6702), .Y(_abc_17692_n6703) );
  OR2X2 OR2X2_2127 ( .A(_abc_17692_n6706), .B(_abc_17692_n6707), .Y(_abc_17692_n6708) );
  OR2X2 OR2X2_2128 ( .A(_abc_17692_n6713), .B(_abc_17692_n6712), .Y(_abc_17692_n6714) );
  OR2X2 OR2X2_2129 ( .A(_abc_17692_n6711), .B(_abc_17692_n6714), .Y(_abc_17692_n6715) );
  OR2X2 OR2X2_213 ( .A(_abc_17692_n1031), .B(_abc_17692_n1025_1), .Y(_abc_17692_n1061) );
  OR2X2 OR2X2_2130 ( .A(_abc_17692_n5836), .B(_abc_17692_n6718), .Y(_abc_17692_n6719) );
  OR2X2 OR2X2_2131 ( .A(_abc_17692_n6721), .B(_abc_17692_n6709), .Y(_abc_17692_n6724) );
  OR2X2 OR2X2_2132 ( .A(_abc_17692_n6725), .B(_abc_17692_n4047_bF_buf3), .Y(_abc_17692_n6726) );
  OR2X2 OR2X2_2133 ( .A(sum_24_), .B(\key_in[24] ), .Y(_abc_17692_n6729) );
  OR2X2 OR2X2_2134 ( .A(_abc_17692_n6731), .B(_abc_17692_n6551), .Y(_abc_17692_n6732) );
  OR2X2 OR2X2_2135 ( .A(_abc_17692_n6295), .B(_abc_17692_n6735), .Y(_abc_17692_n6736) );
  OR2X2 OR2X2_2136 ( .A(_abc_17692_n6737), .B(_abc_17692_n6732), .Y(_abc_17692_n6738) );
  OR2X2 OR2X2_2137 ( .A(_abc_17692_n6742), .B(_abc_17692_n6743), .Y(_abc_17692_n6744) );
  OR2X2 OR2X2_2138 ( .A(_abc_17692_n6745), .B(_abc_17692_n6740), .Y(_abc_17692_n6746) );
  OR2X2 OR2X2_2139 ( .A(_abc_17692_n6747), .B(_abc_17692_n6681), .Y(_abc_17692_n6748) );
  OR2X2 OR2X2_214 ( .A(_abc_17692_n1062), .B(_abc_17692_n1052), .Y(_abc_17692_n1063) );
  OR2X2 OR2X2_2140 ( .A(_abc_17692_n6702), .B(_abc_17692_n6746), .Y(_abc_17692_n6749) );
  OR2X2 OR2X2_2141 ( .A(_abc_17692_n6752), .B(_abc_17692_n6753), .Y(_abc_17692_n6754) );
  OR2X2 OR2X2_2142 ( .A(_abc_17692_n5925), .B(_abc_17692_n6758), .Y(_abc_17692_n6759) );
  OR2X2 OR2X2_2143 ( .A(_abc_17692_n5922), .B(_abc_17692_n6758), .Y(_abc_17692_n6760) );
  OR2X2 OR2X2_2144 ( .A(_abc_17692_n6763), .B(_abc_17692_n6762), .Y(_abc_17692_n6764) );
  OR2X2 OR2X2_2145 ( .A(_abc_17692_n6761), .B(_abc_17692_n6764), .Y(_abc_17692_n6765) );
  OR2X2 OR2X2_2146 ( .A(_abc_17692_n6769), .B(_abc_17692_n6755), .Y(_abc_17692_n6770) );
  OR2X2 OR2X2_2147 ( .A(sum_24_), .B(\key_in[88] ), .Y(_abc_17692_n6777) );
  OR2X2 OR2X2_2148 ( .A(_abc_17692_n6779), .B(_abc_17692_n6486), .Y(_abc_17692_n6780) );
  OR2X2 OR2X2_2149 ( .A(_abc_17692_n6784), .B(_abc_17692_n6780), .Y(_abc_17692_n6785) );
  OR2X2 OR2X2_215 ( .A(_abc_17692_n1064), .B(_abc_17692_n1051), .Y(_abc_17692_n1065) );
  OR2X2 OR2X2_2150 ( .A(_abc_17692_n6783), .B(_abc_17692_n6786), .Y(_abc_17692_n6787) );
  OR2X2 OR2X2_2151 ( .A(_abc_17692_n6789), .B(_abc_17692_n6791), .Y(_abc_17692_n6792) );
  OR2X2 OR2X2_2152 ( .A(_abc_17692_n6793), .B(_abc_17692_n6681), .Y(_abc_17692_n6794) );
  OR2X2 OR2X2_2153 ( .A(_abc_17692_n6792), .B(_abc_17692_n6702), .Y(_abc_17692_n6795) );
  OR2X2 OR2X2_2154 ( .A(_abc_17692_n6798), .B(_abc_17692_n6799), .Y(_abc_17692_n6800) );
  OR2X2 OR2X2_2155 ( .A(_abc_17692_n5875), .B(_abc_17692_n6804), .Y(_abc_17692_n6805) );
  OR2X2 OR2X2_2156 ( .A(_abc_17692_n6809), .B(_abc_17692_n6808), .Y(_abc_17692_n6810) );
  OR2X2 OR2X2_2157 ( .A(_abc_17692_n6814), .B(_abc_17692_n6803), .Y(_abc_17692_n6815) );
  OR2X2 OR2X2_2158 ( .A(_abc_17692_n6815), .B(_abc_17692_n6800), .Y(_abc_17692_n6818) );
  OR2X2 OR2X2_2159 ( .A(sum_24_), .B(\key_in[56] ), .Y(_abc_17692_n6823) );
  OR2X2 OR2X2_216 ( .A(_abc_17692_n1067), .B(_abc_17692_n1060), .Y(_abc_17692_n1068) );
  OR2X2 OR2X2_2160 ( .A(_abc_17692_n6825), .B(_abc_17692_n6520), .Y(_abc_17692_n6826) );
  OR2X2 OR2X2_2161 ( .A(_abc_17692_n6333), .B(_abc_17692_n6829), .Y(_abc_17692_n6830) );
  OR2X2 OR2X2_2162 ( .A(_abc_17692_n6831), .B(_abc_17692_n6826), .Y(_abc_17692_n6832) );
  OR2X2 OR2X2_2163 ( .A(_abc_17692_n6836), .B(_abc_17692_n6837), .Y(_abc_17692_n6838) );
  OR2X2 OR2X2_2164 ( .A(_abc_17692_n6839), .B(_abc_17692_n6834), .Y(_abc_17692_n6840) );
  OR2X2 OR2X2_2165 ( .A(_abc_17692_n6841), .B(_abc_17692_n6681), .Y(_abc_17692_n6842) );
  OR2X2 OR2X2_2166 ( .A(_abc_17692_n6702), .B(_abc_17692_n6840), .Y(_abc_17692_n6843) );
  OR2X2 OR2X2_2167 ( .A(_abc_17692_n6846), .B(_abc_17692_n6847), .Y(_abc_17692_n6848) );
  OR2X2 OR2X2_2168 ( .A(_abc_17692_n6540), .B(_abc_17692_n6357), .Y(_abc_17692_n6850) );
  OR2X2 OR2X2_2169 ( .A(_abc_17692_n6850), .B(_abc_17692_n6363), .Y(_abc_17692_n6851) );
  OR2X2 OR2X2_217 ( .A(_abc_17692_n1068), .B(_abc_17692_n1059), .Y(sum_6__FF_INPUT) );
  OR2X2 OR2X2_2170 ( .A(_abc_17692_n5971), .B(_abc_17692_n6851), .Y(_abc_17692_n6852) );
  OR2X2 OR2X2_2171 ( .A(_abc_17692_n6851), .B(_abc_17692_n5967), .Y(_abc_17692_n6853) );
  OR2X2 OR2X2_2172 ( .A(_abc_17692_n6362), .B(_abc_17692_n6850), .Y(_abc_17692_n6854) );
  OR2X2 OR2X2_2173 ( .A(_abc_17692_n6540), .B(_abc_17692_n6542), .Y(_abc_17692_n6857) );
  OR2X2 OR2X2_2174 ( .A(_abc_17692_n6862), .B(_abc_17692_n6849), .Y(_abc_17692_n6865) );
  OR2X2 OR2X2_2175 ( .A(_abc_17692_n6867), .B(_abc_17692_n1863_bF_buf6), .Y(_abc_17692_n6868) );
  OR2X2 OR2X2_2176 ( .A(_abc_17692_n6820), .B(_abc_17692_n6868), .Y(_abc_17692_n6869) );
  OR2X2 OR2X2_2177 ( .A(_abc_17692_n6869), .B(_abc_17692_n6774), .Y(_abc_17692_n6870) );
  OR2X2 OR2X2_2178 ( .A(_abc_17692_n6880), .B(_abc_17692_n6604), .Y(_abc_17692_n6881) );
  OR2X2 OR2X2_2179 ( .A(_abc_17692_n6879), .B(_abc_17692_n6882), .Y(_abc_17692_n6883) );
  OR2X2 OR2X2_218 ( .A(_abc_17692_n1070), .B(delta_7_), .Y(_abc_17692_n1072) );
  OR2X2 OR2X2_2180 ( .A(_abc_17692_n6883), .B(_abc_17692_n6876), .Y(_abc_17692_n6884) );
  OR2X2 OR2X2_2181 ( .A(_abc_17692_n6885), .B(_abc_17692_n6884), .Y(_abc_17692_n6886) );
  OR2X2 OR2X2_2182 ( .A(_abc_17692_n6886), .B(_abc_17692_n6708), .Y(_abc_17692_n6887) );
  OR2X2 OR2X2_2183 ( .A(_abc_17692_n6510), .B(_abc_17692_n6281), .Y(_abc_17692_n6892) );
  OR2X2 OR2X2_2184 ( .A(_abc_17692_n6892), .B(_abc_17692_n6421), .Y(_abc_17692_n6893) );
  OR2X2 OR2X2_2185 ( .A(_abc_17692_n6012), .B(_abc_17692_n6893), .Y(_abc_17692_n6894) );
  OR2X2 OR2X2_2186 ( .A(_abc_17692_n6893), .B(_abc_17692_n6007), .Y(_abc_17692_n6895) );
  OR2X2 OR2X2_2187 ( .A(_abc_17692_n6892), .B(_abc_17692_n6426), .Y(_abc_17692_n6896) );
  OR2X2 OR2X2_2188 ( .A(_abc_17692_n6504), .B(_abc_17692_n6626), .Y(_abc_17692_n6898) );
  OR2X2 OR2X2_2189 ( .A(_abc_17692_n6903), .B(_abc_17692_n6800), .Y(_abc_17692_n6904) );
  OR2X2 OR2X2_219 ( .A(_abc_17692_n1073), .B(_abc_17692_n1071), .Y(_abc_17692_n1074) );
  OR2X2 OR2X2_2190 ( .A(_abc_17692_n6906), .B(_abc_17692_n6905), .Y(_abc_17692_n6907) );
  OR2X2 OR2X2_2191 ( .A(_abc_17692_n6914), .B(_abc_17692_n6633), .Y(_abc_17692_n6915) );
  OR2X2 OR2X2_2192 ( .A(_abc_17692_n6913), .B(_abc_17692_n6916), .Y(_abc_17692_n6917) );
  OR2X2 OR2X2_2193 ( .A(_abc_17692_n6917), .B(_abc_17692_n6912), .Y(_abc_17692_n6918) );
  OR2X2 OR2X2_2194 ( .A(_abc_17692_n6919), .B(_abc_17692_n6918), .Y(_abc_17692_n6920) );
  OR2X2 OR2X2_2195 ( .A(_abc_17692_n6920), .B(_abc_17692_n6848), .Y(_abc_17692_n6921) );
  OR2X2 OR2X2_2196 ( .A(_abc_17692_n6931), .B(_abc_17692_n6930), .Y(_abc_17692_n6932) );
  OR2X2 OR2X2_2197 ( .A(_abc_17692_n6929), .B(_abc_17692_n6932), .Y(_abc_17692_n6933) );
  OR2X2 OR2X2_2198 ( .A(_abc_17692_n6933), .B(_abc_17692_n6928), .Y(_abc_17692_n6934) );
  OR2X2 OR2X2_2199 ( .A(_abc_17692_n6934), .B(_abc_17692_n6936), .Y(_abc_17692_n6937) );
  OR2X2 OR2X2_22 ( .A(state_8_bF_buf9), .B(delta_27_), .Y(delta_27__FF_INPUT) );
  OR2X2 OR2X2_220 ( .A(_abc_17692_n1078), .B(_abc_17692_n1075), .Y(_abc_17692_n1079) );
  OR2X2 OR2X2_2200 ( .A(_abc_17692_n6937), .B(_abc_17692_n6754), .Y(_abc_17692_n6940) );
  OR2X2 OR2X2_2201 ( .A(_abc_17692_n6925), .B(_abc_17692_n6942), .Y(_abc_17692_n6943) );
  OR2X2 OR2X2_2202 ( .A(_abc_17692_n6943), .B(_abc_17692_n6909), .Y(_abc_17692_n6944) );
  OR2X2 OR2X2_2203 ( .A(_abc_17692_n6944), .B(_abc_17692_n6891), .Y(_abc_17692_n6945) );
  OR2X2 OR2X2_2204 ( .A(_abc_17692_n6947), .B(_abc_17692_n6948), .Y(_abc_17692_n6949) );
  OR2X2 OR2X2_2205 ( .A(_abc_17692_n6946), .B(_abc_17692_n6949), .Y(_abc_17692_n6950) );
  OR2X2 OR2X2_2206 ( .A(_abc_17692_n6872), .B(_abc_17692_n6950), .Y(workunit2_24__FF_INPUT) );
  OR2X2 OR2X2_2207 ( .A(_abc_17692_n6676), .B(_abc_17692_n6663), .Y(_abc_17692_n6953) );
  OR2X2 OR2X2_2208 ( .A(_abc_17692_n4926), .B(workunit1_30_), .Y(_abc_17692_n6955) );
  OR2X2 OR2X2_2209 ( .A(_abc_17692_n6956), .B(workunit1_21_), .Y(_abc_17692_n6957) );
  OR2X2 OR2X2_221 ( .A(_abc_17692_n1080), .B(_abc_17692_n1074), .Y(_abc_17692_n1081) );
  OR2X2 OR2X2_2210 ( .A(_abc_17692_n6954), .B(_abc_17692_n6964), .Y(_abc_17692_n6967) );
  OR2X2 OR2X2_2211 ( .A(_abc_17692_n6695), .B(_abc_17692_n6682), .Y(_abc_17692_n6969) );
  OR2X2 OR2X2_2212 ( .A(sum_25_), .B(\key_in[121] ), .Y(_abc_17692_n6973) );
  OR2X2 OR2X2_2213 ( .A(_abc_17692_n6970), .B(_abc_17692_n6974), .Y(_abc_17692_n6976) );
  OR2X2 OR2X2_2214 ( .A(_abc_17692_n6977), .B(_abc_17692_n6975), .Y(_abc_17692_n6978) );
  OR2X2 OR2X2_2215 ( .A(_abc_17692_n6978), .B(_abc_17692_n6968), .Y(_abc_17692_n6979) );
  OR2X2 OR2X2_2216 ( .A(_abc_17692_n6980), .B(_abc_17692_n6965), .Y(_abc_17692_n6981) );
  OR2X2 OR2X2_2217 ( .A(_abc_17692_n6983), .B(_abc_17692_n6981), .Y(_abc_17692_n6984) );
  OR2X2 OR2X2_2218 ( .A(_abc_17692_n6985), .B(_abc_17692_n6952), .Y(_abc_17692_n6986) );
  OR2X2 OR2X2_2219 ( .A(_abc_17692_n6995), .B(_abc_17692_n4047_bF_buf2), .Y(_abc_17692_n6996) );
  OR2X2 OR2X2_222 ( .A(_abc_17692_n1075), .B(_abc_17692_n1050), .Y(_abc_17692_n1085) );
  OR2X2 OR2X2_2220 ( .A(_abc_17692_n6996), .B(_abc_17692_n6993), .Y(_abc_17692_n6997) );
  OR2X2 OR2X2_2221 ( .A(_abc_17692_n6789), .B(_abc_17692_n6775), .Y(_abc_17692_n6998) );
  OR2X2 OR2X2_2222 ( .A(sum_25_), .B(\key_in[89] ), .Y(_abc_17692_n7001) );
  OR2X2 OR2X2_2223 ( .A(_abc_17692_n6998), .B(_abc_17692_n7003), .Y(_abc_17692_n7004) );
  OR2X2 OR2X2_2224 ( .A(_abc_17692_n7007), .B(_abc_17692_n6968), .Y(_abc_17692_n7008) );
  OR2X2 OR2X2_2225 ( .A(_abc_17692_n7009), .B(_abc_17692_n7005), .Y(_abc_17692_n7010) );
  OR2X2 OR2X2_2226 ( .A(_abc_17692_n7010), .B(_abc_17692_n6981), .Y(_abc_17692_n7011) );
  OR2X2 OR2X2_2227 ( .A(_abc_17692_n7015), .B(_abc_17692_n7013), .Y(_abc_17692_n7016) );
  OR2X2 OR2X2_2228 ( .A(_abc_17692_n7020), .B(_abc_17692_n7017), .Y(_abc_17692_n7021) );
  OR2X2 OR2X2_2229 ( .A(_abc_17692_n7022), .B(_abc_17692_n7016), .Y(_abc_17692_n7023) );
  OR2X2 OR2X2_223 ( .A(_abc_17692_n1056), .B(_abc_17692_n1085), .Y(_abc_17692_n1086) );
  OR2X2 OR2X2_2230 ( .A(_abc_17692_n6740), .B(_abc_17692_n6727), .Y(_abc_17692_n7026) );
  OR2X2 OR2X2_2231 ( .A(sum_25_), .B(\key_in[25] ), .Y(_abc_17692_n7030) );
  OR2X2 OR2X2_2232 ( .A(_abc_17692_n7027), .B(_abc_17692_n7031), .Y(_abc_17692_n7034) );
  OR2X2 OR2X2_2233 ( .A(_abc_17692_n6968), .B(_abc_17692_n7035), .Y(_abc_17692_n7036) );
  OR2X2 OR2X2_2234 ( .A(_abc_17692_n7037), .B(_abc_17692_n7032), .Y(_abc_17692_n7038) );
  OR2X2 OR2X2_2235 ( .A(_abc_17692_n6981), .B(_abc_17692_n7038), .Y(_abc_17692_n7039) );
  OR2X2 OR2X2_2236 ( .A(_abc_17692_n7050), .B(_abc_17692_n7047), .Y(_abc_17692_n7051) );
  OR2X2 OR2X2_2237 ( .A(_abc_17692_n7049), .B(_abc_17692_n7046), .Y(_abc_17692_n7052) );
  OR2X2 OR2X2_2238 ( .A(_abc_17692_n6834), .B(_abc_17692_n6821), .Y(_abc_17692_n7055) );
  OR2X2 OR2X2_2239 ( .A(sum_25_), .B(\key_in[57] ), .Y(_abc_17692_n7059) );
  OR2X2 OR2X2_224 ( .A(_abc_17692_n1093), .B(_abc_17692_n1084), .Y(_abc_17692_n1094) );
  OR2X2 OR2X2_2240 ( .A(_abc_17692_n7056), .B(_abc_17692_n7060), .Y(_abc_17692_n7063) );
  OR2X2 OR2X2_2241 ( .A(_abc_17692_n7066), .B(_abc_17692_n7067), .Y(_abc_17692_n7068) );
  OR2X2 OR2X2_2242 ( .A(_abc_17692_n7068), .B(_abc_17692_n6952), .Y(_abc_17692_n7069) );
  OR2X2 OR2X2_2243 ( .A(_abc_17692_n6968), .B(_abc_17692_n7064), .Y(_abc_17692_n7070) );
  OR2X2 OR2X2_2244 ( .A(_abc_17692_n6981), .B(_abc_17692_n7065), .Y(_abc_17692_n7071) );
  OR2X2 OR2X2_2245 ( .A(_abc_17692_n7072), .B(workunit2_25_), .Y(_abc_17692_n7073) );
  OR2X2 OR2X2_2246 ( .A(_abc_17692_n7078), .B(_abc_17692_n7075), .Y(_abc_17692_n7079) );
  OR2X2 OR2X2_2247 ( .A(_abc_17692_n7077), .B(_abc_17692_n7074), .Y(_abc_17692_n7080) );
  OR2X2 OR2X2_2248 ( .A(_abc_17692_n7082), .B(_abc_17692_n1863_bF_buf4), .Y(_abc_17692_n7083) );
  OR2X2 OR2X2_2249 ( .A(_abc_17692_n7083), .B(_abc_17692_n7054), .Y(_abc_17692_n7084) );
  OR2X2 OR2X2_225 ( .A(_abc_17692_n1083), .B(_abc_17692_n1094), .Y(sum_7__FF_INPUT) );
  OR2X2 OR2X2_2250 ( .A(_abc_17692_n7084), .B(_abc_17692_n7025), .Y(_abc_17692_n7085) );
  OR2X2 OR2X2_2251 ( .A(_abc_17692_n7091), .B(_abc_17692_n6989), .Y(_abc_17692_n7092) );
  OR2X2 OR2X2_2252 ( .A(_abc_17692_n7090), .B(_abc_17692_n6994), .Y(_abc_17692_n7093) );
  OR2X2 OR2X2_2253 ( .A(_abc_17692_n7099), .B(_abc_17692_n7100), .Y(_abc_17692_n7101) );
  OR2X2 OR2X2_2254 ( .A(_abc_17692_n7106), .B(_abc_17692_n7074), .Y(_abc_17692_n7107) );
  OR2X2 OR2X2_2255 ( .A(_abc_17692_n7105), .B(_abc_17692_n7075), .Y(_abc_17692_n7108) );
  OR2X2 OR2X2_2256 ( .A(_abc_17692_n7113), .B(_abc_17692_n7047), .Y(_abc_17692_n7114) );
  OR2X2 OR2X2_2257 ( .A(_abc_17692_n7115), .B(_abc_17692_n7046), .Y(_abc_17692_n7116) );
  OR2X2 OR2X2_2258 ( .A(_abc_17692_n7118), .B(_abc_17692_n7110), .Y(_abc_17692_n7119) );
  OR2X2 OR2X2_2259 ( .A(_abc_17692_n7119), .B(_abc_17692_n7102), .Y(_abc_17692_n7120) );
  OR2X2 OR2X2_226 ( .A(_abc_17692_n1099), .B(_abc_17692_n1096), .Y(_abc_17692_n1100) );
  OR2X2 OR2X2_2260 ( .A(_abc_17692_n7120), .B(_abc_17692_n7095), .Y(_abc_17692_n7121) );
  OR2X2 OR2X2_2261 ( .A(_abc_17692_n7123), .B(_abc_17692_n7124), .Y(_abc_17692_n7125) );
  OR2X2 OR2X2_2262 ( .A(_abc_17692_n7122), .B(_abc_17692_n7125), .Y(_abc_17692_n7126) );
  OR2X2 OR2X2_2263 ( .A(_abc_17692_n7087), .B(_abc_17692_n7126), .Y(workunit2_25__FF_INPUT) );
  OR2X2 OR2X2_2264 ( .A(_abc_17692_n7131), .B(_abc_17692_n6960), .Y(_abc_17692_n7132) );
  OR2X2 OR2X2_2265 ( .A(_abc_17692_n7130), .B(_abc_17692_n7132), .Y(_abc_17692_n7133) );
  OR2X2 OR2X2_2266 ( .A(_abc_17692_n5205), .B(workunit1_31_), .Y(_abc_17692_n7134) );
  OR2X2 OR2X2_2267 ( .A(_abc_17692_n7135), .B(workunit1_22_), .Y(_abc_17692_n7136) );
  OR2X2 OR2X2_2268 ( .A(_abc_17692_n7139), .B(_abc_17692_n7140), .Y(_abc_17692_n7141) );
  OR2X2 OR2X2_2269 ( .A(_abc_17692_n6679), .B(_abc_17692_n7144), .Y(_abc_17692_n7145) );
  OR2X2 OR2X2_227 ( .A(_abc_17692_n1105), .B(_abc_17692_n1101), .Y(_abc_17692_n1106) );
  OR2X2 OR2X2_2270 ( .A(_abc_17692_n7148), .B(_abc_17692_n7143), .Y(_abc_17692_n7149) );
  OR2X2 OR2X2_2271 ( .A(_abc_17692_n7153), .B(_abc_17692_n7028), .Y(_abc_17692_n7154) );
  OR2X2 OR2X2_2272 ( .A(_abc_17692_n7152), .B(_abc_17692_n7154), .Y(_abc_17692_n7155) );
  OR2X2 OR2X2_2273 ( .A(sum_26_), .B(\key_in[26] ), .Y(_abc_17692_n7158) );
  OR2X2 OR2X2_2274 ( .A(_abc_17692_n7165), .B(_abc_17692_n7160), .Y(_abc_17692_n7166) );
  OR2X2 OR2X2_2275 ( .A(_abc_17692_n7167), .B(_abc_17692_n7169), .Y(_abc_17692_n7170) );
  OR2X2 OR2X2_2276 ( .A(_abc_17692_n7171), .B(_abc_17692_n7128), .Y(_abc_17692_n7172) );
  OR2X2 OR2X2_2277 ( .A(_abc_17692_n7170), .B(workunit2_26_), .Y(_abc_17692_n7173) );
  OR2X2 OR2X2_2278 ( .A(_abc_17692_n7046), .B(_abc_17692_n7048), .Y(_abc_17692_n7178) );
  OR2X2 OR2X2_2279 ( .A(_abc_17692_n7046), .B(_abc_17692_n6754), .Y(_abc_17692_n7181) );
  OR2X2 OR2X2_228 ( .A(_abc_17692_n1104_1), .B(_abc_17692_n1100), .Y(_abc_17692_n1107_1) );
  OR2X2 OR2X2_2280 ( .A(_abc_17692_n7183), .B(_abc_17692_n7180), .Y(_abc_17692_n7184) );
  OR2X2 OR2X2_2281 ( .A(_abc_17692_n7184), .B(_abc_17692_n7175), .Y(_abc_17692_n7185) );
  OR2X2 OR2X2_2282 ( .A(_abc_17692_n6787), .B(_abc_17692_n7191), .Y(_abc_17692_n7192) );
  OR2X2 OR2X2_2283 ( .A(_abc_17692_n7193), .B(_abc_17692_n6999), .Y(_abc_17692_n7194) );
  OR2X2 OR2X2_2284 ( .A(sum_26_), .B(\key_in[90] ), .Y(_abc_17692_n7200) );
  OR2X2 OR2X2_2285 ( .A(_abc_17692_n7202), .B(_abc_17692_n7204), .Y(_abc_17692_n7205) );
  OR2X2 OR2X2_2286 ( .A(_abc_17692_n7206), .B(_abc_17692_n7149), .Y(_abc_17692_n7207) );
  OR2X2 OR2X2_2287 ( .A(_abc_17692_n7205), .B(_abc_17692_n7150), .Y(_abc_17692_n7208) );
  OR2X2 OR2X2_2288 ( .A(_abc_17692_n7209), .B(workunit2_26_), .Y(_abc_17692_n7212) );
  OR2X2 OR2X2_2289 ( .A(_abc_17692_n7215), .B(_abc_17692_n7214), .Y(_abc_17692_n7216) );
  OR2X2 OR2X2_229 ( .A(_abc_17692_n1089), .B(_abc_17692_n1073), .Y(_abc_17692_n1110) );
  OR2X2 OR2X2_2290 ( .A(_abc_17692_n7218), .B(_abc_17692_n7216), .Y(_abc_17692_n7219) );
  OR2X2 OR2X2_2291 ( .A(_abc_17692_n7219), .B(_abc_17692_n7213), .Y(_abc_17692_n7222) );
  OR2X2 OR2X2_2292 ( .A(_abc_17692_n7227), .B(_abc_17692_n7057), .Y(_abc_17692_n7228) );
  OR2X2 OR2X2_2293 ( .A(_abc_17692_n7226), .B(_abc_17692_n7228), .Y(_abc_17692_n7229) );
  OR2X2 OR2X2_2294 ( .A(sum_26_), .B(\key_in[58] ), .Y(_abc_17692_n7232) );
  OR2X2 OR2X2_2295 ( .A(_abc_17692_n7229), .B(_abc_17692_n7233), .Y(_abc_17692_n7236) );
  OR2X2 OR2X2_2296 ( .A(_abc_17692_n7149), .B(_abc_17692_n7237), .Y(_abc_17692_n7238) );
  OR2X2 OR2X2_2297 ( .A(_abc_17692_n7150), .B(_abc_17692_n7239), .Y(_abc_17692_n7240) );
  OR2X2 OR2X2_2298 ( .A(_abc_17692_n7241), .B(_abc_17692_n7128), .Y(_abc_17692_n7242) );
  OR2X2 OR2X2_2299 ( .A(_abc_17692_n7243), .B(workunit2_26_), .Y(_abc_17692_n7244) );
  OR2X2 OR2X2_23 ( .A(state_8_bF_buf8), .B(delta_28_), .Y(delta_28__FF_INPUT) );
  OR2X2 OR2X2_230 ( .A(_abc_17692_n1087), .B(_abc_17692_n1110), .Y(_abc_17692_n1111) );
  OR2X2 OR2X2_2300 ( .A(_abc_17692_n7074), .B(_abc_17692_n7076), .Y(_abc_17692_n7249) );
  OR2X2 OR2X2_2301 ( .A(_abc_17692_n7074), .B(_abc_17692_n6848), .Y(_abc_17692_n7251) );
  OR2X2 OR2X2_2302 ( .A(_abc_17692_n6861), .B(_abc_17692_n7251), .Y(_abc_17692_n7252) );
  OR2X2 OR2X2_2303 ( .A(_abc_17692_n7254), .B(_abc_17692_n7246), .Y(_abc_17692_n7255) );
  OR2X2 OR2X2_2304 ( .A(_abc_17692_n7253), .B(_abc_17692_n7245), .Y(_abc_17692_n7256) );
  OR2X2 OR2X2_2305 ( .A(_abc_17692_n7258), .B(_abc_17692_n1863_bF_buf2), .Y(_abc_17692_n7259) );
  OR2X2 OR2X2_2306 ( .A(_abc_17692_n7224), .B(_abc_17692_n7259), .Y(_abc_17692_n7260) );
  OR2X2 OR2X2_2307 ( .A(_abc_17692_n7260), .B(_abc_17692_n7189), .Y(_abc_17692_n7261) );
  OR2X2 OR2X2_2308 ( .A(_abc_17692_n7264), .B(_abc_17692_n6971), .Y(_abc_17692_n7265) );
  OR2X2 OR2X2_2309 ( .A(_abc_17692_n7263), .B(_abc_17692_n7265), .Y(_abc_17692_n7266) );
  OR2X2 OR2X2_231 ( .A(_abc_17692_n1111), .B(_abc_17692_n1100), .Y(_abc_17692_n1112) );
  OR2X2 OR2X2_2310 ( .A(sum_26_), .B(\key_in[122] ), .Y(_abc_17692_n7269) );
  OR2X2 OR2X2_2311 ( .A(_abc_17692_n7266), .B(_abc_17692_n7270), .Y(_abc_17692_n7273) );
  OR2X2 OR2X2_2312 ( .A(_abc_17692_n7274), .B(_abc_17692_n7149), .Y(_abc_17692_n7275) );
  OR2X2 OR2X2_2313 ( .A(_abc_17692_n7276), .B(_abc_17692_n7150), .Y(_abc_17692_n7277) );
  OR2X2 OR2X2_2314 ( .A(_abc_17692_n7278), .B(_abc_17692_n7128), .Y(_abc_17692_n7279) );
  OR2X2 OR2X2_2315 ( .A(_abc_17692_n7280), .B(workunit2_26_), .Y(_abc_17692_n7281) );
  OR2X2 OR2X2_2316 ( .A(_abc_17692_n7284), .B(_abc_17692_n7283), .Y(_abc_17692_n7285) );
  OR2X2 OR2X2_2317 ( .A(_abc_17692_n6720), .B(_abc_17692_n7288), .Y(_abc_17692_n7289) );
  OR2X2 OR2X2_2318 ( .A(_abc_17692_n7290), .B(_abc_17692_n7282), .Y(_abc_17692_n7291) );
  OR2X2 OR2X2_2319 ( .A(_abc_17692_n7293), .B(_abc_17692_n7292), .Y(_abc_17692_n7294) );
  OR2X2 OR2X2_232 ( .A(_abc_17692_n1117), .B(state_8_bF_buf5), .Y(_abc_17692_n1118) );
  OR2X2 OR2X2_2320 ( .A(_abc_17692_n7295), .B(_abc_17692_n4047_bF_buf1), .Y(_abc_17692_n7296) );
  OR2X2 OR2X2_2321 ( .A(_abc_17692_n7299), .B(_abc_17692_n6987), .Y(_abc_17692_n7300) );
  OR2X2 OR2X2_2322 ( .A(_abc_17692_n7303), .B(_abc_17692_n7301), .Y(_abc_17692_n7304) );
  OR2X2 OR2X2_2323 ( .A(_abc_17692_n7304), .B(_abc_17692_n7282), .Y(_abc_17692_n7307) );
  OR2X2 OR2X2_2324 ( .A(_abc_17692_n7013), .B(_abc_17692_n6798), .Y(_abc_17692_n7311) );
  OR2X2 OR2X2_2325 ( .A(_abc_17692_n7312), .B(_abc_17692_n7015), .Y(_abc_17692_n7313) );
  OR2X2 OR2X2_2326 ( .A(_abc_17692_n7016), .B(_abc_17692_n6800), .Y(_abc_17692_n7315) );
  OR2X2 OR2X2_2327 ( .A(_abc_17692_n7317), .B(_abc_17692_n7314), .Y(_abc_17692_n7318) );
  OR2X2 OR2X2_2328 ( .A(_abc_17692_n7318), .B(_abc_17692_n7310), .Y(_abc_17692_n7321) );
  OR2X2 OR2X2_2329 ( .A(_abc_17692_n7324), .B(_abc_17692_n7103), .Y(_abc_17692_n7325) );
  OR2X2 OR2X2_233 ( .A(_abc_17692_n1116), .B(_abc_17692_n1118), .Y(_abc_17692_n1119) );
  OR2X2 OR2X2_2330 ( .A(_abc_17692_n7328), .B(_abc_17692_n7326), .Y(_abc_17692_n7329) );
  OR2X2 OR2X2_2331 ( .A(_abc_17692_n7329), .B(_abc_17692_n7245), .Y(_abc_17692_n7332) );
  OR2X2 OR2X2_2332 ( .A(_abc_17692_n7041), .B(_abc_17692_n7111), .Y(_abc_17692_n7335) );
  OR2X2 OR2X2_2333 ( .A(_abc_17692_n7338), .B(_abc_17692_n7336), .Y(_abc_17692_n7339) );
  OR2X2 OR2X2_2334 ( .A(_abc_17692_n7339), .B(_abc_17692_n7174), .Y(_abc_17692_n7342) );
  OR2X2 OR2X2_2335 ( .A(_abc_17692_n7334), .B(_abc_17692_n7344), .Y(_abc_17692_n7345) );
  OR2X2 OR2X2_2336 ( .A(_abc_17692_n7323), .B(_abc_17692_n7345), .Y(_abc_17692_n7346) );
  OR2X2 OR2X2_2337 ( .A(_abc_17692_n7346), .B(_abc_17692_n7309), .Y(_abc_17692_n7347) );
  OR2X2 OR2X2_2338 ( .A(_abc_17692_n7349), .B(_abc_17692_n7350), .Y(_abc_17692_n7351) );
  OR2X2 OR2X2_2339 ( .A(_abc_17692_n7348), .B(_abc_17692_n7351), .Y(_abc_17692_n7352) );
  OR2X2 OR2X2_234 ( .A(_abc_17692_n1119), .B(_abc_17692_n1109), .Y(sum_8__FF_INPUT) );
  OR2X2 OR2X2_2340 ( .A(_abc_17692_n7298), .B(_abc_17692_n7352), .Y(workunit2_26__FF_INPUT) );
  OR2X2 OR2X2_2341 ( .A(_abc_17692_n7147), .B(_abc_17692_n7141), .Y(_abc_17692_n7355) );
  OR2X2 OR2X2_2342 ( .A(_abc_17692_n7358), .B(_abc_17692_n7357), .Y(_abc_17692_n7359) );
  OR2X2 OR2X2_2343 ( .A(_abc_17692_n7356), .B(_abc_17692_n7360), .Y(_abc_17692_n7361) );
  OR2X2 OR2X2_2344 ( .A(_abc_17692_n7143), .B(_abc_17692_n7139), .Y(_abc_17692_n7362) );
  OR2X2 OR2X2_2345 ( .A(_abc_17692_n7362), .B(_abc_17692_n7359), .Y(_abc_17692_n7363) );
  OR2X2 OR2X2_2346 ( .A(_abc_17692_n7271), .B(_abc_17692_n7267), .Y(_abc_17692_n7365) );
  OR2X2 OR2X2_2347 ( .A(sum_27_), .B(\key_in[123] ), .Y(_abc_17692_n7368) );
  OR2X2 OR2X2_2348 ( .A(_abc_17692_n7365), .B(_abc_17692_n7370), .Y(_abc_17692_n7371) );
  OR2X2 OR2X2_2349 ( .A(_abc_17692_n7374), .B(_abc_17692_n7364), .Y(_abc_17692_n7375) );
  OR2X2 OR2X2_235 ( .A(_abc_17692_n1130), .B(_abc_17692_n1127_1), .Y(_abc_17692_n1131) );
  OR2X2 OR2X2_2350 ( .A(_abc_17692_n7377), .B(_abc_17692_n7376), .Y(_abc_17692_n7378) );
  OR2X2 OR2X2_2351 ( .A(_abc_17692_n7380), .B(_abc_17692_n7372), .Y(_abc_17692_n7381) );
  OR2X2 OR2X2_2352 ( .A(_abc_17692_n7381), .B(_abc_17692_n7378), .Y(_abc_17692_n7382) );
  OR2X2 OR2X2_2353 ( .A(_abc_17692_n7381), .B(_abc_17692_n7364), .Y(_abc_17692_n7386) );
  OR2X2 OR2X2_2354 ( .A(_abc_17692_n7374), .B(_abc_17692_n7378), .Y(_abc_17692_n7387) );
  OR2X2 OR2X2_2355 ( .A(_abc_17692_n7384), .B(_abc_17692_n7389), .Y(_abc_17692_n7390) );
  OR2X2 OR2X2_2356 ( .A(_abc_17692_n7305), .B(_abc_17692_n7391), .Y(_abc_17692_n7392) );
  OR2X2 OR2X2_2357 ( .A(_abc_17692_n7393), .B(_abc_17692_n7390), .Y(_abc_17692_n7394) );
  OR2X2 OR2X2_2358 ( .A(_abc_17692_n7388), .B(_abc_17692_n7385), .Y(_abc_17692_n7395) );
  OR2X2 OR2X2_2359 ( .A(_abc_17692_n7383), .B(workunit2_27_), .Y(_abc_17692_n7396) );
  OR2X2 OR2X2_236 ( .A(_abc_17692_n1129), .B(_abc_17692_n1132), .Y(_abc_17692_n1133) );
  OR2X2 OR2X2_2360 ( .A(_abc_17692_n7392), .B(_abc_17692_n7397), .Y(_abc_17692_n7398) );
  OR2X2 OR2X2_2361 ( .A(_abc_17692_n7196), .B(_abc_17692_n7203), .Y(_abc_17692_n7401) );
  OR2X2 OR2X2_2362 ( .A(sum_27_), .B(\key_in[91] ), .Y(_abc_17692_n7405) );
  OR2X2 OR2X2_2363 ( .A(_abc_17692_n7402), .B(_abc_17692_n7406), .Y(_abc_17692_n7409) );
  OR2X2 OR2X2_2364 ( .A(_abc_17692_n7410), .B(_abc_17692_n7364), .Y(_abc_17692_n7411) );
  OR2X2 OR2X2_2365 ( .A(_abc_17692_n7414), .B(_abc_17692_n7407), .Y(_abc_17692_n7415) );
  OR2X2 OR2X2_2366 ( .A(_abc_17692_n7415), .B(_abc_17692_n7378), .Y(_abc_17692_n7416) );
  OR2X2 OR2X2_2367 ( .A(_abc_17692_n7415), .B(_abc_17692_n7364), .Y(_abc_17692_n7419) );
  OR2X2 OR2X2_2368 ( .A(_abc_17692_n7410), .B(_abc_17692_n7378), .Y(_abc_17692_n7420) );
  OR2X2 OR2X2_2369 ( .A(_abc_17692_n7418), .B(_abc_17692_n7422), .Y(_abc_17692_n7423) );
  OR2X2 OR2X2_237 ( .A(_abc_17692_n1132), .B(_abc_17692_n1138_1), .Y(_abc_17692_n1139) );
  OR2X2 OR2X2_2370 ( .A(_abc_17692_n7429), .B(_abc_17692_n7424), .Y(_abc_17692_n7430) );
  OR2X2 OR2X2_2371 ( .A(_abc_17692_n7428), .B(_abc_17692_n7423), .Y(_abc_17692_n7431) );
  OR2X2 OR2X2_2372 ( .A(sum_27_), .B(\key_in[59] ), .Y(_abc_17692_n7437) );
  OR2X2 OR2X2_2373 ( .A(_abc_17692_n7234), .B(_abc_17692_n7230), .Y(_abc_17692_n7440) );
  OR2X2 OR2X2_2374 ( .A(_abc_17692_n7439), .B(_abc_17692_n7442), .Y(_abc_17692_n7443) );
  OR2X2 OR2X2_2375 ( .A(_abc_17692_n7364), .B(_abc_17692_n7443), .Y(_abc_17692_n7444) );
  OR2X2 OR2X2_2376 ( .A(_abc_17692_n7440), .B(_abc_17692_n7441), .Y(_abc_17692_n7445) );
  OR2X2 OR2X2_2377 ( .A(_abc_17692_n7378), .B(_abc_17692_n7447), .Y(_abc_17692_n7448) );
  OR2X2 OR2X2_2378 ( .A(_abc_17692_n7449), .B(_abc_17692_n7385), .Y(_abc_17692_n7450) );
  OR2X2 OR2X2_2379 ( .A(_abc_17692_n7364), .B(_abc_17692_n7447), .Y(_abc_17692_n7451) );
  OR2X2 OR2X2_238 ( .A(_abc_17692_n1113), .B(_abc_17692_n1139), .Y(_abc_17692_n1140) );
  OR2X2 OR2X2_2380 ( .A(_abc_17692_n7378), .B(_abc_17692_n7443), .Y(_abc_17692_n7452) );
  OR2X2 OR2X2_2381 ( .A(_abc_17692_n7453), .B(workunit2_27_), .Y(_abc_17692_n7454) );
  OR2X2 OR2X2_2382 ( .A(_abc_17692_n7457), .B(_abc_17692_n7455), .Y(_abc_17692_n7458) );
  OR2X2 OR2X2_2383 ( .A(_abc_17692_n7456), .B(_abc_17692_n7459), .Y(_abc_17692_n7460) );
  OR2X2 OR2X2_2384 ( .A(sum_27_), .B(\key_in[27] ), .Y(_abc_17692_n7467) );
  OR2X2 OR2X2_2385 ( .A(_abc_17692_n7160), .B(_abc_17692_n7156), .Y(_abc_17692_n7470) );
  OR2X2 OR2X2_2386 ( .A(_abc_17692_n7469), .B(_abc_17692_n7472), .Y(_abc_17692_n7473) );
  OR2X2 OR2X2_2387 ( .A(_abc_17692_n7364), .B(_abc_17692_n7473), .Y(_abc_17692_n7474) );
  OR2X2 OR2X2_2388 ( .A(_abc_17692_n7470), .B(_abc_17692_n7471), .Y(_abc_17692_n7475) );
  OR2X2 OR2X2_2389 ( .A(_abc_17692_n7378), .B(_abc_17692_n7477), .Y(_abc_17692_n7478) );
  OR2X2 OR2X2_239 ( .A(_abc_17692_n1146), .B(state_8_bF_buf4), .Y(_abc_17692_n1147) );
  OR2X2 OR2X2_2390 ( .A(_abc_17692_n7479), .B(_abc_17692_n7385), .Y(_abc_17692_n7480) );
  OR2X2 OR2X2_2391 ( .A(_abc_17692_n7364), .B(_abc_17692_n7477), .Y(_abc_17692_n7481) );
  OR2X2 OR2X2_2392 ( .A(_abc_17692_n7378), .B(_abc_17692_n7473), .Y(_abc_17692_n7482) );
  OR2X2 OR2X2_2393 ( .A(_abc_17692_n7483), .B(workunit2_27_), .Y(_abc_17692_n7484) );
  OR2X2 OR2X2_2394 ( .A(_abc_17692_n7487), .B(_abc_17692_n7486), .Y(_abc_17692_n7488) );
  OR2X2 OR2X2_2395 ( .A(_abc_17692_n7489), .B(_abc_17692_n7485), .Y(_abc_17692_n7490) );
  OR2X2 OR2X2_2396 ( .A(_abc_17692_n7492), .B(_abc_17692_n7462), .Y(_abc_17692_n7493) );
  OR2X2 OR2X2_2397 ( .A(_abc_17692_n7493), .B(_abc_17692_n7433), .Y(_abc_17692_n7494) );
  OR2X2 OR2X2_2398 ( .A(_abc_17692_n7494), .B(_abc_17692_n7400), .Y(_abc_17692_n7495) );
  OR2X2 OR2X2_2399 ( .A(_abc_17692_n7280), .B(_abc_17692_n7128), .Y(_abc_17692_n7497) );
  OR2X2 OR2X2_24 ( .A(state_8_bF_buf7), .B(delta_31_), .Y(delta_31__FF_INPUT) );
  OR2X2 OR2X2_240 ( .A(_abc_17692_n1145), .B(_abc_17692_n1147), .Y(_abc_17692_n1148) );
  OR2X2 OR2X2_2400 ( .A(_abc_17692_n7501), .B(_abc_17692_n4047_bF_buf0), .Y(_abc_17692_n7502) );
  OR2X2 OR2X2_2401 ( .A(_abc_17692_n7502), .B(_abc_17692_n7500), .Y(_abc_17692_n7503) );
  OR2X2 OR2X2_2402 ( .A(_abc_17692_n7220), .B(_abc_17692_n7210), .Y(_abc_17692_n7504) );
  OR2X2 OR2X2_2403 ( .A(_abc_17692_n7505), .B(_abc_17692_n7424), .Y(_abc_17692_n7506) );
  OR2X2 OR2X2_2404 ( .A(_abc_17692_n7504), .B(_abc_17692_n7423), .Y(_abc_17692_n7507) );
  OR2X2 OR2X2_2405 ( .A(_abc_17692_n7186), .B(_abc_17692_n7510), .Y(_abc_17692_n7511) );
  OR2X2 OR2X2_2406 ( .A(_abc_17692_n7512), .B(_abc_17692_n7485), .Y(_abc_17692_n7513) );
  OR2X2 OR2X2_2407 ( .A(_abc_17692_n7511), .B(_abc_17692_n7486), .Y(_abc_17692_n7514) );
  OR2X2 OR2X2_2408 ( .A(_abc_17692_n7520), .B(_abc_17692_n7459), .Y(_abc_17692_n7521) );
  OR2X2 OR2X2_2409 ( .A(_abc_17692_n7519), .B(_abc_17692_n7455), .Y(_abc_17692_n7522) );
  OR2X2 OR2X2_241 ( .A(_abc_17692_n1135), .B(_abc_17692_n1148), .Y(sum_9__FF_INPUT) );
  OR2X2 OR2X2_2410 ( .A(_abc_17692_n7524), .B(_abc_17692_n1863_bF_buf10), .Y(_abc_17692_n7525) );
  OR2X2 OR2X2_2411 ( .A(_abc_17692_n7516), .B(_abc_17692_n7525), .Y(_abc_17692_n7526) );
  OR2X2 OR2X2_2412 ( .A(_abc_17692_n7526), .B(_abc_17692_n7509), .Y(_abc_17692_n7527) );
  OR2X2 OR2X2_2413 ( .A(_abc_17692_n7530), .B(_abc_17692_n7531), .Y(_abc_17692_n7532) );
  OR2X2 OR2X2_2414 ( .A(_abc_17692_n7529), .B(_abc_17692_n7532), .Y(_abc_17692_n7533) );
  OR2X2 OR2X2_2415 ( .A(_abc_17692_n7533), .B(_abc_17692_n7496), .Y(workunit2_27__FF_INPUT) );
  OR2X2 OR2X2_2416 ( .A(_abc_17692_n7539), .B(_abc_17692_n7357), .Y(_abc_17692_n7540) );
  OR2X2 OR2X2_2417 ( .A(_abc_17692_n7538), .B(_abc_17692_n7540), .Y(_abc_17692_n7541) );
  OR2X2 OR2X2_2418 ( .A(_abc_17692_n7537), .B(_abc_17692_n7541), .Y(_abc_17692_n7542) );
  OR2X2 OR2X2_2419 ( .A(_abc_17692_n7544), .B(_abc_17692_n7543), .Y(_abc_17692_n7545) );
  OR2X2 OR2X2_242 ( .A(_abc_17692_n1153), .B(_abc_17692_n1150), .Y(_abc_17692_n1154) );
  OR2X2 OR2X2_2420 ( .A(_abc_17692_n7542), .B(_abc_17692_n7546), .Y(_abc_17692_n7549) );
  OR2X2 OR2X2_2421 ( .A(sum_28_), .B(\key_in[124] ), .Y(_abc_17692_n7553) );
  OR2X2 OR2X2_2422 ( .A(_abc_17692_n7271), .B(_abc_17692_n7556), .Y(_abc_17692_n7557) );
  OR2X2 OR2X2_2423 ( .A(_abc_17692_n7562), .B(_abc_17692_n7559), .Y(_abc_17692_n7563) );
  OR2X2 OR2X2_2424 ( .A(_abc_17692_n7567), .B(_abc_17692_n7564), .Y(_abc_17692_n7568) );
  OR2X2 OR2X2_2425 ( .A(_abc_17692_n7568), .B(_abc_17692_n7535), .Y(_abc_17692_n7569) );
  OR2X2 OR2X2_2426 ( .A(_abc_17692_n7570), .B(workunit2_28_), .Y(_abc_17692_n7571) );
  OR2X2 OR2X2_2427 ( .A(_abc_17692_n6720), .B(_abc_17692_n7575), .Y(_abc_17692_n7576) );
  OR2X2 OR2X2_2428 ( .A(_abc_17692_n7397), .B(_abc_17692_n7497), .Y(_abc_17692_n7581) );
  OR2X2 OR2X2_2429 ( .A(_abc_17692_n7585), .B(_abc_17692_n7572), .Y(_abc_17692_n7586) );
  OR2X2 OR2X2_243 ( .A(_abc_17692_n1107_1), .B(_abc_17692_n1132), .Y(_abc_17692_n1156) );
  OR2X2 OR2X2_2430 ( .A(_abc_17692_n7584), .B(_abc_17692_n7587), .Y(_abc_17692_n7588) );
  OR2X2 OR2X2_2431 ( .A(_abc_17692_n7589), .B(_abc_17692_n4047_bF_buf4), .Y(_abc_17692_n7590) );
  OR2X2 OR2X2_2432 ( .A(sum_28_), .B(\key_in[28] ), .Y(_abc_17692_n7593) );
  OR2X2 OR2X2_2433 ( .A(_abc_17692_n7160), .B(_abc_17692_n7596), .Y(_abc_17692_n7597) );
  OR2X2 OR2X2_2434 ( .A(_abc_17692_n7602), .B(_abc_17692_n7599), .Y(_abc_17692_n7603) );
  OR2X2 OR2X2_2435 ( .A(_abc_17692_n7606), .B(_abc_17692_n7604), .Y(_abc_17692_n7607) );
  OR2X2 OR2X2_2436 ( .A(_abc_17692_n7608), .B(_abc_17692_n7535), .Y(_abc_17692_n7609) );
  OR2X2 OR2X2_2437 ( .A(_abc_17692_n7607), .B(workunit2_28_), .Y(_abc_17692_n7610) );
  OR2X2 OR2X2_2438 ( .A(_abc_17692_n6768), .B(_abc_17692_n7615), .Y(_abc_17692_n7616) );
  OR2X2 OR2X2_2439 ( .A(_abc_17692_n7617), .B(_abc_17692_n7179), .Y(_abc_17692_n7618) );
  OR2X2 OR2X2_244 ( .A(_abc_17692_n1157), .B(_abc_17692_n1125), .Y(_abc_17692_n1158) );
  OR2X2 OR2X2_2440 ( .A(_abc_17692_n7620), .B(_abc_17692_n7619), .Y(_abc_17692_n7621) );
  OR2X2 OR2X2_2441 ( .A(_abc_17692_n7625), .B(_abc_17692_n7612), .Y(_abc_17692_n7626) );
  OR2X2 OR2X2_2442 ( .A(sum_28_), .B(\key_in[92] ), .Y(_abc_17692_n7633) );
  OR2X2 OR2X2_2443 ( .A(_abc_17692_n7637), .B(_abc_17692_n7635), .Y(_abc_17692_n7638) );
  OR2X2 OR2X2_2444 ( .A(_abc_17692_n7640), .B(_abc_17692_n7642), .Y(_abc_17692_n7643) );
  OR2X2 OR2X2_2445 ( .A(_abc_17692_n7644), .B(_abc_17692_n7565), .Y(_abc_17692_n7645) );
  OR2X2 OR2X2_2446 ( .A(_abc_17692_n7643), .B(_abc_17692_n7550), .Y(_abc_17692_n7646) );
  OR2X2 OR2X2_2447 ( .A(_abc_17692_n7647), .B(workunit2_28_), .Y(_abc_17692_n7650) );
  OR2X2 OR2X2_2448 ( .A(_abc_17692_n7424), .B(_abc_17692_n7310), .Y(_abc_17692_n7653) );
  OR2X2 OR2X2_2449 ( .A(_abc_17692_n7653), .B(_abc_17692_n7652), .Y(_abc_17692_n7654) );
  OR2X2 OR2X2_245 ( .A(_abc_17692_n1160), .B(_abc_17692_n1155), .Y(_abc_17692_n1163) );
  OR2X2 OR2X2_2450 ( .A(_abc_17692_n7657), .B(_abc_17692_n7653), .Y(_abc_17692_n7658) );
  OR2X2 OR2X2_2451 ( .A(_abc_17692_n7660), .B(_abc_17692_n7659), .Y(_abc_17692_n7661) );
  OR2X2 OR2X2_2452 ( .A(_abc_17692_n7664), .B(_abc_17692_n7656), .Y(_abc_17692_n7665) );
  OR2X2 OR2X2_2453 ( .A(_abc_17692_n7665), .B(_abc_17692_n7651), .Y(_abc_17692_n7668) );
  OR2X2 OR2X2_2454 ( .A(sum_28_), .B(\key_in[60] ), .Y(_abc_17692_n7673) );
  OR2X2 OR2X2_2455 ( .A(_abc_17692_n7234), .B(_abc_17692_n7676), .Y(_abc_17692_n7677) );
  OR2X2 OR2X2_2456 ( .A(_abc_17692_n7682), .B(_abc_17692_n7679), .Y(_abc_17692_n7683) );
  OR2X2 OR2X2_2457 ( .A(_abc_17692_n7686), .B(_abc_17692_n7684), .Y(_abc_17692_n7687) );
  OR2X2 OR2X2_2458 ( .A(_abc_17692_n7688), .B(_abc_17692_n7535), .Y(_abc_17692_n7689) );
  OR2X2 OR2X2_2459 ( .A(_abc_17692_n7687), .B(workunit2_28_), .Y(_abc_17692_n7690) );
  OR2X2 OR2X2_246 ( .A(_abc_17692_n1141), .B(_abc_17692_n1166), .Y(_abc_17692_n1167) );
  OR2X2 OR2X2_2460 ( .A(_abc_17692_n7455), .B(_abc_17692_n7245), .Y(_abc_17692_n7693) );
  OR2X2 OR2X2_2461 ( .A(_abc_17692_n7693), .B(_abc_17692_n7251), .Y(_abc_17692_n7694) );
  OR2X2 OR2X2_2462 ( .A(_abc_17692_n6861), .B(_abc_17692_n7694), .Y(_abc_17692_n7695) );
  OR2X2 OR2X2_2463 ( .A(_abc_17692_n7693), .B(_abc_17692_n7250), .Y(_abc_17692_n7696) );
  OR2X2 OR2X2_2464 ( .A(_abc_17692_n7455), .B(_abc_17692_n7518), .Y(_abc_17692_n7699) );
  OR2X2 OR2X2_2465 ( .A(_abc_17692_n7703), .B(_abc_17692_n7692), .Y(_abc_17692_n7706) );
  OR2X2 OR2X2_2466 ( .A(_abc_17692_n7708), .B(_abc_17692_n1863_bF_buf9), .Y(_abc_17692_n7709) );
  OR2X2 OR2X2_2467 ( .A(_abc_17692_n7670), .B(_abc_17692_n7709), .Y(_abc_17692_n7710) );
  OR2X2 OR2X2_2468 ( .A(_abc_17692_n7710), .B(_abc_17692_n7630), .Y(_abc_17692_n7711) );
  OR2X2 OR2X2_2469 ( .A(_abc_17692_n7718), .B(_abc_17692_n7384), .Y(_abc_17692_n7719) );
  OR2X2 OR2X2_247 ( .A(_abc_17692_n1170), .B(_abc_17692_n1154), .Y(_abc_17692_n1173) );
  OR2X2 OR2X2_2470 ( .A(_abc_17692_n7717), .B(_abc_17692_n7719), .Y(_abc_17692_n7720) );
  OR2X2 OR2X2_2471 ( .A(_abc_17692_n7716), .B(_abc_17692_n7720), .Y(_abc_17692_n7721) );
  OR2X2 OR2X2_2472 ( .A(_abc_17692_n7721), .B(_abc_17692_n7587), .Y(_abc_17692_n7722) );
  OR2X2 OR2X2_2473 ( .A(_abc_17692_n7423), .B(_abc_17692_n7213), .Y(_abc_17692_n7728) );
  OR2X2 OR2X2_2474 ( .A(_abc_17692_n7728), .B(_abc_17692_n7315), .Y(_abc_17692_n7729) );
  OR2X2 OR2X2_2475 ( .A(_abc_17692_n6903), .B(_abc_17692_n7729), .Y(_abc_17692_n7730) );
  OR2X2 OR2X2_2476 ( .A(_abc_17692_n7728), .B(_abc_17692_n7313), .Y(_abc_17692_n7731) );
  OR2X2 OR2X2_2477 ( .A(_abc_17692_n7418), .B(_abc_17692_n7426), .Y(_abc_17692_n7733) );
  OR2X2 OR2X2_2478 ( .A(_abc_17692_n7738), .B(_abc_17692_n7727), .Y(_abc_17692_n7741) );
  OR2X2 OR2X2_2479 ( .A(_abc_17692_n7749), .B(_abc_17692_n7748), .Y(_abc_17692_n7750) );
  OR2X2 OR2X2_248 ( .A(_abc_17692_n1176), .B(state_8_bF_buf3), .Y(_abc_17692_n1177) );
  OR2X2 OR2X2_2480 ( .A(_abc_17692_n7747), .B(_abc_17692_n7751), .Y(_abc_17692_n7752) );
  OR2X2 OR2X2_2481 ( .A(_abc_17692_n7746), .B(_abc_17692_n7752), .Y(_abc_17692_n7753) );
  OR2X2 OR2X2_2482 ( .A(_abc_17692_n7753), .B(_abc_17692_n7691), .Y(_abc_17692_n7754) );
  OR2X2 OR2X2_2483 ( .A(_abc_17692_n7765), .B(_abc_17692_n7763), .Y(_abc_17692_n7766) );
  OR2X2 OR2X2_2484 ( .A(_abc_17692_n7762), .B(_abc_17692_n7766), .Y(_abc_17692_n7767) );
  OR2X2 OR2X2_2485 ( .A(_abc_17692_n7761), .B(_abc_17692_n7767), .Y(_abc_17692_n7768) );
  OR2X2 OR2X2_2486 ( .A(_abc_17692_n7768), .B(_abc_17692_n7611), .Y(_abc_17692_n7771) );
  OR2X2 OR2X2_2487 ( .A(_abc_17692_n7758), .B(_abc_17692_n7773), .Y(_abc_17692_n7774) );
  OR2X2 OR2X2_2488 ( .A(_abc_17692_n7774), .B(_abc_17692_n7743), .Y(_abc_17692_n7775) );
  OR2X2 OR2X2_2489 ( .A(_abc_17692_n7775), .B(_abc_17692_n7726), .Y(_abc_17692_n7776) );
  OR2X2 OR2X2_249 ( .A(_abc_17692_n1175), .B(_abc_17692_n1177), .Y(_abc_17692_n1178) );
  OR2X2 OR2X2_2490 ( .A(_abc_17692_n7778), .B(_abc_17692_n7779), .Y(_abc_17692_n7780) );
  OR2X2 OR2X2_2491 ( .A(_abc_17692_n7777), .B(_abc_17692_n7780), .Y(_abc_17692_n7781) );
  OR2X2 OR2X2_2492 ( .A(_abc_17692_n7713), .B(_abc_17692_n7781), .Y(workunit2_28__FF_INPUT) );
  OR2X2 OR2X2_2493 ( .A(_abc_17692_n7547), .B(_abc_17692_n7543), .Y(_abc_17692_n7783) );
  OR2X2 OR2X2_2494 ( .A(_abc_17692_n7783), .B(_abc_17692_n7788), .Y(_abc_17692_n7789) );
  OR2X2 OR2X2_2495 ( .A(_abc_17692_n7638), .B(_abc_17692_n7641), .Y(_abc_17692_n7793) );
  OR2X2 OR2X2_2496 ( .A(sum_29_), .B(\key_in[93] ), .Y(_abc_17692_n7797) );
  OR2X2 OR2X2_2497 ( .A(_abc_17692_n7794), .B(_abc_17692_n7799), .Y(_abc_17692_n7802) );
  OR2X2 OR2X2_2498 ( .A(_abc_17692_n7803), .B(_abc_17692_n7792), .Y(_abc_17692_n7804) );
  OR2X2 OR2X2_2499 ( .A(_abc_17692_n7807), .B(_abc_17692_n7800), .Y(_abc_17692_n7808) );
  OR2X2 OR2X2_25 ( .A(_abc_17692_n629), .B(x_0_), .Y(_abc_17692_n669) );
  OR2X2 OR2X2_250 ( .A(_abc_17692_n1178), .B(_abc_17692_n1165), .Y(sum_10__FF_INPUT) );
  OR2X2 OR2X2_2500 ( .A(_abc_17692_n7808), .B(_abc_17692_n7805), .Y(_abc_17692_n7809) );
  OR2X2 OR2X2_2501 ( .A(_abc_17692_n7813), .B(_abc_17692_n7814), .Y(_abc_17692_n7815) );
  OR2X2 OR2X2_2502 ( .A(_abc_17692_n7811), .B(_abc_17692_n7816), .Y(_abc_17692_n7817) );
  OR2X2 OR2X2_2503 ( .A(_abc_17692_n7819), .B(_abc_17692_n7818), .Y(_abc_17692_n7820) );
  OR2X2 OR2X2_2504 ( .A(_abc_17692_n7821), .B(_abc_17692_n7817), .Y(_abc_17692_n7822) );
  OR2X2 OR2X2_2505 ( .A(_abc_17692_n7599), .B(_abc_17692_n7591), .Y(_abc_17692_n7825) );
  OR2X2 OR2X2_2506 ( .A(sum_29_), .B(\key_in[29] ), .Y(_abc_17692_n7829) );
  OR2X2 OR2X2_2507 ( .A(_abc_17692_n7832), .B(_abc_17692_n7833), .Y(_abc_17692_n7834) );
  OR2X2 OR2X2_2508 ( .A(_abc_17692_n7825), .B(_abc_17692_n7830), .Y(_abc_17692_n7836) );
  OR2X2 OR2X2_2509 ( .A(_abc_17692_n7835), .B(_abc_17692_n7839), .Y(_abc_17692_n7840) );
  OR2X2 OR2X2_251 ( .A(_abc_17692_n1180), .B(delta_11_), .Y(_abc_17692_n1183) );
  OR2X2 OR2X2_2510 ( .A(_abc_17692_n7840), .B(_abc_17692_n7812), .Y(_abc_17692_n7841) );
  OR2X2 OR2X2_2511 ( .A(_abc_17692_n7838), .B(_abc_17692_n7792), .Y(_abc_17692_n7842) );
  OR2X2 OR2X2_2512 ( .A(_abc_17692_n7834), .B(_abc_17692_n7805), .Y(_abc_17692_n7843) );
  OR2X2 OR2X2_2513 ( .A(_abc_17692_n7844), .B(workunit2_29_), .Y(_abc_17692_n7845) );
  OR2X2 OR2X2_2514 ( .A(_abc_17692_n7851), .B(_abc_17692_n7847), .Y(_abc_17692_n7852) );
  OR2X2 OR2X2_2515 ( .A(_abc_17692_n7850), .B(_abc_17692_n7846), .Y(_abc_17692_n7853) );
  OR2X2 OR2X2_2516 ( .A(_abc_17692_n7679), .B(_abc_17692_n7671), .Y(_abc_17692_n7856) );
  OR2X2 OR2X2_2517 ( .A(sum_29_), .B(\key_in[61] ), .Y(_abc_17692_n7860) );
  OR2X2 OR2X2_2518 ( .A(_abc_17692_n7863), .B(_abc_17692_n7864), .Y(_abc_17692_n7865) );
  OR2X2 OR2X2_2519 ( .A(_abc_17692_n7856), .B(_abc_17692_n7861), .Y(_abc_17692_n7867) );
  OR2X2 OR2X2_252 ( .A(_abc_17692_n1188), .B(_abc_17692_n1185), .Y(_abc_17692_n1189) );
  OR2X2 OR2X2_2520 ( .A(_abc_17692_n7866), .B(_abc_17692_n7870), .Y(_abc_17692_n7871) );
  OR2X2 OR2X2_2521 ( .A(_abc_17692_n7871), .B(_abc_17692_n7812), .Y(_abc_17692_n7872) );
  OR2X2 OR2X2_2522 ( .A(_abc_17692_n7869), .B(_abc_17692_n7792), .Y(_abc_17692_n7873) );
  OR2X2 OR2X2_2523 ( .A(_abc_17692_n7865), .B(_abc_17692_n7805), .Y(_abc_17692_n7874) );
  OR2X2 OR2X2_2524 ( .A(_abc_17692_n7875), .B(workunit2_29_), .Y(_abc_17692_n7876) );
  OR2X2 OR2X2_2525 ( .A(_abc_17692_n7880), .B(_abc_17692_n7877), .Y(_abc_17692_n7881) );
  OR2X2 OR2X2_2526 ( .A(_abc_17692_n7883), .B(_abc_17692_n7882), .Y(_abc_17692_n7884) );
  OR2X2 OR2X2_2527 ( .A(_abc_17692_n7886), .B(_abc_17692_n1863_bF_buf7), .Y(_abc_17692_n7887) );
  OR2X2 OR2X2_2528 ( .A(_abc_17692_n7887), .B(_abc_17692_n7855), .Y(_abc_17692_n7888) );
  OR2X2 OR2X2_2529 ( .A(_abc_17692_n7888), .B(_abc_17692_n7824), .Y(_abc_17692_n7889) );
  OR2X2 OR2X2_253 ( .A(_abc_17692_n1187), .B(_abc_17692_n1184), .Y(_abc_17692_n1190) );
  OR2X2 OR2X2_2530 ( .A(_abc_17692_n7559), .B(_abc_17692_n7551), .Y(_abc_17692_n7890) );
  OR2X2 OR2X2_2531 ( .A(sum_29_), .B(\key_in[125] ), .Y(_abc_17692_n7893) );
  OR2X2 OR2X2_2532 ( .A(_abc_17692_n7890), .B(_abc_17692_n7894), .Y(_abc_17692_n7895) );
  OR2X2 OR2X2_2533 ( .A(_abc_17692_n7896), .B(_abc_17692_n7897), .Y(_abc_17692_n7898) );
  OR2X2 OR2X2_2534 ( .A(_abc_17692_n7899), .B(_abc_17692_n7902), .Y(_abc_17692_n7903) );
  OR2X2 OR2X2_2535 ( .A(_abc_17692_n7903), .B(_abc_17692_n7812), .Y(_abc_17692_n7904) );
  OR2X2 OR2X2_2536 ( .A(_abc_17692_n7901), .B(_abc_17692_n7792), .Y(_abc_17692_n7905) );
  OR2X2 OR2X2_2537 ( .A(_abc_17692_n7898), .B(_abc_17692_n7805), .Y(_abc_17692_n7906) );
  OR2X2 OR2X2_2538 ( .A(_abc_17692_n7907), .B(workunit2_29_), .Y(_abc_17692_n7908) );
  OR2X2 OR2X2_2539 ( .A(_abc_17692_n7913), .B(_abc_17692_n7914), .Y(_abc_17692_n7915) );
  OR2X2 OR2X2_254 ( .A(_abc_17692_n1196), .B(_abc_17692_n1185), .Y(_abc_17692_n1197) );
  OR2X2 OR2X2_2540 ( .A(_abc_17692_n7916), .B(_abc_17692_n4047_bF_buf3), .Y(_abc_17692_n7917) );
  OR2X2 OR2X2_2541 ( .A(_abc_17692_n7917), .B(_abc_17692_n7912), .Y(_abc_17692_n7918) );
  OR2X2 OR2X2_2542 ( .A(_abc_17692_n7739), .B(_abc_17692_n7922), .Y(_abc_17692_n7923) );
  OR2X2 OR2X2_2543 ( .A(_abc_17692_n7926), .B(_abc_17692_n7924), .Y(_abc_17692_n7927) );
  OR2X2 OR2X2_2544 ( .A(_abc_17692_n7570), .B(_abc_17692_n7535), .Y(_abc_17692_n7929) );
  OR2X2 OR2X2_2545 ( .A(_abc_17692_n7723), .B(_abc_17692_n7930), .Y(_abc_17692_n7931) );
  OR2X2 OR2X2_2546 ( .A(_abc_17692_n7932), .B(_abc_17692_n7915), .Y(_abc_17692_n7933) );
  OR2X2 OR2X2_2547 ( .A(_abc_17692_n7931), .B(_abc_17692_n7909), .Y(_abc_17692_n7934) );
  OR2X2 OR2X2_2548 ( .A(_abc_17692_n7769), .B(_abc_17692_n7937), .Y(_abc_17692_n7938) );
  OR2X2 OR2X2_2549 ( .A(_abc_17692_n7939), .B(_abc_17692_n7847), .Y(_abc_17692_n7940) );
  OR2X2 OR2X2_255 ( .A(_abc_17692_n1198), .B(_abc_17692_n1184), .Y(_abc_17692_n1199) );
  OR2X2 OR2X2_2550 ( .A(_abc_17692_n7938), .B(_abc_17692_n7846), .Y(_abc_17692_n7941) );
  OR2X2 OR2X2_2551 ( .A(_abc_17692_n7755), .B(_abc_17692_n7944), .Y(_abc_17692_n7945) );
  OR2X2 OR2X2_2552 ( .A(_abc_17692_n7946), .B(_abc_17692_n7882), .Y(_abc_17692_n7947) );
  OR2X2 OR2X2_2553 ( .A(_abc_17692_n7945), .B(_abc_17692_n7877), .Y(_abc_17692_n7948) );
  OR2X2 OR2X2_2554 ( .A(_abc_17692_n7950), .B(_abc_17692_n7943), .Y(_abc_17692_n7951) );
  OR2X2 OR2X2_2555 ( .A(_abc_17692_n7936), .B(_abc_17692_n7951), .Y(_abc_17692_n7952) );
  OR2X2 OR2X2_2556 ( .A(_abc_17692_n7952), .B(_abc_17692_n7928), .Y(_abc_17692_n7953) );
  OR2X2 OR2X2_2557 ( .A(_abc_17692_n7955), .B(_abc_17692_n7956), .Y(_abc_17692_n7957) );
  OR2X2 OR2X2_2558 ( .A(_abc_17692_n7954), .B(_abc_17692_n7957), .Y(_abc_17692_n7958) );
  OR2X2 OR2X2_2559 ( .A(_abc_17692_n7958), .B(_abc_17692_n7920), .Y(workunit2_29__FF_INPUT) );
  OR2X2 OR2X2_256 ( .A(_abc_17692_n1201), .B(_abc_17692_n1193), .Y(_abc_17692_n1202) );
  OR2X2 OR2X2_2560 ( .A(_abc_17692_n7846), .B(_abc_17692_n7611), .Y(_abc_17692_n7960) );
  OR2X2 OR2X2_2561 ( .A(_abc_17692_n7624), .B(_abc_17692_n7960), .Y(_abc_17692_n7961) );
  OR2X2 OR2X2_2562 ( .A(_abc_17692_n7963), .B(_abc_17692_n7962), .Y(_abc_17692_n7964) );
  OR2X2 OR2X2_2563 ( .A(_abc_17692_n7970), .B(_abc_17692_n7969), .Y(_abc_17692_n7971) );
  OR2X2 OR2X2_2564 ( .A(_abc_17692_n7973), .B(_abc_17692_n7784), .Y(_abc_17692_n7974) );
  OR2X2 OR2X2_2565 ( .A(_abc_17692_n7974), .B(_abc_17692_n7972), .Y(_abc_17692_n7977) );
  OR2X2 OR2X2_2566 ( .A(sum_30_), .B(\key_in[30] ), .Y(_abc_17692_n7981) );
  OR2X2 OR2X2_2567 ( .A(_abc_17692_n7985), .B(_abc_17692_n7984), .Y(_abc_17692_n7986) );
  OR2X2 OR2X2_2568 ( .A(_abc_17692_n7986), .B(_abc_17692_n7983), .Y(_abc_17692_n7989) );
  OR2X2 OR2X2_2569 ( .A(_abc_17692_n7990), .B(_abc_17692_n7978), .Y(_abc_17692_n7991) );
  OR2X2 OR2X2_257 ( .A(_abc_17692_n1202), .B(_abc_17692_n1192_1), .Y(sum_11__FF_INPUT) );
  OR2X2 OR2X2_2570 ( .A(_abc_17692_n7992), .B(_abc_17692_n7993), .Y(_abc_17692_n7994) );
  OR2X2 OR2X2_2571 ( .A(_abc_17692_n7994), .B(_abc_17692_n7968), .Y(_abc_17692_n7995) );
  OR2X2 OR2X2_2572 ( .A(_abc_17692_n7997), .B(workunit2_30_), .Y(_abc_17692_n7998) );
  OR2X2 OR2X2_2573 ( .A(_abc_17692_n7967), .B(_abc_17692_n8000), .Y(_abc_17692_n8001) );
  OR2X2 OR2X2_2574 ( .A(_abc_17692_n7966), .B(_abc_17692_n7999), .Y(_abc_17692_n8002) );
  OR2X2 OR2X2_2575 ( .A(_abc_17692_n8008), .B(_abc_17692_n8007), .Y(_abc_17692_n8009) );
  OR2X2 OR2X2_2576 ( .A(_abc_17692_n8006), .B(_abc_17692_n8009), .Y(_abc_17692_n8010) );
  OR2X2 OR2X2_2577 ( .A(sum_30_), .B(\key_in[94] ), .Y(_abc_17692_n8014) );
  OR2X2 OR2X2_2578 ( .A(_abc_17692_n8018), .B(_abc_17692_n8017), .Y(_abc_17692_n8019) );
  OR2X2 OR2X2_2579 ( .A(_abc_17692_n8019), .B(_abc_17692_n8016), .Y(_abc_17692_n8022) );
  OR2X2 OR2X2_258 ( .A(_abc_17692_n1207), .B(_abc_17692_n1204), .Y(_abc_17692_n1208) );
  OR2X2 OR2X2_2580 ( .A(_abc_17692_n8025), .B(_abc_17692_n8026), .Y(_abc_17692_n8027) );
  OR2X2 OR2X2_2581 ( .A(_abc_17692_n8027), .B(workunit2_30_), .Y(_abc_17692_n8028) );
  OR2X2 OR2X2_2582 ( .A(_abc_17692_n8029), .B(_abc_17692_n7968), .Y(_abc_17692_n8030) );
  OR2X2 OR2X2_2583 ( .A(_abc_17692_n8010), .B(_abc_17692_n8031), .Y(_abc_17692_n8032) );
  OR2X2 OR2X2_2584 ( .A(_abc_17692_n7877), .B(_abc_17692_n7691), .Y(_abc_17692_n8037) );
  OR2X2 OR2X2_2585 ( .A(_abc_17692_n7702), .B(_abc_17692_n8037), .Y(_abc_17692_n8038) );
  OR2X2 OR2X2_2586 ( .A(_abc_17692_n7877), .B(_abc_17692_n7879), .Y(_abc_17692_n8041) );
  OR2X2 OR2X2_2587 ( .A(sum_30_), .B(\key_in[62] ), .Y(_abc_17692_n8047) );
  OR2X2 OR2X2_2588 ( .A(_abc_17692_n8051), .B(_abc_17692_n8050), .Y(_abc_17692_n8052) );
  OR2X2 OR2X2_2589 ( .A(_abc_17692_n8052), .B(_abc_17692_n8049), .Y(_abc_17692_n8055) );
  OR2X2 OR2X2_259 ( .A(_abc_17692_n1156), .B(_abc_17692_n1211), .Y(_abc_17692_n1212) );
  OR2X2 OR2X2_2590 ( .A(_abc_17692_n8056), .B(_abc_17692_n8011), .Y(_abc_17692_n8057) );
  OR2X2 OR2X2_2591 ( .A(_abc_17692_n8058), .B(_abc_17692_n7978), .Y(_abc_17692_n8059) );
  OR2X2 OR2X2_2592 ( .A(_abc_17692_n8060), .B(_abc_17692_n7968), .Y(_abc_17692_n8061) );
  OR2X2 OR2X2_2593 ( .A(_abc_17692_n8058), .B(_abc_17692_n8011), .Y(_abc_17692_n8062) );
  OR2X2 OR2X2_2594 ( .A(_abc_17692_n8056), .B(_abc_17692_n7978), .Y(_abc_17692_n8063) );
  OR2X2 OR2X2_2595 ( .A(_abc_17692_n8064), .B(workunit2_30_), .Y(_abc_17692_n8065) );
  OR2X2 OR2X2_2596 ( .A(_abc_17692_n8044), .B(_abc_17692_n8067), .Y(_abc_17692_n8068) );
  OR2X2 OR2X2_2597 ( .A(_abc_17692_n8043), .B(_abc_17692_n8066), .Y(_abc_17692_n8069) );
  OR2X2 OR2X2_2598 ( .A(_abc_17692_n8071), .B(_abc_17692_n1863_bF_buf5), .Y(_abc_17692_n8072) );
  OR2X2 OR2X2_2599 ( .A(_abc_17692_n8036), .B(_abc_17692_n8072), .Y(_abc_17692_n8073) );
  OR2X2 OR2X2_26 ( .A(_abc_17692_n667), .B(x_1_), .Y(_abc_17692_n673) );
  OR2X2 OR2X2_260 ( .A(_abc_17692_n1211), .B(_abc_17692_n1158), .Y(_abc_17692_n1213) );
  OR2X2 OR2X2_2600 ( .A(_abc_17692_n8073), .B(_abc_17692_n8004), .Y(_abc_17692_n8074) );
  OR2X2 OR2X2_2601 ( .A(_abc_17692_n7584), .B(_abc_17692_n8076), .Y(_abc_17692_n8077) );
  OR2X2 OR2X2_2602 ( .A(_abc_17692_n7909), .B(_abc_17692_n7569), .Y(_abc_17692_n8080) );
  OR2X2 OR2X2_2603 ( .A(sum_30_), .B(\key_in[126] ), .Y(_abc_17692_n8086) );
  OR2X2 OR2X2_2604 ( .A(_abc_17692_n7890), .B(_abc_17692_n7891), .Y(_abc_17692_n8089) );
  OR2X2 OR2X2_2605 ( .A(_abc_17692_n8092), .B(_abc_17692_n8093), .Y(_abc_17692_n8094) );
  OR2X2 OR2X2_2606 ( .A(_abc_17692_n8097), .B(_abc_17692_n8095), .Y(_abc_17692_n8098) );
  OR2X2 OR2X2_2607 ( .A(_abc_17692_n8099), .B(_abc_17692_n7968), .Y(_abc_17692_n8100) );
  OR2X2 OR2X2_2608 ( .A(_abc_17692_n8098), .B(workunit2_30_), .Y(_abc_17692_n8101) );
  OR2X2 OR2X2_2609 ( .A(_abc_17692_n8083), .B(_abc_17692_n8102), .Y(_abc_17692_n8103) );
  OR2X2 OR2X2_261 ( .A(_abc_17692_n1214), .B(_abc_17692_n1215), .Y(_abc_17692_n1216) );
  OR2X2 OR2X2_2610 ( .A(_abc_17692_n8098), .B(_abc_17692_n7968), .Y(_abc_17692_n8104) );
  OR2X2 OR2X2_2611 ( .A(_abc_17692_n8099), .B(workunit2_30_), .Y(_abc_17692_n8105) );
  OR2X2 OR2X2_2612 ( .A(_abc_17692_n8082), .B(_abc_17692_n8106), .Y(_abc_17692_n8107) );
  OR2X2 OR2X2_2613 ( .A(_abc_17692_n8108), .B(_abc_17692_n4047_bF_buf2), .Y(_abc_17692_n8109) );
  OR2X2 OR2X2_2614 ( .A(_abc_17692_n8114), .B(_abc_17692_n7914), .Y(_abc_17692_n8115) );
  OR2X2 OR2X2_2615 ( .A(_abc_17692_n8113), .B(_abc_17692_n8116), .Y(_abc_17692_n8117) );
  OR2X2 OR2X2_2616 ( .A(_abc_17692_n8117), .B(_abc_17692_n8106), .Y(_abc_17692_n8118) );
  OR2X2 OR2X2_2617 ( .A(_abc_17692_n6605), .B(_abc_17692_n6398), .Y(_abc_17692_n8126) );
  OR2X2 OR2X2_2618 ( .A(_abc_17692_n8126), .B(_abc_17692_n8125), .Y(_abc_17692_n8127) );
  OR2X2 OR2X2_2619 ( .A(_abc_17692_n8127), .B(_abc_17692_n8124), .Y(_abc_17692_n8128) );
  OR2X2 OR2X2_262 ( .A(_abc_17692_n1220), .B(_abc_17692_n1209), .Y(_abc_17692_n1221) );
  OR2X2 OR2X2_2620 ( .A(_abc_17692_n8128), .B(_abc_17692_n8123), .Y(_abc_17692_n8129) );
  OR2X2 OR2X2_2621 ( .A(_abc_17692_n7390), .B(_abc_17692_n7292), .Y(_abc_17692_n8132) );
  OR2X2 OR2X2_2622 ( .A(_abc_17692_n8132), .B(_abc_17692_n8131), .Y(_abc_17692_n8133) );
  OR2X2 OR2X2_2623 ( .A(_abc_17692_n8130), .B(_abc_17692_n8133), .Y(_abc_17692_n8134) );
  OR2X2 OR2X2_2624 ( .A(_abc_17692_n8132), .B(_abc_17692_n7300), .Y(_abc_17692_n8135) );
  OR2X2 OR2X2_2625 ( .A(_abc_17692_n7915), .B(_abc_17692_n7572), .Y(_abc_17692_n8139) );
  OR2X2 OR2X2_2626 ( .A(_abc_17692_n8138), .B(_abc_17692_n8139), .Y(_abc_17692_n8140) );
  OR2X2 OR2X2_2627 ( .A(_abc_17692_n8141), .B(_abc_17692_n8102), .Y(_abc_17692_n8142) );
  OR2X2 OR2X2_2628 ( .A(_abc_17692_n7817), .B(_abc_17692_n7651), .Y(_abc_17692_n8146) );
  OR2X2 OR2X2_2629 ( .A(_abc_17692_n7737), .B(_abc_17692_n8146), .Y(_abc_17692_n8147) );
  OR2X2 OR2X2_263 ( .A(_abc_17692_n1219), .B(_abc_17692_n1208), .Y(_abc_17692_n1222) );
  OR2X2 OR2X2_2630 ( .A(_abc_17692_n7811), .B(_abc_17692_n7922), .Y(_abc_17692_n8149) );
  OR2X2 OR2X2_2631 ( .A(_abc_17692_n8153), .B(_abc_17692_n8145), .Y(_abc_17692_n8154) );
  OR2X2 OR2X2_2632 ( .A(_abc_17692_n8152), .B(_abc_17692_n8031), .Y(_abc_17692_n8155) );
  OR2X2 OR2X2_2633 ( .A(_abc_17692_n8161), .B(_abc_17692_n8160), .Y(_abc_17692_n8162) );
  OR2X2 OR2X2_2634 ( .A(_abc_17692_n8159), .B(_abc_17692_n8162), .Y(_abc_17692_n8163) );
  OR2X2 OR2X2_2635 ( .A(_abc_17692_n8163), .B(_abc_17692_n8066), .Y(_abc_17692_n8166) );
  OR2X2 OR2X2_2636 ( .A(_abc_17692_n8172), .B(_abc_17692_n8171), .Y(_abc_17692_n8173) );
  OR2X2 OR2X2_2637 ( .A(_abc_17692_n8170), .B(_abc_17692_n8173), .Y(_abc_17692_n8174) );
  OR2X2 OR2X2_2638 ( .A(_abc_17692_n8174), .B(_abc_17692_n7999), .Y(_abc_17692_n8177) );
  OR2X2 OR2X2_2639 ( .A(_abc_17692_n8168), .B(_abc_17692_n8179), .Y(_abc_17692_n8180) );
  OR2X2 OR2X2_264 ( .A(_abc_17692_n1185), .B(_abc_17692_n1195_1), .Y(_abc_17692_n1228) );
  OR2X2 OR2X2_2640 ( .A(_abc_17692_n8180), .B(_abc_17692_n8157), .Y(_abc_17692_n8181) );
  OR2X2 OR2X2_2641 ( .A(_abc_17692_n8181), .B(_abc_17692_n8144), .Y(_abc_17692_n8182) );
  OR2X2 OR2X2_2642 ( .A(_abc_17692_n8184), .B(_abc_17692_n8185), .Y(_abc_17692_n8186) );
  OR2X2 OR2X2_2643 ( .A(_abc_17692_n8183), .B(_abc_17692_n8186), .Y(_abc_17692_n8187) );
  OR2X2 OR2X2_2644 ( .A(_abc_17692_n8111), .B(_abc_17692_n8187), .Y(workunit2_30__FF_INPUT) );
  OR2X2 OR2X2_2645 ( .A(_abc_17692_n1792), .B(\key_in[127] ), .Y(_abc_17692_n8193) );
  OR2X2 OR2X2_2646 ( .A(_abc_17692_n8194), .B(sum_31_), .Y(_abc_17692_n8195) );
  OR2X2 OR2X2_2647 ( .A(_abc_17692_n8192), .B(_abc_17692_n8197), .Y(_abc_17692_n8200) );
  OR2X2 OR2X2_2648 ( .A(_abc_17692_n7975), .B(_abc_17692_n7969), .Y(_abc_17692_n8203) );
  OR2X2 OR2X2_2649 ( .A(_abc_17692_n8206), .B(_abc_17692_n8205), .Y(_abc_17692_n8207) );
  OR2X2 OR2X2_265 ( .A(_abc_17692_n1234), .B(_abc_17692_n1208), .Y(_abc_17692_n1237) );
  OR2X2 OR2X2_2650 ( .A(_abc_17692_n8204), .B(_abc_17692_n8207), .Y(_abc_17692_n8210) );
  OR2X2 OR2X2_2651 ( .A(_abc_17692_n8211), .B(_abc_17692_n8202), .Y(_abc_17692_n8213) );
  OR2X2 OR2X2_2652 ( .A(_abc_17692_n8214), .B(_abc_17692_n8212), .Y(_abc_17692_n8215) );
  OR2X2 OR2X2_2653 ( .A(_abc_17692_n8201), .B(_abc_17692_n8215), .Y(_abc_17692_n8216) );
  OR2X2 OR2X2_2654 ( .A(_abc_17692_n8217), .B(_abc_17692_n8218), .Y(_abc_17692_n8219) );
  OR2X2 OR2X2_2655 ( .A(_abc_17692_n8223), .B(_abc_17692_n4047_bF_buf1), .Y(_abc_17692_n8224) );
  OR2X2 OR2X2_2656 ( .A(_abc_17692_n8224), .B(_abc_17692_n8222), .Y(_abc_17692_n8225) );
  OR2X2 OR2X2_2657 ( .A(_abc_17692_n8033), .B(_abc_17692_n8226), .Y(_abc_17692_n8227) );
  OR2X2 OR2X2_2658 ( .A(_abc_17692_n1792), .B(\key_in[95] ), .Y(_abc_17692_n8230) );
  OR2X2 OR2X2_2659 ( .A(_abc_17692_n8231), .B(sum_31_), .Y(_abc_17692_n8232) );
  OR2X2 OR2X2_266 ( .A(_abc_17692_n1240), .B(state_8_bF_buf2), .Y(_abc_17692_n1241_1) );
  OR2X2 OR2X2_2660 ( .A(_abc_17692_n8229), .B(_abc_17692_n8234), .Y(_abc_17692_n8237) );
  OR2X2 OR2X2_2661 ( .A(_abc_17692_n8215), .B(_abc_17692_n8238), .Y(_abc_17692_n8239) );
  OR2X2 OR2X2_2662 ( .A(_abc_17692_n8218), .B(_abc_17692_n8240), .Y(_abc_17692_n8241) );
  OR2X2 OR2X2_2663 ( .A(_abc_17692_n8228), .B(_abc_17692_n8243), .Y(_abc_17692_n8244) );
  OR2X2 OR2X2_2664 ( .A(_abc_17692_n8227), .B(_abc_17692_n8242), .Y(_abc_17692_n8245) );
  OR2X2 OR2X2_2665 ( .A(_abc_17692_n1792), .B(\key_in[31] ), .Y(_abc_17692_n8253) );
  OR2X2 OR2X2_2666 ( .A(_abc_17692_n8254), .B(sum_31_), .Y(_abc_17692_n8255) );
  OR2X2 OR2X2_2667 ( .A(_abc_17692_n8252), .B(_abc_17692_n8257), .Y(_abc_17692_n8260) );
  OR2X2 OR2X2_2668 ( .A(_abc_17692_n8218), .B(_abc_17692_n8261), .Y(_abc_17692_n8262) );
  OR2X2 OR2X2_2669 ( .A(_abc_17692_n8215), .B(_abc_17692_n8263), .Y(_abc_17692_n8264) );
  OR2X2 OR2X2_267 ( .A(_abc_17692_n1239), .B(_abc_17692_n1241_1), .Y(_abc_17692_n1242) );
  OR2X2 OR2X2_2670 ( .A(_abc_17692_n8251), .B(_abc_17692_n8266), .Y(_abc_17692_n8267) );
  OR2X2 OR2X2_2671 ( .A(_abc_17692_n8250), .B(_abc_17692_n8265), .Y(_abc_17692_n8268) );
  OR2X2 OR2X2_2672 ( .A(_abc_17692_n1792), .B(\key_in[63] ), .Y(_abc_17692_n8276) );
  OR2X2 OR2X2_2673 ( .A(_abc_17692_n8277), .B(sum_31_), .Y(_abc_17692_n8278) );
  OR2X2 OR2X2_2674 ( .A(_abc_17692_n8275), .B(_abc_17692_n8280), .Y(_abc_17692_n8283) );
  OR2X2 OR2X2_2675 ( .A(_abc_17692_n8218), .B(_abc_17692_n8284), .Y(_abc_17692_n8285) );
  OR2X2 OR2X2_2676 ( .A(_abc_17692_n8215), .B(_abc_17692_n8286), .Y(_abc_17692_n8287) );
  OR2X2 OR2X2_2677 ( .A(_abc_17692_n8274), .B(_abc_17692_n8289), .Y(_abc_17692_n8290) );
  OR2X2 OR2X2_2678 ( .A(_abc_17692_n8273), .B(_abc_17692_n8288), .Y(_abc_17692_n8291) );
  OR2X2 OR2X2_2679 ( .A(_abc_17692_n8293), .B(_abc_17692_n1863_bF_buf3), .Y(_abc_17692_n8294) );
  OR2X2 OR2X2_268 ( .A(_abc_17692_n1242), .B(_abc_17692_n1224), .Y(sum_12__FF_INPUT) );
  OR2X2 OR2X2_2680 ( .A(_abc_17692_n8294), .B(_abc_17692_n8270), .Y(_abc_17692_n8295) );
  OR2X2 OR2X2_2681 ( .A(_abc_17692_n8295), .B(_abc_17692_n8247), .Y(_abc_17692_n8296) );
  OR2X2 OR2X2_2682 ( .A(_abc_17692_n8302), .B(_abc_17692_n8301), .Y(_abc_17692_n8303) );
  OR2X2 OR2X2_2683 ( .A(_abc_17692_n8300), .B(_abc_17692_n8304), .Y(_abc_17692_n8305) );
  OR2X2 OR2X2_2684 ( .A(_abc_17692_n8310), .B(_abc_17692_n8243), .Y(_abc_17692_n8311) );
  OR2X2 OR2X2_2685 ( .A(_abc_17692_n8309), .B(_abc_17692_n8242), .Y(_abc_17692_n8312) );
  OR2X2 OR2X2_2686 ( .A(_abc_17692_n8164), .B(_abc_17692_n8315), .Y(_abc_17692_n8316) );
  OR2X2 OR2X2_2687 ( .A(_abc_17692_n8317), .B(_abc_17692_n8289), .Y(_abc_17692_n8318) );
  OR2X2 OR2X2_2688 ( .A(_abc_17692_n8316), .B(_abc_17692_n8288), .Y(_abc_17692_n8319) );
  OR2X2 OR2X2_2689 ( .A(_abc_17692_n8175), .B(_abc_17692_n8322), .Y(_abc_17692_n8323) );
  OR2X2 OR2X2_269 ( .A(_abc_17692_n1253), .B(_abc_17692_n1251), .Y(_abc_17692_n1254) );
  OR2X2 OR2X2_2690 ( .A(_abc_17692_n8324), .B(_abc_17692_n8266), .Y(_abc_17692_n8325) );
  OR2X2 OR2X2_2691 ( .A(_abc_17692_n8323), .B(_abc_17692_n8265), .Y(_abc_17692_n8326) );
  OR2X2 OR2X2_2692 ( .A(_abc_17692_n8321), .B(_abc_17692_n8328), .Y(_abc_17692_n8329) );
  OR2X2 OR2X2_2693 ( .A(_abc_17692_n8329), .B(_abc_17692_n8314), .Y(_abc_17692_n8330) );
  OR2X2 OR2X2_2694 ( .A(_abc_17692_n8330), .B(_abc_17692_n8306), .Y(_abc_17692_n8331) );
  OR2X2 OR2X2_2695 ( .A(_abc_17692_n8333), .B(_abc_17692_n8334), .Y(_abc_17692_n8335) );
  OR2X2 OR2X2_2696 ( .A(_abc_17692_n8332), .B(_abc_17692_n8335), .Y(_abc_17692_n8336) );
  OR2X2 OR2X2_2697 ( .A(_abc_17692_n8336), .B(_abc_17692_n8298), .Y(workunit2_31__FF_INPUT) );
  OR2X2 OR2X2_2698 ( .A(_abc_17692_n8340), .B(_abc_17692_n8339), .Y(_abc_17692_n8341) );
  OR2X2 OR2X2_2699 ( .A(_abc_17692_n8344), .B(_abc_17692_n8342), .Y(_abc_17692_n8345) );
  OR2X2 OR2X2_27 ( .A(_abc_17692_n671), .B(x_2_), .Y(_abc_17692_n677_1) );
  OR2X2 OR2X2_270 ( .A(_abc_17692_n1255), .B(_abc_17692_n1250), .Y(_abc_17692_n1256) );
  OR2X2 OR2X2_2700 ( .A(_abc_17692_n8346), .B(workunit1_0_), .Y(_abc_17692_n8349) );
  OR2X2 OR2X2_2701 ( .A(_abc_17692_n8353), .B(_abc_17692_n8352), .Y(_abc_17692_n8354) );
  OR2X2 OR2X2_2702 ( .A(_abc_17692_n8355), .B(workunit1_0_), .Y(_abc_17692_n8356) );
  OR2X2 OR2X2_2703 ( .A(_abc_17692_n8360), .B(_abc_17692_n8351), .Y(_abc_17692_n8361) );
  OR2X2 OR2X2_2704 ( .A(_abc_17692_n8363), .B(_abc_17692_n8362), .Y(_abc_17692_n8364) );
  OR2X2 OR2X2_2705 ( .A(_abc_17692_n8365), .B(workunit1_0_), .Y(_abc_17692_n8368) );
  OR2X2 OR2X2_2706 ( .A(_abc_17692_n8372), .B(_abc_17692_n8371), .Y(_abc_17692_n8373) );
  OR2X2 OR2X2_2707 ( .A(_abc_17692_n8374), .B(workunit1_0_), .Y(_abc_17692_n8375) );
  OR2X2 OR2X2_2708 ( .A(_abc_17692_n8379), .B(_abc_17692_n8370), .Y(_abc_17692_n8380) );
  OR2X2 OR2X2_2709 ( .A(_abc_17692_n8361), .B(_abc_17692_n8380), .Y(_abc_17692_n8381) );
  OR2X2 OR2X2_271 ( .A(_abc_17692_n1251), .B(_abc_17692_n1259), .Y(_abc_17692_n1260) );
  OR2X2 OR2X2_2710 ( .A(_abc_17692_n8384), .B(_abc_17692_n8385), .Y(_abc_17692_n8386) );
  OR2X2 OR2X2_2711 ( .A(_abc_17692_n8382), .B(_abc_17692_n8386), .Y(workunit1_0__FF_INPUT) );
  OR2X2 OR2X2_2712 ( .A(workunit2_1_bF_buf3), .B(workunit2_6_), .Y(_abc_17692_n8392) );
  OR2X2 OR2X2_2713 ( .A(_abc_17692_n8396), .B(_abc_17692_n8390), .Y(_abc_17692_n8397) );
  OR2X2 OR2X2_2714 ( .A(_abc_17692_n8398), .B(_abc_17692_n8394), .Y(_abc_17692_n8399) );
  OR2X2 OR2X2_2715 ( .A(_abc_17692_n8397), .B(_abc_17692_n8395), .Y(_abc_17692_n8401) );
  OR2X2 OR2X2_2716 ( .A(_abc_17692_n8393), .B(_abc_17692_n8339), .Y(_abc_17692_n8402) );
  OR2X2 OR2X2_2717 ( .A(_abc_17692_n8400), .B(_abc_17692_n8404), .Y(_abc_17692_n8405) );
  OR2X2 OR2X2_2718 ( .A(_abc_17692_n8405), .B(workunit1_1_bF_buf0), .Y(_abc_17692_n8408) );
  OR2X2 OR2X2_2719 ( .A(_abc_17692_n8410), .B(_abc_17692_n8389), .Y(_abc_17692_n8413) );
  OR2X2 OR2X2_272 ( .A(_abc_17692_n1235), .B(_abc_17692_n1260), .Y(_abc_17692_n1261) );
  OR2X2 OR2X2_2720 ( .A(_abc_17692_n1915), .B(_abc_17692_n8403), .Y(_abc_17692_n8416) );
  OR2X2 OR2X2_2721 ( .A(_abc_17692_n1908), .B(_abc_17692_n8399), .Y(_abc_17692_n8417) );
  OR2X2 OR2X2_2722 ( .A(_abc_17692_n1908), .B(_abc_17692_n8403), .Y(_abc_17692_n8420) );
  OR2X2 OR2X2_2723 ( .A(_abc_17692_n1915), .B(_abc_17692_n8399), .Y(_abc_17692_n8421) );
  OR2X2 OR2X2_2724 ( .A(_abc_17692_n8419), .B(_abc_17692_n8423), .Y(_abc_17692_n8424) );
  OR2X2 OR2X2_2725 ( .A(_abc_17692_n8424), .B(_abc_17692_n8426), .Y(_abc_17692_n8427) );
  OR2X2 OR2X2_2726 ( .A(_abc_17692_n8434), .B(_abc_17692_n8435), .Y(_abc_17692_n8436) );
  OR2X2 OR2X2_2727 ( .A(_abc_17692_n8436), .B(workunit1_1_bF_buf1), .Y(_abc_17692_n8439) );
  OR2X2 OR2X2_2728 ( .A(_abc_17692_n8441), .B(_abc_17692_n8433), .Y(_abc_17692_n8442) );
  OR2X2 OR2X2_2729 ( .A(_abc_17692_n8440), .B(_abc_17692_n8432), .Y(_abc_17692_n8443) );
  OR2X2 OR2X2_273 ( .A(_abc_17692_n1270), .B(state_8_bF_buf1), .Y(_abc_17692_n1271) );
  OR2X2 OR2X2_2730 ( .A(_abc_17692_n8431), .B(_abc_17692_n8445), .Y(_abc_17692_n8446) );
  OR2X2 OR2X2_2731 ( .A(_abc_17692_n8446), .B(_abc_17692_n8415), .Y(_abc_17692_n8447) );
  OR2X2 OR2X2_2732 ( .A(_abc_17692_n2007), .B(_abc_17692_n8403), .Y(_abc_17692_n8450) );
  OR2X2 OR2X2_2733 ( .A(_abc_17692_n8453), .B(_abc_17692_n2637), .Y(_abc_17692_n8454) );
  OR2X2 OR2X2_2734 ( .A(_abc_17692_n8455), .B(_abc_17692_n8451), .Y(_abc_17692_n8456) );
  OR2X2 OR2X2_2735 ( .A(_abc_17692_n8456), .B(workunit1_1_bF_buf0), .Y(_abc_17692_n8457) );
  OR2X2 OR2X2_2736 ( .A(_abc_17692_n8459), .B(_abc_17692_n8449), .Y(_abc_17692_n8462) );
  OR2X2 OR2X2_2737 ( .A(_abc_17692_n8447), .B(_abc_17692_n8464), .Y(_abc_17692_n8465) );
  OR2X2 OR2X2_2738 ( .A(_abc_17692_n8467), .B(_abc_17692_n8376), .Y(_abc_17692_n8468) );
  OR2X2 OR2X2_2739 ( .A(_abc_17692_n8424), .B(_abc_17692_n8377), .Y(_abc_17692_n8469) );
  OR2X2 OR2X2_274 ( .A(_abc_17692_n1269), .B(_abc_17692_n1271), .Y(_abc_17692_n1272) );
  OR2X2 OR2X2_2740 ( .A(_abc_17692_n8409), .B(_abc_17692_n8347), .Y(_abc_17692_n8474) );
  OR2X2 OR2X2_2741 ( .A(_abc_17692_n8476), .B(_abc_17692_n8471), .Y(_abc_17692_n8477) );
  OR2X2 OR2X2_2742 ( .A(_abc_17692_n8458), .B(_abc_17692_n8366), .Y(_abc_17692_n8480) );
  OR2X2 OR2X2_2743 ( .A(_abc_17692_n8440), .B(_abc_17692_n8357), .Y(_abc_17692_n8485) );
  OR2X2 OR2X2_2744 ( .A(_abc_17692_n8482), .B(_abc_17692_n8487), .Y(_abc_17692_n8488) );
  OR2X2 OR2X2_2745 ( .A(_abc_17692_n8477), .B(_abc_17692_n8488), .Y(_abc_17692_n8489) );
  OR2X2 OR2X2_2746 ( .A(_abc_17692_n8491), .B(_abc_17692_n8492), .Y(_abc_17692_n8493) );
  OR2X2 OR2X2_2747 ( .A(_abc_17692_n8490), .B(_abc_17692_n8493), .Y(_abc_17692_n8494) );
  OR2X2 OR2X2_2748 ( .A(_abc_17692_n8466), .B(_abc_17692_n8494), .Y(workunit1_1__FF_INPUT) );
  OR2X2 OR2X2_2749 ( .A(_abc_17692_n8498), .B(_abc_17692_n8497), .Y(_abc_17692_n8499) );
  OR2X2 OR2X2_275 ( .A(_abc_17692_n1258_1), .B(_abc_17692_n1272), .Y(sum_13__FF_INPUT) );
  OR2X2 OR2X2_2750 ( .A(_abc_17692_n8496), .B(_abc_17692_n8499), .Y(_abc_17692_n8500) );
  OR2X2 OR2X2_2751 ( .A(_abc_17692_n8394), .B(_abc_17692_n8390), .Y(_abc_17692_n8501) );
  OR2X2 OR2X2_2752 ( .A(_abc_17692_n8501), .B(_abc_17692_n8502), .Y(_abc_17692_n8503) );
  OR2X2 OR2X2_2753 ( .A(_abc_17692_n2087_1), .B(_abc_17692_n8504), .Y(_abc_17692_n8505) );
  OR2X2 OR2X2_2754 ( .A(_abc_17692_n8507), .B(_abc_17692_n8506), .Y(_abc_17692_n8508) );
  OR2X2 OR2X2_2755 ( .A(_abc_17692_n2080), .B(_abc_17692_n8508), .Y(_abc_17692_n8509) );
  OR2X2 OR2X2_2756 ( .A(_abc_17692_n8510), .B(workunit1_2_), .Y(_abc_17692_n8511) );
  OR2X2 OR2X2_2757 ( .A(_abc_17692_n2087_1), .B(_abc_17692_n8508), .Y(_abc_17692_n8512) );
  OR2X2 OR2X2_2758 ( .A(_abc_17692_n2080), .B(_abc_17692_n8504), .Y(_abc_17692_n8513) );
  OR2X2 OR2X2_2759 ( .A(_abc_17692_n8514), .B(_abc_17692_n2062_1), .Y(_abc_17692_n8515) );
  OR2X2 OR2X2_276 ( .A(_abc_17692_n1274), .B(delta_14_), .Y(_abc_17692_n1276) );
  OR2X2 OR2X2_2760 ( .A(_abc_17692_n8428), .B(_abc_17692_n8517), .Y(_abc_17692_n8518) );
  OR2X2 OR2X2_2761 ( .A(_abc_17692_n8518), .B(_abc_17692_n8516), .Y(_abc_17692_n8521) );
  OR2X2 OR2X2_2762 ( .A(_abc_17692_n8528), .B(_abc_17692_n2062_1), .Y(_abc_17692_n8529) );
  OR2X2 OR2X2_2763 ( .A(_abc_17692_n8524), .B(_abc_17692_n8526), .Y(_abc_17692_n8530) );
  OR2X2 OR2X2_2764 ( .A(_abc_17692_n8530), .B(workunit1_2_), .Y(_abc_17692_n8531) );
  OR2X2 OR2X2_2765 ( .A(_abc_17692_n8540), .B(_abc_17692_n8533), .Y(_abc_17692_n8541) );
  OR2X2 OR2X2_2766 ( .A(_abc_17692_n8539), .B(_abc_17692_n8532), .Y(_abc_17692_n8542) );
  OR2X2 OR2X2_2767 ( .A(_abc_17692_n8545), .B(_abc_17692_n8546), .Y(_abc_17692_n8547) );
  OR2X2 OR2X2_2768 ( .A(_abc_17692_n8547), .B(workunit1_2_), .Y(_abc_17692_n8550) );
  OR2X2 OR2X2_2769 ( .A(_abc_17692_n8411), .B(_abc_17692_n8554), .Y(_abc_17692_n8555) );
  OR2X2 OR2X2_277 ( .A(_abc_17692_n1277), .B(_abc_17692_n1275), .Y(_abc_17692_n1278) );
  OR2X2 OR2X2_2770 ( .A(_abc_17692_n8552), .B(_abc_17692_n8555), .Y(_abc_17692_n8558) );
  OR2X2 OR2X2_2771 ( .A(_abc_17692_n8560), .B(_abc_17692_n8544), .Y(_abc_17692_n8561) );
  OR2X2 OR2X2_2772 ( .A(_abc_17692_n8561), .B(_abc_17692_n8523), .Y(_abc_17692_n8562) );
  OR2X2 OR2X2_2773 ( .A(_abc_17692_n2182), .B(_abc_17692_n8504), .Y(_abc_17692_n8563) );
  OR2X2 OR2X2_2774 ( .A(_abc_17692_n2177), .B(_abc_17692_n8508), .Y(_abc_17692_n8564) );
  OR2X2 OR2X2_2775 ( .A(_abc_17692_n8565), .B(_abc_17692_n2062_1), .Y(_abc_17692_n8566) );
  OR2X2 OR2X2_2776 ( .A(_abc_17692_n2177), .B(_abc_17692_n8504), .Y(_abc_17692_n8567) );
  OR2X2 OR2X2_2777 ( .A(_abc_17692_n2182), .B(_abc_17692_n8508), .Y(_abc_17692_n8568) );
  OR2X2 OR2X2_2778 ( .A(_abc_17692_n8569), .B(workunit1_2_), .Y(_abc_17692_n8570) );
  OR2X2 OR2X2_2779 ( .A(_abc_17692_n8460), .B(_abc_17692_n8573), .Y(_abc_17692_n8574) );
  OR2X2 OR2X2_278 ( .A(_abc_17692_n1222), .B(_abc_17692_n1251), .Y(_abc_17692_n1279) );
  OR2X2 OR2X2_2780 ( .A(_abc_17692_n8574), .B(_abc_17692_n8572), .Y(_abc_17692_n8577) );
  OR2X2 OR2X2_2781 ( .A(_abc_17692_n8562), .B(_abc_17692_n8579), .Y(_abc_17692_n8580) );
  OR2X2 OR2X2_2782 ( .A(_abc_17692_n8585), .B(_abc_17692_n8582), .Y(_abc_17692_n8586) );
  OR2X2 OR2X2_2783 ( .A(_abc_17692_n8584), .B(_abc_17692_n8516), .Y(_abc_17692_n8587) );
  OR2X2 OR2X2_2784 ( .A(_abc_17692_n8472), .B(_abc_17692_n8406), .Y(_abc_17692_n8590) );
  OR2X2 OR2X2_2785 ( .A(_abc_17692_n8551), .B(_abc_17692_n8590), .Y(_abc_17692_n8593) );
  OR2X2 OR2X2_2786 ( .A(_abc_17692_n8595), .B(_abc_17692_n8589), .Y(_abc_17692_n8596) );
  OR2X2 OR2X2_2787 ( .A(_abc_17692_n8478), .B(_abc_17692_n8597), .Y(_abc_17692_n8598) );
  OR2X2 OR2X2_2788 ( .A(_abc_17692_n8598), .B(_abc_17692_n8571), .Y(_abc_17692_n8601) );
  OR2X2 OR2X2_2789 ( .A(_abc_17692_n8483), .B(_abc_17692_n8437), .Y(_abc_17692_n8604) );
  OR2X2 OR2X2_279 ( .A(_abc_17692_n1280), .B(_abc_17692_n1248), .Y(_abc_17692_n1281) );
  OR2X2 OR2X2_2790 ( .A(_abc_17692_n8604), .B(_abc_17692_n8532), .Y(_abc_17692_n8607) );
  OR2X2 OR2X2_2791 ( .A(_abc_17692_n8603), .B(_abc_17692_n8609), .Y(_abc_17692_n8610) );
  OR2X2 OR2X2_2792 ( .A(_abc_17692_n8596), .B(_abc_17692_n8610), .Y(_abc_17692_n8611) );
  OR2X2 OR2X2_2793 ( .A(_abc_17692_n8613), .B(_abc_17692_n8614), .Y(_abc_17692_n8615) );
  OR2X2 OR2X2_2794 ( .A(_abc_17692_n8612), .B(_abc_17692_n8615), .Y(_abc_17692_n8616) );
  OR2X2 OR2X2_2795 ( .A(_abc_17692_n8581), .B(_abc_17692_n8616), .Y(workunit1_2__FF_INPUT) );
  OR2X2 OR2X2_2796 ( .A(_abc_17692_n8619), .B(_abc_17692_n8618), .Y(_abc_17692_n8620) );
  OR2X2 OR2X2_2797 ( .A(_abc_17692_n8506), .B(_abc_17692_n8497), .Y(_abc_17692_n8625) );
  OR2X2 OR2X2_2798 ( .A(_abc_17692_n8623), .B(_abc_17692_n8626), .Y(_abc_17692_n8627) );
  OR2X2 OR2X2_2799 ( .A(_abc_17692_n2302), .B(_abc_17692_n8627), .Y(_abc_17692_n8628) );
  OR2X2 OR2X2_28 ( .A(_abc_17692_n675), .B(x_3_), .Y(_abc_17692_n681) );
  OR2X2 OR2X2_280 ( .A(_abc_17692_n1283), .B(_abc_17692_n1278), .Y(_abc_17692_n1284) );
  OR2X2 OR2X2_2800 ( .A(_abc_17692_n8625), .B(_abc_17692_n8624), .Y(_abc_17692_n8629) );
  OR2X2 OR2X2_2801 ( .A(_abc_17692_n8631), .B(_abc_17692_n2306), .Y(_abc_17692_n8632) );
  OR2X2 OR2X2_2802 ( .A(_abc_17692_n8633), .B(_abc_17692_n2249), .Y(_abc_17692_n8634) );
  OR2X2 OR2X2_2803 ( .A(_abc_17692_n8631), .B(_abc_17692_n2302), .Y(_abc_17692_n8635) );
  OR2X2 OR2X2_2804 ( .A(_abc_17692_n2306), .B(_abc_17692_n8627), .Y(_abc_17692_n8636) );
  OR2X2 OR2X2_2805 ( .A(_abc_17692_n8637), .B(workunit1_3_), .Y(_abc_17692_n8638) );
  OR2X2 OR2X2_2806 ( .A(_abc_17692_n8519), .B(_abc_17692_n8640), .Y(_abc_17692_n8641) );
  OR2X2 OR2X2_2807 ( .A(_abc_17692_n8639), .B(_abc_17692_n8641), .Y(_abc_17692_n8644) );
  OR2X2 OR2X2_2808 ( .A(_abc_17692_n8631), .B(_abc_17692_n2268), .Y(_abc_17692_n8647) );
  OR2X2 OR2X2_2809 ( .A(_abc_17692_n2275), .B(_abc_17692_n8627), .Y(_abc_17692_n8648) );
  OR2X2 OR2X2_281 ( .A(_abc_17692_n1265), .B(_abc_17692_n1291), .Y(_abc_17692_n1292) );
  OR2X2 OR2X2_2810 ( .A(_abc_17692_n8649), .B(_abc_17692_n2249), .Y(_abc_17692_n8650) );
  OR2X2 OR2X2_2811 ( .A(_abc_17692_n2268), .B(_abc_17692_n8627), .Y(_abc_17692_n8651) );
  OR2X2 OR2X2_2812 ( .A(_abc_17692_n8631), .B(_abc_17692_n2275), .Y(_abc_17692_n8652) );
  OR2X2 OR2X2_2813 ( .A(_abc_17692_n8653), .B(workunit1_3_), .Y(_abc_17692_n8654) );
  OR2X2 OR2X2_2814 ( .A(_abc_17692_n8660), .B(_abc_17692_n8656), .Y(_abc_17692_n8661) );
  OR2X2 OR2X2_2815 ( .A(_abc_17692_n8659), .B(_abc_17692_n8655), .Y(_abc_17692_n8662) );
  OR2X2 OR2X2_2816 ( .A(_abc_17692_n2335), .B(_abc_17692_n8631), .Y(_abc_17692_n8665) );
  OR2X2 OR2X2_2817 ( .A(_abc_17692_n2331), .B(_abc_17692_n8627), .Y(_abc_17692_n8666) );
  OR2X2 OR2X2_2818 ( .A(_abc_17692_n8668), .B(_abc_17692_n2249), .Y(_abc_17692_n8669) );
  OR2X2 OR2X2_2819 ( .A(_abc_17692_n8667), .B(workunit1_3_), .Y(_abc_17692_n8670) );
  OR2X2 OR2X2_282 ( .A(_abc_17692_n1295), .B(_abc_17692_n1290), .Y(_abc_17692_n1298) );
  OR2X2 OR2X2_2820 ( .A(_abc_17692_n8547), .B(_abc_17692_n2062_1), .Y(_abc_17692_n8672) );
  OR2X2 OR2X2_2821 ( .A(_abc_17692_n8556), .B(_abc_17692_n8673), .Y(_abc_17692_n8674) );
  OR2X2 OR2X2_2822 ( .A(_abc_17692_n8674), .B(_abc_17692_n8671), .Y(_abc_17692_n8677) );
  OR2X2 OR2X2_2823 ( .A(_abc_17692_n8679), .B(_abc_17692_n8664), .Y(_abc_17692_n8680) );
  OR2X2 OR2X2_2824 ( .A(_abc_17692_n8680), .B(_abc_17692_n8646), .Y(_abc_17692_n8681) );
  OR2X2 OR2X2_2825 ( .A(_abc_17692_n2366), .B(_abc_17692_n8631), .Y(_abc_17692_n8682) );
  OR2X2 OR2X2_2826 ( .A(_abc_17692_n2370), .B(_abc_17692_n8627), .Y(_abc_17692_n8683) );
  OR2X2 OR2X2_2827 ( .A(_abc_17692_n8684), .B(_abc_17692_n2249), .Y(_abc_17692_n8685) );
  OR2X2 OR2X2_2828 ( .A(_abc_17692_n2366), .B(_abc_17692_n8627), .Y(_abc_17692_n8686) );
  OR2X2 OR2X2_2829 ( .A(_abc_17692_n2370), .B(_abc_17692_n8631), .Y(_abc_17692_n8687) );
  OR2X2 OR2X2_283 ( .A(_abc_17692_n1300), .B(_abc_17692_n1289), .Y(_abc_17692_n1301) );
  OR2X2 OR2X2_2830 ( .A(_abc_17692_n8688), .B(workunit1_3_), .Y(_abc_17692_n8689) );
  OR2X2 OR2X2_2831 ( .A(_abc_17692_n8569), .B(_abc_17692_n2062_1), .Y(_abc_17692_n8692) );
  OR2X2 OR2X2_2832 ( .A(_abc_17692_n8694), .B(_abc_17692_n8691), .Y(_abc_17692_n8695) );
  OR2X2 OR2X2_2833 ( .A(_abc_17692_n8681), .B(_abc_17692_n8699), .Y(_abc_17692_n8700) );
  OR2X2 OR2X2_2834 ( .A(_abc_17692_n8510), .B(_abc_17692_n2062_1), .Y(_abc_17692_n8703) );
  OR2X2 OR2X2_2835 ( .A(_abc_17692_n8705), .B(_abc_17692_n8702), .Y(_abc_17692_n8706) );
  OR2X2 OR2X2_2836 ( .A(_abc_17692_n8704), .B(_abc_17692_n8639), .Y(_abc_17692_n8707) );
  OR2X2 OR2X2_2837 ( .A(_abc_17692_n8667), .B(_abc_17692_n2249), .Y(_abc_17692_n8710) );
  OR2X2 OR2X2_2838 ( .A(_abc_17692_n8668), .B(workunit1_3_), .Y(_abc_17692_n8711) );
  OR2X2 OR2X2_2839 ( .A(_abc_17692_n8591), .B(_abc_17692_n8548), .Y(_abc_17692_n8713) );
  OR2X2 OR2X2_284 ( .A(_abc_17692_n1288), .B(_abc_17692_n1301), .Y(sum_14__FF_INPUT) );
  OR2X2 OR2X2_2840 ( .A(_abc_17692_n8712), .B(_abc_17692_n8713), .Y(_abc_17692_n8716) );
  OR2X2 OR2X2_2841 ( .A(_abc_17692_n8718), .B(_abc_17692_n8709), .Y(_abc_17692_n8719) );
  OR2X2 OR2X2_2842 ( .A(_abc_17692_n8599), .B(_abc_17692_n8720), .Y(_abc_17692_n8721) );
  OR2X2 OR2X2_2843 ( .A(_abc_17692_n8721), .B(_abc_17692_n8690), .Y(_abc_17692_n8724) );
  OR2X2 OR2X2_2844 ( .A(_abc_17692_n8605), .B(_abc_17692_n8727), .Y(_abc_17692_n8728) );
  OR2X2 OR2X2_2845 ( .A(_abc_17692_n8728), .B(_abc_17692_n8655), .Y(_abc_17692_n8731) );
  OR2X2 OR2X2_2846 ( .A(_abc_17692_n8726), .B(_abc_17692_n8733), .Y(_abc_17692_n8734) );
  OR2X2 OR2X2_2847 ( .A(_abc_17692_n8719), .B(_abc_17692_n8734), .Y(_abc_17692_n8735) );
  OR2X2 OR2X2_2848 ( .A(_abc_17692_n8737), .B(_abc_17692_n8738), .Y(_abc_17692_n8739) );
  OR2X2 OR2X2_2849 ( .A(_abc_17692_n8736), .B(_abc_17692_n8739), .Y(_abc_17692_n8740) );
  OR2X2 OR2X2_285 ( .A(_abc_17692_n1303), .B(delta_15_), .Y(_abc_17692_n1306) );
  OR2X2 OR2X2_2850 ( .A(_abc_17692_n8701), .B(_abc_17692_n8740), .Y(workunit1_3__FF_INPUT) );
  OR2X2 OR2X2_2851 ( .A(_abc_17692_n1814), .B(workunit2_9_), .Y(_abc_17692_n8742) );
  OR2X2 OR2X2_2852 ( .A(_abc_17692_n3471), .B(workunit2_0_), .Y(_abc_17692_n8743) );
  OR2X2 OR2X2_2853 ( .A(_abc_17692_n8744), .B(_abc_17692_n2482), .Y(_abc_17692_n8745) );
  OR2X2 OR2X2_2854 ( .A(_abc_17692_n8746), .B(_abc_17692_n8747), .Y(_abc_17692_n8748) );
  OR2X2 OR2X2_2855 ( .A(_abc_17692_n8748), .B(workunit2_4_), .Y(_abc_17692_n8749) );
  OR2X2 OR2X2_2856 ( .A(_abc_17692_n8499), .B(_abc_17692_n8620), .Y(_abc_17692_n8751) );
  OR2X2 OR2X2_2857 ( .A(_abc_17692_n8754), .B(_abc_17692_n8618), .Y(_abc_17692_n8755) );
  OR2X2 OR2X2_2858 ( .A(_abc_17692_n8753), .B(_abc_17692_n8755), .Y(_abc_17692_n8756) );
  OR2X2 OR2X2_2859 ( .A(_abc_17692_n8758), .B(_abc_17692_n8759), .Y(_abc_17692_n8760) );
  OR2X2 OR2X2_286 ( .A(_abc_17692_n1310), .B(_abc_17692_n1307), .Y(_abc_17692_n1311_1) );
  OR2X2 OR2X2_2860 ( .A(_abc_17692_n8496), .B(_abc_17692_n8751), .Y(_abc_17692_n8761) );
  OR2X2 OR2X2_2861 ( .A(_abc_17692_n8764), .B(_abc_17692_n8757), .Y(_abc_17692_n8765) );
  OR2X2 OR2X2_2862 ( .A(_abc_17692_n8766), .B(_abc_17692_n8768), .Y(_abc_17692_n8769) );
  OR2X2 OR2X2_2863 ( .A(_abc_17692_n8772), .B(_abc_17692_n8770), .Y(_abc_17692_n8773) );
  OR2X2 OR2X2_2864 ( .A(_abc_17692_n8675), .B(_abc_17692_n8774), .Y(_abc_17692_n8775) );
  OR2X2 OR2X2_2865 ( .A(_abc_17692_n8775), .B(_abc_17692_n8773), .Y(_abc_17692_n8778) );
  OR2X2 OR2X2_2866 ( .A(_abc_17692_n8781), .B(_abc_17692_n8782), .Y(_abc_17692_n8783) );
  OR2X2 OR2X2_2867 ( .A(_abc_17692_n8784), .B(workunit1_4_), .Y(_abc_17692_n8785) );
  OR2X2 OR2X2_2868 ( .A(_abc_17692_n8783), .B(_abc_17692_n2433), .Y(_abc_17692_n8786) );
  OR2X2 OR2X2_2869 ( .A(_abc_17692_n8642), .B(_abc_17692_n8788), .Y(_abc_17692_n8789) );
  OR2X2 OR2X2_287 ( .A(_abc_17692_n1313), .B(_abc_17692_n1312), .Y(_abc_17692_n1314) );
  OR2X2 OR2X2_2870 ( .A(_abc_17692_n8789), .B(_abc_17692_n8787), .Y(_abc_17692_n8790) );
  OR2X2 OR2X2_2871 ( .A(_abc_17692_n8796), .B(_abc_17692_n8795), .Y(_abc_17692_n8797) );
  OR2X2 OR2X2_2872 ( .A(_abc_17692_n8800), .B(_abc_17692_n8798), .Y(_abc_17692_n8801) );
  OR2X2 OR2X2_2873 ( .A(_abc_17692_n8805), .B(_abc_17692_n8801), .Y(_abc_17692_n8808) );
  OR2X2 OR2X2_2874 ( .A(_abc_17692_n8810), .B(_abc_17692_n8794), .Y(_abc_17692_n8811) );
  OR2X2 OR2X2_2875 ( .A(_abc_17692_n8811), .B(_abc_17692_n8780), .Y(_abc_17692_n8812) );
  OR2X2 OR2X2_2876 ( .A(_abc_17692_n2572), .B(_abc_17692_n8767), .Y(_abc_17692_n8813) );
  OR2X2 OR2X2_2877 ( .A(_abc_17692_n2567), .B(_abc_17692_n8765), .Y(_abc_17692_n8814) );
  OR2X2 OR2X2_2878 ( .A(_abc_17692_n8815), .B(_abc_17692_n2433), .Y(_abc_17692_n8816) );
  OR2X2 OR2X2_2879 ( .A(_abc_17692_n2572), .B(_abc_17692_n8765), .Y(_abc_17692_n8817) );
  OR2X2 OR2X2_288 ( .A(_abc_17692_n1319), .B(_abc_17692_n1307), .Y(_abc_17692_n1320_1) );
  OR2X2 OR2X2_2880 ( .A(_abc_17692_n2567), .B(_abc_17692_n8767), .Y(_abc_17692_n8818) );
  OR2X2 OR2X2_2881 ( .A(_abc_17692_n8819), .B(workunit1_4_), .Y(_abc_17692_n8820) );
  OR2X2 OR2X2_2882 ( .A(_abc_17692_n8688), .B(_abc_17692_n2249), .Y(_abc_17692_n8823) );
  OR2X2 OR2X2_2883 ( .A(_abc_17692_n8696), .B(_abc_17692_n8824), .Y(_abc_17692_n8825) );
  OR2X2 OR2X2_2884 ( .A(_abc_17692_n8825), .B(_abc_17692_n8822), .Y(_abc_17692_n8828) );
  OR2X2 OR2X2_2885 ( .A(_abc_17692_n8812), .B(_abc_17692_n8830), .Y(_abc_17692_n8831) );
  OR2X2 OR2X2_2886 ( .A(_abc_17692_n8637), .B(_abc_17692_n2249), .Y(_abc_17692_n8834) );
  OR2X2 OR2X2_2887 ( .A(_abc_17692_n8836), .B(_abc_17692_n8833), .Y(_abc_17692_n8837) );
  OR2X2 OR2X2_2888 ( .A(_abc_17692_n8835), .B(_abc_17692_n8787), .Y(_abc_17692_n8838) );
  OR2X2 OR2X2_2889 ( .A(_abc_17692_n8714), .B(_abc_17692_n8842), .Y(_abc_17692_n8843) );
  OR2X2 OR2X2_289 ( .A(_abc_17692_n1318), .B(_abc_17692_n1312), .Y(_abc_17692_n1321) );
  OR2X2 OR2X2_2890 ( .A(_abc_17692_n8843), .B(_abc_17692_n8841), .Y(_abc_17692_n8846) );
  OR2X2 OR2X2_2891 ( .A(_abc_17692_n8848), .B(_abc_17692_n8840), .Y(_abc_17692_n8849) );
  OR2X2 OR2X2_2892 ( .A(_abc_17692_n8722), .B(_abc_17692_n8850), .Y(_abc_17692_n8851) );
  OR2X2 OR2X2_2893 ( .A(_abc_17692_n8851), .B(_abc_17692_n8821), .Y(_abc_17692_n8854) );
  OR2X2 OR2X2_2894 ( .A(_abc_17692_n8729), .B(_abc_17692_n8858), .Y(_abc_17692_n8859) );
  OR2X2 OR2X2_2895 ( .A(_abc_17692_n8859), .B(_abc_17692_n8857), .Y(_abc_17692_n8862) );
  OR2X2 OR2X2_2896 ( .A(_abc_17692_n8856), .B(_abc_17692_n8864), .Y(_abc_17692_n8865) );
  OR2X2 OR2X2_2897 ( .A(_abc_17692_n8849), .B(_abc_17692_n8865), .Y(_abc_17692_n8866) );
  OR2X2 OR2X2_2898 ( .A(_abc_17692_n8868), .B(_abc_17692_n8869), .Y(_abc_17692_n8870) );
  OR2X2 OR2X2_2899 ( .A(_abc_17692_n8867), .B(_abc_17692_n8870), .Y(_abc_17692_n8871) );
  OR2X2 OR2X2_29 ( .A(_abc_17692_n679), .B(x_4_), .Y(_abc_17692_n685) );
  OR2X2 OR2X2_290 ( .A(_abc_17692_n1323), .B(_abc_17692_n1317), .Y(_abc_17692_n1324) );
  OR2X2 OR2X2_2900 ( .A(_abc_17692_n8832), .B(_abc_17692_n8871), .Y(workunit1_4__FF_INPUT) );
  OR2X2 OR2X2_2901 ( .A(_abc_17692_n8763), .B(_abc_17692_n8760), .Y(_abc_17692_n8873) );
  OR2X2 OR2X2_2902 ( .A(_abc_17692_n8876), .B(_abc_17692_n8875), .Y(_abc_17692_n8877) );
  OR2X2 OR2X2_2903 ( .A(_abc_17692_n8877), .B(_abc_17692_n2633), .Y(_abc_17692_n8878) );
  OR2X2 OR2X2_2904 ( .A(workunit2_1_bF_buf1), .B(workunit2_10_bF_buf2), .Y(_abc_17692_n8880) );
  OR2X2 OR2X2_2905 ( .A(_abc_17692_n8881), .B(workunit2_5_), .Y(_abc_17692_n8882) );
  OR2X2 OR2X2_2906 ( .A(_abc_17692_n8757), .B(_abc_17692_n8758), .Y(_abc_17692_n8885) );
  OR2X2 OR2X2_2907 ( .A(_abc_17692_n8887), .B(_abc_17692_n8886), .Y(_abc_17692_n8888) );
  OR2X2 OR2X2_2908 ( .A(_abc_17692_n8884), .B(_abc_17692_n8889), .Y(_abc_17692_n8890) );
  OR2X2 OR2X2_2909 ( .A(_abc_17692_n8885), .B(_abc_17692_n8888), .Y(_abc_17692_n8892) );
  OR2X2 OR2X2_291 ( .A(_abc_17692_n1316), .B(_abc_17692_n1324), .Y(sum_15__FF_INPUT) );
  OR2X2 OR2X2_2910 ( .A(_abc_17692_n8891), .B(_abc_17692_n8895), .Y(_abc_17692_n8896) );
  OR2X2 OR2X2_2911 ( .A(_abc_17692_n8897), .B(_abc_17692_n1817), .Y(_abc_17692_n8898) );
  OR2X2 OR2X2_2912 ( .A(_abc_17692_n8896), .B(workunit1_5_), .Y(_abc_17692_n8899) );
  OR2X2 OR2X2_2913 ( .A(_abc_17692_n8791), .B(_abc_17692_n8901), .Y(_abc_17692_n8902) );
  OR2X2 OR2X2_2914 ( .A(_abc_17692_n8902), .B(_abc_17692_n8900), .Y(_abc_17692_n8905) );
  OR2X2 OR2X2_2915 ( .A(_abc_17692_n2691), .B(_abc_17692_n8894), .Y(_abc_17692_n8908) );
  OR2X2 OR2X2_2916 ( .A(_abc_17692_n2693), .B(_abc_17692_n8890), .Y(_abc_17692_n8909) );
  OR2X2 OR2X2_2917 ( .A(_abc_17692_n8911), .B(workunit1_5_), .Y(_abc_17692_n8914) );
  OR2X2 OR2X2_2918 ( .A(_abc_17692_n8776), .B(_abc_17692_n8916), .Y(_abc_17692_n8917) );
  OR2X2 OR2X2_2919 ( .A(_abc_17692_n8917), .B(_abc_17692_n8915), .Y(_abc_17692_n8920) );
  OR2X2 OR2X2_292 ( .A(_abc_17692_n1329), .B(_abc_17692_n1326), .Y(_abc_17692_n1330) );
  OR2X2 OR2X2_2920 ( .A(_abc_17692_n8924), .B(_abc_17692_n8923), .Y(_abc_17692_n8925) );
  OR2X2 OR2X2_2921 ( .A(_abc_17692_n8925), .B(_abc_17692_n1817), .Y(_abc_17692_n8926) );
  OR2X2 OR2X2_2922 ( .A(_abc_17692_n8894), .B(_abc_17692_n2724), .Y(_abc_17692_n8927) );
  OR2X2 OR2X2_2923 ( .A(_abc_17692_n8890), .B(_abc_17692_n2720), .Y(_abc_17692_n8928) );
  OR2X2 OR2X2_2924 ( .A(_abc_17692_n8929), .B(workunit1_5_), .Y(_abc_17692_n8930) );
  OR2X2 OR2X2_2925 ( .A(_abc_17692_n8806), .B(_abc_17692_n8933), .Y(_abc_17692_n8934) );
  OR2X2 OR2X2_2926 ( .A(_abc_17692_n8934), .B(_abc_17692_n8932), .Y(_abc_17692_n8935) );
  OR2X2 OR2X2_2927 ( .A(_abc_17692_n8939), .B(_abc_17692_n8922), .Y(_abc_17692_n8940) );
  OR2X2 OR2X2_2928 ( .A(_abc_17692_n8940), .B(_abc_17692_n8907), .Y(_abc_17692_n8941) );
  OR2X2 OR2X2_2929 ( .A(_abc_17692_n2752), .B(_abc_17692_n8894), .Y(_abc_17692_n8942) );
  OR2X2 OR2X2_293 ( .A(_abc_17692_n1333), .B(_abc_17692_n1281), .Y(_abc_17692_n1334) );
  OR2X2 OR2X2_2930 ( .A(_abc_17692_n2756), .B(_abc_17692_n8890), .Y(_abc_17692_n8943) );
  OR2X2 OR2X2_2931 ( .A(_abc_17692_n8944), .B(_abc_17692_n1817), .Y(_abc_17692_n8945) );
  OR2X2 OR2X2_2932 ( .A(_abc_17692_n2756), .B(_abc_17692_n8894), .Y(_abc_17692_n8946) );
  OR2X2 OR2X2_2933 ( .A(_abc_17692_n2752), .B(_abc_17692_n8890), .Y(_abc_17692_n8947) );
  OR2X2 OR2X2_2934 ( .A(_abc_17692_n8948), .B(workunit1_5_), .Y(_abc_17692_n8949) );
  OR2X2 OR2X2_2935 ( .A(_abc_17692_n8819), .B(_abc_17692_n2433), .Y(_abc_17692_n8952) );
  OR2X2 OR2X2_2936 ( .A(_abc_17692_n8826), .B(_abc_17692_n8953), .Y(_abc_17692_n8954) );
  OR2X2 OR2X2_2937 ( .A(_abc_17692_n8954), .B(_abc_17692_n8951), .Y(_abc_17692_n8957) );
  OR2X2 OR2X2_2938 ( .A(_abc_17692_n8941), .B(_abc_17692_n8959), .Y(_abc_17692_n8960) );
  OR2X2 OR2X2_2939 ( .A(_abc_17692_n8966), .B(_abc_17692_n8962), .Y(_abc_17692_n8967) );
  OR2X2 OR2X2_294 ( .A(_abc_17692_n1335), .B(_abc_17692_n1336), .Y(_abc_17692_n1337) );
  OR2X2 OR2X2_2940 ( .A(_abc_17692_n8965), .B(_abc_17692_n8900), .Y(_abc_17692_n8968) );
  OR2X2 OR2X2_2941 ( .A(_abc_17692_n8844), .B(_abc_17692_n8770), .Y(_abc_17692_n8972) );
  OR2X2 OR2X2_2942 ( .A(_abc_17692_n8972), .B(_abc_17692_n8971), .Y(_abc_17692_n8975) );
  OR2X2 OR2X2_2943 ( .A(_abc_17692_n8977), .B(_abc_17692_n8970), .Y(_abc_17692_n8978) );
  OR2X2 OR2X2_2944 ( .A(_abc_17692_n8852), .B(_abc_17692_n8979), .Y(_abc_17692_n8980) );
  OR2X2 OR2X2_2945 ( .A(_abc_17692_n8980), .B(_abc_17692_n8950), .Y(_abc_17692_n8983) );
  OR2X2 OR2X2_2946 ( .A(_abc_17692_n8860), .B(_abc_17692_n8798), .Y(_abc_17692_n8986) );
  OR2X2 OR2X2_2947 ( .A(_abc_17692_n8986), .B(_abc_17692_n8931), .Y(_abc_17692_n8989) );
  OR2X2 OR2X2_2948 ( .A(_abc_17692_n8985), .B(_abc_17692_n8991), .Y(_abc_17692_n8992) );
  OR2X2 OR2X2_2949 ( .A(_abc_17692_n8978), .B(_abc_17692_n8992), .Y(_abc_17692_n8993) );
  OR2X2 OR2X2_295 ( .A(_abc_17692_n1279), .B(_abc_17692_n1333), .Y(_abc_17692_n1340) );
  OR2X2 OR2X2_2950 ( .A(_abc_17692_n8995), .B(_abc_17692_n8996), .Y(_abc_17692_n8997) );
  OR2X2 OR2X2_2951 ( .A(_abc_17692_n8994), .B(_abc_17692_n8997), .Y(_abc_17692_n8998) );
  OR2X2 OR2X2_2952 ( .A(_abc_17692_n8961), .B(_abc_17692_n8998), .Y(workunit1_5__FF_INPUT) );
  OR2X2 OR2X2_2953 ( .A(_abc_17692_n8760), .B(_abc_17692_n8888), .Y(_abc_17692_n9000) );
  OR2X2 OR2X2_2954 ( .A(_abc_17692_n8763), .B(_abc_17692_n9000), .Y(_abc_17692_n9001) );
  OR2X2 OR2X2_2955 ( .A(_abc_17692_n8745), .B(_abc_17692_n8887), .Y(_abc_17692_n9002) );
  OR2X2 OR2X2_2956 ( .A(workunit2_2_), .B(workunit2_11_), .Y(_abc_17692_n9007) );
  OR2X2 OR2X2_2957 ( .A(_abc_17692_n9010), .B(_abc_17692_n9005), .Y(_abc_17692_n9011) );
  OR2X2 OR2X2_2958 ( .A(_abc_17692_n9012), .B(_abc_17692_n9009), .Y(_abc_17692_n9013) );
  OR2X2 OR2X2_2959 ( .A(_abc_17692_n8758), .B(_abc_17692_n8886), .Y(_abc_17692_n9017) );
  OR2X2 OR2X2_296 ( .A(_abc_17692_n1342), .B(_abc_17692_n1331_1), .Y(_abc_17692_n1343_1) );
  OR2X2 OR2X2_2960 ( .A(_abc_17692_n9016), .B(_abc_17692_n9018), .Y(_abc_17692_n9019) );
  OR2X2 OR2X2_2961 ( .A(_abc_17692_n9011), .B(_abc_17692_n2862), .Y(_abc_17692_n9020) );
  OR2X2 OR2X2_2962 ( .A(_abc_17692_n9008), .B(workunit2_6_), .Y(_abc_17692_n9021) );
  OR2X2 OR2X2_2963 ( .A(_abc_17692_n9014), .B(_abc_17692_n9023), .Y(_abc_17692_n9024) );
  OR2X2 OR2X2_2964 ( .A(_abc_17692_n9025), .B(_abc_17692_n9027), .Y(_abc_17692_n9028) );
  OR2X2 OR2X2_2965 ( .A(_abc_17692_n9031), .B(_abc_17692_n9029), .Y(_abc_17692_n9032) );
  OR2X2 OR2X2_2966 ( .A(_abc_17692_n8918), .B(_abc_17692_n8912), .Y(_abc_17692_n9033) );
  OR2X2 OR2X2_2967 ( .A(_abc_17692_n9033), .B(_abc_17692_n9032), .Y(_abc_17692_n9036) );
  OR2X2 OR2X2_2968 ( .A(_abc_17692_n9040), .B(_abc_17692_n9039), .Y(_abc_17692_n9041) );
  OR2X2 OR2X2_2969 ( .A(_abc_17692_n9044), .B(_abc_17692_n9042), .Y(_abc_17692_n9045) );
  OR2X2 OR2X2_297 ( .A(_abc_17692_n1312), .B(_abc_17692_n1276), .Y(_abc_17692_n1354) );
  OR2X2 OR2X2_2970 ( .A(_abc_17692_n8903), .B(_abc_17692_n9046), .Y(_abc_17692_n9047) );
  OR2X2 OR2X2_2971 ( .A(_abc_17692_n9047), .B(_abc_17692_n9045), .Y(_abc_17692_n9048) );
  OR2X2 OR2X2_2972 ( .A(_abc_17692_n9054), .B(_abc_17692_n9053), .Y(_abc_17692_n9055) );
  OR2X2 OR2X2_2973 ( .A(_abc_17692_n9057), .B(_abc_17692_n9058), .Y(_abc_17692_n9059) );
  OR2X2 OR2X2_2974 ( .A(_abc_17692_n8931), .B(_abc_17692_n8857), .Y(_abc_17692_n9061) );
  OR2X2 OR2X2_2975 ( .A(_abc_17692_n9061), .B(_abc_17692_n8804), .Y(_abc_17692_n9062) );
  OR2X2 OR2X2_2976 ( .A(_abc_17692_n8931), .B(_abc_17692_n9065), .Y(_abc_17692_n9066) );
  OR2X2 OR2X2_2977 ( .A(_abc_17692_n9069), .B(_abc_17692_n9060), .Y(_abc_17692_n9070) );
  OR2X2 OR2X2_2978 ( .A(_abc_17692_n9052), .B(_abc_17692_n9074), .Y(_abc_17692_n9075) );
  OR2X2 OR2X2_2979 ( .A(_abc_17692_n9075), .B(_abc_17692_n9038), .Y(_abc_17692_n9076) );
  OR2X2 OR2X2_298 ( .A(_abc_17692_n1353), .B(_abc_17692_n1356), .Y(_abc_17692_n1357) );
  OR2X2 OR2X2_2980 ( .A(_abc_17692_n9078), .B(_abc_17692_n9077), .Y(_abc_17692_n9079) );
  OR2X2 OR2X2_2981 ( .A(_abc_17692_n9079), .B(_abc_17692_n2821), .Y(_abc_17692_n9080) );
  OR2X2 OR2X2_2982 ( .A(_abc_17692_n9081), .B(workunit1_6_), .Y(_abc_17692_n9082) );
  OR2X2 OR2X2_2983 ( .A(_abc_17692_n8948), .B(_abc_17692_n1817), .Y(_abc_17692_n9084) );
  OR2X2 OR2X2_2984 ( .A(_abc_17692_n8955), .B(_abc_17692_n9085), .Y(_abc_17692_n9086) );
  OR2X2 OR2X2_2985 ( .A(_abc_17692_n9086), .B(_abc_17692_n9083), .Y(_abc_17692_n9087) );
  OR2X2 OR2X2_2986 ( .A(_abc_17692_n9076), .B(_abc_17692_n9091), .Y(_abc_17692_n9092) );
  OR2X2 OR2X2_2987 ( .A(_abc_17692_n8911), .B(_abc_17692_n1817), .Y(_abc_17692_n9095) );
  OR2X2 OR2X2_2988 ( .A(_abc_17692_n8973), .B(_abc_17692_n9096), .Y(_abc_17692_n9097) );
  OR2X2 OR2X2_2989 ( .A(_abc_17692_n9097), .B(_abc_17692_n9094), .Y(_abc_17692_n9100) );
  OR2X2 OR2X2_299 ( .A(_abc_17692_n1351), .B(_abc_17692_n1357), .Y(_abc_17692_n1358) );
  OR2X2 OR2X2_2990 ( .A(_abc_17692_n8987), .B(_abc_17692_n9103), .Y(_abc_17692_n9104) );
  OR2X2 OR2X2_2991 ( .A(_abc_17692_n9104), .B(_abc_17692_n9059), .Y(_abc_17692_n9105) );
  OR2X2 OR2X2_2992 ( .A(_abc_17692_n9109), .B(_abc_17692_n9102), .Y(_abc_17692_n9110) );
  OR2X2 OR2X2_2993 ( .A(_abc_17692_n8981), .B(_abc_17692_n9112), .Y(_abc_17692_n9113) );
  OR2X2 OR2X2_2994 ( .A(_abc_17692_n9113), .B(_abc_17692_n9111), .Y(_abc_17692_n9116) );
  OR2X2 OR2X2_2995 ( .A(_abc_17692_n9121), .B(_abc_17692_n9045), .Y(_abc_17692_n9122) );
  OR2X2 OR2X2_2996 ( .A(_abc_17692_n9124), .B(_abc_17692_n9123), .Y(_abc_17692_n9125) );
  OR2X2 OR2X2_2997 ( .A(_abc_17692_n9127), .B(_abc_17692_n9118), .Y(_abc_17692_n9128) );
  OR2X2 OR2X2_2998 ( .A(_abc_17692_n9110), .B(_abc_17692_n9128), .Y(_abc_17692_n9129) );
  OR2X2 OR2X2_2999 ( .A(_abc_17692_n9131), .B(_abc_17692_n9132), .Y(_abc_17692_n9133) );
  OR2X2 OR2X2_3 ( .A(state_8_bF_buf8), .B(modereg), .Y(_abc_17692_n631) );
  OR2X2 OR2X2_30 ( .A(_abc_17692_n683), .B(x_5_), .Y(_abc_17692_n687) );
  OR2X2 OR2X2_300 ( .A(_abc_17692_n1358), .B(_abc_17692_n1349), .Y(_abc_17692_n1359) );
  OR2X2 OR2X2_3000 ( .A(_abc_17692_n9130), .B(_abc_17692_n9133), .Y(_abc_17692_n9134) );
  OR2X2 OR2X2_3001 ( .A(_abc_17692_n9134), .B(_abc_17692_n9093), .Y(workunit1_6__FF_INPUT) );
  OR2X2 OR2X2_3002 ( .A(_abc_17692_n9004), .B(_abc_17692_n9013), .Y(_abc_17692_n9136) );
  OR2X2 OR2X2_3003 ( .A(workunit2_3_), .B(workunit2_12_bF_buf0), .Y(_abc_17692_n9140) );
  OR2X2 OR2X2_3004 ( .A(_abc_17692_n2246), .B(workunit2_12_bF_buf3), .Y(_abc_17692_n9143) );
  OR2X2 OR2X2_3005 ( .A(_abc_17692_n4120), .B(workunit2_3_), .Y(_abc_17692_n9144) );
  OR2X2 OR2X2_3006 ( .A(_abc_17692_n9146), .B(_abc_17692_n9142), .Y(_abc_17692_n9147) );
  OR2X2 OR2X2_3007 ( .A(_abc_17692_n9023), .B(_abc_17692_n9009), .Y(_abc_17692_n9149) );
  OR2X2 OR2X2_3008 ( .A(_abc_17692_n9145), .B(_abc_17692_n3060), .Y(_abc_17692_n9150) );
  OR2X2 OR2X2_3009 ( .A(_abc_17692_n9141), .B(workunit2_7_), .Y(_abc_17692_n9151) );
  OR2X2 OR2X2_301 ( .A(_abc_17692_n1359), .B(_abc_17692_n1330), .Y(_abc_17692_n1362) );
  OR2X2 OR2X2_3010 ( .A(_abc_17692_n9148), .B(_abc_17692_n9153), .Y(_abc_17692_n9154) );
  OR2X2 OR2X2_3011 ( .A(_abc_17692_n9154), .B(_abc_17692_n3108), .Y(_abc_17692_n9155) );
  OR2X2 OR2X2_3012 ( .A(_abc_17692_n9149), .B(_abc_17692_n9152), .Y(_abc_17692_n9156) );
  OR2X2 OR2X2_3013 ( .A(_abc_17692_n9137), .B(_abc_17692_n9147), .Y(_abc_17692_n9157) );
  OR2X2 OR2X2_3014 ( .A(_abc_17692_n9158), .B(_abc_17692_n3112), .Y(_abc_17692_n9159) );
  OR2X2 OR2X2_3015 ( .A(_abc_17692_n9160), .B(_abc_17692_n2063), .Y(_abc_17692_n9161) );
  OR2X2 OR2X2_3016 ( .A(_abc_17692_n9158), .B(_abc_17692_n3108), .Y(_abc_17692_n9162) );
  OR2X2 OR2X2_3017 ( .A(_abc_17692_n9154), .B(_abc_17692_n3112), .Y(_abc_17692_n9163) );
  OR2X2 OR2X2_3018 ( .A(_abc_17692_n9164), .B(workunit1_7_), .Y(_abc_17692_n9165) );
  OR2X2 OR2X2_3019 ( .A(_abc_17692_n9170), .B(_abc_17692_n9167), .Y(_abc_17692_n9171) );
  OR2X2 OR2X2_302 ( .A(_abc_17692_n1365), .B(state_8_bF_buf0), .Y(_abc_17692_n1366) );
  OR2X2 OR2X2_3020 ( .A(_abc_17692_n9169), .B(_abc_17692_n9166), .Y(_abc_17692_n9172) );
  OR2X2 OR2X2_3021 ( .A(_abc_17692_n9176), .B(_abc_17692_n9175), .Y(_abc_17692_n9177) );
  OR2X2 OR2X2_3022 ( .A(_abc_17692_n9179), .B(_abc_17692_n9180), .Y(_abc_17692_n9181) );
  OR2X2 OR2X2_3023 ( .A(_abc_17692_n9049), .B(_abc_17692_n9182), .Y(_abc_17692_n9183) );
  OR2X2 OR2X2_3024 ( .A(_abc_17692_n9183), .B(_abc_17692_n9181), .Y(_abc_17692_n9186) );
  OR2X2 OR2X2_3025 ( .A(_abc_17692_n9190), .B(_abc_17692_n9191), .Y(_abc_17692_n9192) );
  OR2X2 OR2X2_3026 ( .A(_abc_17692_n9194), .B(_abc_17692_n9195), .Y(_abc_17692_n9196) );
  OR2X2 OR2X2_3027 ( .A(_abc_17692_n9196), .B(_abc_17692_n9189), .Y(_abc_17692_n9197) );
  OR2X2 OR2X2_3028 ( .A(_abc_17692_n9034), .B(_abc_17692_n9197), .Y(_abc_17692_n9198) );
  OR2X2 OR2X2_3029 ( .A(_abc_17692_n9205), .B(_abc_17692_n9188), .Y(_abc_17692_n9206) );
  OR2X2 OR2X2_303 ( .A(_abc_17692_n1364), .B(_abc_17692_n1366), .Y(_abc_17692_n1367) );
  OR2X2 OR2X2_3030 ( .A(_abc_17692_n9206), .B(_abc_17692_n9174), .Y(_abc_17692_n9207) );
  OR2X2 OR2X2_3031 ( .A(_abc_17692_n9209), .B(_abc_17692_n9208), .Y(_abc_17692_n9210) );
  OR2X2 OR2X2_3032 ( .A(_abc_17692_n9212), .B(_abc_17692_n9213), .Y(_abc_17692_n9214) );
  OR2X2 OR2X2_3033 ( .A(_abc_17692_n9088), .B(_abc_17692_n9216), .Y(_abc_17692_n9217) );
  OR2X2 OR2X2_3034 ( .A(_abc_17692_n9217), .B(_abc_17692_n9215), .Y(_abc_17692_n9218) );
  OR2X2 OR2X2_3035 ( .A(_abc_17692_n9207), .B(_abc_17692_n9222), .Y(_abc_17692_n9223) );
  OR2X2 OR2X2_3036 ( .A(_abc_17692_n9226), .B(_abc_17692_n9196), .Y(_abc_17692_n9227) );
  OR2X2 OR2X2_3037 ( .A(_abc_17692_n9231), .B(_abc_17692_n9230), .Y(_abc_17692_n9232) );
  OR2X2 OR2X2_3038 ( .A(_abc_17692_n9238), .B(_abc_17692_n9166), .Y(_abc_17692_n9239) );
  OR2X2 OR2X2_3039 ( .A(_abc_17692_n9237), .B(_abc_17692_n9167), .Y(_abc_17692_n9240) );
  OR2X2 OR2X2_304 ( .A(_abc_17692_n1347), .B(_abc_17692_n1367), .Y(sum_16__FF_INPUT) );
  OR2X2 OR2X2_3040 ( .A(_abc_17692_n9234), .B(_abc_17692_n9242), .Y(_abc_17692_n9243) );
  OR2X2 OR2X2_3041 ( .A(_abc_17692_n9081), .B(_abc_17692_n2821), .Y(_abc_17692_n9244) );
  OR2X2 OR2X2_3042 ( .A(_abc_17692_n9114), .B(_abc_17692_n9245), .Y(_abc_17692_n9246) );
  OR2X2 OR2X2_3043 ( .A(_abc_17692_n9246), .B(_abc_17692_n9214), .Y(_abc_17692_n9247) );
  OR2X2 OR2X2_3044 ( .A(_abc_17692_n9253), .B(_abc_17692_n9042), .Y(_abc_17692_n9254) );
  OR2X2 OR2X2_3045 ( .A(_abc_17692_n9252), .B(_abc_17692_n9254), .Y(_abc_17692_n9255) );
  OR2X2 OR2X2_3046 ( .A(_abc_17692_n9122), .B(_abc_17692_n9181), .Y(_abc_17692_n9256) );
  OR2X2 OR2X2_3047 ( .A(_abc_17692_n9181), .B(_abc_17692_n9257), .Y(_abc_17692_n9258) );
  OR2X2 OR2X2_3048 ( .A(_abc_17692_n9251), .B(_abc_17692_n9261), .Y(_abc_17692_n9262) );
  OR2X2 OR2X2_3049 ( .A(_abc_17692_n9243), .B(_abc_17692_n9262), .Y(_abc_17692_n9263) );
  OR2X2 OR2X2_305 ( .A(_abc_17692_n1378), .B(_abc_17692_n1375), .Y(_abc_17692_n1379) );
  OR2X2 OR2X2_3050 ( .A(_abc_17692_n9265), .B(_abc_17692_n9266), .Y(_abc_17692_n9267) );
  OR2X2 OR2X2_3051 ( .A(_abc_17692_n9264), .B(_abc_17692_n9267), .Y(_abc_17692_n9268) );
  OR2X2 OR2X2_3052 ( .A(_abc_17692_n9268), .B(_abc_17692_n9224), .Y(workunit1_7__FF_INPUT) );
  OR2X2 OR2X2_3053 ( .A(_abc_17692_n9274), .B(_abc_17692_n9146), .Y(_abc_17692_n9275) );
  OR2X2 OR2X2_3054 ( .A(_abc_17692_n9273), .B(_abc_17692_n9276), .Y(_abc_17692_n9277) );
  OR2X2 OR2X2_3055 ( .A(_abc_17692_n9277), .B(_abc_17692_n9272), .Y(_abc_17692_n9278) );
  OR2X2 OR2X2_3056 ( .A(_abc_17692_n9279), .B(_abc_17692_n9280), .Y(_abc_17692_n9281) );
  OR2X2 OR2X2_3057 ( .A(_abc_17692_n2482), .B(workunit2_13_), .Y(_abc_17692_n9283) );
  OR2X2 OR2X2_3058 ( .A(_abc_17692_n4351), .B(workunit2_4_), .Y(_abc_17692_n9284) );
  OR2X2 OR2X2_3059 ( .A(_abc_17692_n9282), .B(_abc_17692_n9286), .Y(_abc_17692_n9287) );
  OR2X2 OR2X2_306 ( .A(_abc_17692_n1377), .B(_abc_17692_n1380), .Y(_abc_17692_n1381) );
  OR2X2 OR2X2_3060 ( .A(_abc_17692_n9013), .B(_abc_17692_n9147), .Y(_abc_17692_n9290) );
  OR2X2 OR2X2_3061 ( .A(_abc_17692_n9000), .B(_abc_17692_n9290), .Y(_abc_17692_n9291) );
  OR2X2 OR2X2_3062 ( .A(_abc_17692_n9291), .B(_abc_17692_n8763), .Y(_abc_17692_n9292) );
  OR2X2 OR2X2_3063 ( .A(_abc_17692_n9290), .B(_abc_17692_n9003), .Y(_abc_17692_n9293) );
  OR2X2 OR2X2_3064 ( .A(_abc_17692_n9296), .B(_abc_17692_n9289), .Y(_abc_17692_n9297) );
  OR2X2 OR2X2_3065 ( .A(_abc_17692_n3366_1), .B(_abc_17692_n9298), .Y(_abc_17692_n9299) );
  OR2X2 OR2X2_3066 ( .A(_abc_17692_n3368), .B(_abc_17692_n9297), .Y(_abc_17692_n9300) );
  OR2X2 OR2X2_3067 ( .A(_abc_17692_n9301), .B(workunit1_8_bF_buf1), .Y(_abc_17692_n9304) );
  OR2X2 OR2X2_3068 ( .A(_abc_17692_n9219), .B(_abc_17692_n9213), .Y(_abc_17692_n9307) );
  OR2X2 OR2X2_3069 ( .A(_abc_17692_n9308), .B(_abc_17692_n9306), .Y(_abc_17692_n9309) );
  OR2X2 OR2X2_307 ( .A(_abc_17692_n1380), .B(_abc_17692_n1384), .Y(_abc_17692_n1385) );
  OR2X2 OR2X2_3070 ( .A(_abc_17692_n9307), .B(_abc_17692_n9305), .Y(_abc_17692_n9310) );
  OR2X2 OR2X2_3071 ( .A(_abc_17692_n9311), .B(_abc_17692_n4047_bF_buf0), .Y(_abc_17692_n9312) );
  OR2X2 OR2X2_3072 ( .A(_abc_17692_n9298), .B(_abc_17692_n3245), .Y(_abc_17692_n9313) );
  OR2X2 OR2X2_3073 ( .A(_abc_17692_n3246), .B(_abc_17692_n9297), .Y(_abc_17692_n9314) );
  OR2X2 OR2X2_3074 ( .A(_abc_17692_n9317), .B(_abc_17692_n9318), .Y(_abc_17692_n9319) );
  OR2X2 OR2X2_3075 ( .A(_abc_17692_n9184), .B(_abc_17692_n9321), .Y(_abc_17692_n9322) );
  OR2X2 OR2X2_3076 ( .A(_abc_17692_n9322), .B(_abc_17692_n9320), .Y(_abc_17692_n9323) );
  OR2X2 OR2X2_3077 ( .A(_abc_17692_n9298), .B(_abc_17692_n3323), .Y(_abc_17692_n9328) );
  OR2X2 OR2X2_3078 ( .A(_abc_17692_n3324), .B(_abc_17692_n9297), .Y(_abc_17692_n9329) );
  OR2X2 OR2X2_3079 ( .A(_abc_17692_n9330), .B(workunit1_8_bF_buf2), .Y(_abc_17692_n9333) );
  OR2X2 OR2X2_308 ( .A(_abc_17692_n1360), .B(_abc_17692_n1385), .Y(_abc_17692_n1386) );
  OR2X2 OR2X2_3080 ( .A(_abc_17692_n9201), .B(_abc_17692_n9335), .Y(_abc_17692_n9336) );
  OR2X2 OR2X2_3081 ( .A(_abc_17692_n9199), .B(_abc_17692_n9336), .Y(_abc_17692_n9337) );
  OR2X2 OR2X2_3082 ( .A(_abc_17692_n9337), .B(_abc_17692_n9334), .Y(_abc_17692_n9338) );
  OR2X2 OR2X2_3083 ( .A(_abc_17692_n9298), .B(_abc_17692_n3290), .Y(_abc_17692_n9343) );
  OR2X2 OR2X2_3084 ( .A(_abc_17692_n3291), .B(_abc_17692_n9297), .Y(_abc_17692_n9344) );
  OR2X2 OR2X2_3085 ( .A(_abc_17692_n9345), .B(workunit1_8_bF_buf0), .Y(_abc_17692_n9348) );
  OR2X2 OR2X2_3086 ( .A(_abc_17692_n9166), .B(_abc_17692_n9168), .Y(_abc_17692_n9350) );
  OR2X2 OR2X2_3087 ( .A(_abc_17692_n9166), .B(_abc_17692_n9059), .Y(_abc_17692_n9354) );
  OR2X2 OR2X2_3088 ( .A(_abc_17692_n9068), .B(_abc_17692_n9354), .Y(_abc_17692_n9355) );
  OR2X2 OR2X2_3089 ( .A(_abc_17692_n9357), .B(_abc_17692_n9349), .Y(_abc_17692_n9358) );
  OR2X2 OR2X2_309 ( .A(_abc_17692_n1394), .B(state_8_bF_buf9), .Y(_abc_17692_n1395) );
  OR2X2 OR2X2_3090 ( .A(_abc_17692_n9362), .B(_abc_17692_n1863_bF_buf8), .Y(_abc_17692_n9363) );
  OR2X2 OR2X2_3091 ( .A(_abc_17692_n9342), .B(_abc_17692_n9363), .Y(_abc_17692_n9364) );
  OR2X2 OR2X2_3092 ( .A(_abc_17692_n9364), .B(_abc_17692_n9327), .Y(_abc_17692_n9365) );
  OR2X2 OR2X2_3093 ( .A(_abc_17692_n9248), .B(_abc_17692_n9368), .Y(_abc_17692_n9369) );
  OR2X2 OR2X2_3094 ( .A(_abc_17692_n9369), .B(_abc_17692_n9306), .Y(_abc_17692_n9370) );
  OR2X2 OR2X2_3095 ( .A(_abc_17692_n9378), .B(_abc_17692_n9319), .Y(_abc_17692_n9381) );
  OR2X2 OR2X2_3096 ( .A(_abc_17692_n9386), .B(_abc_17692_n9385), .Y(_abc_17692_n9387) );
  OR2X2 OR2X2_3097 ( .A(_abc_17692_n9389), .B(_abc_17692_n9387), .Y(_abc_17692_n9390) );
  OR2X2 OR2X2_3098 ( .A(_abc_17692_n9390), .B(_abc_17692_n9384), .Y(_abc_17692_n9391) );
  OR2X2 OR2X2_3099 ( .A(_abc_17692_n9397), .B(_abc_17692_n9194), .Y(_abc_17692_n9398) );
  OR2X2 OR2X2_31 ( .A(_abc_17692_n688), .B(x_6_), .Y(_abc_17692_n691) );
  OR2X2 OR2X2_310 ( .A(_abc_17692_n1393), .B(_abc_17692_n1395), .Y(_abc_17692_n1396) );
  OR2X2 OR2X2_3100 ( .A(_abc_17692_n9196), .B(_abc_17692_n9032), .Y(_abc_17692_n9399) );
  OR2X2 OR2X2_3101 ( .A(_abc_17692_n9401), .B(_abc_17692_n9398), .Y(_abc_17692_n9402) );
  OR2X2 OR2X2_3102 ( .A(_abc_17692_n9402), .B(_abc_17692_n9396), .Y(_abc_17692_n9405) );
  OR2X2 OR2X2_3103 ( .A(_abc_17692_n9407), .B(_abc_17692_n9395), .Y(_abc_17692_n9408) );
  OR2X2 OR2X2_3104 ( .A(_abc_17692_n9408), .B(_abc_17692_n9383), .Y(_abc_17692_n9409) );
  OR2X2 OR2X2_3105 ( .A(_abc_17692_n9409), .B(_abc_17692_n9374), .Y(_abc_17692_n9410) );
  OR2X2 OR2X2_3106 ( .A(_abc_17692_n9412), .B(_abc_17692_n9413), .Y(_abc_17692_n9414) );
  OR2X2 OR2X2_3107 ( .A(_abc_17692_n9411), .B(_abc_17692_n9414), .Y(_abc_17692_n9415) );
  OR2X2 OR2X2_3108 ( .A(_abc_17692_n9367), .B(_abc_17692_n9415), .Y(workunit1_8__FF_INPUT) );
  OR2X2 OR2X2_3109 ( .A(_abc_17692_n9289), .B(_abc_17692_n9282), .Y(_abc_17692_n9419) );
  OR2X2 OR2X2_311 ( .A(_abc_17692_n1383), .B(_abc_17692_n1396), .Y(sum_17__FF_INPUT) );
  OR2X2 OR2X2_3110 ( .A(workunit2_5_), .B(workunit2_14_bF_buf0), .Y(_abc_17692_n9423) );
  OR2X2 OR2X2_3111 ( .A(_abc_17692_n9426), .B(_abc_17692_n9421), .Y(_abc_17692_n9427) );
  OR2X2 OR2X2_3112 ( .A(_abc_17692_n9428), .B(_abc_17692_n9425), .Y(_abc_17692_n9429) );
  OR2X2 OR2X2_3113 ( .A(_abc_17692_n9431), .B(_abc_17692_n9432), .Y(_abc_17692_n9433) );
  OR2X2 OR2X2_3114 ( .A(_abc_17692_n9434), .B(_abc_17692_n3466), .Y(_abc_17692_n9435) );
  OR2X2 OR2X2_3115 ( .A(_abc_17692_n9433), .B(_abc_17692_n3463), .Y(_abc_17692_n9436) );
  OR2X2 OR2X2_3116 ( .A(_abc_17692_n9440), .B(_abc_17692_n9438), .Y(_abc_17692_n9441) );
  OR2X2 OR2X2_3117 ( .A(_abc_17692_n9445), .B(_abc_17692_n9442), .Y(_abc_17692_n9446) );
  OR2X2 OR2X2_3118 ( .A(_abc_17692_n9434), .B(_abc_17692_n3491), .Y(_abc_17692_n9450) );
  OR2X2 OR2X2_3119 ( .A(_abc_17692_n3494), .B(_abc_17692_n9433), .Y(_abc_17692_n9451) );
  OR2X2 OR2X2_312 ( .A(_abc_17692_n1401), .B(_abc_17692_n1398), .Y(_abc_17692_n1402) );
  OR2X2 OR2X2_3120 ( .A(_abc_17692_n9452), .B(_abc_17692_n2435), .Y(_abc_17692_n9453) );
  OR2X2 OR2X2_3121 ( .A(_abc_17692_n9434), .B(_abc_17692_n3494), .Y(_abc_17692_n9454) );
  OR2X2 OR2X2_3122 ( .A(_abc_17692_n3491), .B(_abc_17692_n9433), .Y(_abc_17692_n9455) );
  OR2X2 OR2X2_3123 ( .A(_abc_17692_n9456), .B(workunit1_9_), .Y(_abc_17692_n9457) );
  OR2X2 OR2X2_3124 ( .A(_abc_17692_n9449), .B(_abc_17692_n9459), .Y(_abc_17692_n9460) );
  OR2X2 OR2X2_3125 ( .A(_abc_17692_n9448), .B(_abc_17692_n9458), .Y(_abc_17692_n9461) );
  OR2X2 OR2X2_3126 ( .A(_abc_17692_n9434), .B(_abc_17692_n3519), .Y(_abc_17692_n9466) );
  OR2X2 OR2X2_3127 ( .A(_abc_17692_n3521), .B(_abc_17692_n9433), .Y(_abc_17692_n9467) );
  OR2X2 OR2X2_3128 ( .A(_abc_17692_n9468), .B(workunit1_9_), .Y(_abc_17692_n9471) );
  OR2X2 OR2X2_3129 ( .A(_abc_17692_n9465), .B(_abc_17692_n9473), .Y(_abc_17692_n9474) );
  OR2X2 OR2X2_313 ( .A(_abc_17692_n1341), .B(_abc_17692_n1405), .Y(_abc_17692_n1406) );
  OR2X2 OR2X2_3130 ( .A(_abc_17692_n9464), .B(_abc_17692_n9472), .Y(_abc_17692_n9475) );
  OR2X2 OR2X2_3131 ( .A(_abc_17692_n9477), .B(_abc_17692_n9463), .Y(_abc_17692_n9478) );
  OR2X2 OR2X2_3132 ( .A(_abc_17692_n9478), .B(_abc_17692_n9447), .Y(_abc_17692_n9479) );
  OR2X2 OR2X2_3133 ( .A(_abc_17692_n3545), .B(_abc_17692_n9434), .Y(_abc_17692_n9481) );
  OR2X2 OR2X2_3134 ( .A(_abc_17692_n3547), .B(_abc_17692_n9433), .Y(_abc_17692_n9482) );
  OR2X2 OR2X2_3135 ( .A(_abc_17692_n9493), .B(_abc_17692_n9491), .Y(_abc_17692_n9494) );
  OR2X2 OR2X2_3136 ( .A(_abc_17692_n9495), .B(_abc_17692_n9479), .Y(_abc_17692_n9496) );
  OR2X2 OR2X2_3137 ( .A(_abc_17692_n9503), .B(_abc_17692_n9504), .Y(_abc_17692_n9505) );
  OR2X2 OR2X2_3138 ( .A(_abc_17692_n9510), .B(_abc_17692_n9444), .Y(_abc_17692_n9511) );
  OR2X2 OR2X2_3139 ( .A(_abc_17692_n9509), .B(_abc_17692_n9441), .Y(_abc_17692_n9512) );
  OR2X2 OR2X2_314 ( .A(_abc_17692_n1407), .B(_abc_17692_n1373), .Y(_abc_17692_n1408) );
  OR2X2 OR2X2_3140 ( .A(_abc_17692_n9518), .B(_abc_17692_n9473), .Y(_abc_17692_n9519) );
  OR2X2 OR2X2_3141 ( .A(_abc_17692_n9520), .B(_abc_17692_n9472), .Y(_abc_17692_n9521) );
  OR2X2 OR2X2_3142 ( .A(_abc_17692_n9528), .B(_abc_17692_n9458), .Y(_abc_17692_n9529) );
  OR2X2 OR2X2_3143 ( .A(_abc_17692_n9527), .B(_abc_17692_n9459), .Y(_abc_17692_n9530) );
  OR2X2 OR2X2_3144 ( .A(_abc_17692_n9523), .B(_abc_17692_n9532), .Y(_abc_17692_n9533) );
  OR2X2 OR2X2_3145 ( .A(_abc_17692_n9533), .B(_abc_17692_n9514), .Y(_abc_17692_n9534) );
  OR2X2 OR2X2_3146 ( .A(_abc_17692_n9534), .B(_abc_17692_n9506), .Y(_abc_17692_n9535) );
  OR2X2 OR2X2_3147 ( .A(_abc_17692_n9537), .B(_abc_17692_n9538), .Y(_abc_17692_n9539) );
  OR2X2 OR2X2_3148 ( .A(_abc_17692_n9536), .B(_abc_17692_n9539), .Y(_abc_17692_n9540) );
  OR2X2 OR2X2_3149 ( .A(_abc_17692_n9540), .B(_abc_17692_n9497), .Y(workunit1_9__FF_INPUT) );
  OR2X2 OR2X2_315 ( .A(_abc_17692_n1410), .B(_abc_17692_n1403_1), .Y(_abc_17692_n1411) );
  OR2X2 OR2X2_3150 ( .A(_abc_17692_n9429), .B(_abc_17692_n9287), .Y(_abc_17692_n9542) );
  OR2X2 OR2X2_3151 ( .A(_abc_17692_n9295), .B(_abc_17692_n9542), .Y(_abc_17692_n9543) );
  OR2X2 OR2X2_3152 ( .A(_abc_17692_n9285), .B(_abc_17692_n3198), .Y(_abc_17692_n9545) );
  OR2X2 OR2X2_3153 ( .A(_abc_17692_n9428), .B(_abc_17692_n9545), .Y(_abc_17692_n9546) );
  OR2X2 OR2X2_3154 ( .A(_abc_17692_n9549), .B(_abc_17692_n9550), .Y(_abc_17692_n9551) );
  OR2X2 OR2X2_3155 ( .A(_abc_17692_n2862), .B(workunit2_15_), .Y(_abc_17692_n9553) );
  OR2X2 OR2X2_3156 ( .A(_abc_17692_n4765), .B(workunit2_6_), .Y(_abc_17692_n9554) );
  OR2X2 OR2X2_3157 ( .A(_abc_17692_n9552), .B(_abc_17692_n9556), .Y(_abc_17692_n9557) );
  OR2X2 OR2X2_3158 ( .A(_abc_17692_n9282), .B(_abc_17692_n9425), .Y(_abc_17692_n9562) );
  OR2X2 OR2X2_3159 ( .A(_abc_17692_n9560), .B(_abc_17692_n9563), .Y(_abc_17692_n9564) );
  OR2X2 OR2X2_316 ( .A(_abc_17692_n1420), .B(_abc_17692_n1402), .Y(_abc_17692_n1423) );
  OR2X2 OR2X2_3160 ( .A(_abc_17692_n9555), .B(_abc_17692_n3751), .Y(_abc_17692_n9565) );
  OR2X2 OR2X2_3161 ( .A(_abc_17692_n9551), .B(workunit2_10_bF_buf0), .Y(_abc_17692_n9566) );
  OR2X2 OR2X2_3162 ( .A(_abc_17692_n9558), .B(_abc_17692_n9568), .Y(_abc_17692_n9569) );
  OR2X2 OR2X2_3163 ( .A(_abc_17692_n9570), .B(_abc_17692_n9572), .Y(_abc_17692_n9573) );
  OR2X2 OR2X2_3164 ( .A(_abc_17692_n9574), .B(_abc_17692_n2638), .Y(_abc_17692_n9575) );
  OR2X2 OR2X2_3165 ( .A(_abc_17692_n9573), .B(workunit1_10_), .Y(_abc_17692_n9576) );
  OR2X2 OR2X2_3166 ( .A(_abc_17692_n9580), .B(_abc_17692_n9579), .Y(_abc_17692_n9581) );
  OR2X2 OR2X2_3167 ( .A(_abc_17692_n9587), .B(_abc_17692_n9578), .Y(_abc_17692_n9590) );
  OR2X2 OR2X2_3168 ( .A(_abc_17692_n9591), .B(_abc_17692_n4047_bF_buf4), .Y(_abc_17692_n9592) );
  OR2X2 OR2X2_3169 ( .A(_abc_17692_n9571), .B(_abc_17692_n3650_1), .Y(_abc_17692_n9593) );
  OR2X2 OR2X2_317 ( .A(_abc_17692_n1426), .B(state_8_bF_buf8), .Y(_abc_17692_n1427) );
  OR2X2 OR2X2_3170 ( .A(_abc_17692_n3651), .B(_abc_17692_n9569), .Y(_abc_17692_n9594) );
  OR2X2 OR2X2_3171 ( .A(_abc_17692_n9598), .B(_abc_17692_n9596), .Y(_abc_17692_n9599) );
  OR2X2 OR2X2_3172 ( .A(_abc_17692_n9604), .B(_abc_17692_n9603), .Y(_abc_17692_n9605) );
  OR2X2 OR2X2_3173 ( .A(_abc_17692_n9602), .B(_abc_17692_n9605), .Y(_abc_17692_n9606) );
  OR2X2 OR2X2_3174 ( .A(_abc_17692_n9606), .B(_abc_17692_n9600), .Y(_abc_17692_n9609) );
  OR2X2 OR2X2_3175 ( .A(_abc_17692_n9612), .B(_abc_17692_n9613), .Y(_abc_17692_n9614) );
  OR2X2 OR2X2_3176 ( .A(_abc_17692_n9615), .B(_abc_17692_n2638), .Y(_abc_17692_n9616) );
  OR2X2 OR2X2_3177 ( .A(_abc_17692_n9614), .B(workunit1_10_), .Y(_abc_17692_n9617) );
  OR2X2 OR2X2_3178 ( .A(_abc_17692_n9620), .B(_abc_17692_n9622), .Y(_abc_17692_n9623) );
  OR2X2 OR2X2_3179 ( .A(_abc_17692_n9626), .B(_abc_17692_n9625), .Y(_abc_17692_n9627) );
  OR2X2 OR2X2_318 ( .A(_abc_17692_n1425), .B(_abc_17692_n1427), .Y(_abc_17692_n1428) );
  OR2X2 OR2X2_3180 ( .A(_abc_17692_n9630), .B(_abc_17692_n9619), .Y(_abc_17692_n9633) );
  OR2X2 OR2X2_3181 ( .A(_abc_17692_n9637), .B(_abc_17692_n9636), .Y(_abc_17692_n9638) );
  OR2X2 OR2X2_3182 ( .A(_abc_17692_n9639), .B(_abc_17692_n2638), .Y(_abc_17692_n9640) );
  OR2X2 OR2X2_3183 ( .A(_abc_17692_n9638), .B(workunit1_10_), .Y(_abc_17692_n9641) );
  OR2X2 OR2X2_3184 ( .A(_abc_17692_n9458), .B(_abc_17692_n9384), .Y(_abc_17692_n9644) );
  OR2X2 OR2X2_3185 ( .A(_abc_17692_n9356), .B(_abc_17692_n9644), .Y(_abc_17692_n9645) );
  OR2X2 OR2X2_3186 ( .A(_abc_17692_n9458), .B(_abc_17692_n9347), .Y(_abc_17692_n9648) );
  OR2X2 OR2X2_3187 ( .A(_abc_17692_n9651), .B(_abc_17692_n9643), .Y(_abc_17692_n9654) );
  OR2X2 OR2X2_3188 ( .A(_abc_17692_n9656), .B(_abc_17692_n1863_bF_buf4), .Y(_abc_17692_n9657) );
  OR2X2 OR2X2_3189 ( .A(_abc_17692_n9635), .B(_abc_17692_n9657), .Y(_abc_17692_n9658) );
  OR2X2 OR2X2_319 ( .A(_abc_17692_n1415), .B(_abc_17692_n1428), .Y(sum_18__FF_INPUT) );
  OR2X2 OR2X2_3190 ( .A(_abc_17692_n9658), .B(_abc_17692_n9611), .Y(_abc_17692_n9659) );
  OR2X2 OR2X2_3191 ( .A(_abc_17692_n9484), .B(_abc_17692_n9499), .Y(_abc_17692_n9664) );
  OR2X2 OR2X2_3192 ( .A(_abc_17692_n9663), .B(_abc_17692_n9665), .Y(_abc_17692_n9666) );
  OR2X2 OR2X2_3193 ( .A(_abc_17692_n9666), .B(_abc_17692_n9577), .Y(_abc_17692_n9667) );
  OR2X2 OR2X2_3194 ( .A(_abc_17692_n9377), .B(_abc_17692_n9673), .Y(_abc_17692_n9674) );
  OR2X2 OR2X2_3195 ( .A(_abc_17692_n9440), .B(_abc_17692_n9508), .Y(_abc_17692_n9676) );
  OR2X2 OR2X2_3196 ( .A(_abc_17692_n9679), .B(_abc_17692_n9599), .Y(_abc_17692_n9682) );
  OR2X2 OR2X2_3197 ( .A(_abc_17692_n9687), .B(_abc_17692_n9525), .Y(_abc_17692_n9688) );
  OR2X2 OR2X2_3198 ( .A(_abc_17692_n9686), .B(_abc_17692_n9689), .Y(_abc_17692_n9690) );
  OR2X2 OR2X2_3199 ( .A(_abc_17692_n9690), .B(_abc_17692_n9642), .Y(_abc_17692_n9691) );
  OR2X2 OR2X2_32 ( .A(_abc_17692_n692_1), .B(x_7_), .Y(_abc_17692_n695) );
  OR2X2 OR2X2_320 ( .A(_abc_17692_n1412), .B(_abc_17692_n1398), .Y(_abc_17692_n1438) );
  OR2X2 OR2X2_3200 ( .A(_abc_17692_n9469), .B(_abc_17692_n9516), .Y(_abc_17692_n9698) );
  OR2X2 OR2X2_3201 ( .A(_abc_17692_n9697), .B(_abc_17692_n9699), .Y(_abc_17692_n9700) );
  OR2X2 OR2X2_3202 ( .A(_abc_17692_n9700), .B(_abc_17692_n9618), .Y(_abc_17692_n9703) );
  OR2X2 OR2X2_3203 ( .A(_abc_17692_n9705), .B(_abc_17692_n9695), .Y(_abc_17692_n9706) );
  OR2X2 OR2X2_3204 ( .A(_abc_17692_n9706), .B(_abc_17692_n9684), .Y(_abc_17692_n9707) );
  OR2X2 OR2X2_3205 ( .A(_abc_17692_n9707), .B(_abc_17692_n9671), .Y(_abc_17692_n9708) );
  OR2X2 OR2X2_3206 ( .A(_abc_17692_n9710), .B(_abc_17692_n9711), .Y(_abc_17692_n9712) );
  OR2X2 OR2X2_3207 ( .A(_abc_17692_n9709), .B(_abc_17692_n9712), .Y(_abc_17692_n9713) );
  OR2X2 OR2X2_3208 ( .A(_abc_17692_n9661), .B(_abc_17692_n9713), .Y(workunit1_10__FF_INPUT) );
  OR2X2 OR2X2_3209 ( .A(_abc_17692_n9568), .B(_abc_17692_n9552), .Y(_abc_17692_n9715) );
  OR2X2 OR2X2_321 ( .A(_abc_17692_n1439), .B(_abc_17692_n1437), .Y(_abc_17692_n1440) );
  OR2X2 OR2X2_3210 ( .A(_abc_17692_n3060), .B(workunit2_16_bF_buf1), .Y(_abc_17692_n9716) );
  OR2X2 OR2X2_3211 ( .A(_abc_17692_n9717), .B(workunit2_7_), .Y(_abc_17692_n9718) );
  OR2X2 OR2X2_3212 ( .A(_abc_17692_n9719), .B(_abc_17692_n3905), .Y(_abc_17692_n9720) );
  OR2X2 OR2X2_3213 ( .A(_abc_17692_n9721), .B(_abc_17692_n9722), .Y(_abc_17692_n9723) );
  OR2X2 OR2X2_3214 ( .A(_abc_17692_n9723), .B(workunit2_11_), .Y(_abc_17692_n9724) );
  OR2X2 OR2X2_3215 ( .A(_abc_17692_n9715), .B(_abc_17692_n9725), .Y(_abc_17692_n9726) );
  OR2X2 OR2X2_3216 ( .A(_abc_17692_n9548), .B(_abc_17692_n9557), .Y(_abc_17692_n9727) );
  OR2X2 OR2X2_3217 ( .A(_abc_17692_n9729), .B(_abc_17692_n9730), .Y(_abc_17692_n9731) );
  OR2X2 OR2X2_3218 ( .A(_abc_17692_n9728), .B(_abc_17692_n9731), .Y(_abc_17692_n9732) );
  OR2X2 OR2X2_3219 ( .A(_abc_17692_n3901), .B(_abc_17692_n9733), .Y(_abc_17692_n9734) );
  OR2X2 OR2X2_322 ( .A(_abc_17692_n1438), .B(_abc_17692_n1436), .Y(_abc_17692_n1441_1) );
  OR2X2 OR2X2_3220 ( .A(_abc_17692_n9735), .B(_abc_17692_n9736), .Y(_abc_17692_n9737) );
  OR2X2 OR2X2_3221 ( .A(_abc_17692_n3896), .B(_abc_17692_n9737), .Y(_abc_17692_n9738) );
  OR2X2 OR2X2_3222 ( .A(_abc_17692_n9742), .B(_abc_17692_n9743), .Y(_abc_17692_n9744) );
  OR2X2 OR2X2_3223 ( .A(_abc_17692_n9750), .B(_abc_17692_n9748), .Y(_abc_17692_n9751) );
  OR2X2 OR2X2_3224 ( .A(_abc_17692_n9752), .B(_abc_17692_n9747), .Y(_abc_17692_n9753) );
  OR2X2 OR2X2_3225 ( .A(_abc_17692_n9737), .B(_abc_17692_n3930_1), .Y(_abc_17692_n9756) );
  OR2X2 OR2X2_3226 ( .A(_abc_17692_n9733), .B(_abc_17692_n3934), .Y(_abc_17692_n9757) );
  OR2X2 OR2X2_3227 ( .A(_abc_17692_n9758), .B(_abc_17692_n2823), .Y(_abc_17692_n9759) );
  OR2X2 OR2X2_3228 ( .A(_abc_17692_n9733), .B(_abc_17692_n3930_1), .Y(_abc_17692_n9760) );
  OR2X2 OR2X2_3229 ( .A(_abc_17692_n9737), .B(_abc_17692_n3934), .Y(_abc_17692_n9761) );
  OR2X2 OR2X2_323 ( .A(_abc_17692_n1447), .B(_abc_17692_n1437), .Y(_abc_17692_n1448) );
  OR2X2 OR2X2_3230 ( .A(_abc_17692_n9762), .B(workunit1_11_bF_buf3), .Y(_abc_17692_n9763) );
  OR2X2 OR2X2_3231 ( .A(_abc_17692_n9769), .B(_abc_17692_n9765), .Y(_abc_17692_n9770) );
  OR2X2 OR2X2_3232 ( .A(_abc_17692_n9768), .B(_abc_17692_n9764), .Y(_abc_17692_n9771) );
  OR2X2 OR2X2_3233 ( .A(_abc_17692_n3959), .B(_abc_17692_n9733), .Y(_abc_17692_n9774) );
  OR2X2 OR2X2_3234 ( .A(_abc_17692_n3961), .B(_abc_17692_n9737), .Y(_abc_17692_n9775) );
  OR2X2 OR2X2_3235 ( .A(_abc_17692_n9778), .B(_abc_17692_n9779), .Y(_abc_17692_n9780) );
  OR2X2 OR2X2_3236 ( .A(_abc_17692_n9777), .B(_abc_17692_n9781), .Y(_abc_17692_n9782) );
  OR2X2 OR2X2_3237 ( .A(_abc_17692_n9786), .B(_abc_17692_n9782), .Y(_abc_17692_n9787) );
  OR2X2 OR2X2_3238 ( .A(_abc_17692_n9776), .B(workunit1_11_bF_buf1), .Y(_abc_17692_n9789) );
  OR2X2 OR2X2_3239 ( .A(_abc_17692_n9785), .B(_abc_17692_n9790), .Y(_abc_17692_n9791) );
  OR2X2 OR2X2_324 ( .A(_abc_17692_n1446), .B(_abc_17692_n1436), .Y(_abc_17692_n1449) );
  OR2X2 OR2X2_3240 ( .A(_abc_17692_n9793), .B(_abc_17692_n9773), .Y(_abc_17692_n9794) );
  OR2X2 OR2X2_3241 ( .A(_abc_17692_n9794), .B(_abc_17692_n9755), .Y(_abc_17692_n9795) );
  OR2X2 OR2X2_3242 ( .A(_abc_17692_n3989), .B(_abc_17692_n9737), .Y(_abc_17692_n9796) );
  OR2X2 OR2X2_3243 ( .A(_abc_17692_n3993), .B(_abc_17692_n9733), .Y(_abc_17692_n9797) );
  OR2X2 OR2X2_3244 ( .A(_abc_17692_n9798), .B(_abc_17692_n2823), .Y(_abc_17692_n9799) );
  OR2X2 OR2X2_3245 ( .A(_abc_17692_n3989), .B(_abc_17692_n9733), .Y(_abc_17692_n9800) );
  OR2X2 OR2X2_3246 ( .A(_abc_17692_n3993), .B(_abc_17692_n9737), .Y(_abc_17692_n9801) );
  OR2X2 OR2X2_3247 ( .A(_abc_17692_n9802), .B(workunit1_11_bF_buf0), .Y(_abc_17692_n9803) );
  OR2X2 OR2X2_3248 ( .A(_abc_17692_n9811), .B(_abc_17692_n9809), .Y(_abc_17692_n9812) );
  OR2X2 OR2X2_3249 ( .A(_abc_17692_n9813), .B(_abc_17692_n9795), .Y(_abc_17692_n9814) );
  OR2X2 OR2X2_325 ( .A(_abc_17692_n1452), .B(state_8_bF_buf7), .Y(_abc_17692_n1453) );
  OR2X2 OR2X2_3250 ( .A(_abc_17692_n9818), .B(_abc_17692_n9819), .Y(_abc_17692_n9820) );
  OR2X2 OR2X2_3251 ( .A(_abc_17692_n9825), .B(_abc_17692_n9748), .Y(_abc_17692_n9826) );
  OR2X2 OR2X2_3252 ( .A(_abc_17692_n9824), .B(_abc_17692_n9747), .Y(_abc_17692_n9827) );
  OR2X2 OR2X2_3253 ( .A(_abc_17692_n9831), .B(_abc_17692_n9764), .Y(_abc_17692_n9832) );
  OR2X2 OR2X2_3254 ( .A(_abc_17692_n9830), .B(_abc_17692_n9765), .Y(_abc_17692_n9833) );
  OR2X2 OR2X2_3255 ( .A(_abc_17692_n9837), .B(_abc_17692_n9790), .Y(_abc_17692_n9838) );
  OR2X2 OR2X2_3256 ( .A(_abc_17692_n9836), .B(_abc_17692_n9782), .Y(_abc_17692_n9839) );
  OR2X2 OR2X2_3257 ( .A(_abc_17692_n9841), .B(_abc_17692_n9835), .Y(_abc_17692_n9842) );
  OR2X2 OR2X2_3258 ( .A(_abc_17692_n9842), .B(_abc_17692_n9829), .Y(_abc_17692_n9843) );
  OR2X2 OR2X2_3259 ( .A(_abc_17692_n9843), .B(_abc_17692_n9821), .Y(_abc_17692_n9844) );
  OR2X2 OR2X2_326 ( .A(_abc_17692_n1451), .B(_abc_17692_n1453), .Y(_abc_17692_n1454) );
  OR2X2 OR2X2_3260 ( .A(_abc_17692_n9846), .B(_abc_17692_n9847), .Y(_abc_17692_n9848) );
  OR2X2 OR2X2_3261 ( .A(_abc_17692_n9845), .B(_abc_17692_n9848), .Y(_abc_17692_n9849) );
  OR2X2 OR2X2_3262 ( .A(_abc_17692_n9815), .B(_abc_17692_n9849), .Y(workunit1_11__FF_INPUT) );
  OR2X2 OR2X2_3263 ( .A(_abc_17692_n9853), .B(_abc_17692_n9730), .Y(_abc_17692_n9854) );
  OR2X2 OR2X2_3264 ( .A(_abc_17692_n9852), .B(_abc_17692_n9855), .Y(_abc_17692_n9856) );
  OR2X2 OR2X2_3265 ( .A(_abc_17692_n9557), .B(_abc_17692_n9731), .Y(_abc_17692_n9857) );
  OR2X2 OR2X2_3266 ( .A(_abc_17692_n9542), .B(_abc_17692_n9857), .Y(_abc_17692_n9858) );
  OR2X2 OR2X2_3267 ( .A(_abc_17692_n9860), .B(_abc_17692_n9856), .Y(_abc_17692_n9861) );
  OR2X2 OR2X2_3268 ( .A(_abc_17692_n9862), .B(_abc_17692_n9863), .Y(_abc_17692_n9864) );
  OR2X2 OR2X2_3269 ( .A(_abc_17692_n9864), .B(workunit2_12_bF_buf1), .Y(_abc_17692_n9867) );
  OR2X2 OR2X2_327 ( .A(_abc_17692_n1443), .B(_abc_17692_n1454), .Y(sum_19__FF_INPUT) );
  OR2X2 OR2X2_3270 ( .A(_abc_17692_n9857), .B(_abc_17692_n9547), .Y(_abc_17692_n9870) );
  OR2X2 OR2X2_3271 ( .A(_abc_17692_n9295), .B(_abc_17692_n9858), .Y(_abc_17692_n9872) );
  OR2X2 OR2X2_3272 ( .A(_abc_17692_n9874), .B(_abc_17692_n9865), .Y(_abc_17692_n9875) );
  OR2X2 OR2X2_3273 ( .A(_abc_17692_n9876), .B(_abc_17692_n9869), .Y(_abc_17692_n9877) );
  OR2X2 OR2X2_3274 ( .A(_abc_17692_n9878), .B(_abc_17692_n4137), .Y(_abc_17692_n9879) );
  OR2X2 OR2X2_3275 ( .A(_abc_17692_n4138), .B(_abc_17692_n9877), .Y(_abc_17692_n9880) );
  OR2X2 OR2X2_3276 ( .A(_abc_17692_n9883), .B(_abc_17692_n9884), .Y(_abc_17692_n9885) );
  OR2X2 OR2X2_3277 ( .A(_abc_17692_n9889), .B(_abc_17692_n9740), .Y(_abc_17692_n9890) );
  OR2X2 OR2X2_3278 ( .A(_abc_17692_n9892), .B(_abc_17692_n9891), .Y(_abc_17692_n9893) );
  OR2X2 OR2X2_3279 ( .A(_abc_17692_n9888), .B(_abc_17692_n9893), .Y(_abc_17692_n9894) );
  OR2X2 OR2X2_328 ( .A(_abc_17692_n1456), .B(delta_20_), .Y(_abc_17692_n1458) );
  OR2X2 OR2X2_3280 ( .A(_abc_17692_n9899), .B(_abc_17692_n9897), .Y(_abc_17692_n9900) );
  OR2X2 OR2X2_3281 ( .A(_abc_17692_n9900), .B(_abc_17692_n9896), .Y(_abc_17692_n9901) );
  OR2X2 OR2X2_3282 ( .A(_abc_17692_n9878), .B(_abc_17692_n4221), .Y(_abc_17692_n9902) );
  OR2X2 OR2X2_3283 ( .A(_abc_17692_n4222), .B(_abc_17692_n9877), .Y(_abc_17692_n9903) );
  OR2X2 OR2X2_3284 ( .A(_abc_17692_n9904), .B(workunit1_12_bF_buf2), .Y(_abc_17692_n9907) );
  OR2X2 OR2X2_3285 ( .A(_abc_17692_n9764), .B(_abc_17692_n9642), .Y(_abc_17692_n9909) );
  OR2X2 OR2X2_3286 ( .A(_abc_17692_n9645), .B(_abc_17692_n9909), .Y(_abc_17692_n9910) );
  OR2X2 OR2X2_3287 ( .A(_abc_17692_n9909), .B(_abc_17692_n9649), .Y(_abc_17692_n9911) );
  OR2X2 OR2X2_3288 ( .A(_abc_17692_n9764), .B(_abc_17692_n9767), .Y(_abc_17692_n9914) );
  OR2X2 OR2X2_3289 ( .A(_abc_17692_n9922), .B(_abc_17692_n9920), .Y(_abc_17692_n9923) );
  OR2X2 OR2X2_329 ( .A(_abc_17692_n1459_1), .B(_abc_17692_n1457), .Y(_abc_17692_n1460) );
  OR2X2 OR2X2_3290 ( .A(_abc_17692_n9923), .B(_abc_17692_n9919), .Y(_abc_17692_n9924) );
  OR2X2 OR2X2_3291 ( .A(_abc_17692_n9878), .B(_abc_17692_n4177), .Y(_abc_17692_n9925) );
  OR2X2 OR2X2_3292 ( .A(_abc_17692_n4178), .B(_abc_17692_n9877), .Y(_abc_17692_n9926) );
  OR2X2 OR2X2_3293 ( .A(_abc_17692_n9927), .B(workunit1_12_bF_buf0), .Y(_abc_17692_n9930) );
  OR2X2 OR2X2_3294 ( .A(_abc_17692_n9937), .B(_abc_17692_n9938), .Y(_abc_17692_n9939) );
  OR2X2 OR2X2_3295 ( .A(_abc_17692_n9936), .B(_abc_17692_n9939), .Y(_abc_17692_n9940) );
  OR2X2 OR2X2_3296 ( .A(_abc_17692_n9935), .B(_abc_17692_n9940), .Y(_abc_17692_n9941) );
  OR2X2 OR2X2_3297 ( .A(_abc_17692_n9945), .B(_abc_17692_n9944), .Y(_abc_17692_n9946) );
  OR2X2 OR2X2_3298 ( .A(_abc_17692_n9946), .B(_abc_17692_n9943), .Y(_abc_17692_n9947) );
  OR2X2 OR2X2_3299 ( .A(_abc_17692_n4093), .B(_abc_17692_n9878), .Y(_abc_17692_n9950) );
  OR2X2 OR2X2_33 ( .A(_abc_17692_n704), .B(_abc_17692_n699), .Y(_abc_17692_n705) );
  OR2X2 OR2X2_330 ( .A(_abc_17692_n1462), .B(_abc_17692_n1408), .Y(_abc_17692_n1463) );
  OR2X2 OR2X2_3300 ( .A(_abc_17692_n4094), .B(_abc_17692_n9877), .Y(_abc_17692_n9951) );
  OR2X2 OR2X2_3301 ( .A(_abc_17692_n9952), .B(workunit1_12_bF_buf2), .Y(_abc_17692_n9955) );
  OR2X2 OR2X2_3302 ( .A(_abc_17692_n9961), .B(_abc_17692_n9962), .Y(_abc_17692_n9963) );
  OR2X2 OR2X2_3303 ( .A(_abc_17692_n9960), .B(_abc_17692_n9963), .Y(_abc_17692_n9964) );
  OR2X2 OR2X2_3304 ( .A(_abc_17692_n9959), .B(_abc_17692_n9964), .Y(_abc_17692_n9965) );
  OR2X2 OR2X2_3305 ( .A(_abc_17692_n9968), .B(_abc_17692_n4047_bF_buf3), .Y(_abc_17692_n9969) );
  OR2X2 OR2X2_3306 ( .A(_abc_17692_n9969), .B(_abc_17692_n9967), .Y(_abc_17692_n9970) );
  OR2X2 OR2X2_3307 ( .A(_abc_17692_n9971), .B(_abc_17692_n627), .Y(_abc_17692_n9972) );
  OR2X2 OR2X2_3308 ( .A(_abc_17692_n9978), .B(_abc_17692_n9976), .Y(_abc_17692_n9979) );
  OR2X2 OR2X2_3309 ( .A(_abc_17692_n9980), .B(_abc_17692_n9979), .Y(_abc_17692_n9981) );
  OR2X2 OR2X2_331 ( .A(_abc_17692_n1464), .B(_abc_17692_n1430), .Y(_abc_17692_n1465) );
  OR2X2 OR2X2_3310 ( .A(_abc_17692_n9975), .B(_abc_17692_n9981), .Y(_abc_17692_n9982) );
  OR2X2 OR2X2_3311 ( .A(_abc_17692_n9985), .B(_abc_17692_n4047_bF_buf2), .Y(_abc_17692_n9986) );
  OR2X2 OR2X2_3312 ( .A(_abc_17692_n9986), .B(_abc_17692_n9983), .Y(_abc_17692_n9987) );
  OR2X2 OR2X2_3313 ( .A(_abc_17692_n9747), .B(_abc_17692_n9600), .Y(_abc_17692_n9988) );
  OR2X2 OR2X2_3314 ( .A(_abc_17692_n9988), .B(_abc_17692_n9677), .Y(_abc_17692_n9993) );
  OR2X2 OR2X2_3315 ( .A(_abc_17692_n9747), .B(_abc_17692_n9823), .Y(_abc_17692_n9996) );
  OR2X2 OR2X2_3316 ( .A(_abc_17692_n10001), .B(_abc_17692_n9991), .Y(_abc_17692_n10002) );
  OR2X2 OR2X2_3317 ( .A(_abc_17692_n10003), .B(_abc_17692_n9897), .Y(_abc_17692_n10004) );
  OR2X2 OR2X2_3318 ( .A(_abc_17692_n10004), .B(_abc_17692_n10000), .Y(_abc_17692_n10005) );
  OR2X2 OR2X2_3319 ( .A(_abc_17692_n10009), .B(_abc_17692_n10007), .Y(_abc_17692_n10010) );
  OR2X2 OR2X2_332 ( .A(_abc_17692_n1406), .B(_abc_17692_n1462), .Y(_abc_17692_n1468) );
  OR2X2 OR2X2_3320 ( .A(_abc_17692_n10006), .B(_abc_17692_n10010), .Y(_abc_17692_n10011) );
  OR2X2 OR2X2_3321 ( .A(_abc_17692_n10013), .B(_abc_17692_n10012), .Y(_abc_17692_n10014) );
  OR2X2 OR2X2_3322 ( .A(_abc_17692_n10009), .B(_abc_17692_n10017), .Y(_abc_17692_n10018) );
  OR2X2 OR2X2_3323 ( .A(_abc_17692_n10015), .B(_abc_17692_n9689), .Y(_abc_17692_n10022) );
  OR2X2 OR2X2_3324 ( .A(_abc_17692_n9686), .B(_abc_17692_n10022), .Y(_abc_17692_n10023) );
  OR2X2 OR2X2_3325 ( .A(_abc_17692_n10015), .B(_abc_17692_n10008), .Y(_abc_17692_n10024) );
  OR2X2 OR2X2_3326 ( .A(_abc_17692_n10026), .B(_abc_17692_n9920), .Y(_abc_17692_n10027) );
  OR2X2 OR2X2_3327 ( .A(_abc_17692_n10027), .B(_abc_17692_n10021), .Y(_abc_17692_n10028) );
  OR2X2 OR2X2_3328 ( .A(_abc_17692_n9781), .B(_abc_17692_n9616), .Y(_abc_17692_n10032) );
  OR2X2 OR2X2_3329 ( .A(_abc_17692_n10035), .B(_abc_17692_n10034), .Y(_abc_17692_n10036) );
  OR2X2 OR2X2_333 ( .A(_abc_17692_n1470), .B(_abc_17692_n1460), .Y(_abc_17692_n1471) );
  OR2X2 OR2X2_3330 ( .A(_abc_17692_n10036), .B(_abc_17692_n10031), .Y(_abc_17692_n10037) );
  OR2X2 OR2X2_3331 ( .A(_abc_17692_n10041), .B(_abc_17692_n9399), .Y(_abc_17692_n10042) );
  OR2X2 OR2X2_3332 ( .A(_abc_17692_n9782), .B(_abc_17692_n9619), .Y(_abc_17692_n10045) );
  OR2X2 OR2X2_3333 ( .A(_abc_17692_n10045), .B(_abc_17692_n10044), .Y(_abc_17692_n10046) );
  OR2X2 OR2X2_3334 ( .A(_abc_17692_n10043), .B(_abc_17692_n10046), .Y(_abc_17692_n10047) );
  OR2X2 OR2X2_3335 ( .A(_abc_17692_n10045), .B(_abc_17692_n10048), .Y(_abc_17692_n10049) );
  OR2X2 OR2X2_3336 ( .A(_abc_17692_n10052), .B(_abc_17692_n9944), .Y(_abc_17692_n10053) );
  OR2X2 OR2X2_3337 ( .A(_abc_17692_n10053), .B(_abc_17692_n10038), .Y(_abc_17692_n10054) );
  OR2X2 OR2X2_3338 ( .A(_abc_17692_n10057), .B(_abc_17692_n712), .Y(_abc_17692_n10058) );
  OR2X2 OR2X2_3339 ( .A(_abc_17692_n10059), .B(_abc_17692_n3026), .Y(_abc_17692_n10060) );
  OR2X2 OR2X2_334 ( .A(_abc_17692_n1482), .B(_abc_17692_n1483), .Y(_abc_17692_n1484) );
  OR2X2 OR2X2_3340 ( .A(_abc_17692_n9869), .B(_abc_17692_n9865), .Y(_abc_17692_n10067) );
  OR2X2 OR2X2_3341 ( .A(_abc_17692_n10068), .B(_abc_17692_n10069), .Y(_abc_17692_n10070) );
  OR2X2 OR2X2_3342 ( .A(_abc_17692_n10070), .B(workunit2_13_), .Y(_abc_17692_n10072) );
  OR2X2 OR2X2_3343 ( .A(_abc_17692_n10073), .B(_abc_17692_n10071), .Y(_abc_17692_n10074) );
  OR2X2 OR2X2_3344 ( .A(_abc_17692_n10067), .B(_abc_17692_n10074), .Y(_abc_17692_n10077) );
  OR2X2 OR2X2_3345 ( .A(_abc_17692_n4426), .B(_abc_17692_n10078), .Y(_abc_17692_n10079) );
  OR2X2 OR2X2_3346 ( .A(_abc_17692_n4428), .B(_abc_17692_n10080), .Y(_abc_17692_n10081) );
  OR2X2 OR2X2_3347 ( .A(_abc_17692_n10085), .B(_abc_17692_n10083), .Y(_abc_17692_n10086) );
  OR2X2 OR2X2_3348 ( .A(_abc_17692_n9968), .B(_abc_17692_n9953), .Y(_abc_17692_n10088) );
  OR2X2 OR2X2_3349 ( .A(_abc_17692_n10091), .B(_abc_17692_n4047_bF_buf1), .Y(_abc_17692_n10092) );
  OR2X2 OR2X2_335 ( .A(_abc_17692_n1481), .B(_abc_17692_n1484), .Y(_abc_17692_n1485) );
  OR2X2 OR2X2_3350 ( .A(_abc_17692_n10092), .B(_abc_17692_n10089), .Y(_abc_17692_n10093) );
  OR2X2 OR2X2_3351 ( .A(_abc_17692_n4346), .B(_abc_17692_n10078), .Y(_abc_17692_n10094) );
  OR2X2 OR2X2_3352 ( .A(_abc_17692_n10080), .B(_abc_17692_n4344_1), .Y(_abc_17692_n10095) );
  OR2X2 OR2X2_3353 ( .A(_abc_17692_n10099), .B(_abc_17692_n10097), .Y(_abc_17692_n10100) );
  OR2X2 OR2X2_3354 ( .A(_abc_17692_n9899), .B(_abc_17692_n9884), .Y(_abc_17692_n10102) );
  OR2X2 OR2X2_3355 ( .A(_abc_17692_n10103), .B(_abc_17692_n10101), .Y(_abc_17692_n10104) );
  OR2X2 OR2X2_3356 ( .A(_abc_17692_n10102), .B(_abc_17692_n10100), .Y(_abc_17692_n10105) );
  OR2X2 OR2X2_3357 ( .A(_abc_17692_n10078), .B(_abc_17692_n4399), .Y(_abc_17692_n10108) );
  OR2X2 OR2X2_3358 ( .A(_abc_17692_n10080), .B(_abc_17692_n4401), .Y(_abc_17692_n10109) );
  OR2X2 OR2X2_3359 ( .A(_abc_17692_n10110), .B(workunit1_13_bF_buf1), .Y(_abc_17692_n10113) );
  OR2X2 OR2X2_336 ( .A(_abc_17692_n1479), .B(_abc_17692_n1485), .Y(_abc_17692_n1486) );
  OR2X2 OR2X2_3360 ( .A(_abc_17692_n9945), .B(_abc_17692_n9928), .Y(_abc_17692_n10116) );
  OR2X2 OR2X2_3361 ( .A(_abc_17692_n10116), .B(_abc_17692_n10115), .Y(_abc_17692_n10117) );
  OR2X2 OR2X2_3362 ( .A(_abc_17692_n10118), .B(_abc_17692_n10114), .Y(_abc_17692_n10119) );
  OR2X2 OR2X2_3363 ( .A(_abc_17692_n4371), .B(_abc_17692_n10078), .Y(_abc_17692_n10122) );
  OR2X2 OR2X2_3364 ( .A(_abc_17692_n10080), .B(_abc_17692_n4374), .Y(_abc_17692_n10123) );
  OR2X2 OR2X2_3365 ( .A(_abc_17692_n10124), .B(_abc_17692_n3208), .Y(_abc_17692_n10125) );
  OR2X2 OR2X2_3366 ( .A(_abc_17692_n4374), .B(_abc_17692_n10078), .Y(_abc_17692_n10126) );
  OR2X2 OR2X2_3367 ( .A(_abc_17692_n4371), .B(_abc_17692_n10080), .Y(_abc_17692_n10127) );
  OR2X2 OR2X2_3368 ( .A(_abc_17692_n10128), .B(workunit1_13_bF_buf0), .Y(_abc_17692_n10129) );
  OR2X2 OR2X2_3369 ( .A(_abc_17692_n10134), .B(_abc_17692_n10131), .Y(_abc_17692_n10135) );
  OR2X2 OR2X2_337 ( .A(_abc_17692_n1486), .B(_abc_17692_n1477), .Y(_abc_17692_n1489) );
  OR2X2 OR2X2_3370 ( .A(_abc_17692_n10133), .B(_abc_17692_n10130), .Y(_abc_17692_n10136) );
  OR2X2 OR2X2_3371 ( .A(_abc_17692_n10138), .B(_abc_17692_n1863_bF_buf0), .Y(_abc_17692_n10139) );
  OR2X2 OR2X2_3372 ( .A(_abc_17692_n10121), .B(_abc_17692_n10139), .Y(_abc_17692_n10140) );
  OR2X2 OR2X2_3373 ( .A(_abc_17692_n10140), .B(_abc_17692_n10107), .Y(_abc_17692_n10141) );
  OR2X2 OR2X2_3374 ( .A(_abc_17692_n9983), .B(_abc_17692_n10145), .Y(_abc_17692_n10146) );
  OR2X2 OR2X2_3375 ( .A(_abc_17692_n10149), .B(_abc_17692_n10147), .Y(_abc_17692_n10150) );
  OR2X2 OR2X2_3376 ( .A(_abc_17692_n10003), .B(_abc_17692_n10152), .Y(_abc_17692_n10153) );
  OR2X2 OR2X2_3377 ( .A(_abc_17692_n10153), .B(_abc_17692_n10101), .Y(_abc_17692_n10154) );
  OR2X2 OR2X2_3378 ( .A(_abc_17692_n10155), .B(_abc_17692_n10100), .Y(_abc_17692_n10156) );
  OR2X2 OR2X2_3379 ( .A(_abc_17692_n10038), .B(_abc_17692_n10160), .Y(_abc_17692_n10161) );
  OR2X2 OR2X2_338 ( .A(_abc_17692_n1491), .B(_abc_17692_n1476), .Y(_abc_17692_n1492) );
  OR2X2 OR2X2_3380 ( .A(_abc_17692_n10162), .B(_abc_17692_n10115), .Y(_abc_17692_n10163) );
  OR2X2 OR2X2_3381 ( .A(_abc_17692_n10161), .B(_abc_17692_n10114), .Y(_abc_17692_n10164) );
  OR2X2 OR2X2_3382 ( .A(_abc_17692_n10026), .B(_abc_17692_n10168), .Y(_abc_17692_n10169) );
  OR2X2 OR2X2_3383 ( .A(_abc_17692_n10172), .B(_abc_17692_n10170), .Y(_abc_17692_n10173) );
  OR2X2 OR2X2_3384 ( .A(_abc_17692_n10174), .B(_abc_17692_n10166), .Y(_abc_17692_n10175) );
  OR2X2 OR2X2_3385 ( .A(_abc_17692_n10175), .B(_abc_17692_n10158), .Y(_abc_17692_n10176) );
  OR2X2 OR2X2_3386 ( .A(_abc_17692_n10176), .B(_abc_17692_n10151), .Y(_abc_17692_n10177) );
  OR2X2 OR2X2_3387 ( .A(_abc_17692_n10179), .B(_abc_17692_n10180), .Y(_abc_17692_n10181) );
  OR2X2 OR2X2_3388 ( .A(_abc_17692_n10178), .B(_abc_17692_n10181), .Y(_abc_17692_n10182) );
  OR2X2 OR2X2_3389 ( .A(_abc_17692_n10182), .B(_abc_17692_n10143), .Y(workunit1_13__FF_INPUT) );
  OR2X2 OR2X2_339 ( .A(_abc_17692_n1475), .B(_abc_17692_n1492), .Y(sum_20__FF_INPUT) );
  OR2X2 OR2X2_3390 ( .A(_abc_17692_n9873), .B(_abc_17692_n10187), .Y(_abc_17692_n10188) );
  OR2X2 OR2X2_3391 ( .A(_abc_17692_n9865), .B(_abc_17692_n10071), .Y(_abc_17692_n10189) );
  OR2X2 OR2X2_3392 ( .A(_abc_17692_n10193), .B(_abc_17692_n10194), .Y(_abc_17692_n10195) );
  OR2X2 OR2X2_3393 ( .A(_abc_17692_n10195), .B(workunit2_14_bF_buf2), .Y(_abc_17692_n10197) );
  OR2X2 OR2X2_3394 ( .A(_abc_17692_n10198), .B(_abc_17692_n10196), .Y(_abc_17692_n10199) );
  OR2X2 OR2X2_3395 ( .A(_abc_17692_n10201), .B(_abc_17692_n10190), .Y(_abc_17692_n10202) );
  OR2X2 OR2X2_3396 ( .A(_abc_17692_n10200), .B(_abc_17692_n10205), .Y(_abc_17692_n10206) );
  OR2X2 OR2X2_3397 ( .A(_abc_17692_n10207), .B(_abc_17692_n10209), .Y(_abc_17692_n10210) );
  OR2X2 OR2X2_3398 ( .A(_abc_17692_n10211), .B(_abc_17692_n5376), .Y(_abc_17692_n10212) );
  OR2X2 OR2X2_3399 ( .A(_abc_17692_n10210), .B(workunit1_14_bF_buf0), .Y(_abc_17692_n10213) );
  OR2X2 OR2X2_34 ( .A(while_flag), .B(state_4_), .Y(_abc_17692_n706) );
  OR2X2 OR2X2_340 ( .A(_abc_17692_n1504), .B(_abc_17692_n1500), .Y(_abc_17692_n1505) );
  OR2X2 OR2X2_3400 ( .A(_abc_17692_n10083), .B(_abc_17692_n10145), .Y(_abc_17692_n10216) );
  OR2X2 OR2X2_3401 ( .A(_abc_17692_n10219), .B(_abc_17692_n10217), .Y(_abc_17692_n10220) );
  OR2X2 OR2X2_3402 ( .A(_abc_17692_n10220), .B(_abc_17692_n10214), .Y(_abc_17692_n10221) );
  OR2X2 OR2X2_3403 ( .A(_abc_17692_n10208), .B(_abc_17692_n4565), .Y(_abc_17692_n10226) );
  OR2X2 OR2X2_3404 ( .A(_abc_17692_n4566), .B(_abc_17692_n10206), .Y(_abc_17692_n10227) );
  OR2X2 OR2X2_3405 ( .A(_abc_17692_n10228), .B(workunit1_14_bF_buf2), .Y(_abc_17692_n10231) );
  OR2X2 OR2X2_3406 ( .A(_abc_17692_n10097), .B(_abc_17692_n10152), .Y(_abc_17692_n10235) );
  OR2X2 OR2X2_3407 ( .A(_abc_17692_n10238), .B(_abc_17692_n10236), .Y(_abc_17692_n10239) );
  OR2X2 OR2X2_3408 ( .A(_abc_17692_n10239), .B(_abc_17692_n10233), .Y(_abc_17692_n10242) );
  OR2X2 OR2X2_3409 ( .A(_abc_17692_n10246), .B(_abc_17692_n10245), .Y(_abc_17692_n10247) );
  OR2X2 OR2X2_341 ( .A(_abc_17692_n1503), .B(_abc_17692_n1506), .Y(_abc_17692_n1507) );
  OR2X2 OR2X2_3410 ( .A(_abc_17692_n10248), .B(_abc_17692_n5376), .Y(_abc_17692_n10249) );
  OR2X2 OR2X2_3411 ( .A(_abc_17692_n10247), .B(workunit1_14_bF_buf1), .Y(_abc_17692_n10250) );
  OR2X2 OR2X2_3412 ( .A(_abc_17692_n10252), .B(_abc_17692_n10168), .Y(_abc_17692_n10253) );
  OR2X2 OR2X2_3413 ( .A(_abc_17692_n10256), .B(_abc_17692_n10254), .Y(_abc_17692_n10257) );
  OR2X2 OR2X2_3414 ( .A(_abc_17692_n10257), .B(_abc_17692_n10251), .Y(_abc_17692_n10260) );
  OR2X2 OR2X2_3415 ( .A(_abc_17692_n10263), .B(_abc_17692_n10264), .Y(_abc_17692_n10265) );
  OR2X2 OR2X2_3416 ( .A(_abc_17692_n10266), .B(_abc_17692_n5376), .Y(_abc_17692_n10267) );
  OR2X2 OR2X2_3417 ( .A(_abc_17692_n10265), .B(workunit1_14_bF_buf0), .Y(_abc_17692_n10268) );
  OR2X2 OR2X2_3418 ( .A(_abc_17692_n10111), .B(_abc_17692_n10160), .Y(_abc_17692_n10270) );
  OR2X2 OR2X2_3419 ( .A(_abc_17692_n10273), .B(_abc_17692_n10271), .Y(_abc_17692_n10274) );
  OR2X2 OR2X2_342 ( .A(_abc_17692_n1506), .B(_abc_17692_n1459_1), .Y(_abc_17692_n1510) );
  OR2X2 OR2X2_3420 ( .A(_abc_17692_n10274), .B(_abc_17692_n10269), .Y(_abc_17692_n10277) );
  OR2X2 OR2X2_3421 ( .A(_abc_17692_n10262), .B(_abc_17692_n10279), .Y(_abc_17692_n10280) );
  OR2X2 OR2X2_3422 ( .A(_abc_17692_n10280), .B(_abc_17692_n10244), .Y(_abc_17692_n10281) );
  OR2X2 OR2X2_3423 ( .A(_abc_17692_n10281), .B(_abc_17692_n10225), .Y(_abc_17692_n10282) );
  OR2X2 OR2X2_3424 ( .A(_abc_17692_n10285), .B(_abc_17692_n10284), .Y(_abc_17692_n10286) );
  OR2X2 OR2X2_3425 ( .A(_abc_17692_n10288), .B(_abc_17692_n10286), .Y(_abc_17692_n10289) );
  OR2X2 OR2X2_3426 ( .A(_abc_17692_n10289), .B(_abc_17692_n10232), .Y(_abc_17692_n10292) );
  OR2X2 OR2X2_3427 ( .A(_abc_17692_n10130), .B(_abc_17692_n9906), .Y(_abc_17692_n10298) );
  OR2X2 OR2X2_3428 ( .A(_abc_17692_n10130), .B(_abc_17692_n9921), .Y(_abc_17692_n10301) );
  OR2X2 OR2X2_3429 ( .A(_abc_17692_n10303), .B(_abc_17692_n10300), .Y(_abc_17692_n10304) );
  OR2X2 OR2X2_343 ( .A(_abc_17692_n1487), .B(_abc_17692_n1510), .Y(_abc_17692_n1511) );
  OR2X2 OR2X2_3430 ( .A(_abc_17692_n10304), .B(_abc_17692_n10295), .Y(_abc_17692_n10307) );
  OR2X2 OR2X2_3431 ( .A(_abc_17692_n10313), .B(_abc_17692_n10312), .Y(_abc_17692_n10314) );
  OR2X2 OR2X2_3432 ( .A(_abc_17692_n10316), .B(_abc_17692_n10314), .Y(_abc_17692_n10317) );
  OR2X2 OR2X2_3433 ( .A(_abc_17692_n10317), .B(_abc_17692_n10310), .Y(_abc_17692_n10320) );
  OR2X2 OR2X2_3434 ( .A(_abc_17692_n10322), .B(_abc_17692_n10309), .Y(_abc_17692_n10323) );
  OR2X2 OR2X2_3435 ( .A(_abc_17692_n10323), .B(_abc_17692_n10294), .Y(_abc_17692_n10324) );
  OR2X2 OR2X2_3436 ( .A(_abc_17692_n10327), .B(_abc_17692_n10326), .Y(_abc_17692_n10328) );
  OR2X2 OR2X2_3437 ( .A(_abc_17692_n10330), .B(_abc_17692_n10328), .Y(_abc_17692_n10331) );
  OR2X2 OR2X2_3438 ( .A(_abc_17692_n10331), .B(_abc_17692_n10325), .Y(_abc_17692_n10334) );
  OR2X2 OR2X2_3439 ( .A(_abc_17692_n10336), .B(_abc_17692_n10324), .Y(_abc_17692_n10337) );
  OR2X2 OR2X2_344 ( .A(_abc_17692_n1520_1), .B(state_8_bF_buf6), .Y(_abc_17692_n1521) );
  OR2X2 OR2X2_3440 ( .A(_abc_17692_n10339), .B(_abc_17692_n10340), .Y(_abc_17692_n10341) );
  OR2X2 OR2X2_3441 ( .A(_abc_17692_n10338), .B(_abc_17692_n10341), .Y(_abc_17692_n10342) );
  OR2X2 OR2X2_3442 ( .A(_abc_17692_n10342), .B(_abc_17692_n10283), .Y(workunit1_14__FF_INPUT) );
  OR2X2 OR2X2_3443 ( .A(_abc_17692_n10205), .B(_abc_17692_n10196), .Y(_abc_17692_n10344) );
  OR2X2 OR2X2_3444 ( .A(_abc_17692_n10345), .B(_abc_17692_n10346), .Y(_abc_17692_n10347) );
  OR2X2 OR2X2_3445 ( .A(_abc_17692_n10347), .B(workunit2_15_), .Y(_abc_17692_n10350) );
  OR2X2 OR2X2_3446 ( .A(_abc_17692_n10344), .B(_abc_17692_n10351), .Y(_abc_17692_n10352) );
  OR2X2 OR2X2_3447 ( .A(_abc_17692_n10192), .B(_abc_17692_n10199), .Y(_abc_17692_n10353) );
  OR2X2 OR2X2_3448 ( .A(_abc_17692_n10355), .B(_abc_17692_n10348), .Y(_abc_17692_n10356) );
  OR2X2 OR2X2_3449 ( .A(_abc_17692_n10354), .B(_abc_17692_n10356), .Y(_abc_17692_n10357) );
  OR2X2 OR2X2_345 ( .A(_abc_17692_n1519), .B(_abc_17692_n1521), .Y(_abc_17692_n1522) );
  OR2X2 OR2X2_3450 ( .A(_abc_17692_n4761), .B(_abc_17692_n10358), .Y(_abc_17692_n10359) );
  OR2X2 OR2X2_3451 ( .A(_abc_17692_n10360), .B(_abc_17692_n10361), .Y(_abc_17692_n10362) );
  OR2X2 OR2X2_3452 ( .A(_abc_17692_n4756), .B(_abc_17692_n10362), .Y(_abc_17692_n10363) );
  OR2X2 OR2X2_3453 ( .A(_abc_17692_n10365), .B(workunit1_15_), .Y(_abc_17692_n10366) );
  OR2X2 OR2X2_3454 ( .A(_abc_17692_n10364), .B(_abc_17692_n3614), .Y(_abc_17692_n10367) );
  OR2X2 OR2X2_3455 ( .A(_abc_17692_n10376), .B(_abc_17692_n10374), .Y(_abc_17692_n10377) );
  OR2X2 OR2X2_3456 ( .A(_abc_17692_n4850), .B(_abc_17692_n10362), .Y(_abc_17692_n10379) );
  OR2X2 OR2X2_3457 ( .A(_abc_17692_n4854), .B(_abc_17692_n10358), .Y(_abc_17692_n10380) );
  OR2X2 OR2X2_3458 ( .A(_abc_17692_n10381), .B(_abc_17692_n3614), .Y(_abc_17692_n10382) );
  OR2X2 OR2X2_3459 ( .A(_abc_17692_n4850), .B(_abc_17692_n10358), .Y(_abc_17692_n10383) );
  OR2X2 OR2X2_346 ( .A(_abc_17692_n1509), .B(_abc_17692_n1522), .Y(sum_21__FF_INPUT) );
  OR2X2 OR2X2_3460 ( .A(_abc_17692_n4854), .B(_abc_17692_n10362), .Y(_abc_17692_n10384) );
  OR2X2 OR2X2_3461 ( .A(_abc_17692_n10385), .B(workunit1_15_), .Y(_abc_17692_n10386) );
  OR2X2 OR2X2_3462 ( .A(_abc_17692_n10389), .B(_abc_17692_n10387), .Y(_abc_17692_n10390) );
  OR2X2 OR2X2_3463 ( .A(_abc_17692_n10388), .B(_abc_17692_n10391), .Y(_abc_17692_n10392) );
  OR2X2 OR2X2_3464 ( .A(_abc_17692_n10362), .B(_abc_17692_n4815), .Y(_abc_17692_n10395) );
  OR2X2 OR2X2_3465 ( .A(_abc_17692_n10358), .B(_abc_17692_n4819), .Y(_abc_17692_n10396) );
  OR2X2 OR2X2_3466 ( .A(_abc_17692_n10397), .B(_abc_17692_n3614), .Y(_abc_17692_n10398) );
  OR2X2 OR2X2_3467 ( .A(_abc_17692_n10358), .B(_abc_17692_n4815), .Y(_abc_17692_n10399) );
  OR2X2 OR2X2_3468 ( .A(_abc_17692_n10362), .B(_abc_17692_n4819), .Y(_abc_17692_n10400) );
  OR2X2 OR2X2_3469 ( .A(_abc_17692_n10401), .B(workunit1_15_), .Y(_abc_17692_n10402) );
  OR2X2 OR2X2_347 ( .A(_abc_17692_n1527), .B(_abc_17692_n1524), .Y(_abc_17692_n1528) );
  OR2X2 OR2X2_3470 ( .A(_abc_17692_n10405), .B(_abc_17692_n10403), .Y(_abc_17692_n10406) );
  OR2X2 OR2X2_3471 ( .A(_abc_17692_n10404), .B(_abc_17692_n10407), .Y(_abc_17692_n10408) );
  OR2X2 OR2X2_3472 ( .A(_abc_17692_n4787), .B(_abc_17692_n10358), .Y(_abc_17692_n10411) );
  OR2X2 OR2X2_3473 ( .A(_abc_17692_n4789_1), .B(_abc_17692_n10362), .Y(_abc_17692_n10412) );
  OR2X2 OR2X2_3474 ( .A(_abc_17692_n10415), .B(_abc_17692_n10416), .Y(_abc_17692_n10417) );
  OR2X2 OR2X2_3475 ( .A(_abc_17692_n10414), .B(_abc_17692_n10418), .Y(_abc_17692_n10419) );
  OR2X2 OR2X2_3476 ( .A(_abc_17692_n10420), .B(_abc_17692_n10419), .Y(_abc_17692_n10421) );
  OR2X2 OR2X2_3477 ( .A(_abc_17692_n10425), .B(_abc_17692_n10424), .Y(_abc_17692_n10426) );
  OR2X2 OR2X2_3478 ( .A(_abc_17692_n10428), .B(_abc_17692_n10410), .Y(_abc_17692_n10429) );
  OR2X2 OR2X2_3479 ( .A(_abc_17692_n10429), .B(_abc_17692_n10394), .Y(_abc_17692_n10430) );
  OR2X2 OR2X2_348 ( .A(_abc_17692_n1530), .B(_abc_17692_n1498), .Y(_abc_17692_n1531) );
  OR2X2 OR2X2_3480 ( .A(_abc_17692_n10430), .B(_abc_17692_n10378), .Y(_abc_17692_n10431) );
  OR2X2 OR2X2_3481 ( .A(_abc_17692_n10433), .B(_abc_17692_n10369), .Y(_abc_17692_n10434) );
  OR2X2 OR2X2_3482 ( .A(_abc_17692_n10435), .B(_abc_17692_n10368), .Y(_abc_17692_n10436) );
  OR2X2 OR2X2_3483 ( .A(_abc_17692_n10442), .B(_abc_17692_n10419), .Y(_abc_17692_n10443) );
  OR2X2 OR2X2_3484 ( .A(_abc_17692_n10441), .B(_abc_17692_n10424), .Y(_abc_17692_n10444) );
  OR2X2 OR2X2_3485 ( .A(_abc_17692_n10450), .B(_abc_17692_n10407), .Y(_abc_17692_n10451) );
  OR2X2 OR2X2_3486 ( .A(_abc_17692_n10449), .B(_abc_17692_n10403), .Y(_abc_17692_n10452) );
  OR2X2 OR2X2_3487 ( .A(_abc_17692_n10446), .B(_abc_17692_n10454), .Y(_abc_17692_n10455) );
  OR2X2 OR2X2_3488 ( .A(_abc_17692_n10455), .B(_abc_17692_n10438), .Y(_abc_17692_n10456) );
  OR2X2 OR2X2_3489 ( .A(_abc_17692_n10460), .B(_abc_17692_n10391), .Y(_abc_17692_n10461) );
  OR2X2 OR2X2_349 ( .A(_abc_17692_n1534), .B(_abc_17692_n1532), .Y(_abc_17692_n1535) );
  OR2X2 OR2X2_3490 ( .A(_abc_17692_n10459), .B(_abc_17692_n10387), .Y(_abc_17692_n10462) );
  OR2X2 OR2X2_3491 ( .A(_abc_17692_n10464), .B(_abc_17692_n10456), .Y(_abc_17692_n10465) );
  OR2X2 OR2X2_3492 ( .A(_abc_17692_n10467), .B(_abc_17692_n10468), .Y(_abc_17692_n10469) );
  OR2X2 OR2X2_3493 ( .A(_abc_17692_n10466), .B(_abc_17692_n10469), .Y(_abc_17692_n10470) );
  OR2X2 OR2X2_3494 ( .A(_abc_17692_n10470), .B(_abc_17692_n10432), .Y(workunit1_15__FF_INPUT) );
  OR2X2 OR2X2_3495 ( .A(_abc_17692_n10474), .B(_abc_17692_n9858), .Y(_abc_17692_n10475) );
  OR2X2 OR2X2_3496 ( .A(_abc_17692_n9295), .B(_abc_17692_n10475), .Y(_abc_17692_n10476) );
  OR2X2 OR2X2_3497 ( .A(_abc_17692_n9871), .B(_abc_17692_n10474), .Y(_abc_17692_n10477) );
  OR2X2 OR2X2_3498 ( .A(_abc_17692_n10479), .B(_abc_17692_n10348), .Y(_abc_17692_n10480) );
  OR2X2 OR2X2_3499 ( .A(_abc_17692_n10478), .B(_abc_17692_n10480), .Y(_abc_17692_n10481) );
  OR2X2 OR2X2_35 ( .A(state_13_), .B(state_12_), .Y(_abc_17692_n708) );
  OR2X2 OR2X2_350 ( .A(_abc_17692_n1535), .B(_abc_17692_n1529), .Y(_abc_17692_n1536) );
  OR2X2 OR2X2_3500 ( .A(_abc_17692_n4120), .B(workunit2_21_), .Y(_abc_17692_n10485) );
  OR2X2 OR2X2_3501 ( .A(_abc_17692_n6095), .B(workunit2_12_bF_buf0), .Y(_abc_17692_n10486) );
  OR2X2 OR2X2_3502 ( .A(_abc_17692_n10489), .B(_abc_17692_n10490), .Y(_abc_17692_n10491) );
  OR2X2 OR2X2_3503 ( .A(_abc_17692_n10495), .B(_abc_17692_n10481), .Y(_abc_17692_n10496) );
  OR2X2 OR2X2_3504 ( .A(_abc_17692_n10496), .B(_abc_17692_n10494), .Y(_abc_17692_n10497) );
  OR2X2 OR2X2_3505 ( .A(_abc_17692_n10492), .B(_abc_17692_n10499), .Y(_abc_17692_n10500) );
  OR2X2 OR2X2_3506 ( .A(_abc_17692_n10501), .B(_abc_17692_n4964), .Y(_abc_17692_n10502) );
  OR2X2 OR2X2_3507 ( .A(_abc_17692_n4965), .B(_abc_17692_n10500), .Y(_abc_17692_n10503) );
  OR2X2 OR2X2_3508 ( .A(_abc_17692_n10504), .B(workunit1_16_bF_buf0), .Y(_abc_17692_n10507) );
  OR2X2 OR2X2_3509 ( .A(_abc_17692_n10512), .B(_abc_17692_n10511), .Y(_abc_17692_n10513) );
  OR2X2 OR2X2_351 ( .A(_abc_17692_n1515), .B(_abc_17692_n1541), .Y(_abc_17692_n1542) );
  OR2X2 OR2X2_3510 ( .A(_abc_17692_n10510), .B(_abc_17692_n10513), .Y(_abc_17692_n10514) );
  OR2X2 OR2X2_3511 ( .A(_abc_17692_n10516), .B(_abc_17692_n10514), .Y(_abc_17692_n10517) );
  OR2X2 OR2X2_3512 ( .A(_abc_17692_n10517), .B(_abc_17692_n10508), .Y(_abc_17692_n10520) );
  OR2X2 OR2X2_3513 ( .A(_abc_17692_n10501), .B(_abc_17692_n5010), .Y(_abc_17692_n10523) );
  OR2X2 OR2X2_3514 ( .A(_abc_17692_n5011), .B(_abc_17692_n10500), .Y(_abc_17692_n10524) );
  OR2X2 OR2X2_3515 ( .A(_abc_17692_n10525), .B(workunit1_16_bF_buf2), .Y(_abc_17692_n10528) );
  OR2X2 OR2X2_3516 ( .A(_abc_17692_n10403), .B(_abc_17692_n10251), .Y(_abc_17692_n10530) );
  OR2X2 OR2X2_3517 ( .A(_abc_17692_n10530), .B(_abc_17692_n10299), .Y(_abc_17692_n10531) );
  OR2X2 OR2X2_3518 ( .A(_abc_17692_n10403), .B(_abc_17692_n10448), .Y(_abc_17692_n10534) );
  OR2X2 OR2X2_3519 ( .A(_abc_17692_n10530), .B(_abc_17692_n10301), .Y(_abc_17692_n10537) );
  OR2X2 OR2X2_352 ( .A(_abc_17692_n1545), .B(_abc_17692_n1528), .Y(_abc_17692_n1548) );
  OR2X2 OR2X2_3520 ( .A(_abc_17692_n10537), .B(_abc_17692_n9917), .Y(_abc_17692_n10538) );
  OR2X2 OR2X2_3521 ( .A(_abc_17692_n10540), .B(_abc_17692_n10529), .Y(_abc_17692_n10541) );
  OR2X2 OR2X2_3522 ( .A(_abc_17692_n10501), .B(_abc_17692_n5056), .Y(_abc_17692_n10546) );
  OR2X2 OR2X2_3523 ( .A(_abc_17692_n5057), .B(_abc_17692_n10500), .Y(_abc_17692_n10547) );
  OR2X2 OR2X2_3524 ( .A(_abc_17692_n10548), .B(workunit1_16_bF_buf0), .Y(_abc_17692_n10551) );
  OR2X2 OR2X2_3525 ( .A(_abc_17692_n10555), .B(_abc_17692_n10556), .Y(_abc_17692_n10557) );
  OR2X2 OR2X2_3526 ( .A(_abc_17692_n10557), .B(_abc_17692_n10554), .Y(_abc_17692_n10558) );
  OR2X2 OR2X2_3527 ( .A(_abc_17692_n10560), .B(_abc_17692_n10558), .Y(_abc_17692_n10561) );
  OR2X2 OR2X2_3528 ( .A(_abc_17692_n10561), .B(_abc_17692_n10552), .Y(_abc_17692_n10562) );
  OR2X2 OR2X2_3529 ( .A(_abc_17692_n10566), .B(_abc_17692_n10545), .Y(_abc_17692_n10567) );
  OR2X2 OR2X2_353 ( .A(_abc_17692_n1551), .B(state_8_bF_buf5), .Y(_abc_17692_n1552) );
  OR2X2 OR2X2_3530 ( .A(_abc_17692_n10567), .B(_abc_17692_n10522), .Y(_abc_17692_n10568) );
  OR2X2 OR2X2_3531 ( .A(_abc_17692_n5103), .B(_abc_17692_n10501), .Y(_abc_17692_n10569) );
  OR2X2 OR2X2_3532 ( .A(_abc_17692_n5104), .B(_abc_17692_n10500), .Y(_abc_17692_n10570) );
  OR2X2 OR2X2_3533 ( .A(_abc_17692_n10571), .B(workunit1_16_bF_buf2), .Y(_abc_17692_n10574) );
  OR2X2 OR2X2_3534 ( .A(_abc_17692_n10578), .B(_abc_17692_n10579), .Y(_abc_17692_n10580) );
  OR2X2 OR2X2_3535 ( .A(_abc_17692_n10580), .B(_abc_17692_n10577), .Y(_abc_17692_n10581) );
  OR2X2 OR2X2_3536 ( .A(_abc_17692_n10583), .B(_abc_17692_n10581), .Y(_abc_17692_n10584) );
  OR2X2 OR2X2_3537 ( .A(_abc_17692_n10584), .B(_abc_17692_n10575), .Y(_abc_17692_n10585) );
  OR2X2 OR2X2_3538 ( .A(_abc_17692_n10589), .B(_abc_17692_n10568), .Y(_abc_17692_n10590) );
  OR2X2 OR2X2_3539 ( .A(_abc_17692_n10596), .B(_abc_17692_n10595), .Y(_abc_17692_n10597) );
  OR2X2 OR2X2_354 ( .A(_abc_17692_n1550_1), .B(_abc_17692_n1552), .Y(_abc_17692_n1553) );
  OR2X2 OR2X2_3540 ( .A(_abc_17692_n10594), .B(_abc_17692_n10598), .Y(_abc_17692_n10599) );
  OR2X2 OR2X2_3541 ( .A(_abc_17692_n10601), .B(_abc_17692_n10599), .Y(_abc_17692_n10602) );
  OR2X2 OR2X2_3542 ( .A(_abc_17692_n10602), .B(_abc_17692_n10592), .Y(_abc_17692_n10603) );
  OR2X2 OR2X2_3543 ( .A(_abc_17692_n10368), .B(_abc_17692_n10232), .Y(_abc_17692_n10610) );
  OR2X2 OR2X2_3544 ( .A(_abc_17692_n10610), .B(_abc_17692_n10609), .Y(_abc_17692_n10611) );
  OR2X2 OR2X2_3545 ( .A(_abc_17692_n10368), .B(_abc_17692_n10372), .Y(_abc_17692_n10614) );
  OR2X2 OR2X2_3546 ( .A(_abc_17692_n10610), .B(_abc_17692_n10618), .Y(_abc_17692_n10619) );
  OR2X2 OR2X2_3547 ( .A(_abc_17692_n10621), .B(_abc_17692_n10617), .Y(_abc_17692_n10622) );
  OR2X2 OR2X2_3548 ( .A(_abc_17692_n10622), .B(_abc_17692_n10608), .Y(_abc_17692_n10625) );
  OR2X2 OR2X2_3549 ( .A(_abc_17692_n10418), .B(_abc_17692_n10267), .Y(_abc_17692_n10631) );
  OR2X2 OR2X2_355 ( .A(_abc_17692_n1540), .B(_abc_17692_n1553), .Y(sum_22__FF_INPUT) );
  OR2X2 OR2X2_3550 ( .A(_abc_17692_n10630), .B(_abc_17692_n10633), .Y(_abc_17692_n10634) );
  OR2X2 OR2X2_3551 ( .A(_abc_17692_n10634), .B(_abc_17692_n10636), .Y(_abc_17692_n10637) );
  OR2X2 OR2X2_3552 ( .A(_abc_17692_n10637), .B(_abc_17692_n10628), .Y(_abc_17692_n10640) );
  OR2X2 OR2X2_3553 ( .A(_abc_17692_n10650), .B(_abc_17692_n10645), .Y(_abc_17692_n10651) );
  OR2X2 OR2X2_3554 ( .A(_abc_17692_n10653), .B(_abc_17692_n10651), .Y(_abc_17692_n10654) );
  OR2X2 OR2X2_3555 ( .A(_abc_17692_n10654), .B(_abc_17692_n10643), .Y(_abc_17692_n10655) );
  OR2X2 OR2X2_3556 ( .A(_abc_17692_n10659), .B(_abc_17692_n10642), .Y(_abc_17692_n10660) );
  OR2X2 OR2X2_3557 ( .A(_abc_17692_n10660), .B(_abc_17692_n10627), .Y(_abc_17692_n10661) );
  OR2X2 OR2X2_3558 ( .A(_abc_17692_n10661), .B(_abc_17692_n10607), .Y(_abc_17692_n10662) );
  OR2X2 OR2X2_3559 ( .A(_abc_17692_n10664), .B(_abc_17692_n10665), .Y(_abc_17692_n10666) );
  OR2X2 OR2X2_356 ( .A(_abc_17692_n1537), .B(_abc_17692_n1524), .Y(_abc_17692_n1563) );
  OR2X2 OR2X2_3560 ( .A(_abc_17692_n10663), .B(_abc_17692_n10666), .Y(_abc_17692_n10667) );
  OR2X2 OR2X2_3561 ( .A(_abc_17692_n10591), .B(_abc_17692_n10667), .Y(workunit1_16__FF_INPUT) );
  OR2X2 OR2X2_3562 ( .A(_abc_17692_n10499), .B(_abc_17692_n10489), .Y(_abc_17692_n10669) );
  OR2X2 OR2X2_3563 ( .A(_abc_17692_n4351), .B(workunit2_22_), .Y(_abc_17692_n10670) );
  OR2X2 OR2X2_3564 ( .A(_abc_17692_n6293), .B(workunit2_13_), .Y(_abc_17692_n10671) );
  OR2X2 OR2X2_3565 ( .A(_abc_17692_n10669), .B(_abc_17692_n10679), .Y(_abc_17692_n10680) );
  OR2X2 OR2X2_3566 ( .A(_abc_17692_n5312), .B(_abc_17692_n10683), .Y(_abc_17692_n10684) );
  OR2X2 OR2X2_3567 ( .A(_abc_17692_n5314), .B(_abc_17692_n10685), .Y(_abc_17692_n10686) );
  OR2X2 OR2X2_3568 ( .A(_abc_17692_n10698), .B(_abc_17692_n4047_bF_buf0), .Y(_abc_17692_n10699) );
  OR2X2 OR2X2_3569 ( .A(_abc_17692_n10699), .B(_abc_17692_n10696), .Y(_abc_17692_n10700) );
  OR2X2 OR2X2_357 ( .A(_abc_17692_n1564), .B(_abc_17692_n1562_1), .Y(_abc_17692_n1565) );
  OR2X2 OR2X2_3570 ( .A(_abc_17692_n5253), .B(_abc_17692_n10683), .Y(_abc_17692_n10701) );
  OR2X2 OR2X2_3571 ( .A(_abc_17692_n5255), .B(_abc_17692_n10685), .Y(_abc_17692_n10702) );
  OR2X2 OR2X2_3572 ( .A(_abc_17692_n10710), .B(_abc_17692_n10709), .Y(_abc_17692_n10711) );
  OR2X2 OR2X2_3573 ( .A(_abc_17692_n10713), .B(_abc_17692_n10712), .Y(_abc_17692_n10714) );
  OR2X2 OR2X2_3574 ( .A(_abc_17692_n5231), .B(_abc_17692_n10683), .Y(_abc_17692_n10717) );
  OR2X2 OR2X2_3575 ( .A(_abc_17692_n10685), .B(_abc_17692_n5228), .Y(_abc_17692_n10718) );
  OR2X2 OR2X2_3576 ( .A(_abc_17692_n10721), .B(_abc_17692_n10722), .Y(_abc_17692_n10723) );
  OR2X2 OR2X2_3577 ( .A(_abc_17692_n10725), .B(_abc_17692_n10723), .Y(_abc_17692_n10726) );
  OR2X2 OR2X2_3578 ( .A(_abc_17692_n10724), .B(_abc_17692_n10727), .Y(_abc_17692_n10728) );
  OR2X2 OR2X2_3579 ( .A(_abc_17692_n10731), .B(_abc_17692_n10732), .Y(_abc_17692_n10733) );
  OR2X2 OR2X2_358 ( .A(_abc_17692_n1563), .B(_abc_17692_n1561), .Y(_abc_17692_n1566) );
  OR2X2 OR2X2_3580 ( .A(_abc_17692_n10733), .B(_abc_17692_n4059), .Y(_abc_17692_n10734) );
  OR2X2 OR2X2_3581 ( .A(_abc_17692_n10735), .B(workunit1_17_), .Y(_abc_17692_n10736) );
  OR2X2 OR2X2_3582 ( .A(_abc_17692_n10738), .B(_abc_17692_n10737), .Y(_abc_17692_n10739) );
  OR2X2 OR2X2_3583 ( .A(_abc_17692_n10741), .B(_abc_17692_n10740), .Y(_abc_17692_n10742) );
  OR2X2 OR2X2_3584 ( .A(_abc_17692_n10744), .B(_abc_17692_n1863_bF_buf3), .Y(_abc_17692_n10745) );
  OR2X2 OR2X2_3585 ( .A(_abc_17692_n10745), .B(_abc_17692_n10730), .Y(_abc_17692_n10746) );
  OR2X2 OR2X2_3586 ( .A(_abc_17692_n10746), .B(_abc_17692_n10716), .Y(_abc_17692_n10747) );
  OR2X2 OR2X2_3587 ( .A(_abc_17692_n10755), .B(_abc_17692_n10756), .Y(_abc_17692_n10757) );
  OR2X2 OR2X2_3588 ( .A(_abc_17692_n10762), .B(_abc_17692_n10712), .Y(_abc_17692_n10763) );
  OR2X2 OR2X2_3589 ( .A(_abc_17692_n10764), .B(_abc_17692_n10709), .Y(_abc_17692_n10765) );
  OR2X2 OR2X2_359 ( .A(_abc_17692_n1571), .B(_abc_17692_n1561), .Y(_abc_17692_n1572) );
  OR2X2 OR2X2_3590 ( .A(_abc_17692_n10772), .B(_abc_17692_n10737), .Y(_abc_17692_n10773) );
  OR2X2 OR2X2_3591 ( .A(_abc_17692_n10771), .B(_abc_17692_n10740), .Y(_abc_17692_n10774) );
  OR2X2 OR2X2_3592 ( .A(_abc_17692_n10780), .B(_abc_17692_n10723), .Y(_abc_17692_n10781) );
  OR2X2 OR2X2_3593 ( .A(_abc_17692_n10782), .B(_abc_17692_n10727), .Y(_abc_17692_n10783) );
  OR2X2 OR2X2_3594 ( .A(_abc_17692_n10785), .B(_abc_17692_n10776), .Y(_abc_17692_n10786) );
  OR2X2 OR2X2_3595 ( .A(_abc_17692_n10786), .B(_abc_17692_n10767), .Y(_abc_17692_n10787) );
  OR2X2 OR2X2_3596 ( .A(_abc_17692_n10787), .B(_abc_17692_n10758), .Y(_abc_17692_n10788) );
  OR2X2 OR2X2_3597 ( .A(_abc_17692_n10790), .B(_abc_17692_n10791), .Y(_abc_17692_n10792) );
  OR2X2 OR2X2_3598 ( .A(_abc_17692_n10789), .B(_abc_17692_n10792), .Y(_abc_17692_n10793) );
  OR2X2 OR2X2_3599 ( .A(_abc_17692_n10793), .B(_abc_17692_n10749), .Y(workunit1_17__FF_INPUT) );
  OR2X2 OR2X2_36 ( .A(state_5_), .B(state_1_), .Y(_abc_17692_n709) );
  OR2X2 OR2X2_360 ( .A(_abc_17692_n1573), .B(_abc_17692_n1562_1), .Y(_abc_17692_n1574) );
  OR2X2 OR2X2_3600 ( .A(_abc_17692_n10795), .B(_abc_17692_n10674), .Y(_abc_17692_n10796) );
  OR2X2 OR2X2_3601 ( .A(_abc_17692_n10798), .B(_abc_17692_n10796), .Y(_abc_17692_n10799) );
  OR2X2 OR2X2_3602 ( .A(_abc_17692_n4623), .B(workunit2_23_), .Y(_abc_17692_n10800) );
  OR2X2 OR2X2_3603 ( .A(_abc_17692_n6505), .B(workunit2_14_bF_buf1), .Y(_abc_17692_n10801) );
  OR2X2 OR2X2_3604 ( .A(_abc_17692_n10804), .B(_abc_17692_n10805), .Y(_abc_17692_n10806) );
  OR2X2 OR2X2_3605 ( .A(_abc_17692_n10810), .B(_abc_17692_n10808), .Y(_abc_17692_n10811) );
  OR2X2 OR2X2_3606 ( .A(_abc_17692_n5521), .B(_abc_17692_n10812), .Y(_abc_17692_n10813) );
  OR2X2 OR2X2_3607 ( .A(_abc_17692_n5522), .B(_abc_17692_n10811), .Y(_abc_17692_n10814) );
  OR2X2 OR2X2_3608 ( .A(_abc_17692_n10817), .B(_abc_17692_n10818), .Y(_abc_17692_n10819) );
  OR2X2 OR2X2_3609 ( .A(_abc_17692_n10688), .B(_abc_17692_n10751), .Y(_abc_17692_n10820) );
  OR2X2 OR2X2_361 ( .A(_abc_17692_n1577), .B(state_8_bF_buf4), .Y(_abc_17692_n1578) );
  OR2X2 OR2X2_3610 ( .A(_abc_17692_n10823), .B(_abc_17692_n10821), .Y(_abc_17692_n10824) );
  OR2X2 OR2X2_3611 ( .A(_abc_17692_n10824), .B(_abc_17692_n10819), .Y(_abc_17692_n10825) );
  OR2X2 OR2X2_3612 ( .A(_abc_17692_n5410), .B(_abc_17692_n10812), .Y(_abc_17692_n10830) );
  OR2X2 OR2X2_3613 ( .A(_abc_17692_n5413), .B(_abc_17692_n10811), .Y(_abc_17692_n10831) );
  OR2X2 OR2X2_3614 ( .A(_abc_17692_n10832), .B(workunit1_18_), .Y(_abc_17692_n10835) );
  OR2X2 OR2X2_3615 ( .A(_abc_17692_n10704), .B(_abc_17692_n10760), .Y(_abc_17692_n10838) );
  OR2X2 OR2X2_3616 ( .A(_abc_17692_n10841), .B(_abc_17692_n10839), .Y(_abc_17692_n10842) );
  OR2X2 OR2X2_3617 ( .A(_abc_17692_n10842), .B(_abc_17692_n10837), .Y(_abc_17692_n10845) );
  OR2X2 OR2X2_3618 ( .A(_abc_17692_n10812), .B(_abc_17692_n5482), .Y(_abc_17692_n10848) );
  OR2X2 OR2X2_3619 ( .A(_abc_17692_n5483), .B(_abc_17692_n10811), .Y(_abc_17692_n10849) );
  OR2X2 OR2X2_362 ( .A(_abc_17692_n1576), .B(_abc_17692_n1578), .Y(_abc_17692_n1579) );
  OR2X2 OR2X2_3620 ( .A(_abc_17692_n10850), .B(_abc_17692_n4322), .Y(_abc_17692_n10851) );
  OR2X2 OR2X2_3621 ( .A(_abc_17692_n10852), .B(workunit1_18_), .Y(_abc_17692_n10853) );
  OR2X2 OR2X2_3622 ( .A(_abc_17692_n10721), .B(_abc_17692_n10778), .Y(_abc_17692_n10856) );
  OR2X2 OR2X2_3623 ( .A(_abc_17692_n10859), .B(_abc_17692_n10857), .Y(_abc_17692_n10860) );
  OR2X2 OR2X2_3624 ( .A(_abc_17692_n10860), .B(_abc_17692_n10854), .Y(_abc_17692_n10863) );
  OR2X2 OR2X2_3625 ( .A(_abc_17692_n10812), .B(_abc_17692_n5444), .Y(_abc_17692_n10866) );
  OR2X2 OR2X2_3626 ( .A(_abc_17692_n5446), .B(_abc_17692_n10811), .Y(_abc_17692_n10867) );
  OR2X2 OR2X2_3627 ( .A(_abc_17692_n10868), .B(workunit1_18_), .Y(_abc_17692_n10869) );
  OR2X2 OR2X2_3628 ( .A(_abc_17692_n10874), .B(_abc_17692_n10875), .Y(_abc_17692_n10876) );
  OR2X2 OR2X2_3629 ( .A(_abc_17692_n10020), .B(_abc_17692_n10878), .Y(_abc_17692_n10879) );
  OR2X2 OR2X2_363 ( .A(_abc_17692_n1568), .B(_abc_17692_n1579), .Y(sum_23__FF_INPUT) );
  OR2X2 OR2X2_3630 ( .A(_abc_17692_n10880), .B(_abc_17692_n10882), .Y(_abc_17692_n10883) );
  OR2X2 OR2X2_3631 ( .A(_abc_17692_n10885), .B(_abc_17692_n10873), .Y(_abc_17692_n10888) );
  OR2X2 OR2X2_3632 ( .A(_abc_17692_n10890), .B(_abc_17692_n10865), .Y(_abc_17692_n10891) );
  OR2X2 OR2X2_3633 ( .A(_abc_17692_n10891), .B(_abc_17692_n10847), .Y(_abc_17692_n10892) );
  OR2X2 OR2X2_3634 ( .A(_abc_17692_n10892), .B(_abc_17692_n10829), .Y(_abc_17692_n10893) );
  OR2X2 OR2X2_3635 ( .A(_abc_17692_n10693), .B(_abc_17692_n10573), .Y(_abc_17692_n10898) );
  OR2X2 OR2X2_3636 ( .A(_abc_17692_n10902), .B(_abc_17692_n10900), .Y(_abc_17692_n10903) );
  OR2X2 OR2X2_3637 ( .A(_abc_17692_n10903), .B(_abc_17692_n10895), .Y(_abc_17692_n10904) );
  OR2X2 OR2X2_3638 ( .A(_abc_17692_n10907), .B(_abc_17692_n4047_bF_buf4), .Y(_abc_17692_n10908) );
  OR2X2 OR2X2_3639 ( .A(_abc_17692_n10910), .B(_abc_17692_n10909), .Y(_abc_17692_n10911) );
  OR2X2 OR2X2_364 ( .A(_abc_17692_n1581), .B(delta_24_), .Y(_abc_17692_n1583) );
  OR2X2 OR2X2_3640 ( .A(_abc_17692_n10913), .B(_abc_17692_n10911), .Y(_abc_17692_n10914) );
  OR2X2 OR2X2_3641 ( .A(_abc_17692_n10914), .B(_abc_17692_n10836), .Y(_abc_17692_n10915) );
  OR2X2 OR2X2_3642 ( .A(_abc_17692_n10922), .B(_abc_17692_n10921), .Y(_abc_17692_n10923) );
  OR2X2 OR2X2_3643 ( .A(_abc_17692_n10925), .B(_abc_17692_n10923), .Y(_abc_17692_n10926) );
  OR2X2 OR2X2_3644 ( .A(_abc_17692_n10926), .B(_abc_17692_n10920), .Y(_abc_17692_n10929) );
  OR2X2 OR2X2_3645 ( .A(_abc_17692_n10737), .B(_abc_17692_n10527), .Y(_abc_17692_n10934) );
  OR2X2 OR2X2_3646 ( .A(_abc_17692_n10938), .B(_abc_17692_n10936), .Y(_abc_17692_n10939) );
  OR2X2 OR2X2_3647 ( .A(_abc_17692_n10939), .B(_abc_17692_n10872), .Y(_abc_17692_n10940) );
  OR2X2 OR2X2_3648 ( .A(_abc_17692_n10944), .B(_abc_17692_n1863_bF_buf0), .Y(_abc_17692_n10945) );
  OR2X2 OR2X2_3649 ( .A(_abc_17692_n10945), .B(_abc_17692_n10931), .Y(_abc_17692_n10946) );
  OR2X2 OR2X2_365 ( .A(_abc_17692_n1584), .B(_abc_17692_n1582), .Y(_abc_17692_n1585) );
  OR2X2 OR2X2_3650 ( .A(_abc_17692_n10946), .B(_abc_17692_n10919), .Y(_abc_17692_n10947) );
  OR2X2 OR2X2_3651 ( .A(_abc_17692_n10950), .B(_abc_17692_n10951), .Y(_abc_17692_n10952) );
  OR2X2 OR2X2_3652 ( .A(_abc_17692_n10949), .B(_abc_17692_n10952), .Y(_abc_17692_n10953) );
  OR2X2 OR2X2_3653 ( .A(_abc_17692_n10953), .B(_abc_17692_n10894), .Y(workunit1_18__FF_INPUT) );
  OR2X2 OR2X2_3654 ( .A(_abc_17692_n10808), .B(_abc_17692_n10804), .Y(_abc_17692_n10955) );
  OR2X2 OR2X2_3655 ( .A(_abc_17692_n4765), .B(workunit2_24_), .Y(_abc_17692_n10957) );
  OR2X2 OR2X2_3656 ( .A(_abc_17692_n6657_1), .B(workunit2_15_), .Y(_abc_17692_n10958) );
  OR2X2 OR2X2_3657 ( .A(_abc_17692_n10971), .B(_abc_17692_n5708), .Y(_abc_17692_n10972) );
  OR2X2 OR2X2_3658 ( .A(_abc_17692_n10967), .B(_abc_17692_n10969), .Y(_abc_17692_n10973) );
  OR2X2 OR2X2_3659 ( .A(_abc_17692_n5711), .B(_abc_17692_n10973), .Y(_abc_17692_n10974) );
  OR2X2 OR2X2_366 ( .A(_abc_17692_n1467), .B(_abc_17692_n1588), .Y(_abc_17692_n1589) );
  OR2X2 OR2X2_3660 ( .A(_abc_17692_n5708), .B(_abc_17692_n10973), .Y(_abc_17692_n10977) );
  OR2X2 OR2X2_3661 ( .A(_abc_17692_n10971), .B(_abc_17692_n5711), .Y(_abc_17692_n10978) );
  OR2X2 OR2X2_3662 ( .A(_abc_17692_n10976), .B(_abc_17692_n10980), .Y(_abc_17692_n10981) );
  OR2X2 OR2X2_3663 ( .A(_abc_17692_n10984), .B(_abc_17692_n10981), .Y(_abc_17692_n10985) );
  OR2X2 OR2X2_3664 ( .A(_abc_17692_n10987), .B(_abc_17692_n10986), .Y(_abc_17692_n10988) );
  OR2X2 OR2X2_3665 ( .A(_abc_17692_n5622), .B(_abc_17692_n10971), .Y(_abc_17692_n10991) );
  OR2X2 OR2X2_3666 ( .A(_abc_17692_n5620), .B(_abc_17692_n10973), .Y(_abc_17692_n10992) );
  OR2X2 OR2X2_3667 ( .A(_abc_17692_n10994), .B(workunit1_19_), .Y(_abc_17692_n10995) );
  OR2X2 OR2X2_3668 ( .A(_abc_17692_n10993), .B(_abc_17692_n4494), .Y(_abc_17692_n10996) );
  OR2X2 OR2X2_3669 ( .A(_abc_17692_n10999), .B(_abc_17692_n10997), .Y(_abc_17692_n11000) );
  OR2X2 OR2X2_367 ( .A(_abc_17692_n1591), .B(_abc_17692_n1555), .Y(_abc_17692_n1592) );
  OR2X2 OR2X2_3670 ( .A(_abc_17692_n10998), .B(_abc_17692_n11001), .Y(_abc_17692_n11002) );
  OR2X2 OR2X2_3671 ( .A(_abc_17692_n5680), .B(_abc_17692_n10973), .Y(_abc_17692_n11005) );
  OR2X2 OR2X2_3672 ( .A(_abc_17692_n10971), .B(_abc_17692_n5683), .Y(_abc_17692_n11006) );
  OR2X2 OR2X2_3673 ( .A(_abc_17692_n11007), .B(workunit1_19_), .Y(_abc_17692_n11008) );
  OR2X2 OR2X2_3674 ( .A(_abc_17692_n10971), .B(_abc_17692_n5680), .Y(_abc_17692_n11009) );
  OR2X2 OR2X2_3675 ( .A(_abc_17692_n5683), .B(_abc_17692_n10973), .Y(_abc_17692_n11010) );
  OR2X2 OR2X2_3676 ( .A(_abc_17692_n11011), .B(_abc_17692_n4494), .Y(_abc_17692_n11012) );
  OR2X2 OR2X2_3677 ( .A(_abc_17692_n11015), .B(_abc_17692_n11013), .Y(_abc_17692_n11016) );
  OR2X2 OR2X2_3678 ( .A(_abc_17692_n11017), .B(_abc_17692_n11018), .Y(_abc_17692_n11019) );
  OR2X2 OR2X2_3679 ( .A(_abc_17692_n11014), .B(_abc_17692_n11019), .Y(_abc_17692_n11020) );
  OR2X2 OR2X2_368 ( .A(_abc_17692_n1590), .B(_abc_17692_n1592), .Y(_abc_17692_n1593) );
  OR2X2 OR2X2_3680 ( .A(_abc_17692_n11004), .B(_abc_17692_n11022), .Y(_abc_17692_n11023) );
  OR2X2 OR2X2_3681 ( .A(_abc_17692_n11023), .B(_abc_17692_n10990), .Y(_abc_17692_n11024) );
  OR2X2 OR2X2_3682 ( .A(_abc_17692_n5651), .B(_abc_17692_n10971), .Y(_abc_17692_n11025) );
  OR2X2 OR2X2_3683 ( .A(_abc_17692_n5648), .B(_abc_17692_n10973), .Y(_abc_17692_n11026) );
  OR2X2 OR2X2_3684 ( .A(_abc_17692_n5651), .B(_abc_17692_n10973), .Y(_abc_17692_n11029) );
  OR2X2 OR2X2_3685 ( .A(_abc_17692_n5648), .B(_abc_17692_n10971), .Y(_abc_17692_n11030) );
  OR2X2 OR2X2_3686 ( .A(_abc_17692_n11028), .B(_abc_17692_n11032), .Y(_abc_17692_n11033) );
  OR2X2 OR2X2_3687 ( .A(_abc_17692_n11031), .B(workunit1_19_), .Y(_abc_17692_n11038) );
  OR2X2 OR2X2_3688 ( .A(_abc_17692_n11027), .B(_abc_17692_n4494), .Y(_abc_17692_n11039) );
  OR2X2 OR2X2_3689 ( .A(_abc_17692_n11037), .B(_abc_17692_n11041), .Y(_abc_17692_n11042) );
  OR2X2 OR2X2_369 ( .A(_abc_17692_n1468), .B(_abc_17692_n1588), .Y(_abc_17692_n1596) );
  OR2X2 OR2X2_3690 ( .A(_abc_17692_n11043), .B(_abc_17692_n11024), .Y(_abc_17692_n11044) );
  OR2X2 OR2X2_3691 ( .A(_abc_17692_n10826), .B(_abc_17692_n11046), .Y(_abc_17692_n11047) );
  OR2X2 OR2X2_3692 ( .A(_abc_17692_n11048), .B(_abc_17692_n11040), .Y(_abc_17692_n11049) );
  OR2X2 OR2X2_3693 ( .A(_abc_17692_n11047), .B(_abc_17692_n11033), .Y(_abc_17692_n11050) );
  OR2X2 OR2X2_3694 ( .A(_abc_17692_n11056), .B(_abc_17692_n10997), .Y(_abc_17692_n11057) );
  OR2X2 OR2X2_3695 ( .A(_abc_17692_n11058), .B(_abc_17692_n11001), .Y(_abc_17692_n11059) );
  OR2X2 OR2X2_3696 ( .A(_abc_17692_n10868), .B(_abc_17692_n4322), .Y(_abc_17692_n11062) );
  OR2X2 OR2X2_3697 ( .A(_abc_17692_n10886), .B(_abc_17692_n11063), .Y(_abc_17692_n11064) );
  OR2X2 OR2X2_3698 ( .A(_abc_17692_n11065), .B(_abc_17692_n11013), .Y(_abc_17692_n11066) );
  OR2X2 OR2X2_3699 ( .A(_abc_17692_n11064), .B(_abc_17692_n11019), .Y(_abc_17692_n11067) );
  OR2X2 OR2X2_37 ( .A(_abc_17692_n708), .B(_abc_17692_n709), .Y(_abc_17692_n710) );
  OR2X2 OR2X2_370 ( .A(_abc_17692_n1598_1), .B(_abc_17692_n1585), .Y(_abc_17692_n1599) );
  OR2X2 OR2X2_3700 ( .A(_abc_17692_n11071), .B(_abc_17692_n10981), .Y(_abc_17692_n11072) );
  OR2X2 OR2X2_3701 ( .A(_abc_17692_n11070), .B(_abc_17692_n10986), .Y(_abc_17692_n11073) );
  OR2X2 OR2X2_3702 ( .A(_abc_17692_n11075), .B(_abc_17692_n11069), .Y(_abc_17692_n11076) );
  OR2X2 OR2X2_3703 ( .A(_abc_17692_n11061), .B(_abc_17692_n11076), .Y(_abc_17692_n11077) );
  OR2X2 OR2X2_3704 ( .A(_abc_17692_n11077), .B(_abc_17692_n11052), .Y(_abc_17692_n11078) );
  OR2X2 OR2X2_3705 ( .A(_abc_17692_n11080), .B(_abc_17692_n11081), .Y(_abc_17692_n11082) );
  OR2X2 OR2X2_3706 ( .A(_abc_17692_n11079), .B(_abc_17692_n11082), .Y(_abc_17692_n11083) );
  OR2X2 OR2X2_3707 ( .A(_abc_17692_n11045), .B(_abc_17692_n11083), .Y(workunit1_19__FF_INPUT) );
  OR2X2 OR2X2_3708 ( .A(_abc_17692_n10484), .B(_abc_17692_n11087), .Y(_abc_17692_n11088) );
  OR2X2 OR2X2_3709 ( .A(_abc_17692_n11092), .B(_abc_17692_n10963), .Y(_abc_17692_n11093) );
  OR2X2 OR2X2_371 ( .A(_abc_17692_n1608), .B(_abc_17692_n1609), .Y(_abc_17692_n1610) );
  OR2X2 OR2X2_3710 ( .A(_abc_17692_n9717), .B(workunit2_25_), .Y(_abc_17692_n11096) );
  OR2X2 OR2X2_3711 ( .A(_abc_17692_n6952), .B(workunit2_16_bF_buf1), .Y(_abc_17692_n11097) );
  OR2X2 OR2X2_3712 ( .A(_abc_17692_n11100), .B(_abc_17692_n11101), .Y(_abc_17692_n11102) );
  OR2X2 OR2X2_3713 ( .A(_abc_17692_n11104), .B(_abc_17692_n11105), .Y(_abc_17692_n11106) );
  OR2X2 OR2X2_3714 ( .A(_abc_17692_n11103), .B(_abc_17692_n11108), .Y(_abc_17692_n11109) );
  OR2X2 OR2X2_3715 ( .A(_abc_17692_n5814), .B(_abc_17692_n11110), .Y(_abc_17692_n11111) );
  OR2X2 OR2X2_3716 ( .A(_abc_17692_n5815), .B(_abc_17692_n11109), .Y(_abc_17692_n11112) );
  OR2X2 OR2X2_3717 ( .A(_abc_17692_n11115), .B(_abc_17692_n11116), .Y(_abc_17692_n11117) );
  OR2X2 OR2X2_3718 ( .A(_abc_17692_n11122), .B(_abc_17692_n10899), .Y(_abc_17692_n11123) );
  OR2X2 OR2X2_3719 ( .A(_abc_17692_n11124), .B(_abc_17692_n11032), .Y(_abc_17692_n11125) );
  OR2X2 OR2X2_372 ( .A(_abc_17692_n1607), .B(_abc_17692_n1610), .Y(_abc_17692_n1611) );
  OR2X2 OR2X2_3720 ( .A(_abc_17692_n11121), .B(_abc_17692_n11128), .Y(_abc_17692_n11129) );
  OR2X2 OR2X2_3721 ( .A(_abc_17692_n11129), .B(_abc_17692_n11118), .Y(_abc_17692_n11132) );
  OR2X2 OR2X2_3722 ( .A(_abc_17692_n11133), .B(_abc_17692_n4047_bF_buf3), .Y(_abc_17692_n11134) );
  OR2X2 OR2X2_3723 ( .A(_abc_17692_n11110), .B(_abc_17692_n5859), .Y(_abc_17692_n11135) );
  OR2X2 OR2X2_3724 ( .A(_abc_17692_n5860), .B(_abc_17692_n11109), .Y(_abc_17692_n11136) );
  OR2X2 OR2X2_3725 ( .A(_abc_17692_n11137), .B(workunit1_20_), .Y(_abc_17692_n11140) );
  OR2X2 OR2X2_3726 ( .A(_abc_17692_n11144), .B(_abc_17692_n10834), .Y(_abc_17692_n11145) );
  OR2X2 OR2X2_3727 ( .A(_abc_17692_n11147), .B(_abc_17692_n11143), .Y(_abc_17692_n11148) );
  OR2X2 OR2X2_3728 ( .A(_abc_17692_n11150), .B(_abc_17692_n11148), .Y(_abc_17692_n11151) );
  OR2X2 OR2X2_3729 ( .A(_abc_17692_n11151), .B(_abc_17692_n11141), .Y(_abc_17692_n11152) );
  OR2X2 OR2X2_373 ( .A(_abc_17692_n1613_1), .B(_abc_17692_n1611), .Y(_abc_17692_n1614) );
  OR2X2 OR2X2_3730 ( .A(_abc_17692_n11110), .B(_abc_17692_n5905), .Y(_abc_17692_n11157) );
  OR2X2 OR2X2_3731 ( .A(_abc_17692_n5906), .B(_abc_17692_n11109), .Y(_abc_17692_n11158) );
  OR2X2 OR2X2_3732 ( .A(_abc_17692_n11161), .B(_abc_17692_n11162), .Y(_abc_17692_n11163) );
  OR2X2 OR2X2_3733 ( .A(_abc_17692_n11167), .B(_abc_17692_n10980), .Y(_abc_17692_n11168) );
  OR2X2 OR2X2_3734 ( .A(_abc_17692_n11168), .B(_abc_17692_n11166), .Y(_abc_17692_n11169) );
  OR2X2 OR2X2_3735 ( .A(_abc_17692_n11171), .B(_abc_17692_n11169), .Y(_abc_17692_n11172) );
  OR2X2 OR2X2_3736 ( .A(_abc_17692_n11172), .B(_abc_17692_n11164), .Y(_abc_17692_n11175) );
  OR2X2 OR2X2_3737 ( .A(_abc_17692_n11110), .B(_abc_17692_n5952), .Y(_abc_17692_n11178) );
  OR2X2 OR2X2_3738 ( .A(_abc_17692_n5953), .B(_abc_17692_n11109), .Y(_abc_17692_n11179) );
  OR2X2 OR2X2_3739 ( .A(_abc_17692_n11182), .B(_abc_17692_n11183), .Y(_abc_17692_n11184) );
  OR2X2 OR2X2_374 ( .A(_abc_17692_n1614), .B(_abc_17692_n1605), .Y(_abc_17692_n1617) );
  OR2X2 OR2X2_3740 ( .A(_abc_17692_n11019), .B(_abc_17692_n10873), .Y(_abc_17692_n11186) );
  OR2X2 OR2X2_3741 ( .A(_abc_17692_n11186), .B(_abc_17692_n10935), .Y(_abc_17692_n11187) );
  OR2X2 OR2X2_3742 ( .A(_abc_17692_n11018), .B(_abc_17692_n10870), .Y(_abc_17692_n11188) );
  OR2X2 OR2X2_3743 ( .A(_abc_17692_n10539), .B(_abc_17692_n11194), .Y(_abc_17692_n11195) );
  OR2X2 OR2X2_3744 ( .A(_abc_17692_n11197), .B(_abc_17692_n11185), .Y(_abc_17692_n11200) );
  OR2X2 OR2X2_3745 ( .A(_abc_17692_n11202), .B(_abc_17692_n1863_bF_buf8), .Y(_abc_17692_n11203) );
  OR2X2 OR2X2_3746 ( .A(_abc_17692_n11177), .B(_abc_17692_n11203), .Y(_abc_17692_n11204) );
  OR2X2 OR2X2_3747 ( .A(_abc_17692_n11204), .B(_abc_17692_n11156), .Y(_abc_17692_n11205) );
  OR2X2 OR2X2_3748 ( .A(_abc_17692_n11210), .B(_abc_17692_n11211), .Y(_abc_17692_n11212) );
  OR2X2 OR2X2_3749 ( .A(_abc_17692_n11212), .B(_abc_17692_n11209), .Y(_abc_17692_n11213) );
  OR2X2 OR2X2_375 ( .A(_abc_17692_n1619), .B(_abc_17692_n1604), .Y(_abc_17692_n1620) );
  OR2X2 OR2X2_3750 ( .A(_abc_17692_n11215), .B(_abc_17692_n11213), .Y(_abc_17692_n11216) );
  OR2X2 OR2X2_3751 ( .A(_abc_17692_n11216), .B(_abc_17692_n11117), .Y(_abc_17692_n11217) );
  OR2X2 OR2X2_3752 ( .A(_abc_17692_n10997), .B(_abc_17692_n10836), .Y(_abc_17692_n11224) );
  OR2X2 OR2X2_3753 ( .A(_abc_17692_n11224), .B(_abc_17692_n11223), .Y(_abc_17692_n11225) );
  OR2X2 OR2X2_3754 ( .A(_abc_17692_n10997), .B(_abc_17692_n11055), .Y(_abc_17692_n11228) );
  OR2X2 OR2X2_3755 ( .A(_abc_17692_n11234), .B(_abc_17692_n11231), .Y(_abc_17692_n11235) );
  OR2X2 OR2X2_3756 ( .A(_abc_17692_n11235), .B(_abc_17692_n11222), .Y(_abc_17692_n11238) );
  OR2X2 OR2X2_3757 ( .A(_abc_17692_n11013), .B(_abc_17692_n10872), .Y(_abc_17692_n11241) );
  OR2X2 OR2X2_3758 ( .A(_abc_17692_n11241), .B(_abc_17692_n10876), .Y(_abc_17692_n11242) );
  OR2X2 OR2X2_3759 ( .A(_abc_17692_n11013), .B(_abc_17692_n11062), .Y(_abc_17692_n11245) );
  OR2X2 OR2X2_376 ( .A(_abc_17692_n1603), .B(_abc_17692_n1620), .Y(sum_24__FF_INPUT) );
  OR2X2 OR2X2_3760 ( .A(_abc_17692_n11241), .B(_abc_17692_n10882), .Y(_abc_17692_n11249) );
  OR2X2 OR2X2_3761 ( .A(_abc_17692_n11251), .B(_abc_17692_n11248), .Y(_abc_17692_n11252) );
  OR2X2 OR2X2_3762 ( .A(_abc_17692_n11252), .B(_abc_17692_n11184), .Y(_abc_17692_n11253) );
  OR2X2 OR2X2_3763 ( .A(_abc_17692_n11262), .B(_abc_17692_n11260), .Y(_abc_17692_n11263) );
  OR2X2 OR2X2_3764 ( .A(_abc_17692_n11263), .B(_abc_17692_n11259), .Y(_abc_17692_n11264) );
  OR2X2 OR2X2_3765 ( .A(_abc_17692_n10419), .B(_abc_17692_n10310), .Y(_abc_17692_n11267) );
  OR2X2 OR2X2_3766 ( .A(_abc_17692_n11267), .B(_abc_17692_n11266), .Y(_abc_17692_n11268) );
  OR2X2 OR2X2_3767 ( .A(_abc_17692_n11267), .B(_abc_17692_n11270), .Y(_abc_17692_n11271) );
  OR2X2 OR2X2_3768 ( .A(_abc_17692_n10051), .B(_abc_17692_n11271), .Y(_abc_17692_n11272) );
  OR2X2 OR2X2_3769 ( .A(_abc_17692_n11273), .B(_abc_17692_n11275), .Y(_abc_17692_n11276) );
  OR2X2 OR2X2_377 ( .A(_abc_17692_n1600), .B(_abc_17692_n1630), .Y(_abc_17692_n1631) );
  OR2X2 OR2X2_3770 ( .A(_abc_17692_n11278), .B(_abc_17692_n11163), .Y(_abc_17692_n11281) );
  OR2X2 OR2X2_3771 ( .A(_abc_17692_n11283), .B(_abc_17692_n11257), .Y(_abc_17692_n11284) );
  OR2X2 OR2X2_3772 ( .A(_abc_17692_n11284), .B(_abc_17692_n11240), .Y(_abc_17692_n11285) );
  OR2X2 OR2X2_3773 ( .A(_abc_17692_n11285), .B(_abc_17692_n11221), .Y(_abc_17692_n11286) );
  OR2X2 OR2X2_3774 ( .A(_abc_17692_n11288), .B(_abc_17692_n11289), .Y(_abc_17692_n11290) );
  OR2X2 OR2X2_3775 ( .A(_abc_17692_n11287), .B(_abc_17692_n11290), .Y(_abc_17692_n11291) );
  OR2X2 OR2X2_3776 ( .A(_abc_17692_n11291), .B(_abc_17692_n11207), .Y(workunit1_20__FF_INPUT) );
  OR2X2 OR2X2_3777 ( .A(_abc_17692_n11108), .B(_abc_17692_n11100), .Y(_abc_17692_n11293) );
  OR2X2 OR2X2_3778 ( .A(_abc_17692_n5260), .B(workunit2_26_), .Y(_abc_17692_n11294) );
  OR2X2 OR2X2_3779 ( .A(_abc_17692_n7128), .B(workunit2_17_), .Y(_abc_17692_n11295) );
  OR2X2 OR2X2_378 ( .A(_abc_17692_n1632), .B(_abc_17692_n1629), .Y(_abc_17692_n1633) );
  OR2X2 OR2X2_3780 ( .A(_abc_17692_n11293), .B(_abc_17692_n11303), .Y(_abc_17692_n11306) );
  OR2X2 OR2X2_3781 ( .A(_abc_17692_n6088), .B(_abc_17692_n11307), .Y(_abc_17692_n11308) );
  OR2X2 OR2X2_3782 ( .A(_abc_17692_n11309), .B(_abc_17692_n6087), .Y(_abc_17692_n11310) );
  OR2X2 OR2X2_3783 ( .A(_abc_17692_n11314), .B(_abc_17692_n11312), .Y(_abc_17692_n11315) );
  OR2X2 OR2X2_3784 ( .A(_abc_17692_n11317), .B(_abc_17692_n11315), .Y(_abc_17692_n11318) );
  OR2X2 OR2X2_3785 ( .A(_abc_17692_n11316), .B(_abc_17692_n11319), .Y(_abc_17692_n11320) );
  OR2X2 OR2X2_3786 ( .A(_abc_17692_n11307), .B(_abc_17692_n6115), .Y(_abc_17692_n11323) );
  OR2X2 OR2X2_3787 ( .A(_abc_17692_n11309), .B(_abc_17692_n6116), .Y(_abc_17692_n11324) );
  OR2X2 OR2X2_3788 ( .A(_abc_17692_n11328), .B(_abc_17692_n11326), .Y(_abc_17692_n11329) );
  OR2X2 OR2X2_3789 ( .A(_abc_17692_n11174), .B(_abc_17692_n11330), .Y(_abc_17692_n11331) );
  OR2X2 OR2X2_379 ( .A(_abc_17692_n1631), .B(_abc_17692_n1628), .Y(_abc_17692_n1634) );
  OR2X2 OR2X2_3790 ( .A(_abc_17692_n11329), .B(_abc_17692_n11162), .Y(_abc_17692_n11335) );
  OR2X2 OR2X2_3791 ( .A(_abc_17692_n11173), .B(_abc_17692_n11335), .Y(_abc_17692_n11336) );
  OR2X2 OR2X2_3792 ( .A(_abc_17692_n6144), .B(_abc_17692_n11307), .Y(_abc_17692_n11339) );
  OR2X2 OR2X2_3793 ( .A(_abc_17692_n11309), .B(_abc_17692_n6143), .Y(_abc_17692_n11340) );
  OR2X2 OR2X2_3794 ( .A(_abc_17692_n11341), .B(_abc_17692_n4926), .Y(_abc_17692_n11342) );
  OR2X2 OR2X2_3795 ( .A(_abc_17692_n6143), .B(_abc_17692_n11307), .Y(_abc_17692_n11343) );
  OR2X2 OR2X2_3796 ( .A(_abc_17692_n6144), .B(_abc_17692_n11309), .Y(_abc_17692_n11344) );
  OR2X2 OR2X2_3797 ( .A(_abc_17692_n11345), .B(workunit1_21_), .Y(_abc_17692_n11346) );
  OR2X2 OR2X2_3798 ( .A(_abc_17692_n11351), .B(_abc_17692_n11348), .Y(_abc_17692_n11352) );
  OR2X2 OR2X2_3799 ( .A(_abc_17692_n11350), .B(_abc_17692_n11347), .Y(_abc_17692_n11353) );
  OR2X2 OR2X2_38 ( .A(state_7_bF_buf3), .B(state_6_bF_buf4), .Y(_abc_17692_n714_1) );
  OR2X2 OR2X2_380 ( .A(_abc_17692_n1629), .B(_abc_17692_n1584), .Y(_abc_17692_n1637) );
  OR2X2 OR2X2_3800 ( .A(_abc_17692_n11338), .B(_abc_17692_n11355), .Y(_abc_17692_n11356) );
  OR2X2 OR2X2_3801 ( .A(_abc_17692_n11356), .B(_abc_17692_n11322), .Y(_abc_17692_n11357) );
  OR2X2 OR2X2_3802 ( .A(_abc_17692_n11358), .B(_abc_17692_n11359), .Y(_abc_17692_n11360) );
  OR2X2 OR2X2_3803 ( .A(_abc_17692_n11362), .B(_abc_17692_n11363), .Y(_abc_17692_n11364) );
  OR2X2 OR2X2_3804 ( .A(_abc_17692_n11370), .B(_abc_17692_n11367), .Y(_abc_17692_n11371) );
  OR2X2 OR2X2_3805 ( .A(_abc_17692_n11372), .B(_abc_17692_n11357), .Y(_abc_17692_n11373) );
  OR2X2 OR2X2_3806 ( .A(_abc_17692_n11218), .B(_abc_17692_n11375), .Y(_abc_17692_n11376) );
  OR2X2 OR2X2_3807 ( .A(_abc_17692_n11379), .B(_abc_17692_n11377), .Y(_abc_17692_n11380) );
  OR2X2 OR2X2_3808 ( .A(_abc_17692_n11386), .B(_abc_17692_n11319), .Y(_abc_17692_n11387) );
  OR2X2 OR2X2_3809 ( .A(_abc_17692_n11385), .B(_abc_17692_n11315), .Y(_abc_17692_n11388) );
  OR2X2 OR2X2_381 ( .A(_abc_17692_n1615), .B(_abc_17692_n1637), .Y(_abc_17692_n1638) );
  OR2X2 OR2X2_3810 ( .A(_abc_17692_n11394), .B(_abc_17692_n11347), .Y(_abc_17692_n11395) );
  OR2X2 OR2X2_3811 ( .A(_abc_17692_n11393), .B(_abc_17692_n11348), .Y(_abc_17692_n11396) );
  OR2X2 OR2X2_3812 ( .A(_abc_17692_n11401), .B(_abc_17692_n11329), .Y(_abc_17692_n11402) );
  OR2X2 OR2X2_3813 ( .A(_abc_17692_n11403), .B(_abc_17692_n11330), .Y(_abc_17692_n11404) );
  OR2X2 OR2X2_3814 ( .A(_abc_17692_n11406), .B(_abc_17692_n11398), .Y(_abc_17692_n11407) );
  OR2X2 OR2X2_3815 ( .A(_abc_17692_n11407), .B(_abc_17692_n11390), .Y(_abc_17692_n11408) );
  OR2X2 OR2X2_3816 ( .A(_abc_17692_n11408), .B(_abc_17692_n11381), .Y(_abc_17692_n11409) );
  OR2X2 OR2X2_3817 ( .A(_abc_17692_n11411), .B(_abc_17692_n11412), .Y(_abc_17692_n11413) );
  OR2X2 OR2X2_3818 ( .A(_abc_17692_n11410), .B(_abc_17692_n11413), .Y(_abc_17692_n11414) );
  OR2X2 OR2X2_3819 ( .A(_abc_17692_n11414), .B(_abc_17692_n11374), .Y(workunit1_21__FF_INPUT) );
  OR2X2 OR2X2_382 ( .A(_abc_17692_n1647), .B(state_8_bF_buf3), .Y(_abc_17692_n1648) );
  OR2X2 OR2X2_3820 ( .A(_abc_17692_n11095), .B(_abc_17692_n11417), .Y(_abc_17692_n11418) );
  OR2X2 OR2X2_3821 ( .A(_abc_17692_n11419), .B(_abc_17692_n11298), .Y(_abc_17692_n11420) );
  OR2X2 OR2X2_3822 ( .A(_abc_17692_n5430), .B(workunit2_27_), .Y(_abc_17692_n11423) );
  OR2X2 OR2X2_3823 ( .A(_abc_17692_n7385), .B(workunit2_18_), .Y(_abc_17692_n11424) );
  OR2X2 OR2X2_3824 ( .A(_abc_17692_n11427), .B(_abc_17692_n11428), .Y(_abc_17692_n11429) );
  OR2X2 OR2X2_3825 ( .A(_abc_17692_n11431), .B(_abc_17692_n11420), .Y(_abc_17692_n11432) );
  OR2X2 OR2X2_3826 ( .A(_abc_17692_n11430), .B(_abc_17692_n11434), .Y(_abc_17692_n11435) );
  OR2X2 OR2X2_3827 ( .A(_abc_17692_n6272), .B(_abc_17692_n11436), .Y(_abc_17692_n11437) );
  OR2X2 OR2X2_3828 ( .A(_abc_17692_n6273), .B(_abc_17692_n11435), .Y(_abc_17692_n11438) );
  OR2X2 OR2X2_3829 ( .A(_abc_17692_n11439), .B(workunit1_22_), .Y(_abc_17692_n11442) );
  OR2X2 OR2X2_383 ( .A(_abc_17692_n1646), .B(_abc_17692_n1648), .Y(_abc_17692_n1649) );
  OR2X2 OR2X2_3830 ( .A(_abc_17692_n11445), .B(_abc_17692_n11444), .Y(_abc_17692_n11446) );
  OR2X2 OR2X2_3831 ( .A(_abc_17692_n11448), .B(_abc_17692_n11446), .Y(_abc_17692_n11449) );
  OR2X2 OR2X2_3832 ( .A(_abc_17692_n11449), .B(_abc_17692_n11443), .Y(_abc_17692_n11452) );
  OR2X2 OR2X2_3833 ( .A(_abc_17692_n11436), .B(_abc_17692_n6349), .Y(_abc_17692_n11455) );
  OR2X2 OR2X2_3834 ( .A(_abc_17692_n6350), .B(_abc_17692_n11435), .Y(_abc_17692_n11456) );
  OR2X2 OR2X2_3835 ( .A(_abc_17692_n11459), .B(_abc_17692_n11460), .Y(_abc_17692_n11461) );
  OR2X2 OR2X2_3836 ( .A(_abc_17692_n11347), .B(_abc_17692_n11349), .Y(_abc_17692_n11464) );
  OR2X2 OR2X2_3837 ( .A(_abc_17692_n11347), .B(_abc_17692_n11184), .Y(_abc_17692_n11467) );
  OR2X2 OR2X2_3838 ( .A(_abc_17692_n11469), .B(_abc_17692_n11466), .Y(_abc_17692_n11470) );
  OR2X2 OR2X2_3839 ( .A(_abc_17692_n11470), .B(_abc_17692_n11461), .Y(_abc_17692_n11473) );
  OR2X2 OR2X2_384 ( .A(_abc_17692_n1636_1), .B(_abc_17692_n1649), .Y(sum_25__FF_INPUT) );
  OR2X2 OR2X2_3840 ( .A(_abc_17692_n11477), .B(_abc_17692_n11476), .Y(_abc_17692_n11478) );
  OR2X2 OR2X2_3841 ( .A(_abc_17692_n11479), .B(_abc_17692_n5205), .Y(_abc_17692_n11480) );
  OR2X2 OR2X2_3842 ( .A(_abc_17692_n11478), .B(workunit1_22_), .Y(_abc_17692_n11481) );
  OR2X2 OR2X2_3843 ( .A(_abc_17692_n11332), .B(_abc_17692_n11484), .Y(_abc_17692_n11485) );
  OR2X2 OR2X2_3844 ( .A(_abc_17692_n11488), .B(_abc_17692_n11483), .Y(_abc_17692_n11489) );
  OR2X2 OR2X2_3845 ( .A(_abc_17692_n11487), .B(_abc_17692_n11482), .Y(_abc_17692_n11490) );
  OR2X2 OR2X2_3846 ( .A(_abc_17692_n11492), .B(_abc_17692_n11475), .Y(_abc_17692_n11493) );
  OR2X2 OR2X2_3847 ( .A(_abc_17692_n11493), .B(_abc_17692_n11454), .Y(_abc_17692_n11494) );
  OR2X2 OR2X2_3848 ( .A(_abc_17692_n11495), .B(_abc_17692_n11496), .Y(_abc_17692_n11497) );
  OR2X2 OR2X2_3849 ( .A(_abc_17692_n11498), .B(_abc_17692_n5205), .Y(_abc_17692_n11499) );
  OR2X2 OR2X2_385 ( .A(_abc_17692_n1654), .B(_abc_17692_n1651), .Y(_abc_17692_n1655) );
  OR2X2 OR2X2_3850 ( .A(_abc_17692_n11497), .B(workunit1_22_), .Y(_abc_17692_n11500) );
  OR2X2 OR2X2_3851 ( .A(_abc_17692_n11504), .B(_abc_17692_n11503), .Y(_abc_17692_n11505) );
  OR2X2 OR2X2_3852 ( .A(_abc_17692_n11507), .B(_abc_17692_n11505), .Y(_abc_17692_n11508) );
  OR2X2 OR2X2_3853 ( .A(_abc_17692_n11508), .B(_abc_17692_n11502), .Y(_abc_17692_n11511) );
  OR2X2 OR2X2_3854 ( .A(_abc_17692_n11494), .B(_abc_17692_n11513), .Y(_abc_17692_n11514) );
  OR2X2 OR2X2_3855 ( .A(_abc_17692_n11362), .B(_abc_17692_n11375), .Y(_abc_17692_n11517) );
  OR2X2 OR2X2_3856 ( .A(_abc_17692_n11364), .B(_abc_17692_n11118), .Y(_abc_17692_n11519) );
  OR2X2 OR2X2_3857 ( .A(_abc_17692_n11521), .B(_abc_17692_n11518), .Y(_abc_17692_n11522) );
  OR2X2 OR2X2_3858 ( .A(_abc_17692_n11522), .B(_abc_17692_n11501), .Y(_abc_17692_n11525) );
  OR2X2 OR2X2_3859 ( .A(_abc_17692_n11315), .B(_abc_17692_n11141), .Y(_abc_17692_n11529) );
  OR2X2 OR2X2_386 ( .A(_abc_17692_n1597), .B(_abc_17692_n1658), .Y(_abc_17692_n1659) );
  OR2X2 OR2X2_3860 ( .A(_abc_17692_n11533), .B(_abc_17692_n11314), .Y(_abc_17692_n11534) );
  OR2X2 OR2X2_3861 ( .A(_abc_17692_n11531), .B(_abc_17692_n11535), .Y(_abc_17692_n11536) );
  OR2X2 OR2X2_3862 ( .A(_abc_17692_n11536), .B(_abc_17692_n11528), .Y(_abc_17692_n11539) );
  OR2X2 OR2X2_3863 ( .A(_abc_17692_n11348), .B(_abc_17692_n11185), .Y(_abc_17692_n11543) );
  OR2X2 OR2X2_3864 ( .A(_abc_17692_n11547), .B(_abc_17692_n11546), .Y(_abc_17692_n11548) );
  OR2X2 OR2X2_3865 ( .A(_abc_17692_n11545), .B(_abc_17692_n11549), .Y(_abc_17692_n11550) );
  OR2X2 OR2X2_3866 ( .A(_abc_17692_n11550), .B(_abc_17692_n11542), .Y(_abc_17692_n11551) );
  OR2X2 OR2X2_3867 ( .A(_abc_17692_n11326), .B(_abc_17692_n11399), .Y(_abc_17692_n11557) );
  OR2X2 OR2X2_3868 ( .A(_abc_17692_n11560), .B(_abc_17692_n11558), .Y(_abc_17692_n11561) );
  OR2X2 OR2X2_3869 ( .A(_abc_17692_n11561), .B(_abc_17692_n11482), .Y(_abc_17692_n11564) );
  OR2X2 OR2X2_387 ( .A(_abc_17692_n1660_1), .B(_abc_17692_n1622), .Y(_abc_17692_n1661) );
  OR2X2 OR2X2_3870 ( .A(_abc_17692_n11566), .B(_abc_17692_n11555), .Y(_abc_17692_n11567) );
  OR2X2 OR2X2_3871 ( .A(_abc_17692_n11567), .B(_abc_17692_n11541), .Y(_abc_17692_n11568) );
  OR2X2 OR2X2_3872 ( .A(_abc_17692_n11568), .B(_abc_17692_n11527), .Y(_abc_17692_n11569) );
  OR2X2 OR2X2_3873 ( .A(_abc_17692_n11571), .B(_abc_17692_n11572), .Y(_abc_17692_n11573) );
  OR2X2 OR2X2_3874 ( .A(_abc_17692_n11570), .B(_abc_17692_n11573), .Y(_abc_17692_n11574) );
  OR2X2 OR2X2_3875 ( .A(_abc_17692_n11515), .B(_abc_17692_n11574), .Y(workunit1_22__FF_INPUT) );
  OR2X2 OR2X2_3876 ( .A(_abc_17692_n11422), .B(_abc_17692_n11429), .Y(_abc_17692_n11577) );
  OR2X2 OR2X2_3877 ( .A(_abc_17692_n5626), .B(workunit2_28_), .Y(_abc_17692_n11579) );
  OR2X2 OR2X2_3878 ( .A(_abc_17692_n7535), .B(workunit2_19_), .Y(_abc_17692_n11580) );
  OR2X2 OR2X2_3879 ( .A(_abc_17692_n11434), .B(_abc_17692_n11427), .Y(_abc_17692_n11590) );
  OR2X2 OR2X2_388 ( .A(_abc_17692_n1664), .B(_abc_17692_n1656), .Y(_abc_17692_n1665) );
  OR2X2 OR2X2_3880 ( .A(_abc_17692_n11589), .B(_abc_17692_n11591), .Y(_abc_17692_n11592) );
  OR2X2 OR2X2_3881 ( .A(_abc_17692_n6501), .B(_abc_17692_n11592), .Y(_abc_17692_n11593) );
  OR2X2 OR2X2_3882 ( .A(_abc_17692_n11590), .B(_abc_17692_n11587), .Y(_abc_17692_n11594) );
  OR2X2 OR2X2_3883 ( .A(_abc_17692_n11578), .B(_abc_17692_n11588), .Y(_abc_17692_n11595) );
  OR2X2 OR2X2_3884 ( .A(_abc_17692_n6493), .B(_abc_17692_n11596), .Y(_abc_17692_n11597) );
  OR2X2 OR2X2_3885 ( .A(_abc_17692_n11598), .B(workunit1_23_), .Y(_abc_17692_n11599) );
  OR2X2 OR2X2_3886 ( .A(_abc_17692_n6501), .B(_abc_17692_n11596), .Y(_abc_17692_n11600) );
  OR2X2 OR2X2_3887 ( .A(_abc_17692_n6493), .B(_abc_17692_n11592), .Y(_abc_17692_n11601) );
  OR2X2 OR2X2_3888 ( .A(_abc_17692_n11602), .B(_abc_17692_n5378), .Y(_abc_17692_n11603) );
  OR2X2 OR2X2_3889 ( .A(_abc_17692_n11606), .B(_abc_17692_n11604), .Y(_abc_17692_n11607) );
  OR2X2 OR2X2_389 ( .A(_abc_17692_n1642), .B(_abc_17692_n1670), .Y(_abc_17692_n1671) );
  OR2X2 OR2X2_3890 ( .A(_abc_17692_n11605), .B(_abc_17692_n11608), .Y(_abc_17692_n11609) );
  OR2X2 OR2X2_3891 ( .A(_abc_17692_n11596), .B(_abc_17692_n6559), .Y(_abc_17692_n11612) );
  OR2X2 OR2X2_3892 ( .A(_abc_17692_n11592), .B(_abc_17692_n6563), .Y(_abc_17692_n11613) );
  OR2X2 OR2X2_3893 ( .A(_abc_17692_n11592), .B(_abc_17692_n6559), .Y(_abc_17692_n11616) );
  OR2X2 OR2X2_3894 ( .A(_abc_17692_n11596), .B(_abc_17692_n6563), .Y(_abc_17692_n11617) );
  OR2X2 OR2X2_3895 ( .A(_abc_17692_n11615), .B(_abc_17692_n11619), .Y(_abc_17692_n11620) );
  OR2X2 OR2X2_3896 ( .A(_abc_17692_n11625), .B(_abc_17692_n11621), .Y(_abc_17692_n11626) );
  OR2X2 OR2X2_3897 ( .A(_abc_17692_n11624), .B(_abc_17692_n11620), .Y(_abc_17692_n11627) );
  OR2X2 OR2X2_3898 ( .A(_abc_17692_n11592), .B(_abc_17692_n6528), .Y(_abc_17692_n11630) );
  OR2X2 OR2X2_3899 ( .A(_abc_17692_n11596), .B(_abc_17692_n6532), .Y(_abc_17692_n11631) );
  OR2X2 OR2X2_39 ( .A(state_4_), .B(state_2_), .Y(_abc_17692_n718) );
  OR2X2 OR2X2_390 ( .A(_abc_17692_n1640), .B(_abc_17692_n1671), .Y(_abc_17692_n1672) );
  OR2X2 OR2X2_3900 ( .A(_abc_17692_n11632), .B(workunit1_23_), .Y(_abc_17692_n11633) );
  OR2X2 OR2X2_3901 ( .A(_abc_17692_n11596), .B(_abc_17692_n6528), .Y(_abc_17692_n11634) );
  OR2X2 OR2X2_3902 ( .A(_abc_17692_n11592), .B(_abc_17692_n6532), .Y(_abc_17692_n11635) );
  OR2X2 OR2X2_3903 ( .A(_abc_17692_n11636), .B(_abc_17692_n5378), .Y(_abc_17692_n11637) );
  OR2X2 OR2X2_3904 ( .A(_abc_17692_n11458), .B(_abc_17692_n5205), .Y(_abc_17692_n11639) );
  OR2X2 OR2X2_3905 ( .A(_abc_17692_n11641), .B(_abc_17692_n11638), .Y(_abc_17692_n11642) );
  OR2X2 OR2X2_3906 ( .A(_abc_17692_n11643), .B(_abc_17692_n11644), .Y(_abc_17692_n11645) );
  OR2X2 OR2X2_3907 ( .A(_abc_17692_n11640), .B(_abc_17692_n11645), .Y(_abc_17692_n11646) );
  OR2X2 OR2X2_3908 ( .A(_abc_17692_n11629), .B(_abc_17692_n11648), .Y(_abc_17692_n11649) );
  OR2X2 OR2X2_3909 ( .A(_abc_17692_n11649), .B(_abc_17692_n11611), .Y(_abc_17692_n11650) );
  OR2X2 OR2X2_391 ( .A(_abc_17692_n1672), .B(_abc_17692_n1655), .Y(_abc_17692_n1675) );
  OR2X2 OR2X2_3910 ( .A(_abc_17692_n6597_1), .B(_abc_17692_n11596), .Y(_abc_17692_n11651) );
  OR2X2 OR2X2_3911 ( .A(_abc_17692_n6592), .B(_abc_17692_n11592), .Y(_abc_17692_n11652) );
  OR2X2 OR2X2_3912 ( .A(_abc_17692_n6597_1), .B(_abc_17692_n11592), .Y(_abc_17692_n11655) );
  OR2X2 OR2X2_3913 ( .A(_abc_17692_n6592), .B(_abc_17692_n11596), .Y(_abc_17692_n11656) );
  OR2X2 OR2X2_3914 ( .A(_abc_17692_n11654), .B(_abc_17692_n11658), .Y(_abc_17692_n11659) );
  OR2X2 OR2X2_3915 ( .A(_abc_17692_n11497), .B(_abc_17692_n5205), .Y(_abc_17692_n11660) );
  OR2X2 OR2X2_3916 ( .A(_abc_17692_n11657), .B(workunit1_23_), .Y(_abc_17692_n11664) );
  OR2X2 OR2X2_3917 ( .A(_abc_17692_n11653), .B(_abc_17692_n5378), .Y(_abc_17692_n11665) );
  OR2X2 OR2X2_3918 ( .A(_abc_17692_n11663), .B(_abc_17692_n11667), .Y(_abc_17692_n11668) );
  OR2X2 OR2X2_3919 ( .A(_abc_17692_n11669), .B(_abc_17692_n11650), .Y(_abc_17692_n11670) );
  OR2X2 OR2X2_392 ( .A(_abc_17692_n1678), .B(state_8_bF_buf2), .Y(_abc_17692_n1679) );
  OR2X2 OR2X2_3920 ( .A(_abc_17692_n11523), .B(_abc_17692_n11672), .Y(_abc_17692_n11673) );
  OR2X2 OR2X2_3921 ( .A(_abc_17692_n11674), .B(_abc_17692_n11666), .Y(_abc_17692_n11675) );
  OR2X2 OR2X2_3922 ( .A(_abc_17692_n11673), .B(_abc_17692_n11659), .Y(_abc_17692_n11676) );
  OR2X2 OR2X2_3923 ( .A(_abc_17692_n11683), .B(_abc_17692_n11608), .Y(_abc_17692_n11684) );
  OR2X2 OR2X2_3924 ( .A(_abc_17692_n11682), .B(_abc_17692_n11604), .Y(_abc_17692_n11685) );
  OR2X2 OR2X2_3925 ( .A(_abc_17692_n11552), .B(_abc_17692_n11459), .Y(_abc_17692_n11688) );
  OR2X2 OR2X2_3926 ( .A(_abc_17692_n11689), .B(_abc_17692_n11638), .Y(_abc_17692_n11690) );
  OR2X2 OR2X2_3927 ( .A(_abc_17692_n11688), .B(_abc_17692_n11645), .Y(_abc_17692_n11691) );
  OR2X2 OR2X2_3928 ( .A(_abc_17692_n11562), .B(_abc_17692_n11694), .Y(_abc_17692_n11695) );
  OR2X2 OR2X2_3929 ( .A(_abc_17692_n11696), .B(_abc_17692_n11621), .Y(_abc_17692_n11697) );
  OR2X2 OR2X2_393 ( .A(_abc_17692_n1677), .B(_abc_17692_n1679), .Y(_abc_17692_n1680) );
  OR2X2 OR2X2_3930 ( .A(_abc_17692_n11695), .B(_abc_17692_n11620), .Y(_abc_17692_n11698) );
  OR2X2 OR2X2_3931 ( .A(_abc_17692_n11700), .B(_abc_17692_n11693), .Y(_abc_17692_n11701) );
  OR2X2 OR2X2_3932 ( .A(_abc_17692_n11701), .B(_abc_17692_n11687), .Y(_abc_17692_n11702) );
  OR2X2 OR2X2_3933 ( .A(_abc_17692_n11702), .B(_abc_17692_n11678), .Y(_abc_17692_n11703) );
  OR2X2 OR2X2_3934 ( .A(_abc_17692_n11705), .B(_abc_17692_n11706), .Y(_abc_17692_n11707) );
  OR2X2 OR2X2_3935 ( .A(_abc_17692_n11704), .B(_abc_17692_n11707), .Y(_abc_17692_n11708) );
  OR2X2 OR2X2_3936 ( .A(_abc_17692_n11671), .B(_abc_17692_n11708), .Y(workunit1_23__FF_INPUT) );
  OR2X2 OR2X2_3937 ( .A(_abc_17692_n5769), .B(workunit2_29_), .Y(_abc_17692_n11710) );
  OR2X2 OR2X2_3938 ( .A(_abc_17692_n7812), .B(workunit2_20_), .Y(_abc_17692_n11711) );
  OR2X2 OR2X2_3939 ( .A(_abc_17692_n11714), .B(_abc_17692_n11715), .Y(_abc_17692_n11716) );
  OR2X2 OR2X2_394 ( .A(_abc_17692_n1669), .B(_abc_17692_n1680), .Y(sum_26__FF_INPUT) );
  OR2X2 OR2X2_3940 ( .A(_abc_17692_n11718), .B(_abc_17692_n11585), .Y(_abc_17692_n11719) );
  OR2X2 OR2X2_3941 ( .A(_abc_17692_n11721), .B(_abc_17692_n11421), .Y(_abc_17692_n11722) );
  OR2X2 OR2X2_3942 ( .A(_abc_17692_n11417), .B(_abc_17692_n11721), .Y(_abc_17692_n11724) );
  OR2X2 OR2X2_3943 ( .A(_abc_17692_n11094), .B(_abc_17692_n11724), .Y(_abc_17692_n11725) );
  OR2X2 OR2X2_3944 ( .A(_abc_17692_n11724), .B(_abc_17692_n11087), .Y(_abc_17692_n11727) );
  OR2X2 OR2X2_3945 ( .A(_abc_17692_n10484), .B(_abc_17692_n11727), .Y(_abc_17692_n11728) );
  OR2X2 OR2X2_3946 ( .A(_abc_17692_n11731), .B(_abc_17692_n11732), .Y(_abc_17692_n11733) );
  OR2X2 OR2X2_3947 ( .A(_abc_17692_n6700), .B(_abc_17692_n11734), .Y(_abc_17692_n11735) );
  OR2X2 OR2X2_3948 ( .A(_abc_17692_n6699), .B(_abc_17692_n11733), .Y(_abc_17692_n11736) );
  OR2X2 OR2X2_3949 ( .A(_abc_17692_n11740), .B(_abc_17692_n11738), .Y(_abc_17692_n11741) );
  OR2X2 OR2X2_395 ( .A(_abc_17692_n1682), .B(delta_27_), .Y(_abc_17692_n1684) );
  OR2X2 OR2X2_3950 ( .A(_abc_17692_n11654), .B(_abc_17692_n11660), .Y(_abc_17692_n11745) );
  OR2X2 OR2X2_3951 ( .A(_abc_17692_n11749), .B(_abc_17692_n11127), .Y(_abc_17692_n11750) );
  OR2X2 OR2X2_3952 ( .A(_abc_17692_n11756), .B(_abc_17692_n11741), .Y(_abc_17692_n11759) );
  OR2X2 OR2X2_3953 ( .A(_abc_17692_n11760), .B(_abc_17692_n4047_bF_buf2), .Y(_abc_17692_n11761) );
  OR2X2 OR2X2_3954 ( .A(_abc_17692_n6793), .B(_abc_17692_n11734), .Y(_abc_17692_n11762) );
  OR2X2 OR2X2_3955 ( .A(_abc_17692_n6792), .B(_abc_17692_n11733), .Y(_abc_17692_n11763) );
  OR2X2 OR2X2_3956 ( .A(_abc_17692_n11764), .B(workunit1_24_), .Y(_abc_17692_n11767) );
  OR2X2 OR2X2_3957 ( .A(_abc_17692_n11775), .B(_abc_17692_n11774), .Y(_abc_17692_n11776) );
  OR2X2 OR2X2_3958 ( .A(_abc_17692_n11773), .B(_abc_17692_n11776), .Y(_abc_17692_n11777) );
  OR2X2 OR2X2_3959 ( .A(_abc_17692_n11778), .B(_abc_17692_n11777), .Y(_abc_17692_n11779) );
  OR2X2 OR2X2_396 ( .A(_abc_17692_n1685_1), .B(_abc_17692_n1683), .Y(_abc_17692_n1686) );
  OR2X2 OR2X2_3960 ( .A(_abc_17692_n11772), .B(_abc_17692_n11779), .Y(_abc_17692_n11780) );
  OR2X2 OR2X2_3961 ( .A(_abc_17692_n11780), .B(_abc_17692_n11769), .Y(_abc_17692_n11781) );
  OR2X2 OR2X2_3962 ( .A(_abc_17692_n6747), .B(_abc_17692_n11734), .Y(_abc_17692_n11786) );
  OR2X2 OR2X2_3963 ( .A(_abc_17692_n6746), .B(_abc_17692_n11733), .Y(_abc_17692_n11787) );
  OR2X2 OR2X2_3964 ( .A(_abc_17692_n11791), .B(_abc_17692_n11789), .Y(_abc_17692_n11792) );
  OR2X2 OR2X2_3965 ( .A(_abc_17692_n11795), .B(_abc_17692_n11619), .Y(_abc_17692_n11796) );
  OR2X2 OR2X2_3966 ( .A(_abc_17692_n11796), .B(_abc_17692_n11794), .Y(_abc_17692_n11797) );
  OR2X2 OR2X2_3967 ( .A(_abc_17692_n11797), .B(_abc_17692_n11800), .Y(_abc_17692_n11801) );
  OR2X2 OR2X2_3968 ( .A(_abc_17692_n11803), .B(_abc_17692_n11801), .Y(_abc_17692_n11804) );
  OR2X2 OR2X2_3969 ( .A(_abc_17692_n11804), .B(_abc_17692_n11792), .Y(_abc_17692_n11807) );
  OR2X2 OR2X2_397 ( .A(_abc_17692_n1686), .B(_abc_17692_n1651), .Y(_abc_17692_n1687) );
  OR2X2 OR2X2_3970 ( .A(_abc_17692_n6841), .B(_abc_17692_n11734), .Y(_abc_17692_n11810) );
  OR2X2 OR2X2_3971 ( .A(_abc_17692_n6840), .B(_abc_17692_n11733), .Y(_abc_17692_n11811) );
  OR2X2 OR2X2_3972 ( .A(_abc_17692_n11815), .B(_abc_17692_n11813), .Y(_abc_17692_n11816) );
  OR2X2 OR2X2_3973 ( .A(_abc_17692_n11645), .B(_abc_17692_n11542), .Y(_abc_17692_n11817) );
  OR2X2 OR2X2_3974 ( .A(_abc_17692_n11817), .B(_abc_17692_n11467), .Y(_abc_17692_n11818) );
  OR2X2 OR2X2_3975 ( .A(_abc_17692_n11195), .B(_abc_17692_n11818), .Y(_abc_17692_n11819) );
  OR2X2 OR2X2_3976 ( .A(_abc_17692_n11818), .B(_abc_17692_n11191), .Y(_abc_17692_n11820) );
  OR2X2 OR2X2_3977 ( .A(_abc_17692_n11817), .B(_abc_17692_n11465), .Y(_abc_17692_n11821) );
  OR2X2 OR2X2_3978 ( .A(_abc_17692_n11643), .B(_abc_17692_n11639), .Y(_abc_17692_n11822) );
  OR2X2 OR2X2_3979 ( .A(_abc_17692_n11827), .B(_abc_17692_n11816), .Y(_abc_17692_n11830) );
  OR2X2 OR2X2_398 ( .A(_abc_17692_n1666), .B(_abc_17692_n1687), .Y(_abc_17692_n1688) );
  OR2X2 OR2X2_3980 ( .A(_abc_17692_n11832), .B(_abc_17692_n1863_bF_buf0), .Y(_abc_17692_n11833) );
  OR2X2 OR2X2_3981 ( .A(_abc_17692_n11833), .B(_abc_17692_n11809), .Y(_abc_17692_n11834) );
  OR2X2 OR2X2_3982 ( .A(_abc_17692_n11834), .B(_abc_17692_n11785), .Y(_abc_17692_n11835) );
  OR2X2 OR2X2_3983 ( .A(_abc_17692_n11844), .B(_abc_17692_n11843), .Y(_abc_17692_n11845) );
  OR2X2 OR2X2_3984 ( .A(_abc_17692_n11845), .B(_abc_17692_n11842), .Y(_abc_17692_n11846) );
  OR2X2 OR2X2_3985 ( .A(_abc_17692_n11846), .B(_abc_17692_n11841), .Y(_abc_17692_n11847) );
  OR2X2 OR2X2_3986 ( .A(_abc_17692_n11847), .B(_abc_17692_n11848), .Y(_abc_17692_n11849) );
  OR2X2 OR2X2_3987 ( .A(_abc_17692_n11849), .B(_abc_17692_n11838), .Y(_abc_17692_n11850) );
  OR2X2 OR2X2_3988 ( .A(_abc_17692_n11604), .B(_abc_17692_n11443), .Y(_abc_17692_n11855) );
  OR2X2 OR2X2_3989 ( .A(_abc_17692_n11855), .B(_abc_17692_n11529), .Y(_abc_17692_n11856) );
  OR2X2 OR2X2_399 ( .A(_abc_17692_n1663), .B(_abc_17692_n1690), .Y(_abc_17692_n1691) );
  OR2X2 OR2X2_3990 ( .A(_abc_17692_n11230), .B(_abc_17692_n11856), .Y(_abc_17692_n11857) );
  OR2X2 OR2X2_3991 ( .A(_abc_17692_n11855), .B(_abc_17692_n11534), .Y(_abc_17692_n11858) );
  OR2X2 OR2X2_3992 ( .A(_abc_17692_n11604), .B(_abc_17692_n11681), .Y(_abc_17692_n11861) );
  OR2X2 OR2X2_3993 ( .A(_abc_17692_n9999), .B(_abc_17692_n10619), .Y(_abc_17692_n11865) );
  OR2X2 OR2X2_3994 ( .A(_abc_17692_n11867), .B(_abc_17692_n11856), .Y(_abc_17692_n11868) );
  OR2X2 OR2X2_3995 ( .A(_abc_17692_n11866), .B(_abc_17692_n11868), .Y(_abc_17692_n11869) );
  OR2X2 OR2X2_3996 ( .A(_abc_17692_n11871), .B(_abc_17692_n11768), .Y(_abc_17692_n11874) );
  OR2X2 OR2X2_3997 ( .A(_abc_17692_n11638), .B(_abc_17692_n11461), .Y(_abc_17692_n11878) );
  OR2X2 OR2X2_3998 ( .A(_abc_17692_n11878), .B(_abc_17692_n11543), .Y(_abc_17692_n11879) );
  OR2X2 OR2X2_3999 ( .A(_abc_17692_n11879), .B(_abc_17692_n11247), .Y(_abc_17692_n11880) );
  OR2X2 OR2X2_4 ( .A(_abc_17692_n632), .B(mode), .Y(_abc_17692_n633) );
  OR2X2 OR2X2_40 ( .A(_abc_17692_n718), .B(state_11_), .Y(_abc_17692_n719) );
  OR2X2 OR2X2_400 ( .A(_abc_17692_n1698), .B(_abc_17692_n1699), .Y(_abc_17692_n1700) );
  OR2X2 OR2X2_4000 ( .A(_abc_17692_n11878), .B(_abc_17692_n11548), .Y(_abc_17692_n11881) );
  OR2X2 OR2X2_4001 ( .A(_abc_17692_n11638), .B(_abc_17692_n11884), .Y(_abc_17692_n11885) );
  OR2X2 OR2X2_4002 ( .A(_abc_17692_n11879), .B(_abc_17692_n11249), .Y(_abc_17692_n11889) );
  OR2X2 OR2X2_4003 ( .A(_abc_17692_n11889), .B(_abc_17692_n10880), .Y(_abc_17692_n11890) );
  OR2X2 OR2X2_4004 ( .A(_abc_17692_n11892), .B(_abc_17692_n11877), .Y(_abc_17692_n11893) );
  OR2X2 OR2X2_4005 ( .A(_abc_17692_n11891), .B(_abc_17692_n11816), .Y(_abc_17692_n11894) );
  OR2X2 OR2X2_4006 ( .A(_abc_17692_n11904), .B(_abc_17692_n11903), .Y(_abc_17692_n11905) );
  OR2X2 OR2X2_4007 ( .A(_abc_17692_n11905), .B(_abc_17692_n11902), .Y(_abc_17692_n11906) );
  OR2X2 OR2X2_4008 ( .A(_abc_17692_n11906), .B(_abc_17692_n11901), .Y(_abc_17692_n11907) );
  OR2X2 OR2X2_4009 ( .A(_abc_17692_n11907), .B(_abc_17692_n11900), .Y(_abc_17692_n11908) );
  OR2X2 OR2X2_401 ( .A(_abc_17692_n1673), .B(_abc_17692_n1700), .Y(_abc_17692_n1701) );
  OR2X2 OR2X2_4010 ( .A(_abc_17692_n11909), .B(_abc_17692_n11792), .Y(_abc_17692_n11910) );
  OR2X2 OR2X2_4011 ( .A(_abc_17692_n11908), .B(_abc_17692_n11911), .Y(_abc_17692_n11912) );
  OR2X2 OR2X2_4012 ( .A(_abc_17692_n11914), .B(_abc_17692_n11896), .Y(_abc_17692_n11915) );
  OR2X2 OR2X2_4013 ( .A(_abc_17692_n11876), .B(_abc_17692_n11915), .Y(_abc_17692_n11916) );
  OR2X2 OR2X2_4014 ( .A(_abc_17692_n11916), .B(_abc_17692_n11854), .Y(_abc_17692_n11917) );
  OR2X2 OR2X2_4015 ( .A(_abc_17692_n11919), .B(_abc_17692_n11920), .Y(_abc_17692_n11921) );
  OR2X2 OR2X2_4016 ( .A(_abc_17692_n11918), .B(_abc_17692_n11921), .Y(_abc_17692_n11922) );
  OR2X2 OR2X2_4017 ( .A(_abc_17692_n11837), .B(_abc_17692_n11922), .Y(workunit1_24__FF_INPUT) );
  OR2X2 OR2X2_4018 ( .A(_abc_17692_n11731), .B(_abc_17692_n11714), .Y(_abc_17692_n11924) );
  OR2X2 OR2X2_4019 ( .A(_abc_17692_n6095), .B(workunit2_30_), .Y(_abc_17692_n11926) );
  OR2X2 OR2X2_402 ( .A(_abc_17692_n1709), .B(_abc_17692_n1697), .Y(_abc_17692_n1710) );
  OR2X2 OR2X2_4020 ( .A(_abc_17692_n7968), .B(workunit2_21_), .Y(_abc_17692_n11927) );
  OR2X2 OR2X2_4021 ( .A(_abc_17692_n11936), .B(_abc_17692_n11937), .Y(_abc_17692_n11938) );
  OR2X2 OR2X2_4022 ( .A(_abc_17692_n7010), .B(_abc_17692_n11938), .Y(_abc_17692_n11939) );
  OR2X2 OR2X2_4023 ( .A(_abc_17692_n7007), .B(_abc_17692_n11940), .Y(_abc_17692_n11941) );
  OR2X2 OR2X2_4024 ( .A(_abc_17692_n11942), .B(workunit1_25_), .Y(_abc_17692_n11943) );
  OR2X2 OR2X2_4025 ( .A(_abc_17692_n7010), .B(_abc_17692_n11940), .Y(_abc_17692_n11944) );
  OR2X2 OR2X2_4026 ( .A(_abc_17692_n7007), .B(_abc_17692_n11938), .Y(_abc_17692_n11945) );
  OR2X2 OR2X2_4027 ( .A(_abc_17692_n11946), .B(_abc_17692_n5782), .Y(_abc_17692_n11947) );
  OR2X2 OR2X2_4028 ( .A(_abc_17692_n11953), .B(_abc_17692_n11949), .Y(_abc_17692_n11954) );
  OR2X2 OR2X2_4029 ( .A(_abc_17692_n11955), .B(_abc_17692_n11948), .Y(_abc_17692_n11956) );
  OR2X2 OR2X2_403 ( .A(_abc_17692_n1696), .B(_abc_17692_n1710), .Y(sum_27__FF_INPUT) );
  OR2X2 OR2X2_4030 ( .A(_abc_17692_n7065), .B(_abc_17692_n11938), .Y(_abc_17692_n11959) );
  OR2X2 OR2X2_4031 ( .A(_abc_17692_n7064), .B(_abc_17692_n11940), .Y(_abc_17692_n11960) );
  OR2X2 OR2X2_4032 ( .A(_abc_17692_n11961), .B(workunit1_25_), .Y(_abc_17692_n11962) );
  OR2X2 OR2X2_4033 ( .A(_abc_17692_n7065), .B(_abc_17692_n11940), .Y(_abc_17692_n11963) );
  OR2X2 OR2X2_4034 ( .A(_abc_17692_n7064), .B(_abc_17692_n11938), .Y(_abc_17692_n11964) );
  OR2X2 OR2X2_4035 ( .A(_abc_17692_n11965), .B(_abc_17692_n5782), .Y(_abc_17692_n11966) );
  OR2X2 OR2X2_4036 ( .A(_abc_17692_n11971), .B(_abc_17692_n11967), .Y(_abc_17692_n11972) );
  OR2X2 OR2X2_4037 ( .A(_abc_17692_n11970), .B(_abc_17692_n11973), .Y(_abc_17692_n11974) );
  OR2X2 OR2X2_4038 ( .A(_abc_17692_n7038), .B(_abc_17692_n11940), .Y(_abc_17692_n11977) );
  OR2X2 OR2X2_4039 ( .A(_abc_17692_n7035), .B(_abc_17692_n11938), .Y(_abc_17692_n11978) );
  OR2X2 OR2X2_404 ( .A(_abc_17692_n1712), .B(delta_28_), .Y(_abc_17692_n1714) );
  OR2X2 OR2X2_4040 ( .A(_abc_17692_n7038), .B(_abc_17692_n11938), .Y(_abc_17692_n11981) );
  OR2X2 OR2X2_4041 ( .A(_abc_17692_n7035), .B(_abc_17692_n11940), .Y(_abc_17692_n11982) );
  OR2X2 OR2X2_4042 ( .A(_abc_17692_n11980), .B(_abc_17692_n11984), .Y(_abc_17692_n11985) );
  OR2X2 OR2X2_4043 ( .A(_abc_17692_n11988), .B(_abc_17692_n11985), .Y(_abc_17692_n11989) );
  OR2X2 OR2X2_4044 ( .A(_abc_17692_n11991), .B(_abc_17692_n11990), .Y(_abc_17692_n11992) );
  OR2X2 OR2X2_4045 ( .A(_abc_17692_n11994), .B(_abc_17692_n11976), .Y(_abc_17692_n11995) );
  OR2X2 OR2X2_4046 ( .A(_abc_17692_n11995), .B(_abc_17692_n11958), .Y(_abc_17692_n11996) );
  OR2X2 OR2X2_4047 ( .A(_abc_17692_n6978), .B(_abc_17692_n11940), .Y(_abc_17692_n11997) );
  OR2X2 OR2X2_4048 ( .A(_abc_17692_n6983), .B(_abc_17692_n11938), .Y(_abc_17692_n11998) );
  OR2X2 OR2X2_4049 ( .A(_abc_17692_n6978), .B(_abc_17692_n11938), .Y(_abc_17692_n12002) );
  OR2X2 OR2X2_405 ( .A(_abc_17692_n1715), .B(_abc_17692_n1713), .Y(_abc_17692_n1716) );
  OR2X2 OR2X2_4050 ( .A(_abc_17692_n6983), .B(_abc_17692_n11940), .Y(_abc_17692_n12003) );
  OR2X2 OR2X2_4051 ( .A(_abc_17692_n12000), .B(_abc_17692_n12005), .Y(_abc_17692_n12012) );
  OR2X2 OR2X2_4052 ( .A(_abc_17692_n12014), .B(_abc_17692_n12011), .Y(_abc_17692_n12015) );
  OR2X2 OR2X2_4053 ( .A(_abc_17692_n12016), .B(_abc_17692_n11996), .Y(_abc_17692_n12017) );
  OR2X2 OR2X2_4054 ( .A(_abc_17692_n12021), .B(_abc_17692_n12012), .Y(_abc_17692_n12022) );
  OR2X2 OR2X2_4055 ( .A(_abc_17692_n12020), .B(_abc_17692_n12007), .Y(_abc_17692_n12023) );
  OR2X2 OR2X2_4056 ( .A(_abc_17692_n12027), .B(_abc_17692_n11949), .Y(_abc_17692_n12028) );
  OR2X2 OR2X2_4057 ( .A(_abc_17692_n12026), .B(_abc_17692_n11948), .Y(_abc_17692_n12029) );
  OR2X2 OR2X2_4058 ( .A(_abc_17692_n12034), .B(_abc_17692_n11973), .Y(_abc_17692_n12035) );
  OR2X2 OR2X2_4059 ( .A(_abc_17692_n12033), .B(_abc_17692_n11967), .Y(_abc_17692_n12036) );
  OR2X2 OR2X2_406 ( .A(_abc_17692_n1692), .B(_abc_17692_n1717), .Y(_abc_17692_n1718) );
  OR2X2 OR2X2_4060 ( .A(_abc_17692_n12043), .B(_abc_17692_n12041), .Y(_abc_17692_n12044) );
  OR2X2 OR2X2_4061 ( .A(_abc_17692_n12045), .B(_abc_17692_n12038), .Y(_abc_17692_n12046) );
  OR2X2 OR2X2_4062 ( .A(_abc_17692_n12046), .B(_abc_17692_n12031), .Y(_abc_17692_n12047) );
  OR2X2 OR2X2_4063 ( .A(_abc_17692_n12047), .B(_abc_17692_n12025), .Y(_abc_17692_n12048) );
  OR2X2 OR2X2_4064 ( .A(_abc_17692_n12050), .B(_abc_17692_n12051), .Y(_abc_17692_n12052) );
  OR2X2 OR2X2_4065 ( .A(_abc_17692_n12049), .B(_abc_17692_n12052), .Y(_abc_17692_n12053) );
  OR2X2 OR2X2_4066 ( .A(_abc_17692_n12018), .B(_abc_17692_n12053), .Y(workunit1_25__FF_INPUT) );
  OR2X2 OR2X2_4067 ( .A(_abc_17692_n11949), .B(_abc_17692_n11952), .Y(_abc_17692_n12057) );
  OR2X2 OR2X2_4068 ( .A(_abc_17692_n12056), .B(_abc_17692_n12059), .Y(_abc_17692_n12060) );
  OR2X2 OR2X2_4069 ( .A(_abc_17692_n11714), .B(_abc_17692_n11930), .Y(_abc_17692_n12063) );
  OR2X2 OR2X2_407 ( .A(_abc_17692_n1721), .B(_abc_17692_n1716), .Y(_abc_17692_n1722) );
  OR2X2 OR2X2_4070 ( .A(_abc_17692_n12062), .B(_abc_17692_n12064), .Y(_abc_17692_n12065) );
  OR2X2 OR2X2_4071 ( .A(_abc_17692_n6293), .B(workunit2_31_), .Y(_abc_17692_n12067) );
  OR2X2 OR2X2_4072 ( .A(_abc_17692_n8202), .B(workunit2_22_), .Y(_abc_17692_n12068) );
  OR2X2 OR2X2_4073 ( .A(_abc_17692_n12071), .B(_abc_17692_n12072), .Y(_abc_17692_n12073) );
  OR2X2 OR2X2_4074 ( .A(_abc_17692_n12074), .B(_abc_17692_n12076), .Y(_abc_17692_n12077) );
  OR2X2 OR2X2_4075 ( .A(_abc_17692_n7205), .B(_abc_17692_n12078), .Y(_abc_17692_n12079) );
  OR2X2 OR2X2_4076 ( .A(_abc_17692_n7206), .B(_abc_17692_n12077), .Y(_abc_17692_n12080) );
  OR2X2 OR2X2_4077 ( .A(_abc_17692_n12081), .B(workunit1_26_), .Y(_abc_17692_n12084) );
  OR2X2 OR2X2_4078 ( .A(_abc_17692_n12060), .B(_abc_17692_n12085), .Y(_abc_17692_n12086) );
  OR2X2 OR2X2_4079 ( .A(_abc_17692_n12091), .B(_abc_17692_n12092), .Y(_abc_17692_n12093) );
  OR2X2 OR2X2_408 ( .A(_abc_17692_n1720), .B(_abc_17692_n1723), .Y(_abc_17692_n1724) );
  OR2X2 OR2X2_4080 ( .A(_abc_17692_n12094), .B(_abc_17692_n6065), .Y(_abc_17692_n12095) );
  OR2X2 OR2X2_4081 ( .A(_abc_17692_n12093), .B(workunit1_26_), .Y(_abc_17692_n12096) );
  OR2X2 OR2X2_4082 ( .A(_abc_17692_n11984), .B(_abc_17692_n11986), .Y(_abc_17692_n12099) );
  OR2X2 OR2X2_4083 ( .A(_abc_17692_n12101), .B(_abc_17692_n11980), .Y(_abc_17692_n12102) );
  OR2X2 OR2X2_4084 ( .A(_abc_17692_n12103), .B(_abc_17692_n12098), .Y(_abc_17692_n12104) );
  OR2X2 OR2X2_4085 ( .A(_abc_17692_n12102), .B(_abc_17692_n12097), .Y(_abc_17692_n12105) );
  OR2X2 OR2X2_4086 ( .A(_abc_17692_n7239), .B(_abc_17692_n12078), .Y(_abc_17692_n12108) );
  OR2X2 OR2X2_4087 ( .A(_abc_17692_n7237), .B(_abc_17692_n12077), .Y(_abc_17692_n12109) );
  OR2X2 OR2X2_4088 ( .A(_abc_17692_n12112), .B(_abc_17692_n12113), .Y(_abc_17692_n12114) );
  OR2X2 OR2X2_4089 ( .A(_abc_17692_n12117), .B(_abc_17692_n12116), .Y(_abc_17692_n12118) );
  OR2X2 OR2X2_409 ( .A(_abc_17692_n1703), .B(_abc_17692_n1729), .Y(_abc_17692_n1730) );
  OR2X2 OR2X2_4090 ( .A(_abc_17692_n12121), .B(_abc_17692_n12119), .Y(_abc_17692_n12122) );
  OR2X2 OR2X2_4091 ( .A(_abc_17692_n12122), .B(_abc_17692_n12115), .Y(_abc_17692_n12125) );
  OR2X2 OR2X2_4092 ( .A(_abc_17692_n12127), .B(_abc_17692_n1863_bF_buf7), .Y(_abc_17692_n12128) );
  OR2X2 OR2X2_4093 ( .A(_abc_17692_n12107), .B(_abc_17692_n12128), .Y(_abc_17692_n12129) );
  OR2X2 OR2X2_4094 ( .A(_abc_17692_n12129), .B(_abc_17692_n12090), .Y(_abc_17692_n12130) );
  OR2X2 OR2X2_4095 ( .A(_abc_17692_n12005), .B(_abc_17692_n12008), .Y(_abc_17692_n12131) );
  OR2X2 OR2X2_4096 ( .A(_abc_17692_n12134), .B(_abc_17692_n12132), .Y(_abc_17692_n12135) );
  OR2X2 OR2X2_4097 ( .A(_abc_17692_n7276), .B(_abc_17692_n12078), .Y(_abc_17692_n12136) );
  OR2X2 OR2X2_4098 ( .A(_abc_17692_n7274), .B(_abc_17692_n12077), .Y(_abc_17692_n12137) );
  OR2X2 OR2X2_4099 ( .A(_abc_17692_n12138), .B(_abc_17692_n6065), .Y(_abc_17692_n12139) );
  OR2X2 OR2X2_41 ( .A(state_3_bF_buf4), .B(state_15_bF_buf4), .Y(_abc_17692_n721) );
  OR2X2 OR2X2_410 ( .A(_abc_17692_n1730), .B(_abc_17692_n1723), .Y(_abc_17692_n1733) );
  OR2X2 OR2X2_4100 ( .A(_abc_17692_n12140), .B(workunit1_26_), .Y(_abc_17692_n12141) );
  OR2X2 OR2X2_4101 ( .A(_abc_17692_n12135), .B(_abc_17692_n12143), .Y(_abc_17692_n12146) );
  OR2X2 OR2X2_4102 ( .A(_abc_17692_n12147), .B(_abc_17692_n4047_bF_buf1), .Y(_abc_17692_n12148) );
  OR2X2 OR2X2_4103 ( .A(_abc_17692_n12152), .B(_abc_17692_n12151), .Y(_abc_17692_n12153) );
  OR2X2 OR2X2_4104 ( .A(_abc_17692_n12155), .B(_abc_17692_n12153), .Y(_abc_17692_n12156) );
  OR2X2 OR2X2_4105 ( .A(_abc_17692_n12156), .B(_abc_17692_n12142), .Y(_abc_17692_n12159) );
  OR2X2 OR2X2_4106 ( .A(_abc_17692_n11948), .B(_abc_17692_n11766), .Y(_abc_17692_n12165) );
  OR2X2 OR2X2_4107 ( .A(_abc_17692_n12169), .B(_abc_17692_n12167), .Y(_abc_17692_n12170) );
  OR2X2 OR2X2_4108 ( .A(_abc_17692_n12170), .B(_abc_17692_n12162), .Y(_abc_17692_n12173) );
  OR2X2 OR2X2_4109 ( .A(_abc_17692_n11967), .B(_abc_17692_n12032), .Y(_abc_17692_n12178) );
  OR2X2 OR2X2_411 ( .A(_abc_17692_n1735), .B(_abc_17692_n1727), .Y(_abc_17692_n1736) );
  OR2X2 OR2X2_4110 ( .A(_abc_17692_n11967), .B(_abc_17692_n11816), .Y(_abc_17692_n12181) );
  OR2X2 OR2X2_4111 ( .A(_abc_17692_n12183), .B(_abc_17692_n12180), .Y(_abc_17692_n12184) );
  OR2X2 OR2X2_4112 ( .A(_abc_17692_n12184), .B(_abc_17692_n12114), .Y(_abc_17692_n12185) );
  OR2X2 OR2X2_4113 ( .A(_abc_17692_n11909), .B(_abc_17692_n12191), .Y(_abc_17692_n12192) );
  OR2X2 OR2X2_4114 ( .A(_abc_17692_n12193), .B(_abc_17692_n12194), .Y(_abc_17692_n12195) );
  OR2X2 OR2X2_4115 ( .A(_abc_17692_n12197), .B(_abc_17692_n12098), .Y(_abc_17692_n12198) );
  OR2X2 OR2X2_4116 ( .A(_abc_17692_n12199), .B(_abc_17692_n12097), .Y(_abc_17692_n12200) );
  OR2X2 OR2X2_4117 ( .A(_abc_17692_n12202), .B(_abc_17692_n12189), .Y(_abc_17692_n12203) );
  OR2X2 OR2X2_4118 ( .A(_abc_17692_n12203), .B(_abc_17692_n12175), .Y(_abc_17692_n12204) );
  OR2X2 OR2X2_4119 ( .A(_abc_17692_n12204), .B(_abc_17692_n12161), .Y(_abc_17692_n12205) );
  OR2X2 OR2X2_412 ( .A(_abc_17692_n1726), .B(_abc_17692_n1736), .Y(sum_28__FF_INPUT) );
  OR2X2 OR2X2_4120 ( .A(_abc_17692_n12207), .B(_abc_17692_n12208), .Y(_abc_17692_n12209) );
  OR2X2 OR2X2_4121 ( .A(_abc_17692_n12206), .B(_abc_17692_n12209), .Y(_abc_17692_n12210) );
  OR2X2 OR2X2_4122 ( .A(_abc_17692_n12150), .B(_abc_17692_n12210), .Y(workunit1_26__FF_INPUT) );
  OR2X2 OR2X2_4123 ( .A(_abc_17692_n12076), .B(_abc_17692_n12071), .Y(_abc_17692_n12212) );
  OR2X2 OR2X2_4124 ( .A(_abc_17692_n12212), .B(_abc_17692_n12218), .Y(_abc_17692_n12221) );
  OR2X2 OR2X2_4125 ( .A(_abc_17692_n7381), .B(_abc_17692_n12222), .Y(_abc_17692_n12223) );
  OR2X2 OR2X2_4126 ( .A(_abc_17692_n7374), .B(_abc_17692_n12224), .Y(_abc_17692_n12225) );
  OR2X2 OR2X2_4127 ( .A(_abc_17692_n12226), .B(workunit1_27_), .Y(_abc_17692_n12227) );
  OR2X2 OR2X2_4128 ( .A(_abc_17692_n7374), .B(_abc_17692_n12222), .Y(_abc_17692_n12228) );
  OR2X2 OR2X2_4129 ( .A(_abc_17692_n7381), .B(_abc_17692_n12224), .Y(_abc_17692_n12229) );
  OR2X2 OR2X2_413 ( .A(_abc_17692_n1749), .B(_abc_17692_n1745), .Y(_abc_17692_n1750) );
  OR2X2 OR2X2_4130 ( .A(_abc_17692_n12230), .B(_abc_17692_n6242), .Y(_abc_17692_n12231) );
  OR2X2 OR2X2_4131 ( .A(_abc_17692_n12140), .B(_abc_17692_n6065), .Y(_abc_17692_n12233) );
  OR2X2 OR2X2_4132 ( .A(_abc_17692_n12144), .B(_abc_17692_n12234), .Y(_abc_17692_n12235) );
  OR2X2 OR2X2_4133 ( .A(_abc_17692_n12238), .B(_abc_17692_n12239), .Y(_abc_17692_n12240) );
  OR2X2 OR2X2_4134 ( .A(_abc_17692_n12241), .B(_abc_17692_n4047_bF_buf0), .Y(_abc_17692_n12242) );
  OR2X2 OR2X2_4135 ( .A(_abc_17692_n12242), .B(_abc_17692_n12237), .Y(_abc_17692_n12243) );
  OR2X2 OR2X2_4136 ( .A(_abc_17692_n7477), .B(_abc_17692_n12222), .Y(_abc_17692_n12244) );
  OR2X2 OR2X2_4137 ( .A(_abc_17692_n7473), .B(_abc_17692_n12224), .Y(_abc_17692_n12245) );
  OR2X2 OR2X2_4138 ( .A(_abc_17692_n7473), .B(_abc_17692_n12222), .Y(_abc_17692_n12248) );
  OR2X2 OR2X2_4139 ( .A(_abc_17692_n7477), .B(_abc_17692_n12224), .Y(_abc_17692_n12249) );
  OR2X2 OR2X2_414 ( .A(_abc_17692_n1748), .B(_abc_17692_n1744), .Y(_abc_17692_n1751) );
  OR2X2 OR2X2_4140 ( .A(_abc_17692_n12247), .B(_abc_17692_n12251), .Y(_abc_17692_n12252) );
  OR2X2 OR2X2_4141 ( .A(_abc_17692_n12257), .B(_abc_17692_n12253), .Y(_abc_17692_n12258) );
  OR2X2 OR2X2_4142 ( .A(_abc_17692_n12256), .B(_abc_17692_n12252), .Y(_abc_17692_n12259) );
  OR2X2 OR2X2_4143 ( .A(_abc_17692_n7415), .B(_abc_17692_n12222), .Y(_abc_17692_n12262) );
  OR2X2 OR2X2_4144 ( .A(_abc_17692_n7410), .B(_abc_17692_n12224), .Y(_abc_17692_n12263) );
  OR2X2 OR2X2_4145 ( .A(_abc_17692_n12264), .B(workunit1_27_), .Y(_abc_17692_n12265) );
  OR2X2 OR2X2_4146 ( .A(_abc_17692_n7410), .B(_abc_17692_n12222), .Y(_abc_17692_n12266) );
  OR2X2 OR2X2_4147 ( .A(_abc_17692_n7415), .B(_abc_17692_n12224), .Y(_abc_17692_n12267) );
  OR2X2 OR2X2_4148 ( .A(_abc_17692_n12268), .B(_abc_17692_n6242), .Y(_abc_17692_n12269) );
  OR2X2 OR2X2_4149 ( .A(_abc_17692_n12272), .B(_abc_17692_n12270), .Y(_abc_17692_n12273) );
  OR2X2 OR2X2_415 ( .A(_abc_17692_n1731), .B(_abc_17692_n1715), .Y(_abc_17692_n1755_1) );
  OR2X2 OR2X2_4150 ( .A(_abc_17692_n12271), .B(_abc_17692_n12274), .Y(_abc_17692_n12275) );
  OR2X2 OR2X2_4151 ( .A(_abc_17692_n7447), .B(_abc_17692_n12222), .Y(_abc_17692_n12278) );
  OR2X2 OR2X2_4152 ( .A(_abc_17692_n7443), .B(_abc_17692_n12224), .Y(_abc_17692_n12279) );
  OR2X2 OR2X2_4153 ( .A(_abc_17692_n7443), .B(_abc_17692_n12222), .Y(_abc_17692_n12282) );
  OR2X2 OR2X2_4154 ( .A(_abc_17692_n7447), .B(_abc_17692_n12224), .Y(_abc_17692_n12283) );
  OR2X2 OR2X2_4155 ( .A(_abc_17692_n12281), .B(_abc_17692_n12285), .Y(_abc_17692_n12286) );
  OR2X2 OR2X2_4156 ( .A(_abc_17692_n12123), .B(_abc_17692_n12113), .Y(_abc_17692_n12287) );
  OR2X2 OR2X2_4157 ( .A(_abc_17692_n12288), .B(_abc_17692_n12286), .Y(_abc_17692_n12289) );
  OR2X2 OR2X2_4158 ( .A(_abc_17692_n12284), .B(workunit1_27_), .Y(_abc_17692_n12290) );
  OR2X2 OR2X2_4159 ( .A(_abc_17692_n12280), .B(_abc_17692_n6242), .Y(_abc_17692_n12291) );
  OR2X2 OR2X2_416 ( .A(_abc_17692_n1755_1), .B(_abc_17692_n1744), .Y(_abc_17692_n1756) );
  OR2X2 OR2X2_4160 ( .A(_abc_17692_n12287), .B(_abc_17692_n12292), .Y(_abc_17692_n12293) );
  OR2X2 OR2X2_4161 ( .A(_abc_17692_n12295), .B(_abc_17692_n1863_bF_buf5), .Y(_abc_17692_n12296) );
  OR2X2 OR2X2_4162 ( .A(_abc_17692_n12277), .B(_abc_17692_n12296), .Y(_abc_17692_n12297) );
  OR2X2 OR2X2_4163 ( .A(_abc_17692_n12297), .B(_abc_17692_n12261), .Y(_abc_17692_n12298) );
  OR2X2 OR2X2_4164 ( .A(_abc_17692_n12302), .B(_abc_17692_n12240), .Y(_abc_17692_n12303) );
  OR2X2 OR2X2_4165 ( .A(_abc_17692_n12301), .B(_abc_17692_n12232), .Y(_abc_17692_n12304) );
  OR2X2 OR2X2_4166 ( .A(_abc_17692_n12311), .B(_abc_17692_n12274), .Y(_abc_17692_n12312) );
  OR2X2 OR2X2_4167 ( .A(_abc_17692_n12310), .B(_abc_17692_n12270), .Y(_abc_17692_n12313) );
  OR2X2 OR2X2_4168 ( .A(_abc_17692_n12319), .B(_abc_17692_n12286), .Y(_abc_17692_n12320) );
  OR2X2 OR2X2_4169 ( .A(_abc_17692_n12318), .B(_abc_17692_n12292), .Y(_abc_17692_n12321) );
  OR2X2 OR2X2_417 ( .A(_abc_17692_n1757), .B(_abc_17692_n1745), .Y(_abc_17692_n1758_1) );
  OR2X2 OR2X2_4170 ( .A(_abc_17692_n12325), .B(_abc_17692_n12252), .Y(_abc_17692_n12326) );
  OR2X2 OR2X2_4171 ( .A(_abc_17692_n12324), .B(_abc_17692_n12253), .Y(_abc_17692_n12327) );
  OR2X2 OR2X2_4172 ( .A(_abc_17692_n12323), .B(_abc_17692_n12329), .Y(_abc_17692_n12330) );
  OR2X2 OR2X2_4173 ( .A(_abc_17692_n12330), .B(_abc_17692_n12315), .Y(_abc_17692_n12331) );
  OR2X2 OR2X2_4174 ( .A(_abc_17692_n12331), .B(_abc_17692_n12306), .Y(_abc_17692_n12332) );
  OR2X2 OR2X2_4175 ( .A(_abc_17692_n12334), .B(_abc_17692_n12335), .Y(_abc_17692_n12336) );
  OR2X2 OR2X2_4176 ( .A(_abc_17692_n12333), .B(_abc_17692_n12336), .Y(_abc_17692_n12337) );
  OR2X2 OR2X2_4177 ( .A(_abc_17692_n12337), .B(_abc_17692_n12300), .Y(workunit1_27__FF_INPUT) );
  OR2X2 OR2X2_4178 ( .A(_abc_17692_n12340), .B(_abc_17692_n12339), .Y(_abc_17692_n12341) );
  OR2X2 OR2X2_4179 ( .A(_abc_17692_n12071), .B(_abc_17692_n12213), .Y(_abc_17692_n12342) );
  OR2X2 OR2X2_418 ( .A(_abc_17692_n1760), .B(_abc_17692_n1754), .Y(_abc_17692_n1761) );
  OR2X2 OR2X2_4180 ( .A(_abc_17692_n12076), .B(_abc_17692_n12342), .Y(_abc_17692_n12343) );
  OR2X2 OR2X2_4181 ( .A(_abc_17692_n12346), .B(_abc_17692_n12348), .Y(_abc_17692_n12349) );
  OR2X2 OR2X2_4182 ( .A(_abc_17692_n7566), .B(_abc_17692_n12350), .Y(_abc_17692_n12351) );
  OR2X2 OR2X2_4183 ( .A(_abc_17692_n7563), .B(_abc_17692_n12349), .Y(_abc_17692_n12352) );
  OR2X2 OR2X2_4184 ( .A(_abc_17692_n12354), .B(_abc_17692_n6468_1), .Y(_abc_17692_n12355) );
  OR2X2 OR2X2_4185 ( .A(_abc_17692_n12353), .B(workunit1_28_), .Y(_abc_17692_n12356) );
  OR2X2 OR2X2_4186 ( .A(_abc_17692_n11755), .B(_abc_17692_n12361), .Y(_abc_17692_n12362) );
  OR2X2 OR2X2_4187 ( .A(_abc_17692_n12239), .B(_abc_17692_n12234), .Y(_abc_17692_n12364) );
  OR2X2 OR2X2_4188 ( .A(_abc_17692_n12363), .B(_abc_17692_n12365), .Y(_abc_17692_n12366) );
  OR2X2 OR2X2_4189 ( .A(_abc_17692_n12369), .B(_abc_17692_n12358), .Y(_abc_17692_n12370) );
  OR2X2 OR2X2_419 ( .A(_abc_17692_n1753), .B(_abc_17692_n1761), .Y(sum_29__FF_INPUT) );
  OR2X2 OR2X2_4190 ( .A(_abc_17692_n12373), .B(_abc_17692_n4047_bF_buf4), .Y(_abc_17692_n12374) );
  OR2X2 OR2X2_4191 ( .A(_abc_17692_n7644), .B(_abc_17692_n12350), .Y(_abc_17692_n12375) );
  OR2X2 OR2X2_4192 ( .A(_abc_17692_n7643), .B(_abc_17692_n12349), .Y(_abc_17692_n12376) );
  OR2X2 OR2X2_4193 ( .A(_abc_17692_n12377), .B(workunit1_28_), .Y(_abc_17692_n12380) );
  OR2X2 OR2X2_4194 ( .A(_abc_17692_n12388), .B(_abc_17692_n12387), .Y(_abc_17692_n12389) );
  OR2X2 OR2X2_4195 ( .A(_abc_17692_n12386), .B(_abc_17692_n12389), .Y(_abc_17692_n12390) );
  OR2X2 OR2X2_4196 ( .A(_abc_17692_n12385), .B(_abc_17692_n12390), .Y(_abc_17692_n12391) );
  OR2X2 OR2X2_4197 ( .A(_abc_17692_n12391), .B(_abc_17692_n12382), .Y(_abc_17692_n12394) );
  OR2X2 OR2X2_4198 ( .A(_abc_17692_n7605), .B(_abc_17692_n12350), .Y(_abc_17692_n12397) );
  OR2X2 OR2X2_4199 ( .A(_abc_17692_n7603), .B(_abc_17692_n12349), .Y(_abc_17692_n12398) );
  OR2X2 OR2X2_42 ( .A(_abc_17692_n725_bF_buf7), .B(_auto_iopadmap_cc_313_execute_30065_0_), .Y(_abc_17692_n726) );
  OR2X2 OR2X2_420 ( .A(_abc_17692_n1766), .B(_abc_17692_n1763), .Y(_abc_17692_n1767) );
  OR2X2 OR2X2_4200 ( .A(_abc_17692_n12400), .B(_abc_17692_n6468_1), .Y(_abc_17692_n12401) );
  OR2X2 OR2X2_4201 ( .A(_abc_17692_n12399), .B(workunit1_28_), .Y(_abc_17692_n12402) );
  OR2X2 OR2X2_4202 ( .A(_abc_17692_n12100), .B(_abc_17692_n11980), .Y(_abc_17692_n12409) );
  OR2X2 OR2X2_4203 ( .A(_abc_17692_n12412), .B(_abc_17692_n12251), .Y(_abc_17692_n12413) );
  OR2X2 OR2X2_4204 ( .A(_abc_17692_n12413), .B(_abc_17692_n12411), .Y(_abc_17692_n12414) );
  OR2X2 OR2X2_4205 ( .A(_abc_17692_n12408), .B(_abc_17692_n12414), .Y(_abc_17692_n12415) );
  OR2X2 OR2X2_4206 ( .A(_abc_17692_n12415), .B(_abc_17692_n12404), .Y(_abc_17692_n12416) );
  OR2X2 OR2X2_4207 ( .A(_abc_17692_n7685), .B(_abc_17692_n12350), .Y(_abc_17692_n12421) );
  OR2X2 OR2X2_4208 ( .A(_abc_17692_n7683), .B(_abc_17692_n12349), .Y(_abc_17692_n12422) );
  OR2X2 OR2X2_4209 ( .A(_abc_17692_n12424), .B(_abc_17692_n6468_1), .Y(_abc_17692_n12425) );
  OR2X2 OR2X2_421 ( .A(_abc_17692_n1748), .B(_abc_17692_n1771), .Y(_abc_17692_n1772) );
  OR2X2 OR2X2_4210 ( .A(_abc_17692_n12423), .B(workunit1_28_), .Y(_abc_17692_n12426) );
  OR2X2 OR2X2_4211 ( .A(_abc_17692_n12286), .B(_abc_17692_n12114), .Y(_abc_17692_n12430) );
  OR2X2 OR2X2_4212 ( .A(_abc_17692_n12430), .B(_abc_17692_n12429), .Y(_abc_17692_n12431) );
  OR2X2 OR2X2_4213 ( .A(_abc_17692_n11826), .B(_abc_17692_n12431), .Y(_abc_17692_n12432) );
  OR2X2 OR2X2_4214 ( .A(_abc_17692_n12430), .B(_abc_17692_n12118), .Y(_abc_17692_n12433) );
  OR2X2 OR2X2_4215 ( .A(_abc_17692_n12285), .B(_abc_17692_n12113), .Y(_abc_17692_n12434) );
  OR2X2 OR2X2_4216 ( .A(_abc_17692_n12439), .B(_abc_17692_n12428), .Y(_abc_17692_n12442) );
  OR2X2 OR2X2_4217 ( .A(_abc_17692_n12444), .B(_abc_17692_n1863_bF_buf3), .Y(_abc_17692_n12445) );
  OR2X2 OR2X2_4218 ( .A(_abc_17692_n12445), .B(_abc_17692_n12420), .Y(_abc_17692_n12446) );
  OR2X2 OR2X2_4219 ( .A(_abc_17692_n12446), .B(_abc_17692_n12396), .Y(_abc_17692_n12447) );
  OR2X2 OR2X2_422 ( .A(_abc_17692_n1774), .B(_abc_17692_n1768), .Y(_abc_17692_n1775_1) );
  OR2X2 OR2X2_4220 ( .A(_abc_17692_n12456), .B(_abc_17692_n12454), .Y(_abc_17692_n12457) );
  OR2X2 OR2X2_4221 ( .A(_abc_17692_n12457), .B(_abc_17692_n12453), .Y(_abc_17692_n12458) );
  OR2X2 OR2X2_4222 ( .A(_abc_17692_n12452), .B(_abc_17692_n12458), .Y(_abc_17692_n12459) );
  OR2X2 OR2X2_4223 ( .A(_abc_17692_n12459), .B(_abc_17692_n12357), .Y(_abc_17692_n12462) );
  OR2X2 OR2X2_4224 ( .A(_abc_17692_n12270), .B(_abc_17692_n12085), .Y(_abc_17692_n12466) );
  OR2X2 OR2X2_4225 ( .A(_abc_17692_n12466), .B(_abc_17692_n12465), .Y(_abc_17692_n12467) );
  OR2X2 OR2X2_4226 ( .A(_abc_17692_n11870), .B(_abc_17692_n12467), .Y(_abc_17692_n12468) );
  OR2X2 OR2X2_4227 ( .A(_abc_17692_n12466), .B(_abc_17692_n12166), .Y(_abc_17692_n12469) );
  OR2X2 OR2X2_4228 ( .A(_abc_17692_n12270), .B(_abc_17692_n12309), .Y(_abc_17692_n12472) );
  OR2X2 OR2X2_4229 ( .A(_abc_17692_n12476), .B(_abc_17692_n12381), .Y(_abc_17692_n12479) );
  OR2X2 OR2X2_423 ( .A(_abc_17692_n1773), .B(_abc_17692_n1767), .Y(_abc_17692_n1776) );
  OR2X2 OR2X2_4230 ( .A(_abc_17692_n12292), .B(_abc_17692_n12115), .Y(_abc_17692_n12482) );
  OR2X2 OR2X2_4231 ( .A(_abc_17692_n12482), .B(_abc_17692_n12181), .Y(_abc_17692_n12483) );
  OR2X2 OR2X2_4232 ( .A(_abc_17692_n11891), .B(_abc_17692_n12483), .Y(_abc_17692_n12484) );
  OR2X2 OR2X2_4233 ( .A(_abc_17692_n12179), .B(_abc_17692_n12482), .Y(_abc_17692_n12485) );
  OR2X2 OR2X2_4234 ( .A(_abc_17692_n12292), .B(_abc_17692_n12317), .Y(_abc_17692_n12488) );
  OR2X2 OR2X2_4235 ( .A(_abc_17692_n12492), .B(_abc_17692_n12427), .Y(_abc_17692_n12493) );
  OR2X2 OR2X2_4236 ( .A(_abc_17692_n12504), .B(_abc_17692_n12502), .Y(_abc_17692_n12505) );
  OR2X2 OR2X2_4237 ( .A(_abc_17692_n12505), .B(_abc_17692_n12501), .Y(_abc_17692_n12506) );
  OR2X2 OR2X2_4238 ( .A(_abc_17692_n12500), .B(_abc_17692_n12506), .Y(_abc_17692_n12507) );
  OR2X2 OR2X2_4239 ( .A(_abc_17692_n12507), .B(_abc_17692_n12403), .Y(_abc_17692_n12510) );
  OR2X2 OR2X2_424 ( .A(_abc_17692_n1779), .B(_abc_17692_n1742), .Y(_abc_17692_n1780) );
  OR2X2 OR2X2_4240 ( .A(_abc_17692_n12497), .B(_abc_17692_n12512), .Y(_abc_17692_n12513) );
  OR2X2 OR2X2_4241 ( .A(_abc_17692_n12513), .B(_abc_17692_n12481), .Y(_abc_17692_n12514) );
  OR2X2 OR2X2_4242 ( .A(_abc_17692_n12514), .B(_abc_17692_n12464), .Y(_abc_17692_n12515) );
  OR2X2 OR2X2_4243 ( .A(_abc_17692_n12517), .B(_abc_17692_n12518), .Y(_abc_17692_n12519) );
  OR2X2 OR2X2_4244 ( .A(_abc_17692_n12516), .B(_abc_17692_n12519), .Y(_abc_17692_n12520) );
  OR2X2 OR2X2_4245 ( .A(_abc_17692_n12520), .B(_abc_17692_n12449), .Y(workunit1_28__FF_INPUT) );
  OR2X2 OR2X2_4246 ( .A(_abc_17692_n12348), .B(_abc_17692_n12339), .Y(_abc_17692_n12522) );
  OR2X2 OR2X2_4247 ( .A(_abc_17692_n12522), .B(_abc_17692_n12528), .Y(_abc_17692_n12531) );
  OR2X2 OR2X2_4248 ( .A(_abc_17692_n7898), .B(_abc_17692_n12532), .Y(_abc_17692_n12533) );
  OR2X2 OR2X2_4249 ( .A(_abc_17692_n7901), .B(_abc_17692_n12534), .Y(_abc_17692_n12535) );
  OR2X2 OR2X2_425 ( .A(_abc_17692_n1780), .B(_abc_17692_n1767), .Y(_abc_17692_n1781) );
  OR2X2 OR2X2_4250 ( .A(_abc_17692_n7901), .B(_abc_17692_n12532), .Y(_abc_17692_n12538) );
  OR2X2 OR2X2_4251 ( .A(_abc_17692_n7898), .B(_abc_17692_n12534), .Y(_abc_17692_n12539) );
  OR2X2 OR2X2_4252 ( .A(_abc_17692_n12537), .B(_abc_17692_n12541), .Y(_abc_17692_n12542) );
  OR2X2 OR2X2_4253 ( .A(_abc_17692_n12353), .B(_abc_17692_n6468_1), .Y(_abc_17692_n12543) );
  OR2X2 OR2X2_4254 ( .A(_abc_17692_n12540), .B(workunit1_29_), .Y(_abc_17692_n12547) );
  OR2X2 OR2X2_4255 ( .A(_abc_17692_n12536), .B(_abc_17692_n6659_1), .Y(_abc_17692_n12548) );
  OR2X2 OR2X2_4256 ( .A(_abc_17692_n12550), .B(_abc_17692_n4047_bF_buf3), .Y(_abc_17692_n12551) );
  OR2X2 OR2X2_4257 ( .A(_abc_17692_n12551), .B(_abc_17692_n12546), .Y(_abc_17692_n12552) );
  OR2X2 OR2X2_4258 ( .A(_abc_17692_n7803), .B(_abc_17692_n12532), .Y(_abc_17692_n12553) );
  OR2X2 OR2X2_4259 ( .A(_abc_17692_n7808), .B(_abc_17692_n12534), .Y(_abc_17692_n12554) );
  OR2X2 OR2X2_426 ( .A(_abc_17692_n1786), .B(state_8_bF_buf1), .Y(_abc_17692_n1787) );
  OR2X2 OR2X2_4260 ( .A(_abc_17692_n12555), .B(workunit1_29_), .Y(_abc_17692_n12556) );
  OR2X2 OR2X2_4261 ( .A(_abc_17692_n7808), .B(_abc_17692_n12532), .Y(_abc_17692_n12557) );
  OR2X2 OR2X2_4262 ( .A(_abc_17692_n7803), .B(_abc_17692_n12534), .Y(_abc_17692_n12558) );
  OR2X2 OR2X2_4263 ( .A(_abc_17692_n12559), .B(_abc_17692_n6659_1), .Y(_abc_17692_n12560) );
  OR2X2 OR2X2_4264 ( .A(_abc_17692_n12392), .B(_abc_17692_n12564), .Y(_abc_17692_n12565) );
  OR2X2 OR2X2_4265 ( .A(_abc_17692_n12566), .B(_abc_17692_n12562), .Y(_abc_17692_n12567) );
  OR2X2 OR2X2_4266 ( .A(_abc_17692_n12565), .B(_abc_17692_n12561), .Y(_abc_17692_n12568) );
  OR2X2 OR2X2_4267 ( .A(_abc_17692_n7834), .B(_abc_17692_n12532), .Y(_abc_17692_n12571) );
  OR2X2 OR2X2_4268 ( .A(_abc_17692_n7838), .B(_abc_17692_n12534), .Y(_abc_17692_n12572) );
  OR2X2 OR2X2_4269 ( .A(_abc_17692_n7838), .B(_abc_17692_n12532), .Y(_abc_17692_n12575) );
  OR2X2 OR2X2_427 ( .A(_abc_17692_n1785), .B(_abc_17692_n1787), .Y(_abc_17692_n1788_1) );
  OR2X2 OR2X2_4270 ( .A(_abc_17692_n7834), .B(_abc_17692_n12534), .Y(_abc_17692_n12576) );
  OR2X2 OR2X2_4271 ( .A(_abc_17692_n12574), .B(_abc_17692_n12578), .Y(_abc_17692_n12579) );
  OR2X2 OR2X2_4272 ( .A(_abc_17692_n12582), .B(_abc_17692_n12579), .Y(_abc_17692_n12583) );
  OR2X2 OR2X2_4273 ( .A(_abc_17692_n12585), .B(_abc_17692_n12584), .Y(_abc_17692_n12586) );
  OR2X2 OR2X2_4274 ( .A(_abc_17692_n7865), .B(_abc_17692_n12532), .Y(_abc_17692_n12589) );
  OR2X2 OR2X2_4275 ( .A(_abc_17692_n7869), .B(_abc_17692_n12534), .Y(_abc_17692_n12590) );
  OR2X2 OR2X2_4276 ( .A(_abc_17692_n7869), .B(_abc_17692_n12532), .Y(_abc_17692_n12593) );
  OR2X2 OR2X2_4277 ( .A(_abc_17692_n7865), .B(_abc_17692_n12534), .Y(_abc_17692_n12594) );
  OR2X2 OR2X2_4278 ( .A(_abc_17692_n12592), .B(_abc_17692_n12596), .Y(_abc_17692_n12597) );
  OR2X2 OR2X2_4279 ( .A(_abc_17692_n12423), .B(_abc_17692_n6468_1), .Y(_abc_17692_n12598) );
  OR2X2 OR2X2_428 ( .A(_abc_17692_n1778), .B(_abc_17692_n1788_1), .Y(sum_30__FF_INPUT) );
  OR2X2 OR2X2_4280 ( .A(_abc_17692_n12440), .B(_abc_17692_n12599), .Y(_abc_17692_n12600) );
  OR2X2 OR2X2_4281 ( .A(_abc_17692_n12601), .B(_abc_17692_n12597), .Y(_abc_17692_n12602) );
  OR2X2 OR2X2_4282 ( .A(_abc_17692_n12595), .B(workunit1_29_), .Y(_abc_17692_n12603) );
  OR2X2 OR2X2_4283 ( .A(_abc_17692_n12591), .B(_abc_17692_n6659_1), .Y(_abc_17692_n12604) );
  OR2X2 OR2X2_4284 ( .A(_abc_17692_n12600), .B(_abc_17692_n12605), .Y(_abc_17692_n12606) );
  OR2X2 OR2X2_4285 ( .A(_abc_17692_n12608), .B(_abc_17692_n1863_bF_buf1), .Y(_abc_17692_n12609) );
  OR2X2 OR2X2_4286 ( .A(_abc_17692_n12609), .B(_abc_17692_n12588), .Y(_abc_17692_n12610) );
  OR2X2 OR2X2_4287 ( .A(_abc_17692_n12610), .B(_abc_17692_n12570), .Y(_abc_17692_n12611) );
  OR2X2 OR2X2_4288 ( .A(_abc_17692_n12615), .B(_abc_17692_n12542), .Y(_abc_17692_n12616) );
  OR2X2 OR2X2_4289 ( .A(_abc_17692_n12614), .B(_abc_17692_n12549), .Y(_abc_17692_n12617) );
  OR2X2 OR2X2_429 ( .A(_abc_17692_n1790), .B(sum_31_), .Y(_abc_17692_n1791) );
  OR2X2 OR2X2_4290 ( .A(_abc_17692_n12621), .B(_abc_17692_n12562), .Y(_abc_17692_n12622) );
  OR2X2 OR2X2_4291 ( .A(_abc_17692_n12620), .B(_abc_17692_n12561), .Y(_abc_17692_n12623) );
  OR2X2 OR2X2_4292 ( .A(_abc_17692_n12626), .B(_abc_17692_n12584), .Y(_abc_17692_n12627) );
  OR2X2 OR2X2_4293 ( .A(_abc_17692_n12628), .B(_abc_17692_n12579), .Y(_abc_17692_n12629) );
  OR2X2 OR2X2_4294 ( .A(_abc_17692_n12633), .B(_abc_17692_n12597), .Y(_abc_17692_n12634) );
  OR2X2 OR2X2_4295 ( .A(_abc_17692_n12632), .B(_abc_17692_n12605), .Y(_abc_17692_n12635) );
  OR2X2 OR2X2_4296 ( .A(_abc_17692_n12631), .B(_abc_17692_n12637), .Y(_abc_17692_n12638) );
  OR2X2 OR2X2_4297 ( .A(_abc_17692_n12638), .B(_abc_17692_n12625), .Y(_abc_17692_n12639) );
  OR2X2 OR2X2_4298 ( .A(_abc_17692_n12639), .B(_abc_17692_n12619), .Y(_abc_17692_n12640) );
  OR2X2 OR2X2_4299 ( .A(_abc_17692_n12642), .B(_abc_17692_n12643), .Y(_abc_17692_n12644) );
  OR2X2 OR2X2_43 ( .A(_abc_17692_n727_bF_buf7), .B(workunit2_0_), .Y(_abc_17692_n728) );
  OR2X2 OR2X2_430 ( .A(_abc_17692_n1792), .B(delta_31_), .Y(_abc_17692_n1793) );
  OR2X2 OR2X2_4300 ( .A(_abc_17692_n12641), .B(_abc_17692_n12644), .Y(_abc_17692_n12645) );
  OR2X2 OR2X2_4301 ( .A(_abc_17692_n12645), .B(_abc_17692_n12613), .Y(workunit1_29__FF_INPUT) );
  OR2X2 OR2X2_4302 ( .A(_abc_17692_n12649), .B(_abc_17692_n12648), .Y(_abc_17692_n12650) );
  OR2X2 OR2X2_4303 ( .A(_abc_17692_n12522), .B(_abc_17692_n12523), .Y(_abc_17692_n12652) );
  OR2X2 OR2X2_4304 ( .A(_abc_17692_n12653), .B(_abc_17692_n12651), .Y(_abc_17692_n12656) );
  OR2X2 OR2X2_4305 ( .A(_abc_17692_n12647), .B(_abc_17692_n12657), .Y(_abc_17692_n12658) );
  OR2X2 OR2X2_4306 ( .A(_abc_17692_n7990), .B(_abc_17692_n12659), .Y(_abc_17692_n12660) );
  OR2X2 OR2X2_4307 ( .A(_abc_17692_n12661), .B(_abc_17692_n6956), .Y(_abc_17692_n12662) );
  OR2X2 OR2X2_4308 ( .A(_abc_17692_n7990), .B(_abc_17692_n12657), .Y(_abc_17692_n12663) );
  OR2X2 OR2X2_4309 ( .A(_abc_17692_n12647), .B(_abc_17692_n12659), .Y(_abc_17692_n12664) );
  OR2X2 OR2X2_431 ( .A(_abc_17692_n1798), .B(_abc_17692_n1795), .Y(_abc_17692_n1799) );
  OR2X2 OR2X2_4310 ( .A(_abc_17692_n12665), .B(workunit1_30_), .Y(_abc_17692_n12666) );
  OR2X2 OR2X2_4311 ( .A(_abc_17692_n12671), .B(_abc_17692_n12578), .Y(_abc_17692_n12672) );
  OR2X2 OR2X2_4312 ( .A(_abc_17692_n12670), .B(_abc_17692_n12672), .Y(_abc_17692_n12673) );
  OR2X2 OR2X2_4313 ( .A(_abc_17692_n12673), .B(_abc_17692_n12668), .Y(_abc_17692_n12674) );
  OR2X2 OR2X2_4314 ( .A(_abc_17692_n12680), .B(_abc_17692_n12679), .Y(_abc_17692_n12681) );
  OR2X2 OR2X2_4315 ( .A(_abc_17692_n12682), .B(workunit1_30_), .Y(_abc_17692_n12683) );
  OR2X2 OR2X2_4316 ( .A(_abc_17692_n12681), .B(_abc_17692_n6956), .Y(_abc_17692_n12684) );
  OR2X2 OR2X2_4317 ( .A(_abc_17692_n12689), .B(_abc_17692_n12688), .Y(_abc_17692_n12690) );
  OR2X2 OR2X2_4318 ( .A(_abc_17692_n12687), .B(_abc_17692_n12690), .Y(_abc_17692_n12691) );
  OR2X2 OR2X2_4319 ( .A(_abc_17692_n12691), .B(_abc_17692_n12685), .Y(_abc_17692_n12694) );
  OR2X2 OR2X2_432 ( .A(_abc_17692_n1797), .B(_abc_17692_n1794), .Y(_abc_17692_n1800) );
  OR2X2 OR2X2_4320 ( .A(_abc_17692_n8058), .B(_abc_17692_n12657), .Y(_abc_17692_n12697) );
  OR2X2 OR2X2_4321 ( .A(_abc_17692_n8056), .B(_abc_17692_n12659), .Y(_abc_17692_n12698) );
  OR2X2 OR2X2_4322 ( .A(_abc_17692_n12699), .B(workunit1_30_), .Y(_abc_17692_n12700) );
  OR2X2 OR2X2_4323 ( .A(_abc_17692_n8056), .B(_abc_17692_n12657), .Y(_abc_17692_n12701) );
  OR2X2 OR2X2_4324 ( .A(_abc_17692_n8058), .B(_abc_17692_n12659), .Y(_abc_17692_n12702) );
  OR2X2 OR2X2_4325 ( .A(_abc_17692_n12703), .B(_abc_17692_n6956), .Y(_abc_17692_n12704) );
  OR2X2 OR2X2_4326 ( .A(_abc_17692_n12597), .B(_abc_17692_n12427), .Y(_abc_17692_n12706) );
  OR2X2 OR2X2_4327 ( .A(_abc_17692_n12438), .B(_abc_17692_n12706), .Y(_abc_17692_n12707) );
  OR2X2 OR2X2_4328 ( .A(_abc_17692_n12592), .B(_abc_17692_n12598), .Y(_abc_17692_n12708) );
  OR2X2 OR2X2_4329 ( .A(_abc_17692_n12711), .B(_abc_17692_n12705), .Y(_abc_17692_n12712) );
  OR2X2 OR2X2_433 ( .A(_abc_17692_n1782), .B(_abc_17692_n1803), .Y(_abc_17692_n1804_1) );
  OR2X2 OR2X2_4330 ( .A(_abc_17692_n12699), .B(_abc_17692_n6956), .Y(_abc_17692_n12713) );
  OR2X2 OR2X2_4331 ( .A(_abc_17692_n12703), .B(workunit1_30_), .Y(_abc_17692_n12714) );
  OR2X2 OR2X2_4332 ( .A(_abc_17692_n12710), .B(_abc_17692_n12715), .Y(_abc_17692_n12716) );
  OR2X2 OR2X2_4333 ( .A(_abc_17692_n12718), .B(_abc_17692_n1863_bF_buf10), .Y(_abc_17692_n12719) );
  OR2X2 OR2X2_4334 ( .A(_abc_17692_n12696), .B(_abc_17692_n12719), .Y(_abc_17692_n12720) );
  OR2X2 OR2X2_4335 ( .A(_abc_17692_n12720), .B(_abc_17692_n12678), .Y(_abc_17692_n12721) );
  OR2X2 OR2X2_4336 ( .A(_abc_17692_n8094), .B(_abc_17692_n12657), .Y(_abc_17692_n12722) );
  OR2X2 OR2X2_4337 ( .A(_abc_17692_n8096), .B(_abc_17692_n12659), .Y(_abc_17692_n12723) );
  OR2X2 OR2X2_4338 ( .A(_abc_17692_n12725), .B(_abc_17692_n6956), .Y(_abc_17692_n12726) );
  OR2X2 OR2X2_4339 ( .A(_abc_17692_n12724), .B(workunit1_30_), .Y(_abc_17692_n12727) );
  OR2X2 OR2X2_434 ( .A(_abc_17692_n1805), .B(_abc_17692_n1795), .Y(_abc_17692_n1806) );
  OR2X2 OR2X2_4340 ( .A(_abc_17692_n12368), .B(_abc_17692_n12730), .Y(_abc_17692_n12731) );
  OR2X2 OR2X2_4341 ( .A(_abc_17692_n12732), .B(_abc_17692_n12537), .Y(_abc_17692_n12733) );
  OR2X2 OR2X2_4342 ( .A(_abc_17692_n12735), .B(_abc_17692_n12728), .Y(_abc_17692_n12736) );
  OR2X2 OR2X2_4343 ( .A(_abc_17692_n12724), .B(_abc_17692_n6956), .Y(_abc_17692_n12737) );
  OR2X2 OR2X2_4344 ( .A(_abc_17692_n12725), .B(workunit1_30_), .Y(_abc_17692_n12738) );
  OR2X2 OR2X2_4345 ( .A(_abc_17692_n12734), .B(_abc_17692_n12739), .Y(_abc_17692_n12740) );
  OR2X2 OR2X2_4346 ( .A(_abc_17692_n12741), .B(_abc_17692_n4047_bF_buf2), .Y(_abc_17692_n12742) );
  OR2X2 OR2X2_4347 ( .A(_abc_17692_n11040), .B(_abc_17692_n12746), .Y(_abc_17692_n12747) );
  OR2X2 OR2X2_4348 ( .A(_abc_17692_n11666), .B(_abc_17692_n11502), .Y(_abc_17692_n12751) );
  OR2X2 OR2X2_4349 ( .A(_abc_17692_n12751), .B(_abc_17692_n11519), .Y(_abc_17692_n12752) );
  OR2X2 OR2X2_435 ( .A(_abc_17692_n1804_1), .B(_abc_17692_n1794), .Y(_abc_17692_n1807) );
  OR2X2 OR2X2_4350 ( .A(_abc_17692_n12750), .B(_abc_17692_n12752), .Y(_abc_17692_n12753) );
  OR2X2 OR2X2_4351 ( .A(_abc_17692_n12751), .B(_abc_17692_n12754), .Y(_abc_17692_n12755) );
  OR2X2 OR2X2_4352 ( .A(_abc_17692_n11666), .B(_abc_17692_n11499), .Y(_abc_17692_n12757) );
  OR2X2 OR2X2_4353 ( .A(_abc_17692_n12752), .B(_abc_17692_n12762), .Y(_abc_17692_n12763) );
  OR2X2 OR2X2_4354 ( .A(_abc_17692_n12763), .B(_abc_17692_n12761), .Y(_abc_17692_n12764) );
  OR2X2 OR2X2_4355 ( .A(_abc_17692_n12232), .B(_abc_17692_n12143), .Y(_abc_17692_n12767) );
  OR2X2 OR2X2_4356 ( .A(_abc_17692_n12767), .B(_abc_17692_n12766), .Y(_abc_17692_n12768) );
  OR2X2 OR2X2_4357 ( .A(_abc_17692_n12765), .B(_abc_17692_n12768), .Y(_abc_17692_n12769) );
  OR2X2 OR2X2_4358 ( .A(_abc_17692_n12772), .B(_abc_17692_n12767), .Y(_abc_17692_n12773) );
  OR2X2 OR2X2_4359 ( .A(_abc_17692_n12232), .B(_abc_17692_n12139), .Y(_abc_17692_n12775) );
  OR2X2 OR2X2_436 ( .A(_abc_17692_n1810), .B(state_8_bF_buf0), .Y(_abc_17692_n1811) );
  OR2X2 OR2X2_4360 ( .A(_abc_17692_n12549), .B(_abc_17692_n12358), .Y(_abc_17692_n12779) );
  OR2X2 OR2X2_4361 ( .A(_abc_17692_n12778), .B(_abc_17692_n12779), .Y(_abc_17692_n12780) );
  OR2X2 OR2X2_4362 ( .A(_abc_17692_n12549), .B(_abc_17692_n12355), .Y(_abc_17692_n12783) );
  OR2X2 OR2X2_4363 ( .A(_abc_17692_n12785), .B(_abc_17692_n12728), .Y(_abc_17692_n12786) );
  OR2X2 OR2X2_4364 ( .A(_abc_17692_n12790), .B(_abc_17692_n12781), .Y(_abc_17692_n12791) );
  OR2X2 OR2X2_4365 ( .A(_abc_17692_n12788), .B(_abc_17692_n12791), .Y(_abc_17692_n12792) );
  OR2X2 OR2X2_4366 ( .A(_abc_17692_n12792), .B(_abc_17692_n12739), .Y(_abc_17692_n12793) );
  OR2X2 OR2X2_4367 ( .A(_abc_17692_n12561), .B(_abc_17692_n12382), .Y(_abc_17692_n12797) );
  OR2X2 OR2X2_4368 ( .A(_abc_17692_n12475), .B(_abc_17692_n12797), .Y(_abc_17692_n12798) );
  OR2X2 OR2X2_4369 ( .A(_abc_17692_n12561), .B(_abc_17692_n12379), .Y(_abc_17692_n12801) );
  OR2X2 OR2X2_437 ( .A(_abc_17692_n1809), .B(_abc_17692_n1811), .Y(_abc_17692_n1812) );
  OR2X2 OR2X2_4370 ( .A(_abc_17692_n12804), .B(_abc_17692_n12796), .Y(_abc_17692_n12805) );
  OR2X2 OR2X2_4371 ( .A(_abc_17692_n12803), .B(_abc_17692_n12685), .Y(_abc_17692_n12806) );
  OR2X2 OR2X2_4372 ( .A(_abc_17692_n12605), .B(_abc_17692_n12428), .Y(_abc_17692_n12809) );
  OR2X2 OR2X2_4373 ( .A(_abc_17692_n12491), .B(_abc_17692_n12809), .Y(_abc_17692_n12810) );
  OR2X2 OR2X2_4374 ( .A(_abc_17692_n12605), .B(_abc_17692_n12425), .Y(_abc_17692_n12813) );
  OR2X2 OR2X2_4375 ( .A(_abc_17692_n12815), .B(_abc_17692_n12705), .Y(_abc_17692_n12816) );
  OR2X2 OR2X2_4376 ( .A(_abc_17692_n12817), .B(_abc_17692_n12715), .Y(_abc_17692_n12818) );
  OR2X2 OR2X2_4377 ( .A(_abc_17692_n12825), .B(_abc_17692_n12823), .Y(_abc_17692_n12826) );
  OR2X2 OR2X2_4378 ( .A(_abc_17692_n12822), .B(_abc_17692_n12826), .Y(_abc_17692_n12827) );
  OR2X2 OR2X2_4379 ( .A(_abc_17692_n12827), .B(_abc_17692_n12667), .Y(_abc_17692_n12830) );
  OR2X2 OR2X2_438 ( .A(_abc_17692_n1802), .B(_abc_17692_n1812), .Y(sum_31__FF_INPUT) );
  OR2X2 OR2X2_4380 ( .A(_abc_17692_n12820), .B(_abc_17692_n12832), .Y(_abc_17692_n12833) );
  OR2X2 OR2X2_4381 ( .A(_abc_17692_n12833), .B(_abc_17692_n12808), .Y(_abc_17692_n12834) );
  OR2X2 OR2X2_4382 ( .A(_abc_17692_n12834), .B(_abc_17692_n12795), .Y(_abc_17692_n12835) );
  OR2X2 OR2X2_4383 ( .A(_abc_17692_n12837), .B(_abc_17692_n12838), .Y(_abc_17692_n12839) );
  OR2X2 OR2X2_4384 ( .A(_abc_17692_n12836), .B(_abc_17692_n12839), .Y(_abc_17692_n12840) );
  OR2X2 OR2X2_4385 ( .A(_abc_17692_n12744), .B(_abc_17692_n12840), .Y(workunit1_30__FF_INPUT) );
  OR2X2 OR2X2_4386 ( .A(_abc_17692_n12654), .B(_abc_17692_n12648), .Y(_abc_17692_n12844) );
  OR2X2 OR2X2_4387 ( .A(_abc_17692_n12845), .B(_abc_17692_n12846), .Y(_abc_17692_n12847) );
  OR2X2 OR2X2_4388 ( .A(_abc_17692_n12851), .B(_abc_17692_n12848), .Y(_abc_17692_n12852) );
  OR2X2 OR2X2_4389 ( .A(_abc_17692_n12852), .B(_abc_17692_n7135), .Y(_abc_17692_n12855) );
  OR2X2 OR2X2_439 ( .A(_abc_17692_n1818), .B(_abc_17692_n1815_1), .Y(_abc_17692_n1819) );
  OR2X2 OR2X2_4390 ( .A(_abc_17692_n12858), .B(_abc_17692_n12859), .Y(_abc_17692_n12860) );
  OR2X2 OR2X2_4391 ( .A(_abc_17692_n12863), .B(_abc_17692_n4047_bF_buf1), .Y(_abc_17692_n12864) );
  OR2X2 OR2X2_4392 ( .A(_abc_17692_n12864), .B(_abc_17692_n12861), .Y(_abc_17692_n12865) );
  OR2X2 OR2X2_4393 ( .A(_abc_17692_n12692), .B(_abc_17692_n12866), .Y(_abc_17692_n12867) );
  OR2X2 OR2X2_4394 ( .A(_abc_17692_n8238), .B(_abc_17692_n12856), .Y(_abc_17692_n12869) );
  OR2X2 OR2X2_4395 ( .A(_abc_17692_n8240), .B(_abc_17692_n12857), .Y(_abc_17692_n12870) );
  OR2X2 OR2X2_4396 ( .A(_abc_17692_n12868), .B(_abc_17692_n12872), .Y(_abc_17692_n12873) );
  OR2X2 OR2X2_4397 ( .A(_abc_17692_n12867), .B(_abc_17692_n12871), .Y(_abc_17692_n12874) );
  OR2X2 OR2X2_4398 ( .A(_abc_17692_n12675), .B(_abc_17692_n12877), .Y(_abc_17692_n12878) );
  OR2X2 OR2X2_4399 ( .A(_abc_17692_n12857), .B(_abc_17692_n8261), .Y(_abc_17692_n12880) );
  OR2X2 OR2X2_44 ( .A(_abc_17692_n725_bF_buf5), .B(_auto_iopadmap_cc_313_execute_30065_1_), .Y(_abc_17692_n730_1) );
  OR2X2 OR2X2_440 ( .A(sum_0_), .B(\key_in[0] ), .Y(_abc_17692_n1822) );
  OR2X2 OR2X2_4400 ( .A(_abc_17692_n8263), .B(_abc_17692_n12856), .Y(_abc_17692_n12881) );
  OR2X2 OR2X2_4401 ( .A(_abc_17692_n12879), .B(_abc_17692_n12882), .Y(_abc_17692_n12883) );
  OR2X2 OR2X2_4402 ( .A(_abc_17692_n12878), .B(_abc_17692_n12884), .Y(_abc_17692_n12885) );
  OR2X2 OR2X2_4403 ( .A(_abc_17692_n12856), .B(_abc_17692_n8284), .Y(_abc_17692_n12890) );
  OR2X2 OR2X2_4404 ( .A(_abc_17692_n12857), .B(_abc_17692_n8286), .Y(_abc_17692_n12891) );
  OR2X2 OR2X2_4405 ( .A(_abc_17692_n12889), .B(_abc_17692_n12892), .Y(_abc_17692_n12893) );
  OR2X2 OR2X2_4406 ( .A(_abc_17692_n12888), .B(_abc_17692_n12894), .Y(_abc_17692_n12895) );
  OR2X2 OR2X2_4407 ( .A(_abc_17692_n12897), .B(_abc_17692_n1863_bF_buf8), .Y(_abc_17692_n12898) );
  OR2X2 OR2X2_4408 ( .A(_abc_17692_n12898), .B(_abc_17692_n12887), .Y(_abc_17692_n12899) );
  OR2X2 OR2X2_4409 ( .A(_abc_17692_n12899), .B(_abc_17692_n12876), .Y(_abc_17692_n12900) );
  OR2X2 OR2X2_441 ( .A(_abc_17692_n1827), .B(_abc_17692_n1825), .Y(_abc_17692_n1828) );
  OR2X2 OR2X2_4410 ( .A(_abc_17692_n12904), .B(_abc_17692_n12903), .Y(_abc_17692_n12905) );
  OR2X2 OR2X2_4411 ( .A(_abc_17692_n12905), .B(_abc_17692_n12860), .Y(_abc_17692_n12906) );
  OR2X2 OR2X2_4412 ( .A(_abc_17692_n12907), .B(_abc_17692_n12862), .Y(_abc_17692_n12908) );
  OR2X2 OR2X2_4413 ( .A(_abc_17692_n12914), .B(_abc_17692_n12872), .Y(_abc_17692_n12915) );
  OR2X2 OR2X2_4414 ( .A(_abc_17692_n12913), .B(_abc_17692_n12871), .Y(_abc_17692_n12916) );
  OR2X2 OR2X2_4415 ( .A(_abc_17692_n12920), .B(_abc_17692_n12894), .Y(_abc_17692_n12921) );
  OR2X2 OR2X2_4416 ( .A(_abc_17692_n12919), .B(_abc_17692_n12892), .Y(_abc_17692_n12922) );
  OR2X2 OR2X2_4417 ( .A(_abc_17692_n12828), .B(_abc_17692_n12925), .Y(_abc_17692_n12926) );
  OR2X2 OR2X2_4418 ( .A(_abc_17692_n12927), .B(_abc_17692_n12884), .Y(_abc_17692_n12928) );
  OR2X2 OR2X2_4419 ( .A(_abc_17692_n12926), .B(_abc_17692_n12882), .Y(_abc_17692_n12929) );
  OR2X2 OR2X2_442 ( .A(_abc_17692_n1828), .B(_abc_17692_n1814), .Y(_abc_17692_n1829) );
  OR2X2 OR2X2_4420 ( .A(_abc_17692_n12931), .B(_abc_17692_n12924), .Y(_abc_17692_n12932) );
  OR2X2 OR2X2_4421 ( .A(_abc_17692_n12932), .B(_abc_17692_n12918), .Y(_abc_17692_n12933) );
  OR2X2 OR2X2_4422 ( .A(_abc_17692_n12933), .B(_abc_17692_n12910), .Y(_abc_17692_n12934) );
  OR2X2 OR2X2_4423 ( .A(_abc_17692_n12936), .B(_abc_17692_n12937), .Y(_abc_17692_n12938) );
  OR2X2 OR2X2_4424 ( .A(_abc_17692_n12935), .B(_abc_17692_n12938), .Y(_abc_17692_n12939) );
  OR2X2 OR2X2_4425 ( .A(_abc_17692_n12939), .B(_abc_17692_n12902), .Y(workunit1_31__FF_INPUT) );
  OR2X2 OR2X2_4426 ( .A(state_12_), .B(state_11_), .Y(_abc_17692_n12942) );
  OR2X2 OR2X2_4427 ( .A(_abc_17692_n12946), .B(_abc_17692_n12947), .Y(_abc_17692_n12948) );
  OR2X2 OR2X2_4428 ( .A(_abc_17692_n12945), .B(_abc_17692_n12948), .Y(selectslice_0__FF_INPUT) );
  OR2X2 OR2X2_4429 ( .A(_abc_17692_n12951), .B(_abc_17692_n12952), .Y(_abc_17692_n12953) );
  OR2X2 OR2X2_443 ( .A(_abc_17692_n1831), .B(workunit2_0_), .Y(_abc_17692_n1832) );
  OR2X2 OR2X2_4430 ( .A(_abc_17692_n12950), .B(_abc_17692_n12953), .Y(selectslice_1__FF_INPUT) );
  OR2X2 OR2X2_444 ( .A(sum_0_), .B(\key_in[32] ), .Y(_abc_17692_n1837) );
  OR2X2 OR2X2_445 ( .A(_abc_17692_n1841), .B(_abc_17692_n1840), .Y(_abc_17692_n1842) );
  OR2X2 OR2X2_446 ( .A(_abc_17692_n1843), .B(workunit2_0_), .Y(_abc_17692_n1844) );
  OR2X2 OR2X2_447 ( .A(_abc_17692_n1842), .B(_abc_17692_n1814), .Y(_abc_17692_n1847) );
  OR2X2 OR2X2_448 ( .A(_abc_17692_n1834), .B(_abc_17692_n1849), .Y(_abc_17692_n1850) );
  OR2X2 OR2X2_449 ( .A(sum_0_), .B(\key_in[96] ), .Y(_abc_17692_n1853) );
  OR2X2 OR2X2_45 ( .A(_abc_17692_n727_bF_buf6), .B(workunit2_1_bF_buf3), .Y(_abc_17692_n731_1) );
  OR2X2 OR2X2_450 ( .A(_abc_17692_n1857), .B(_abc_17692_n1856), .Y(_abc_17692_n1858) );
  OR2X2 OR2X2_451 ( .A(_abc_17692_n1859), .B(workunit2_0_), .Y(_abc_17692_n1864) );
  OR2X2 OR2X2_452 ( .A(sum_0_), .B(\key_in[64] ), .Y(_abc_17692_n1869) );
  OR2X2 OR2X2_453 ( .A(_abc_17692_n1873), .B(_abc_17692_n1872), .Y(_abc_17692_n1874) );
  OR2X2 OR2X2_454 ( .A(_abc_17692_n1875), .B(workunit2_0_), .Y(_abc_17692_n1876) );
  OR2X2 OR2X2_455 ( .A(_abc_17692_n1881), .B(_abc_17692_n1866), .Y(_abc_17692_n1882) );
  OR2X2 OR2X2_456 ( .A(_abc_17692_n1882), .B(_abc_17692_n1850), .Y(_abc_17692_n1883) );
  OR2X2 OR2X2_457 ( .A(_abc_17692_n1886), .B(_abc_17692_n1887), .Y(_abc_17692_n1888) );
  OR2X2 OR2X2_458 ( .A(_abc_17692_n1884_1), .B(_abc_17692_n1888), .Y(workunit2_0__FF_INPUT) );
  OR2X2 OR2X2_459 ( .A(workunit1_1_bF_buf1), .B(workunit1_6_), .Y(_abc_17692_n1892) );
  OR2X2 OR2X2_46 ( .A(_abc_17692_n725_bF_buf4), .B(_auto_iopadmap_cc_313_execute_30065_2_), .Y(_abc_17692_n733) );
  OR2X2 OR2X2_460 ( .A(_abc_17692_n1893), .B(_abc_17692_n1891), .Y(_abc_17692_n1894) );
  OR2X2 OR2X2_461 ( .A(_abc_17692_n1894), .B(_abc_17692_n1890), .Y(_abc_17692_n1895) );
  OR2X2 OR2X2_462 ( .A(_abc_17692_n1897), .B(_abc_17692_n1815_1), .Y(_abc_17692_n1898) );
  OR2X2 OR2X2_463 ( .A(sum_1_), .B(\key_in[65] ), .Y(_abc_17692_n1902) );
  OR2X2 OR2X2_464 ( .A(_abc_17692_n1905), .B(_abc_17692_n1900), .Y(_abc_17692_n1906) );
  OR2X2 OR2X2_465 ( .A(_abc_17692_n1907), .B(_abc_17692_n1904), .Y(_abc_17692_n1908) );
  OR2X2 OR2X2_466 ( .A(_abc_17692_n1911), .B(_abc_17692_n1910), .Y(_abc_17692_n1912) );
  OR2X2 OR2X2_467 ( .A(_abc_17692_n1906), .B(_abc_17692_n1868), .Y(_abc_17692_n1913) );
  OR2X2 OR2X2_468 ( .A(_abc_17692_n1903), .B(_abc_17692_n1867_1), .Y(_abc_17692_n1914) );
  OR2X2 OR2X2_469 ( .A(_abc_17692_n1909), .B(_abc_17692_n1916), .Y(_abc_17692_n1917) );
  OR2X2 OR2X2_47 ( .A(_abc_17692_n727_bF_buf5), .B(workunit2_2_), .Y(_abc_17692_n734) );
  OR2X2 OR2X2_470 ( .A(_abc_17692_n1912), .B(_abc_17692_n1915), .Y(_abc_17692_n1920) );
  OR2X2 OR2X2_471 ( .A(_abc_17692_n1899), .B(_abc_17692_n1908), .Y(_abc_17692_n1921) );
  OR2X2 OR2X2_472 ( .A(_abc_17692_n1918), .B(_abc_17692_n1923), .Y(_abc_17692_n1924) );
  OR2X2 OR2X2_473 ( .A(_abc_17692_n1924), .B(_abc_17692_n1926), .Y(_abc_17692_n1927) );
  OR2X2 OR2X2_474 ( .A(sum_1_), .B(\key_in[1] ), .Y(_abc_17692_n1936) );
  OR2X2 OR2X2_475 ( .A(_abc_17692_n1939), .B(_abc_17692_n1934), .Y(_abc_17692_n1940) );
  OR2X2 OR2X2_476 ( .A(_abc_17692_n1941), .B(_abc_17692_n1938), .Y(_abc_17692_n1942) );
  OR2X2 OR2X2_477 ( .A(_abc_17692_n1940), .B(_abc_17692_n1821), .Y(_abc_17692_n1944) );
  OR2X2 OR2X2_478 ( .A(_abc_17692_n1937), .B(_abc_17692_n1820), .Y(_abc_17692_n1945) );
  OR2X2 OR2X2_479 ( .A(_abc_17692_n1943), .B(_abc_17692_n1947), .Y(_abc_17692_n1948) );
  OR2X2 OR2X2_48 ( .A(_abc_17692_n725_bF_buf3), .B(_auto_iopadmap_cc_313_execute_30065_3_), .Y(_abc_17692_n736) );
  OR2X2 OR2X2_480 ( .A(_abc_17692_n1912), .B(_abc_17692_n1946), .Y(_abc_17692_n1950) );
  OR2X2 OR2X2_481 ( .A(_abc_17692_n1899), .B(_abc_17692_n1942), .Y(_abc_17692_n1951) );
  OR2X2 OR2X2_482 ( .A(_abc_17692_n1949), .B(_abc_17692_n1953), .Y(_abc_17692_n1954) );
  OR2X2 OR2X2_483 ( .A(_abc_17692_n1954), .B(_abc_17692_n1933), .Y(_abc_17692_n1955) );
  OR2X2 OR2X2_484 ( .A(_abc_17692_n1952), .B(_abc_17692_n1919_1), .Y(_abc_17692_n1956) );
  OR2X2 OR2X2_485 ( .A(_abc_17692_n1948), .B(workunit2_1_bF_buf3), .Y(_abc_17692_n1957) );
  OR2X2 OR2X2_486 ( .A(_abc_17692_n1958), .B(_abc_17692_n1932), .Y(_abc_17692_n1959) );
  OR2X2 OR2X2_487 ( .A(sum_1_), .B(\key_in[33] ), .Y(_abc_17692_n1966) );
  OR2X2 OR2X2_488 ( .A(_abc_17692_n1971_1), .B(_abc_17692_n1964), .Y(_abc_17692_n1972) );
  OR2X2 OR2X2_489 ( .A(_abc_17692_n1973), .B(_abc_17692_n1968), .Y(_abc_17692_n1974_1) );
  OR2X2 OR2X2_49 ( .A(_abc_17692_n727_bF_buf4), .B(workunit2_3_), .Y(_abc_17692_n737) );
  OR2X2 OR2X2_490 ( .A(_abc_17692_n1912), .B(_abc_17692_n1974_1), .Y(_abc_17692_n1975) );
  OR2X2 OR2X2_491 ( .A(_abc_17692_n1972), .B(_abc_17692_n1836), .Y(_abc_17692_n1976) );
  OR2X2 OR2X2_492 ( .A(_abc_17692_n1967), .B(_abc_17692_n1835), .Y(_abc_17692_n1977) );
  OR2X2 OR2X2_493 ( .A(_abc_17692_n1899), .B(_abc_17692_n1978), .Y(_abc_17692_n1979) );
  OR2X2 OR2X2_494 ( .A(_abc_17692_n1912), .B(_abc_17692_n1978), .Y(_abc_17692_n1982) );
  OR2X2 OR2X2_495 ( .A(_abc_17692_n1899), .B(_abc_17692_n1974_1), .Y(_abc_17692_n1983) );
  OR2X2 OR2X2_496 ( .A(_abc_17692_n1981_1), .B(_abc_17692_n1985), .Y(_abc_17692_n1986) );
  OR2X2 OR2X2_497 ( .A(_abc_17692_n1986), .B(_abc_17692_n1963), .Y(_abc_17692_n1989) );
  OR2X2 OR2X2_498 ( .A(_abc_17692_n1961), .B(_abc_17692_n1991), .Y(_abc_17692_n1992) );
  OR2X2 OR2X2_499 ( .A(_abc_17692_n1992), .B(_abc_17692_n1931), .Y(_abc_17692_n1993_1) );
  OR2X2 OR2X2_5 ( .A(state_8_bF_buf6), .B(delta_0_), .Y(delta_0__FF_INPUT) );
  OR2X2 OR2X2_50 ( .A(_abc_17692_n725_bF_buf2), .B(_auto_iopadmap_cc_313_execute_30065_4_), .Y(_abc_17692_n739) );
  OR2X2 OR2X2_500 ( .A(sum_1_), .B(\key_in[97] ), .Y(_abc_17692_n1997) );
  OR2X2 OR2X2_501 ( .A(_abc_17692_n1998), .B(_abc_17692_n1851), .Y(_abc_17692_n2001) );
  OR2X2 OR2X2_502 ( .A(_abc_17692_n2002), .B(_abc_17692_n1912), .Y(_abc_17692_n2003) );
  OR2X2 OR2X2_503 ( .A(_abc_17692_n2004_1), .B(_abc_17692_n1995), .Y(_abc_17692_n2005) );
  OR2X2 OR2X2_504 ( .A(_abc_17692_n2006), .B(_abc_17692_n1999), .Y(_abc_17692_n2007) );
  OR2X2 OR2X2_505 ( .A(_abc_17692_n1899), .B(_abc_17692_n2007), .Y(_abc_17692_n2008) );
  OR2X2 OR2X2_506 ( .A(_abc_17692_n2009), .B(_abc_17692_n1919_1), .Y(_abc_17692_n2010) );
  OR2X2 OR2X2_507 ( .A(_abc_17692_n2012), .B(_abc_17692_n2011), .Y(_abc_17692_n2013) );
  OR2X2 OR2X2_508 ( .A(_abc_17692_n2013), .B(workunit2_1_bF_buf1), .Y(_abc_17692_n2014) );
  OR2X2 OR2X2_509 ( .A(_abc_17692_n2015), .B(_abc_17692_n1994), .Y(_abc_17692_n2016_1) );
  OR2X2 OR2X2_51 ( .A(_abc_17692_n727_bF_buf3), .B(workunit2_4_), .Y(_abc_17692_n740) );
  OR2X2 OR2X2_510 ( .A(_abc_17692_n2018), .B(_abc_17692_n2019), .Y(_abc_17692_n2020) );
  OR2X2 OR2X2_511 ( .A(_abc_17692_n2020), .B(_abc_17692_n2017), .Y(_abc_17692_n2021) );
  OR2X2 OR2X2_512 ( .A(_abc_17692_n1993_1), .B(_abc_17692_n2023), .Y(_abc_17692_n2024) );
  OR2X2 OR2X2_513 ( .A(_abc_17692_n1922), .B(_abc_17692_n1919_1), .Y(_abc_17692_n2026) );
  OR2X2 OR2X2_514 ( .A(_abc_17692_n1917), .B(workunit2_1_bF_buf3), .Y(_abc_17692_n2027) );
  OR2X2 OR2X2_515 ( .A(_abc_17692_n2028), .B(_abc_17692_n1878), .Y(_abc_17692_n2029) );
  OR2X2 OR2X2_516 ( .A(_abc_17692_n1924), .B(_abc_17692_n1879), .Y(_abc_17692_n2030) );
  OR2X2 OR2X2_517 ( .A(_abc_17692_n1958), .B(_abc_17692_n2033), .Y(_abc_17692_n2036) );
  OR2X2 OR2X2_518 ( .A(_abc_17692_n2032), .B(_abc_17692_n2038), .Y(_abc_17692_n2039) );
  OR2X2 OR2X2_519 ( .A(_abc_17692_n2020), .B(_abc_17692_n1861), .Y(_abc_17692_n2040) );
  OR2X2 OR2X2_52 ( .A(_abc_17692_n725_bF_buf1), .B(_auto_iopadmap_cc_313_execute_30065_5_), .Y(_abc_17692_n742) );
  OR2X2 OR2X2_520 ( .A(_abc_17692_n2015), .B(_abc_17692_n1860), .Y(_abc_17692_n2041) );
  OR2X2 OR2X2_521 ( .A(_abc_17692_n1986), .B(_abc_17692_n1847), .Y(_abc_17692_n2044) );
  OR2X2 OR2X2_522 ( .A(_abc_17692_n1984), .B(_abc_17692_n1919_1), .Y(_abc_17692_n2046) );
  OR2X2 OR2X2_523 ( .A(_abc_17692_n1980), .B(workunit2_1_bF_buf2), .Y(_abc_17692_n2047) );
  OR2X2 OR2X2_524 ( .A(_abc_17692_n2048), .B(_abc_17692_n2045), .Y(_abc_17692_n2049_1) );
  OR2X2 OR2X2_525 ( .A(_abc_17692_n2043), .B(_abc_17692_n2051), .Y(_abc_17692_n2052_1) );
  OR2X2 OR2X2_526 ( .A(_abc_17692_n2039), .B(_abc_17692_n2052_1), .Y(_abc_17692_n2053) );
  OR2X2 OR2X2_527 ( .A(_abc_17692_n2055), .B(_abc_17692_n2056), .Y(_abc_17692_n2057) );
  OR2X2 OR2X2_528 ( .A(_abc_17692_n2054), .B(_abc_17692_n2057), .Y(_abc_17692_n2058) );
  OR2X2 OR2X2_529 ( .A(_abc_17692_n2058), .B(_abc_17692_n2025), .Y(workunit2_1__FF_INPUT) );
  OR2X2 OR2X2_53 ( .A(_abc_17692_n727_bF_buf2), .B(workunit2_5_), .Y(_abc_17692_n743) );
  OR2X2 OR2X2_530 ( .A(_abc_17692_n1910), .B(_abc_17692_n1891), .Y(_abc_17692_n2060) );
  OR2X2 OR2X2_531 ( .A(_abc_17692_n2064), .B(_abc_17692_n2061), .Y(_abc_17692_n2065) );
  OR2X2 OR2X2_532 ( .A(_abc_17692_n2069), .B(_abc_17692_n2067), .Y(_abc_17692_n2070) );
  OR2X2 OR2X2_533 ( .A(sum_2_), .B(\key_in[66] ), .Y(_abc_17692_n2074) );
  OR2X2 OR2X2_534 ( .A(_abc_17692_n2071), .B(_abc_17692_n2076), .Y(_abc_17692_n2077) );
  OR2X2 OR2X2_535 ( .A(_abc_17692_n1904), .B(_abc_17692_n1900), .Y(_abc_17692_n2078) );
  OR2X2 OR2X2_536 ( .A(_abc_17692_n2078), .B(_abc_17692_n2075), .Y(_abc_17692_n2079) );
  OR2X2 OR2X2_537 ( .A(_abc_17692_n2070), .B(_abc_17692_n2080), .Y(_abc_17692_n2081) );
  OR2X2 OR2X2_538 ( .A(_abc_17692_n2068), .B(_abc_17692_n2065), .Y(_abc_17692_n2082) );
  OR2X2 OR2X2_539 ( .A(_abc_17692_n2060), .B(_abc_17692_n2066), .Y(_abc_17692_n2083) );
  OR2X2 OR2X2_54 ( .A(_abc_17692_n725_bF_buf0), .B(_auto_iopadmap_cc_313_execute_30065_6_), .Y(_abc_17692_n745) );
  OR2X2 OR2X2_540 ( .A(_abc_17692_n2086), .B(_abc_17692_n2085), .Y(_abc_17692_n2087_1) );
  OR2X2 OR2X2_541 ( .A(_abc_17692_n2084), .B(_abc_17692_n2087_1), .Y(_abc_17692_n2088) );
  OR2X2 OR2X2_542 ( .A(_abc_17692_n2089), .B(workunit2_2_), .Y(_abc_17692_n2090) );
  OR2X2 OR2X2_543 ( .A(_abc_17692_n2092), .B(_abc_17692_n2093), .Y(_abc_17692_n2094) );
  OR2X2 OR2X2_544 ( .A(_abc_17692_n2094), .B(_abc_17692_n2091), .Y(_abc_17692_n2095) );
  OR2X2 OR2X2_545 ( .A(_abc_17692_n1928), .B(_abc_17692_n2097), .Y(_abc_17692_n2098) );
  OR2X2 OR2X2_546 ( .A(_abc_17692_n2098), .B(_abc_17692_n2096), .Y(_abc_17692_n2101) );
  OR2X2 OR2X2_547 ( .A(_abc_17692_n1968), .B(_abc_17692_n1964), .Y(_abc_17692_n2104) );
  OR2X2 OR2X2_548 ( .A(sum_2_), .B(\key_in[34] ), .Y(_abc_17692_n2107) );
  OR2X2 OR2X2_549 ( .A(_abc_17692_n2112_1), .B(_abc_17692_n2109), .Y(_abc_17692_n2113) );
  OR2X2 OR2X2_55 ( .A(_abc_17692_n727_bF_buf1), .B(workunit2_6_), .Y(_abc_17692_n746) );
  OR2X2 OR2X2_550 ( .A(_abc_17692_n2070), .B(_abc_17692_n2113), .Y(_abc_17692_n2114) );
  OR2X2 OR2X2_551 ( .A(_abc_17692_n2110), .B(_abc_17692_n2111), .Y(_abc_17692_n2115) );
  OR2X2 OR2X2_552 ( .A(_abc_17692_n2104), .B(_abc_17692_n2108), .Y(_abc_17692_n2116) );
  OR2X2 OR2X2_553 ( .A(_abc_17692_n2084), .B(_abc_17692_n2117), .Y(_abc_17692_n2118) );
  OR2X2 OR2X2_554 ( .A(_abc_17692_n2119), .B(_abc_17692_n2091), .Y(_abc_17692_n2120) );
  OR2X2 OR2X2_555 ( .A(_abc_17692_n2070), .B(_abc_17692_n2117), .Y(_abc_17692_n2121) );
  OR2X2 OR2X2_556 ( .A(_abc_17692_n2084), .B(_abc_17692_n2113), .Y(_abc_17692_n2122) );
  OR2X2 OR2X2_557 ( .A(_abc_17692_n2123), .B(workunit2_2_), .Y(_abc_17692_n2124) );
  OR2X2 OR2X2_558 ( .A(_abc_17692_n1987), .B(_abc_17692_n2126), .Y(_abc_17692_n2127) );
  OR2X2 OR2X2_559 ( .A(_abc_17692_n2127), .B(_abc_17692_n2125), .Y(_abc_17692_n2130) );
  OR2X2 OR2X2_56 ( .A(_abc_17692_n725_bF_buf7), .B(_auto_iopadmap_cc_313_execute_30065_7_), .Y(_abc_17692_n748) );
  OR2X2 OR2X2_560 ( .A(_abc_17692_n1938), .B(_abc_17692_n1934), .Y(_abc_17692_n2133) );
  OR2X2 OR2X2_561 ( .A(sum_2_), .B(\key_in[2] ), .Y(_abc_17692_n2136) );
  OR2X2 OR2X2_562 ( .A(_abc_17692_n2133), .B(_abc_17692_n2137_1), .Y(_abc_17692_n2140) );
  OR2X2 OR2X2_563 ( .A(_abc_17692_n2141), .B(_abc_17692_n2070), .Y(_abc_17692_n2142) );
  OR2X2 OR2X2_564 ( .A(_abc_17692_n2145), .B(_abc_17692_n2138), .Y(_abc_17692_n2146) );
  OR2X2 OR2X2_565 ( .A(_abc_17692_n2084), .B(_abc_17692_n2146), .Y(_abc_17692_n2147) );
  OR2X2 OR2X2_566 ( .A(_abc_17692_n2148), .B(_abc_17692_n2091), .Y(_abc_17692_n2149) );
  OR2X2 OR2X2_567 ( .A(_abc_17692_n2151), .B(_abc_17692_n2150), .Y(_abc_17692_n2152) );
  OR2X2 OR2X2_568 ( .A(_abc_17692_n2152), .B(workunit2_2_), .Y(_abc_17692_n2153) );
  OR2X2 OR2X2_569 ( .A(_abc_17692_n2154), .B(_abc_17692_n2157), .Y(_abc_17692_n2158) );
  OR2X2 OR2X2_57 ( .A(_abc_17692_n727_bF_buf0), .B(workunit2_7_), .Y(_abc_17692_n749) );
  OR2X2 OR2X2_570 ( .A(_abc_17692_n2152), .B(_abc_17692_n2091), .Y(_abc_17692_n2159) );
  OR2X2 OR2X2_571 ( .A(_abc_17692_n2148), .B(workunit2_2_), .Y(_abc_17692_n2160) );
  OR2X2 OR2X2_572 ( .A(_abc_17692_n2162), .B(_abc_17692_n2155), .Y(_abc_17692_n2163) );
  OR2X2 OR2X2_573 ( .A(_abc_17692_n2163), .B(_abc_17692_n2161), .Y(_abc_17692_n2164) );
  OR2X2 OR2X2_574 ( .A(_abc_17692_n2166), .B(_abc_17692_n2132), .Y(_abc_17692_n2167) );
  OR2X2 OR2X2_575 ( .A(_abc_17692_n2167), .B(_abc_17692_n2103), .Y(_abc_17692_n2168) );
  OR2X2 OR2X2_576 ( .A(_abc_17692_n1999), .B(_abc_17692_n1995), .Y(_abc_17692_n2169) );
  OR2X2 OR2X2_577 ( .A(sum_2_), .B(\key_in[98] ), .Y(_abc_17692_n2172) );
  OR2X2 OR2X2_578 ( .A(_abc_17692_n2169), .B(_abc_17692_n2173), .Y(_abc_17692_n2176) );
  OR2X2 OR2X2_579 ( .A(_abc_17692_n2177), .B(_abc_17692_n2070), .Y(_abc_17692_n2178) );
  OR2X2 OR2X2_58 ( .A(_abc_17692_n725_bF_buf6), .B(_auto_iopadmap_cc_313_execute_30065_8_), .Y(_abc_17692_n751_1) );
  OR2X2 OR2X2_580 ( .A(_abc_17692_n2181), .B(_abc_17692_n2174), .Y(_abc_17692_n2182) );
  OR2X2 OR2X2_581 ( .A(_abc_17692_n2182), .B(_abc_17692_n2084), .Y(_abc_17692_n2183) );
  OR2X2 OR2X2_582 ( .A(_abc_17692_n2184), .B(_abc_17692_n2091), .Y(_abc_17692_n2185) );
  OR2X2 OR2X2_583 ( .A(_abc_17692_n2182), .B(_abc_17692_n2070), .Y(_abc_17692_n2186) );
  OR2X2 OR2X2_584 ( .A(_abc_17692_n2177), .B(_abc_17692_n2084), .Y(_abc_17692_n2187) );
  OR2X2 OR2X2_585 ( .A(_abc_17692_n2188), .B(workunit2_2_), .Y(_abc_17692_n2189) );
  OR2X2 OR2X2_586 ( .A(_abc_17692_n2190), .B(_abc_17692_n2193), .Y(_abc_17692_n2194) );
  OR2X2 OR2X2_587 ( .A(_abc_17692_n2188), .B(_abc_17692_n2091), .Y(_abc_17692_n2195) );
  OR2X2 OR2X2_588 ( .A(_abc_17692_n2184), .B(workunit2_2_), .Y(_abc_17692_n2196) );
  OR2X2 OR2X2_589 ( .A(_abc_17692_n2198), .B(_abc_17692_n2197), .Y(_abc_17692_n2199) );
  OR2X2 OR2X2_59 ( .A(_abc_17692_n727_bF_buf7), .B(workunit2_8_bF_buf3), .Y(_abc_17692_n752) );
  OR2X2 OR2X2_590 ( .A(_abc_17692_n2168), .B(_abc_17692_n2201), .Y(_abc_17692_n2202) );
  OR2X2 OR2X2_591 ( .A(_abc_17692_n2089), .B(_abc_17692_n2091), .Y(_abc_17692_n2204) );
  OR2X2 OR2X2_592 ( .A(_abc_17692_n2094), .B(workunit2_2_), .Y(_abc_17692_n2205) );
  OR2X2 OR2X2_593 ( .A(_abc_17692_n2207), .B(_abc_17692_n1918), .Y(_abc_17692_n2208) );
  OR2X2 OR2X2_594 ( .A(_abc_17692_n2206), .B(_abc_17692_n2208), .Y(_abc_17692_n2209) );
  OR2X2 OR2X2_595 ( .A(_abc_17692_n2210), .B(_abc_17692_n2096), .Y(_abc_17692_n2211_1) );
  OR2X2 OR2X2_596 ( .A(_abc_17692_n2034), .B(_abc_17692_n1949), .Y(_abc_17692_n2214_1) );
  OR2X2 OR2X2_597 ( .A(_abc_17692_n2154), .B(_abc_17692_n2214_1), .Y(_abc_17692_n2217) );
  OR2X2 OR2X2_598 ( .A(_abc_17692_n2213), .B(_abc_17692_n2219), .Y(_abc_17692_n2220) );
  OR2X2 OR2X2_599 ( .A(_abc_17692_n2221), .B(_abc_17692_n2197), .Y(_abc_17692_n2222) );
  OR2X2 OR2X2_6 ( .A(state_8_bF_buf5), .B(delta_3_), .Y(delta_3__FF_INPUT) );
  OR2X2 OR2X2_60 ( .A(_abc_17692_n725_bF_buf5), .B(_auto_iopadmap_cc_313_execute_30065_9_), .Y(_abc_17692_n754) );
  OR2X2 OR2X2_600 ( .A(_abc_17692_n2223), .B(_abc_17692_n2018), .Y(_abc_17692_n2224) );
  OR2X2 OR2X2_601 ( .A(_abc_17692_n2190), .B(_abc_17692_n2224), .Y(_abc_17692_n2225) );
  OR2X2 OR2X2_602 ( .A(_abc_17692_n2228), .B(_abc_17692_n2125), .Y(_abc_17692_n2229) );
  OR2X2 OR2X2_603 ( .A(_abc_17692_n2123), .B(_abc_17692_n2091), .Y(_abc_17692_n2230) );
  OR2X2 OR2X2_604 ( .A(_abc_17692_n2119), .B(workunit2_2_), .Y(_abc_17692_n2231) );
  OR2X2 OR2X2_605 ( .A(_abc_17692_n2233), .B(_abc_17692_n1981_1), .Y(_abc_17692_n2234) );
  OR2X2 OR2X2_606 ( .A(_abc_17692_n2232), .B(_abc_17692_n2234), .Y(_abc_17692_n2235) );
  OR2X2 OR2X2_607 ( .A(_abc_17692_n2227), .B(_abc_17692_n2237), .Y(_abc_17692_n2238) );
  OR2X2 OR2X2_608 ( .A(_abc_17692_n2220), .B(_abc_17692_n2238), .Y(_abc_17692_n2239) );
  OR2X2 OR2X2_609 ( .A(_abc_17692_n2241), .B(_abc_17692_n2242_1), .Y(_abc_17692_n2243) );
  OR2X2 OR2X2_61 ( .A(_abc_17692_n727_bF_buf6), .B(workunit2_9_), .Y(_abc_17692_n755) );
  OR2X2 OR2X2_610 ( .A(_abc_17692_n2240), .B(_abc_17692_n2243), .Y(_abc_17692_n2244) );
  OR2X2 OR2X2_611 ( .A(_abc_17692_n2244), .B(_abc_17692_n2203), .Y(workunit2_2__FF_INPUT) );
  OR2X2 OR2X2_612 ( .A(_abc_17692_n2067), .B(_abc_17692_n2061), .Y(_abc_17692_n2247) );
  OR2X2 OR2X2_613 ( .A(_abc_17692_n2251), .B(_abc_17692_n2248), .Y(_abc_17692_n2252) );
  OR2X2 OR2X2_614 ( .A(_abc_17692_n2247), .B(_abc_17692_n2252), .Y(_abc_17692_n2253) );
  OR2X2 OR2X2_615 ( .A(_abc_17692_n2255), .B(_abc_17692_n2256), .Y(_abc_17692_n2257_1) );
  OR2X2 OR2X2_616 ( .A(_abc_17692_n2109), .B(_abc_17692_n2105), .Y(_abc_17692_n2259) );
  OR2X2 OR2X2_617 ( .A(sum_3_), .B(\key_in[35] ), .Y(_abc_17692_n2262) );
  OR2X2 OR2X2_618 ( .A(_abc_17692_n2259), .B(_abc_17692_n2264), .Y(_abc_17692_n2265) );
  OR2X2 OR2X2_619 ( .A(_abc_17692_n2266), .B(_abc_17692_n2263), .Y(_abc_17692_n2267) );
  OR2X2 OR2X2_62 ( .A(_abc_17692_n725_bF_buf4), .B(_auto_iopadmap_cc_313_execute_30065_10_), .Y(_abc_17692_n757) );
  OR2X2 OR2X2_620 ( .A(_abc_17692_n2258), .B(_abc_17692_n2268), .Y(_abc_17692_n2269) );
  OR2X2 OR2X2_621 ( .A(_abc_17692_n2270), .B(_abc_17692_n2271), .Y(_abc_17692_n2272) );
  OR2X2 OR2X2_622 ( .A(_abc_17692_n2273), .B(_abc_17692_n2274), .Y(_abc_17692_n2275) );
  OR2X2 OR2X2_623 ( .A(_abc_17692_n2272), .B(_abc_17692_n2275), .Y(_abc_17692_n2276) );
  OR2X2 OR2X2_624 ( .A(_abc_17692_n2277), .B(_abc_17692_n2246), .Y(_abc_17692_n2278_1) );
  OR2X2 OR2X2_625 ( .A(_abc_17692_n2258), .B(_abc_17692_n2275), .Y(_abc_17692_n2279) );
  OR2X2 OR2X2_626 ( .A(_abc_17692_n2272), .B(_abc_17692_n2268), .Y(_abc_17692_n2280) );
  OR2X2 OR2X2_627 ( .A(_abc_17692_n2281), .B(workunit2_3_), .Y(_abc_17692_n2282) );
  OR2X2 OR2X2_628 ( .A(_abc_17692_n2285), .B(_abc_17692_n2283), .Y(_abc_17692_n2286) );
  OR2X2 OR2X2_629 ( .A(_abc_17692_n2281), .B(_abc_17692_n2246), .Y(_abc_17692_n2287) );
  OR2X2 OR2X2_63 ( .A(_abc_17692_n727_bF_buf5), .B(workunit2_10_bF_buf3), .Y(_abc_17692_n758) );
  OR2X2 OR2X2_630 ( .A(_abc_17692_n2277), .B(workunit2_3_), .Y(_abc_17692_n2288) );
  OR2X2 OR2X2_631 ( .A(_abc_17692_n2284), .B(_abc_17692_n2289), .Y(_abc_17692_n2290) );
  OR2X2 OR2X2_632 ( .A(_abc_17692_n2085), .B(_abc_17692_n2072), .Y(_abc_17692_n2293) );
  OR2X2 OR2X2_633 ( .A(sum_3_), .B(\key_in[67] ), .Y(_abc_17692_n2296) );
  OR2X2 OR2X2_634 ( .A(_abc_17692_n2293), .B(_abc_17692_n2298), .Y(_abc_17692_n2299) );
  OR2X2 OR2X2_635 ( .A(_abc_17692_n2300), .B(_abc_17692_n2297), .Y(_abc_17692_n2301) );
  OR2X2 OR2X2_636 ( .A(_abc_17692_n2258), .B(_abc_17692_n2302), .Y(_abc_17692_n2303) );
  OR2X2 OR2X2_637 ( .A(_abc_17692_n2304), .B(_abc_17692_n2305), .Y(_abc_17692_n2306) );
  OR2X2 OR2X2_638 ( .A(_abc_17692_n2272), .B(_abc_17692_n2306), .Y(_abc_17692_n2307) );
  OR2X2 OR2X2_639 ( .A(_abc_17692_n2308), .B(_abc_17692_n2246), .Y(_abc_17692_n2309) );
  OR2X2 OR2X2_64 ( .A(_abc_17692_n725_bF_buf3), .B(_auto_iopadmap_cc_313_execute_30065_11_), .Y(_abc_17692_n760) );
  OR2X2 OR2X2_640 ( .A(_abc_17692_n2310), .B(_abc_17692_n2311), .Y(_abc_17692_n2312) );
  OR2X2 OR2X2_641 ( .A(_abc_17692_n2312), .B(workunit2_3_), .Y(_abc_17692_n2313) );
  OR2X2 OR2X2_642 ( .A(_abc_17692_n2099), .B(_abc_17692_n2315), .Y(_abc_17692_n2316) );
  OR2X2 OR2X2_643 ( .A(_abc_17692_n2316), .B(_abc_17692_n2314), .Y(_abc_17692_n2319) );
  OR2X2 OR2X2_644 ( .A(sum_3_), .B(\key_in[3] ), .Y(_abc_17692_n2325) );
  OR2X2 OR2X2_645 ( .A(_abc_17692_n2138), .B(_abc_17692_n2134), .Y(_abc_17692_n2328) );
  OR2X2 OR2X2_646 ( .A(_abc_17692_n2327), .B(_abc_17692_n2330), .Y(_abc_17692_n2331) );
  OR2X2 OR2X2_647 ( .A(_abc_17692_n2331), .B(_abc_17692_n2258), .Y(_abc_17692_n2332) );
  OR2X2 OR2X2_648 ( .A(_abc_17692_n2328), .B(_abc_17692_n2329_1), .Y(_abc_17692_n2333) );
  OR2X2 OR2X2_649 ( .A(_abc_17692_n2335), .B(_abc_17692_n2272), .Y(_abc_17692_n2336) );
  OR2X2 OR2X2_65 ( .A(_abc_17692_n727_bF_buf4), .B(workunit2_11_), .Y(_abc_17692_n761) );
  OR2X2 OR2X2_650 ( .A(_abc_17692_n2337), .B(_abc_17692_n2246), .Y(_abc_17692_n2338) );
  OR2X2 OR2X2_651 ( .A(_abc_17692_n2335), .B(_abc_17692_n2258), .Y(_abc_17692_n2339) );
  OR2X2 OR2X2_652 ( .A(_abc_17692_n2331), .B(_abc_17692_n2272), .Y(_abc_17692_n2340_1) );
  OR2X2 OR2X2_653 ( .A(_abc_17692_n2341), .B(workunit2_3_), .Y(_abc_17692_n2342) );
  OR2X2 OR2X2_654 ( .A(_abc_17692_n2344), .B(_abc_17692_n2343), .Y(_abc_17692_n2345) );
  OR2X2 OR2X2_655 ( .A(_abc_17692_n2341), .B(_abc_17692_n2246), .Y(_abc_17692_n2346) );
  OR2X2 OR2X2_656 ( .A(_abc_17692_n2337), .B(workunit2_3_), .Y(_abc_17692_n2347) );
  OR2X2 OR2X2_657 ( .A(_abc_17692_n2350), .B(_abc_17692_n2349), .Y(_abc_17692_n2351) );
  OR2X2 OR2X2_658 ( .A(_abc_17692_n2351), .B(_abc_17692_n2348), .Y(_abc_17692_n2352) );
  OR2X2 OR2X2_659 ( .A(_abc_17692_n2354), .B(_abc_17692_n2321), .Y(_abc_17692_n2355) );
  OR2X2 OR2X2_66 ( .A(_abc_17692_n725_bF_buf2), .B(_auto_iopadmap_cc_313_execute_30065_12_), .Y(_abc_17692_n763) );
  OR2X2 OR2X2_660 ( .A(_abc_17692_n2355), .B(_abc_17692_n2292), .Y(_abc_17692_n2356) );
  OR2X2 OR2X2_661 ( .A(_abc_17692_n2174), .B(_abc_17692_n2170), .Y(_abc_17692_n2357) );
  OR2X2 OR2X2_662 ( .A(sum_3_), .B(\key_in[99] ), .Y(_abc_17692_n2360) );
  OR2X2 OR2X2_663 ( .A(_abc_17692_n2365), .B(_abc_17692_n2362), .Y(_abc_17692_n2366) );
  OR2X2 OR2X2_664 ( .A(_abc_17692_n2366), .B(_abc_17692_n2258), .Y(_abc_17692_n2367) );
  OR2X2 OR2X2_665 ( .A(_abc_17692_n2357), .B(_abc_17692_n2361_1), .Y(_abc_17692_n2369) );
  OR2X2 OR2X2_666 ( .A(_abc_17692_n2370), .B(_abc_17692_n2272), .Y(_abc_17692_n2371) );
  OR2X2 OR2X2_667 ( .A(_abc_17692_n2372), .B(_abc_17692_n2246), .Y(_abc_17692_n2373) );
  OR2X2 OR2X2_668 ( .A(_abc_17692_n2370), .B(_abc_17692_n2258), .Y(_abc_17692_n2374) );
  OR2X2 OR2X2_669 ( .A(_abc_17692_n2366), .B(_abc_17692_n2272), .Y(_abc_17692_n2375) );
  OR2X2 OR2X2_67 ( .A(_abc_17692_n727_bF_buf3), .B(workunit2_12_bF_buf3), .Y(_abc_17692_n764) );
  OR2X2 OR2X2_670 ( .A(_abc_17692_n2376), .B(workunit2_3_), .Y(_abc_17692_n2377) );
  OR2X2 OR2X2_671 ( .A(_abc_17692_n2380_1), .B(_abc_17692_n2378), .Y(_abc_17692_n2381) );
  OR2X2 OR2X2_672 ( .A(_abc_17692_n2376), .B(_abc_17692_n2246), .Y(_abc_17692_n2382) );
  OR2X2 OR2X2_673 ( .A(_abc_17692_n2372), .B(workunit2_3_), .Y(_abc_17692_n2383) );
  OR2X2 OR2X2_674 ( .A(_abc_17692_n2379), .B(_abc_17692_n2384), .Y(_abc_17692_n2385) );
  OR2X2 OR2X2_675 ( .A(_abc_17692_n2356), .B(_abc_17692_n2387), .Y(_abc_17692_n2388) );
  OR2X2 OR2X2_676 ( .A(_abc_17692_n2312), .B(_abc_17692_n2246), .Y(_abc_17692_n2390) );
  OR2X2 OR2X2_677 ( .A(_abc_17692_n2308), .B(workunit2_3_), .Y(_abc_17692_n2391) );
  OR2X2 OR2X2_678 ( .A(_abc_17692_n2394), .B(_abc_17692_n2393), .Y(_abc_17692_n2395) );
  OR2X2 OR2X2_679 ( .A(_abc_17692_n2395), .B(_abc_17692_n2392), .Y(_abc_17692_n2396) );
  OR2X2 OR2X2_68 ( .A(_abc_17692_n725_bF_buf1), .B(_auto_iopadmap_cc_313_execute_30065_13_), .Y(_abc_17692_n766_1) );
  OR2X2 OR2X2_680 ( .A(_abc_17692_n2397), .B(_abc_17692_n2314), .Y(_abc_17692_n2398) );
  OR2X2 OR2X2_681 ( .A(_abc_17692_n2215), .B(_abc_17692_n2401), .Y(_abc_17692_n2402) );
  OR2X2 OR2X2_682 ( .A(_abc_17692_n2402), .B(_abc_17692_n2343), .Y(_abc_17692_n2405) );
  OR2X2 OR2X2_683 ( .A(_abc_17692_n2407), .B(_abc_17692_n2400), .Y(_abc_17692_n2408) );
  OR2X2 OR2X2_684 ( .A(_abc_17692_n2409), .B(_abc_17692_n2378), .Y(_abc_17692_n2410) );
  OR2X2 OR2X2_685 ( .A(_abc_17692_n2412), .B(_abc_17692_n2411), .Y(_abc_17692_n2413) );
  OR2X2 OR2X2_686 ( .A(_abc_17692_n2413), .B(_abc_17692_n2384), .Y(_abc_17692_n2414) );
  OR2X2 OR2X2_687 ( .A(_abc_17692_n2417), .B(_abc_17692_n2283), .Y(_abc_17692_n2418) );
  OR2X2 OR2X2_688 ( .A(_abc_17692_n2420), .B(_abc_17692_n2419), .Y(_abc_17692_n2421) );
  OR2X2 OR2X2_689 ( .A(_abc_17692_n2421), .B(_abc_17692_n2289), .Y(_abc_17692_n2422) );
  OR2X2 OR2X2_69 ( .A(_abc_17692_n727_bF_buf2), .B(workunit2_13_), .Y(_abc_17692_n767) );
  OR2X2 OR2X2_690 ( .A(_abc_17692_n2416), .B(_abc_17692_n2424), .Y(_abc_17692_n2425) );
  OR2X2 OR2X2_691 ( .A(_abc_17692_n2408), .B(_abc_17692_n2425), .Y(_abc_17692_n2426) );
  OR2X2 OR2X2_692 ( .A(_abc_17692_n2428), .B(_abc_17692_n2429), .Y(_abc_17692_n2430) );
  OR2X2 OR2X2_693 ( .A(_abc_17692_n2427), .B(_abc_17692_n2430), .Y(_abc_17692_n2431) );
  OR2X2 OR2X2_694 ( .A(_abc_17692_n2431), .B(_abc_17692_n2389), .Y(workunit2_3__FF_INPUT) );
  OR2X2 OR2X2_695 ( .A(_abc_17692_n1816), .B(workunit1_9_), .Y(_abc_17692_n2434) );
  OR2X2 OR2X2_696 ( .A(_abc_17692_n2435), .B(workunit1_0_), .Y(_abc_17692_n2436) );
  OR2X2 OR2X2_697 ( .A(_abc_17692_n2437), .B(_abc_17692_n2433), .Y(_abc_17692_n2438) );
  OR2X2 OR2X2_698 ( .A(_abc_17692_n2439), .B(_abc_17692_n2440), .Y(_abc_17692_n2441) );
  OR2X2 OR2X2_699 ( .A(_abc_17692_n2441), .B(workunit1_4_), .Y(_abc_17692_n2442) );
  OR2X2 OR2X2_7 ( .A(state_8_bF_buf4), .B(delta_4_), .Y(delta_4__FF_INPUT) );
  OR2X2 OR2X2_70 ( .A(_abc_17692_n725_bF_buf0), .B(_auto_iopadmap_cc_313_execute_30065_14_), .Y(_abc_17692_n769) );
  OR2X2 OR2X2_700 ( .A(_abc_17692_n2444), .B(_abc_17692_n2248), .Y(_abc_17692_n2445) );
  OR2X2 OR2X2_701 ( .A(_abc_17692_n2447), .B(_abc_17692_n2445), .Y(_abc_17692_n2448) );
  OR2X2 OR2X2_702 ( .A(_abc_17692_n2450), .B(_abc_17692_n2451), .Y(_abc_17692_n2452) );
  OR2X2 OR2X2_703 ( .A(_abc_17692_n2068), .B(_abc_17692_n2454), .Y(_abc_17692_n2455) );
  OR2X2 OR2X2_704 ( .A(_abc_17692_n2457), .B(_abc_17692_n2449), .Y(_abc_17692_n2458) );
  OR2X2 OR2X2_705 ( .A(_abc_17692_n2460), .B(_abc_17692_n2323), .Y(_abc_17692_n2461) );
  OR2X2 OR2X2_706 ( .A(_abc_17692_n2463), .B(_abc_17692_n2461), .Y(_abc_17692_n2464) );
  OR2X2 OR2X2_707 ( .A(sum_4_), .B(\key_in[4] ), .Y(_abc_17692_n2467) );
  OR2X2 OR2X2_708 ( .A(_abc_17692_n2143), .B(_abc_17692_n2471), .Y(_abc_17692_n2472) );
  OR2X2 OR2X2_709 ( .A(_abc_17692_n2475), .B(_abc_17692_n2469_1), .Y(_abc_17692_n2476) );
  OR2X2 OR2X2_71 ( .A(_abc_17692_n727_bF_buf1), .B(workunit2_14_bF_buf3), .Y(_abc_17692_n770) );
  OR2X2 OR2X2_710 ( .A(_abc_17692_n2477), .B(_abc_17692_n2479_1), .Y(_abc_17692_n2480) );
  OR2X2 OR2X2_711 ( .A(_abc_17692_n2484), .B(_abc_17692_n2481), .Y(_abc_17692_n2485) );
  OR2X2 OR2X2_712 ( .A(_abc_17692_n2487), .B(_abc_17692_n2486), .Y(_abc_17692_n2488) );
  OR2X2 OR2X2_713 ( .A(_abc_17692_n2490_1), .B(_abc_17692_n2489), .Y(_abc_17692_n2491) );
  OR2X2 OR2X2_714 ( .A(_abc_17692_n2491), .B(_abc_17692_n2485), .Y(_abc_17692_n2492) );
  OR2X2 OR2X2_715 ( .A(sum_4_), .B(\key_in[68] ), .Y(_abc_17692_n2497) );
  OR2X2 OR2X2_716 ( .A(_abc_17692_n2499), .B(_abc_17692_n2294), .Y(_abc_17692_n2500_1) );
  OR2X2 OR2X2_717 ( .A(_abc_17692_n2502), .B(_abc_17692_n2500_1), .Y(_abc_17692_n2503) );
  OR2X2 OR2X2_718 ( .A(_abc_17692_n2507), .B(_abc_17692_n2504), .Y(_abc_17692_n2508) );
  OR2X2 OR2X2_719 ( .A(_abc_17692_n2511), .B(_abc_17692_n2509), .Y(_abc_17692_n2512) );
  OR2X2 OR2X2_72 ( .A(_abc_17692_n725_bF_buf7), .B(_auto_iopadmap_cc_313_execute_30065_15_), .Y(_abc_17692_n772) );
  OR2X2 OR2X2_720 ( .A(_abc_17692_n2512), .B(_abc_17692_n2482), .Y(_abc_17692_n2513) );
  OR2X2 OR2X2_721 ( .A(_abc_17692_n2514), .B(workunit2_4_), .Y(_abc_17692_n2515) );
  OR2X2 OR2X2_722 ( .A(_abc_17692_n2317), .B(_abc_17692_n2518), .Y(_abc_17692_n2519) );
  OR2X2 OR2X2_723 ( .A(_abc_17692_n2519), .B(_abc_17692_n2517), .Y(_abc_17692_n2520) );
  OR2X2 OR2X2_724 ( .A(_abc_17692_n2525), .B(_abc_17692_n2260), .Y(_abc_17692_n2526) );
  OR2X2 OR2X2_725 ( .A(_abc_17692_n2528), .B(_abc_17692_n2526), .Y(_abc_17692_n2529) );
  OR2X2 OR2X2_726 ( .A(sum_4_), .B(\key_in[36] ), .Y(_abc_17692_n2532) );
  OR2X2 OR2X2_727 ( .A(_abc_17692_n2110), .B(_abc_17692_n2536), .Y(_abc_17692_n2537) );
  OR2X2 OR2X2_728 ( .A(_abc_17692_n2540), .B(_abc_17692_n2534), .Y(_abc_17692_n2541) );
  OR2X2 OR2X2_729 ( .A(_abc_17692_n2542), .B(_abc_17692_n2544), .Y(_abc_17692_n2545) );
  OR2X2 OR2X2_73 ( .A(_abc_17692_n727_bF_buf0), .B(workunit2_15_), .Y(_abc_17692_n773) );
  OR2X2 OR2X2_730 ( .A(_abc_17692_n2548), .B(_abc_17692_n2546), .Y(_abc_17692_n2549) );
  OR2X2 OR2X2_731 ( .A(_abc_17692_n2551), .B(_abc_17692_n2549), .Y(_abc_17692_n2554) );
  OR2X2 OR2X2_732 ( .A(_abc_17692_n2556), .B(_abc_17692_n2524), .Y(_abc_17692_n2557) );
  OR2X2 OR2X2_733 ( .A(_abc_17692_n2557), .B(_abc_17692_n2494), .Y(_abc_17692_n2558) );
  OR2X2 OR2X2_734 ( .A(_abc_17692_n2362), .B(_abc_17692_n2358), .Y(_abc_17692_n2559) );
  OR2X2 OR2X2_735 ( .A(sum_4_), .B(\key_in[100] ), .Y(_abc_17692_n2562) );
  OR2X2 OR2X2_736 ( .A(_abc_17692_n2559), .B(_abc_17692_n2563), .Y(_abc_17692_n2566) );
  OR2X2 OR2X2_737 ( .A(_abc_17692_n2567), .B(_abc_17692_n2458), .Y(_abc_17692_n2568) );
  OR2X2 OR2X2_738 ( .A(_abc_17692_n2571), .B(_abc_17692_n2564), .Y(_abc_17692_n2572) );
  OR2X2 OR2X2_739 ( .A(_abc_17692_n2572), .B(_abc_17692_n2459_1), .Y(_abc_17692_n2573) );
  OR2X2 OR2X2_74 ( .A(_abc_17692_n725_bF_buf6), .B(_auto_iopadmap_cc_313_execute_30065_16_), .Y(_abc_17692_n775) );
  OR2X2 OR2X2_740 ( .A(_abc_17692_n2574), .B(_abc_17692_n2482), .Y(_abc_17692_n2575) );
  OR2X2 OR2X2_741 ( .A(_abc_17692_n2572), .B(_abc_17692_n2458), .Y(_abc_17692_n2576) );
  OR2X2 OR2X2_742 ( .A(_abc_17692_n2567), .B(_abc_17692_n2459_1), .Y(_abc_17692_n2577) );
  OR2X2 OR2X2_743 ( .A(_abc_17692_n2578), .B(workunit2_4_), .Y(_abc_17692_n2579) );
  OR2X2 OR2X2_744 ( .A(_abc_17692_n2581_1), .B(_abc_17692_n2580), .Y(_abc_17692_n2582) );
  OR2X2 OR2X2_745 ( .A(_abc_17692_n2578), .B(_abc_17692_n2482), .Y(_abc_17692_n2583) );
  OR2X2 OR2X2_746 ( .A(_abc_17692_n2574), .B(workunit2_4_), .Y(_abc_17692_n2584) );
  OR2X2 OR2X2_747 ( .A(_abc_17692_n2586), .B(_abc_17692_n2585), .Y(_abc_17692_n2587) );
  OR2X2 OR2X2_748 ( .A(_abc_17692_n2558), .B(_abc_17692_n2589), .Y(_abc_17692_n2590) );
  OR2X2 OR2X2_749 ( .A(_abc_17692_n2593), .B(_abc_17692_n2592), .Y(_abc_17692_n2594) );
  OR2X2 OR2X2_75 ( .A(_abc_17692_n727_bF_buf7), .B(workunit2_16_bF_buf3), .Y(_abc_17692_n776) );
  OR2X2 OR2X2_750 ( .A(_abc_17692_n2594), .B(_abc_17692_n2516), .Y(_abc_17692_n2595) );
  OR2X2 OR2X2_751 ( .A(_abc_17692_n2596), .B(_abc_17692_n2517), .Y(_abc_17692_n2597) );
  OR2X2 OR2X2_752 ( .A(_abc_17692_n2403), .B(_abc_17692_n2600), .Y(_abc_17692_n2601) );
  OR2X2 OR2X2_753 ( .A(_abc_17692_n2601), .B(_abc_17692_n2486), .Y(_abc_17692_n2604) );
  OR2X2 OR2X2_754 ( .A(_abc_17692_n2599), .B(_abc_17692_n2606), .Y(_abc_17692_n2607) );
  OR2X2 OR2X2_755 ( .A(_abc_17692_n2608_1), .B(_abc_17692_n2585), .Y(_abc_17692_n2609) );
  OR2X2 OR2X2_756 ( .A(_abc_17692_n2611), .B(_abc_17692_n2610), .Y(_abc_17692_n2612) );
  OR2X2 OR2X2_757 ( .A(_abc_17692_n2612), .B(_abc_17692_n2580), .Y(_abc_17692_n2613) );
  OR2X2 OR2X2_758 ( .A(_abc_17692_n2616), .B(_abc_17692_n2549), .Y(_abc_17692_n2617) );
  OR2X2 OR2X2_759 ( .A(_abc_17692_n2620), .B(_abc_17692_n2619), .Y(_abc_17692_n2621) );
  OR2X2 OR2X2_76 ( .A(_abc_17692_n725_bF_buf5), .B(_auto_iopadmap_cc_313_execute_30065_17_), .Y(_abc_17692_n778) );
  OR2X2 OR2X2_760 ( .A(_abc_17692_n2621), .B(_abc_17692_n2618), .Y(_abc_17692_n2622) );
  OR2X2 OR2X2_761 ( .A(_abc_17692_n2615), .B(_abc_17692_n2624), .Y(_abc_17692_n2625) );
  OR2X2 OR2X2_762 ( .A(_abc_17692_n2607), .B(_abc_17692_n2625), .Y(_abc_17692_n2626) );
  OR2X2 OR2X2_763 ( .A(_abc_17692_n2628), .B(_abc_17692_n2629), .Y(_abc_17692_n2630) );
  OR2X2 OR2X2_764 ( .A(_abc_17692_n2627), .B(_abc_17692_n2630), .Y(_abc_17692_n2631) );
  OR2X2 OR2X2_765 ( .A(_abc_17692_n2591), .B(_abc_17692_n2631), .Y(workunit2_4__FF_INPUT) );
  OR2X2 OR2X2_766 ( .A(_abc_17692_n2456), .B(_abc_17692_n2452), .Y(_abc_17692_n2634_1) );
  OR2X2 OR2X2_767 ( .A(_abc_17692_n2639), .B(_abc_17692_n2636), .Y(_abc_17692_n2640) );
  OR2X2 OR2X2_768 ( .A(_abc_17692_n2640), .B(_abc_17692_n1817), .Y(_abc_17692_n2641) );
  OR2X2 OR2X2_769 ( .A(workunit1_1_bF_buf2), .B(workunit1_10_), .Y(_abc_17692_n2643) );
  OR2X2 OR2X2_77 ( .A(_abc_17692_n727_bF_buf6), .B(workunit2_17_), .Y(_abc_17692_n779) );
  OR2X2 OR2X2_770 ( .A(_abc_17692_n2644), .B(workunit1_5_), .Y(_abc_17692_n2645) );
  OR2X2 OR2X2_771 ( .A(_abc_17692_n2449), .B(_abc_17692_n2450), .Y(_abc_17692_n2648) );
  OR2X2 OR2X2_772 ( .A(_abc_17692_n2650), .B(_abc_17692_n2649), .Y(_abc_17692_n2651) );
  OR2X2 OR2X2_773 ( .A(_abc_17692_n2647), .B(_abc_17692_n2652), .Y(_abc_17692_n2653) );
  OR2X2 OR2X2_774 ( .A(_abc_17692_n2504), .B(_abc_17692_n2495), .Y(_abc_17692_n2654) );
  OR2X2 OR2X2_775 ( .A(sum_5_), .B(\key_in[69] ), .Y(_abc_17692_n2657) );
  OR2X2 OR2X2_776 ( .A(_abc_17692_n2654), .B(_abc_17692_n2659), .Y(_abc_17692_n2660) );
  OR2X2 OR2X2_777 ( .A(_abc_17692_n2648), .B(_abc_17692_n2651), .Y(_abc_17692_n2666) );
  OR2X2 OR2X2_778 ( .A(_abc_17692_n2635), .B(_abc_17692_n2646), .Y(_abc_17692_n2667) );
  OR2X2 OR2X2_779 ( .A(_abc_17692_n2665), .B(_abc_17692_n2669), .Y(_abc_17692_n2670) );
  OR2X2 OR2X2_78 ( .A(_abc_17692_n725_bF_buf4), .B(_auto_iopadmap_cc_313_execute_30065_18_), .Y(_abc_17692_n781) );
  OR2X2 OR2X2_780 ( .A(_abc_17692_n2671), .B(_abc_17692_n2633), .Y(_abc_17692_n2672) );
  OR2X2 OR2X2_781 ( .A(_abc_17692_n2670), .B(workunit2_5_), .Y(_abc_17692_n2673) );
  OR2X2 OR2X2_782 ( .A(_abc_17692_n2514), .B(_abc_17692_n2482), .Y(_abc_17692_n2675) );
  OR2X2 OR2X2_783 ( .A(_abc_17692_n2521), .B(_abc_17692_n2676), .Y(_abc_17692_n2677) );
  OR2X2 OR2X2_784 ( .A(_abc_17692_n2677), .B(_abc_17692_n2674), .Y(_abc_17692_n2680) );
  OR2X2 OR2X2_785 ( .A(_abc_17692_n2469_1), .B(_abc_17692_n2465), .Y(_abc_17692_n2683) );
  OR2X2 OR2X2_786 ( .A(_abc_17692_n2686), .B(_abc_17692_n2684), .Y(_abc_17692_n2687) );
  OR2X2 OR2X2_787 ( .A(_abc_17692_n2683), .B(_abc_17692_n2687), .Y(_abc_17692_n2688) );
  OR2X2 OR2X2_788 ( .A(_abc_17692_n2691), .B(_abc_17692_n2668), .Y(_abc_17692_n2692) );
  OR2X2 OR2X2_789 ( .A(_abc_17692_n2693), .B(_abc_17692_n2653), .Y(_abc_17692_n2694) );
  OR2X2 OR2X2_79 ( .A(_abc_17692_n727_bF_buf5), .B(workunit2_18_), .Y(_abc_17692_n782) );
  OR2X2 OR2X2_790 ( .A(_abc_17692_n2695), .B(_abc_17692_n2633), .Y(_abc_17692_n2696) );
  OR2X2 OR2X2_791 ( .A(_abc_17692_n2697), .B(workunit2_5_), .Y(_abc_17692_n2698) );
  OR2X2 OR2X2_792 ( .A(_abc_17692_n2703), .B(_abc_17692_n2700), .Y(_abc_17692_n2704) );
  OR2X2 OR2X2_793 ( .A(_abc_17692_n2705), .B(_abc_17692_n2701), .Y(_abc_17692_n2706) );
  OR2X2 OR2X2_794 ( .A(_abc_17692_n2706), .B(_abc_17692_n2699), .Y(_abc_17692_n2707) );
  OR2X2 OR2X2_795 ( .A(_abc_17692_n2538_1), .B(_abc_17692_n2539), .Y(_abc_17692_n2710) );
  OR2X2 OR2X2_796 ( .A(_abc_17692_n2714), .B(_abc_17692_n2712), .Y(_abc_17692_n2715) );
  OR2X2 OR2X2_797 ( .A(_abc_17692_n2534), .B(_abc_17692_n2530), .Y(_abc_17692_n2718) );
  OR2X2 OR2X2_798 ( .A(_abc_17692_n2717), .B(_abc_17692_n2719), .Y(_abc_17692_n2720) );
  OR2X2 OR2X2_799 ( .A(_abc_17692_n2668), .B(_abc_17692_n2720), .Y(_abc_17692_n2721) );
  OR2X2 OR2X2_8 ( .A(state_8_bF_buf3), .B(delta_5_), .Y(delta_5__FF_INPUT) );
  OR2X2 OR2X2_80 ( .A(_abc_17692_n725_bF_buf3), .B(_auto_iopadmap_cc_313_execute_30065_19_), .Y(_abc_17692_n784) );
  OR2X2 OR2X2_800 ( .A(_abc_17692_n2718), .B(_abc_17692_n2715), .Y(_abc_17692_n2722) );
  OR2X2 OR2X2_801 ( .A(_abc_17692_n2711), .B(_abc_17692_n2716_1), .Y(_abc_17692_n2723_1) );
  OR2X2 OR2X2_802 ( .A(_abc_17692_n2653), .B(_abc_17692_n2724), .Y(_abc_17692_n2725) );
  OR2X2 OR2X2_803 ( .A(_abc_17692_n2726), .B(_abc_17692_n2633), .Y(_abc_17692_n2727) );
  OR2X2 OR2X2_804 ( .A(_abc_17692_n2668), .B(_abc_17692_n2724), .Y(_abc_17692_n2728) );
  OR2X2 OR2X2_805 ( .A(_abc_17692_n2653), .B(_abc_17692_n2720), .Y(_abc_17692_n2729) );
  OR2X2 OR2X2_806 ( .A(_abc_17692_n2730), .B(workunit2_5_), .Y(_abc_17692_n2731) );
  OR2X2 OR2X2_807 ( .A(_abc_17692_n2552_1), .B(_abc_17692_n2734_1), .Y(_abc_17692_n2735) );
  OR2X2 OR2X2_808 ( .A(_abc_17692_n2735), .B(_abc_17692_n2733), .Y(_abc_17692_n2736) );
  OR2X2 OR2X2_809 ( .A(_abc_17692_n2740), .B(_abc_17692_n2709), .Y(_abc_17692_n2741) );
  OR2X2 OR2X2_81 ( .A(_abc_17692_n727_bF_buf4), .B(workunit2_19_), .Y(_abc_17692_n785) );
  OR2X2 OR2X2_810 ( .A(_abc_17692_n2741), .B(_abc_17692_n2682), .Y(_abc_17692_n2742) );
  OR2X2 OR2X2_811 ( .A(sum_5_), .B(\key_in[101] ), .Y(_abc_17692_n2746) );
  OR2X2 OR2X2_812 ( .A(_abc_17692_n2564), .B(_abc_17692_n2560), .Y(_abc_17692_n2749) );
  OR2X2 OR2X2_813 ( .A(_abc_17692_n2748), .B(_abc_17692_n2751), .Y(_abc_17692_n2752) );
  OR2X2 OR2X2_814 ( .A(_abc_17692_n2752), .B(_abc_17692_n2668), .Y(_abc_17692_n2753) );
  OR2X2 OR2X2_815 ( .A(_abc_17692_n2749), .B(_abc_17692_n2750), .Y(_abc_17692_n2754) );
  OR2X2 OR2X2_816 ( .A(_abc_17692_n2756), .B(_abc_17692_n2653), .Y(_abc_17692_n2757_1) );
  OR2X2 OR2X2_817 ( .A(_abc_17692_n2758), .B(_abc_17692_n2633), .Y(_abc_17692_n2759) );
  OR2X2 OR2X2_818 ( .A(_abc_17692_n2756), .B(_abc_17692_n2668), .Y(_abc_17692_n2760) );
  OR2X2 OR2X2_819 ( .A(_abc_17692_n2752), .B(_abc_17692_n2653), .Y(_abc_17692_n2761) );
  OR2X2 OR2X2_82 ( .A(_abc_17692_n725_bF_buf2), .B(_auto_iopadmap_cc_313_execute_30065_20_), .Y(_abc_17692_n787) );
  OR2X2 OR2X2_820 ( .A(_abc_17692_n2762), .B(workunit2_5_), .Y(_abc_17692_n2763) );
  OR2X2 OR2X2_821 ( .A(_abc_17692_n2765), .B(_abc_17692_n2764), .Y(_abc_17692_n2766) );
  OR2X2 OR2X2_822 ( .A(_abc_17692_n2762), .B(_abc_17692_n2633), .Y(_abc_17692_n2767) );
  OR2X2 OR2X2_823 ( .A(_abc_17692_n2758), .B(workunit2_5_), .Y(_abc_17692_n2768) );
  OR2X2 OR2X2_824 ( .A(_abc_17692_n2770), .B(_abc_17692_n2769), .Y(_abc_17692_n2771) );
  OR2X2 OR2X2_825 ( .A(_abc_17692_n2742), .B(_abc_17692_n2773), .Y(_abc_17692_n2774) );
  OR2X2 OR2X2_826 ( .A(_abc_17692_n2778), .B(_abc_17692_n2777), .Y(_abc_17692_n2779) );
  OR2X2 OR2X2_827 ( .A(_abc_17692_n2779), .B(_abc_17692_n2776), .Y(_abc_17692_n2780) );
  OR2X2 OR2X2_828 ( .A(_abc_17692_n2781), .B(_abc_17692_n2674), .Y(_abc_17692_n2782) );
  OR2X2 OR2X2_829 ( .A(_abc_17692_n2602), .B(_abc_17692_n2481), .Y(_abc_17692_n2785) );
  OR2X2 OR2X2_83 ( .A(_abc_17692_n727_bF_buf3), .B(workunit2_20_), .Y(_abc_17692_n788) );
  OR2X2 OR2X2_830 ( .A(_abc_17692_n2785), .B(_abc_17692_n2700), .Y(_abc_17692_n2788) );
  OR2X2 OR2X2_831 ( .A(_abc_17692_n2784), .B(_abc_17692_n2790), .Y(_abc_17692_n2791) );
  OR2X2 OR2X2_832 ( .A(_abc_17692_n2792), .B(_abc_17692_n2769), .Y(_abc_17692_n2793) );
  OR2X2 OR2X2_833 ( .A(_abc_17692_n2795), .B(_abc_17692_n2794), .Y(_abc_17692_n2796) );
  OR2X2 OR2X2_834 ( .A(_abc_17692_n2796), .B(_abc_17692_n2764), .Y(_abc_17692_n2797_1) );
  OR2X2 OR2X2_835 ( .A(_abc_17692_n2801), .B(_abc_17692_n2733), .Y(_abc_17692_n2802) );
  OR2X2 OR2X2_836 ( .A(_abc_17692_n2803), .B(_abc_17692_n2546), .Y(_abc_17692_n2804) );
  OR2X2 OR2X2_837 ( .A(_abc_17692_n2804), .B(_abc_17692_n2732), .Y(_abc_17692_n2805) );
  OR2X2 OR2X2_838 ( .A(_abc_17692_n2799), .B(_abc_17692_n2807), .Y(_abc_17692_n2808) );
  OR2X2 OR2X2_839 ( .A(_abc_17692_n2791), .B(_abc_17692_n2808), .Y(_abc_17692_n2809) );
  OR2X2 OR2X2_84 ( .A(_abc_17692_n725_bF_buf1), .B(_auto_iopadmap_cc_313_execute_30065_21_), .Y(_abc_17692_n790) );
  OR2X2 OR2X2_840 ( .A(_abc_17692_n2811), .B(_abc_17692_n2812_1), .Y(_abc_17692_n2813) );
  OR2X2 OR2X2_841 ( .A(_abc_17692_n2810), .B(_abc_17692_n2813), .Y(_abc_17692_n2814) );
  OR2X2 OR2X2_842 ( .A(_abc_17692_n2775), .B(_abc_17692_n2814), .Y(workunit2_5__FF_INPUT) );
  OR2X2 OR2X2_843 ( .A(_abc_17692_n2450), .B(_abc_17692_n2649), .Y(_abc_17692_n2818) );
  OR2X2 OR2X2_844 ( .A(_abc_17692_n2817), .B(_abc_17692_n2819), .Y(_abc_17692_n2820) );
  OR2X2 OR2X2_845 ( .A(_abc_17692_n2824), .B(_abc_17692_n2822), .Y(_abc_17692_n2825) );
  OR2X2 OR2X2_846 ( .A(_abc_17692_n2825), .B(_abc_17692_n2821), .Y(_abc_17692_n2826) );
  OR2X2 OR2X2_847 ( .A(workunit1_2_), .B(workunit1_11_bF_buf0), .Y(_abc_17692_n2828) );
  OR2X2 OR2X2_848 ( .A(_abc_17692_n2829), .B(workunit1_6_), .Y(_abc_17692_n2830_1) );
  OR2X2 OR2X2_849 ( .A(_abc_17692_n2438), .B(_abc_17692_n2650), .Y(_abc_17692_n2834) );
  OR2X2 OR2X2_85 ( .A(_abc_17692_n727_bF_buf2), .B(workunit2_21_), .Y(_abc_17692_n791) );
  OR2X2 OR2X2_850 ( .A(_abc_17692_n2838), .B(_abc_17692_n2837), .Y(_abc_17692_n2839) );
  OR2X2 OR2X2_851 ( .A(_abc_17692_n2840), .B(_abc_17692_n2832), .Y(_abc_17692_n2841) );
  OR2X2 OR2X2_852 ( .A(_abc_17692_n2659), .B(_abc_17692_n2496), .Y(_abc_17692_n2845) );
  OR2X2 OR2X2_853 ( .A(_abc_17692_n2844), .B(_abc_17692_n2847), .Y(_abc_17692_n2848) );
  OR2X2 OR2X2_854 ( .A(sum_6_), .B(\key_in[70] ), .Y(_abc_17692_n2851) );
  OR2X2 OR2X2_855 ( .A(_abc_17692_n2848), .B(_abc_17692_n2852), .Y(_abc_17692_n2855) );
  OR2X2 OR2X2_856 ( .A(_abc_17692_n2858), .B(_abc_17692_n2859), .Y(_abc_17692_n2860) );
  OR2X2 OR2X2_857 ( .A(_abc_17692_n2864), .B(_abc_17692_n2861), .Y(_abc_17692_n2865) );
  OR2X2 OR2X2_858 ( .A(_abc_17692_n2678), .B(_abc_17692_n2866), .Y(_abc_17692_n2867_1) );
  OR2X2 OR2X2_859 ( .A(_abc_17692_n2867_1), .B(_abc_17692_n2865), .Y(_abc_17692_n2868) );
  OR2X2 OR2X2_86 ( .A(_abc_17692_n725_bF_buf0), .B(_auto_iopadmap_cc_313_execute_30065_22_), .Y(_abc_17692_n793) );
  OR2X2 OR2X2_860 ( .A(_abc_17692_n2474), .B(_abc_17692_n2687), .Y(_abc_17692_n2873) );
  OR2X2 OR2X2_861 ( .A(_abc_17692_n2465), .B(_abc_17692_n2684), .Y(_abc_17692_n2877) );
  OR2X2 OR2X2_862 ( .A(_abc_17692_n2875), .B(_abc_17692_n2878), .Y(_abc_17692_n2879) );
  OR2X2 OR2X2_863 ( .A(sum_6_), .B(\key_in[6] ), .Y(_abc_17692_n2882) );
  OR2X2 OR2X2_864 ( .A(_abc_17692_n2887), .B(_abc_17692_n2884), .Y(_abc_17692_n2888) );
  OR2X2 OR2X2_865 ( .A(_abc_17692_n2891), .B(_abc_17692_n2889), .Y(_abc_17692_n2892) );
  OR2X2 OR2X2_866 ( .A(_abc_17692_n2892), .B(workunit2_6_), .Y(_abc_17692_n2895) );
  OR2X2 OR2X2_867 ( .A(_abc_17692_n2897), .B(_abc_17692_n2896), .Y(_abc_17692_n2898) );
  OR2X2 OR2X2_868 ( .A(_abc_17692_n2901), .B(_abc_17692_n2900), .Y(_abc_17692_n2902) );
  OR2X2 OR2X2_869 ( .A(_abc_17692_n2902), .B(_abc_17692_n2899), .Y(_abc_17692_n2903) );
  OR2X2 OR2X2_87 ( .A(_abc_17692_n727_bF_buf1), .B(workunit2_22_), .Y(_abc_17692_n794) );
  OR2X2 OR2X2_870 ( .A(_abc_17692_n2530), .B(_abc_17692_n2712), .Y(_abc_17692_n2909) );
  OR2X2 OR2X2_871 ( .A(_abc_17692_n2907), .B(_abc_17692_n2910), .Y(_abc_17692_n2911) );
  OR2X2 OR2X2_872 ( .A(sum_6_), .B(\key_in[38] ), .Y(_abc_17692_n2914) );
  OR2X2 OR2X2_873 ( .A(_abc_17692_n2538_1), .B(_abc_17692_n2917), .Y(_abc_17692_n2918) );
  OR2X2 OR2X2_874 ( .A(_abc_17692_n2922), .B(_abc_17692_n2916_1), .Y(_abc_17692_n2923) );
  OR2X2 OR2X2_875 ( .A(_abc_17692_n2924), .B(_abc_17692_n2926_1), .Y(_abc_17692_n2927) );
  OR2X2 OR2X2_876 ( .A(_abc_17692_n2928), .B(_abc_17692_n2862), .Y(_abc_17692_n2929) );
  OR2X2 OR2X2_877 ( .A(_abc_17692_n2927), .B(workunit2_6_), .Y(_abc_17692_n2930) );
  OR2X2 OR2X2_878 ( .A(_abc_17692_n2732), .B(_abc_17692_n2618), .Y(_abc_17692_n2933) );
  OR2X2 OR2X2_879 ( .A(_abc_17692_n2933), .B(_abc_17692_n2550), .Y(_abc_17692_n2934) );
  OR2X2 OR2X2_88 ( .A(_abc_17692_n725_bF_buf7), .B(_auto_iopadmap_cc_313_execute_30065_23_), .Y(_abc_17692_n796) );
  OR2X2 OR2X2_880 ( .A(_abc_17692_n2732), .B(_abc_17692_n2937), .Y(_abc_17692_n2938_1) );
  OR2X2 OR2X2_881 ( .A(_abc_17692_n2941), .B(_abc_17692_n2932), .Y(_abc_17692_n2942) );
  OR2X2 OR2X2_882 ( .A(_abc_17692_n2905), .B(_abc_17692_n2946), .Y(_abc_17692_n2947) );
  OR2X2 OR2X2_883 ( .A(_abc_17692_n2947), .B(_abc_17692_n2872), .Y(_abc_17692_n2948) );
  OR2X2 OR2X2_884 ( .A(_abc_17692_n2750), .B(_abc_17692_n2561), .Y(_abc_17692_n2951) );
  OR2X2 OR2X2_885 ( .A(_abc_17692_n2950), .B(_abc_17692_n2953), .Y(_abc_17692_n2954) );
  OR2X2 OR2X2_886 ( .A(sum_6_), .B(\key_in[102] ), .Y(_abc_17692_n2957) );
  OR2X2 OR2X2_887 ( .A(_abc_17692_n2954), .B(_abc_17692_n2958), .Y(_abc_17692_n2961) );
  OR2X2 OR2X2_888 ( .A(_abc_17692_n2964), .B(_abc_17692_n2965), .Y(_abc_17692_n2966) );
  OR2X2 OR2X2_889 ( .A(_abc_17692_n2966), .B(_abc_17692_n2862), .Y(_abc_17692_n2967) );
  OR2X2 OR2X2_89 ( .A(_abc_17692_n727_bF_buf0), .B(workunit2_23_), .Y(_abc_17692_n797) );
  OR2X2 OR2X2_890 ( .A(_abc_17692_n2968), .B(workunit2_6_), .Y(_abc_17692_n2969) );
  OR2X2 OR2X2_891 ( .A(_abc_17692_n2972), .B(_abc_17692_n2970), .Y(_abc_17692_n2973) );
  OR2X2 OR2X2_892 ( .A(_abc_17692_n2971), .B(_abc_17692_n2974), .Y(_abc_17692_n2975) );
  OR2X2 OR2X2_893 ( .A(_abc_17692_n2948), .B(_abc_17692_n2977), .Y(_abc_17692_n2978) );
  OR2X2 OR2X2_894 ( .A(_abc_17692_n2697), .B(_abc_17692_n2633), .Y(_abc_17692_n2980) );
  OR2X2 OR2X2_895 ( .A(_abc_17692_n2786), .B(_abc_17692_n2981), .Y(_abc_17692_n2982) );
  OR2X2 OR2X2_896 ( .A(_abc_17692_n2982), .B(_abc_17692_n2896), .Y(_abc_17692_n2985) );
  OR2X2 OR2X2_897 ( .A(_abc_17692_n2989), .B(_abc_17692_n2988), .Y(_abc_17692_n2990) );
  OR2X2 OR2X2_898 ( .A(_abc_17692_n2990), .B(_abc_17692_n2931), .Y(_abc_17692_n2991) );
  OR2X2 OR2X2_899 ( .A(_abc_17692_n2995_1), .B(_abc_17692_n2987), .Y(_abc_17692_n2996) );
  OR2X2 OR2X2_9 ( .A(state_8_bF_buf2), .B(delta_7_), .Y(delta_7__FF_INPUT) );
  OR2X2 OR2X2_90 ( .A(_abc_17692_n725_bF_buf6), .B(_auto_iopadmap_cc_313_execute_30065_24_), .Y(_abc_17692_n799_1) );
  OR2X2 OR2X2_900 ( .A(_abc_17692_n2997), .B(_abc_17692_n2970), .Y(_abc_17692_n2998_1) );
  OR2X2 OR2X2_901 ( .A(_abc_17692_n3000), .B(_abc_17692_n2999), .Y(_abc_17692_n3001) );
  OR2X2 OR2X2_902 ( .A(_abc_17692_n3001), .B(_abc_17692_n2974), .Y(_abc_17692_n3002) );
  OR2X2 OR2X2_903 ( .A(_abc_17692_n2670), .B(_abc_17692_n2633), .Y(_abc_17692_n3005) );
  OR2X2 OR2X2_904 ( .A(_abc_17692_n3006), .B(_abc_17692_n2865), .Y(_abc_17692_n3007) );
  OR2X2 OR2X2_905 ( .A(_abc_17692_n3010), .B(_abc_17692_n3009_1), .Y(_abc_17692_n3011) );
  OR2X2 OR2X2_906 ( .A(_abc_17692_n3011), .B(_abc_17692_n3008), .Y(_abc_17692_n3012) );
  OR2X2 OR2X2_907 ( .A(_abc_17692_n3004), .B(_abc_17692_n3014), .Y(_abc_17692_n3015) );
  OR2X2 OR2X2_908 ( .A(_abc_17692_n2996), .B(_abc_17692_n3015), .Y(_abc_17692_n3016) );
  OR2X2 OR2X2_909 ( .A(_abc_17692_n3018), .B(_abc_17692_n3019), .Y(_abc_17692_n3020) );
  OR2X2 OR2X2_91 ( .A(_abc_17692_n727_bF_buf7), .B(workunit2_24_), .Y(_abc_17692_n800) );
  OR2X2 OR2X2_910 ( .A(_abc_17692_n3017), .B(_abc_17692_n3020), .Y(_abc_17692_n3021) );
  OR2X2 OR2X2_911 ( .A(_abc_17692_n3021), .B(_abc_17692_n2979), .Y(workunit2_6__FF_INPUT) );
  OR2X2 OR2X2_912 ( .A(_abc_17692_n3027), .B(_abc_17692_n3025), .Y(_abc_17692_n3028) );
  OR2X2 OR2X2_913 ( .A(_abc_17692_n3028), .B(_abc_17692_n2063), .Y(_abc_17692_n3029) );
  OR2X2 OR2X2_914 ( .A(workunit1_3_), .B(workunit1_12_bF_buf0), .Y(_abc_17692_n3031) );
  OR2X2 OR2X2_915 ( .A(_abc_17692_n3032), .B(workunit1_7_), .Y(_abc_17692_n3033) );
  OR2X2 OR2X2_916 ( .A(_abc_17692_n2832), .B(_abc_17692_n2837), .Y(_abc_17692_n3036) );
  OR2X2 OR2X2_917 ( .A(_abc_17692_n3038), .B(_abc_17692_n3037), .Y(_abc_17692_n3039) );
  OR2X2 OR2X2_918 ( .A(_abc_17692_n3035), .B(_abc_17692_n3040), .Y(_abc_17692_n3041) );
  OR2X2 OR2X2_919 ( .A(_abc_17692_n2884), .B(_abc_17692_n2880), .Y(_abc_17692_n3042) );
  OR2X2 OR2X2_92 ( .A(_abc_17692_n725_bF_buf5), .B(_auto_iopadmap_cc_313_execute_30065_25_), .Y(_abc_17692_n802) );
  OR2X2 OR2X2_920 ( .A(sum_7_), .B(\key_in[7] ), .Y(_abc_17692_n3046) );
  OR2X2 OR2X2_921 ( .A(_abc_17692_n3048), .B(_abc_17692_n3050), .Y(_abc_17692_n3051) );
  OR2X2 OR2X2_922 ( .A(_abc_17692_n3036), .B(_abc_17692_n3039), .Y(_abc_17692_n3053) );
  OR2X2 OR2X2_923 ( .A(_abc_17692_n3057), .B(_abc_17692_n3052), .Y(_abc_17692_n3058_1) );
  OR2X2 OR2X2_924 ( .A(_abc_17692_n3062), .B(_abc_17692_n3059), .Y(_abc_17692_n3063) );
  OR2X2 OR2X2_925 ( .A(_abc_17692_n2892), .B(_abc_17692_n2862), .Y(_abc_17692_n3065) );
  OR2X2 OR2X2_926 ( .A(_abc_17692_n3067), .B(_abc_17692_n3064), .Y(_abc_17692_n3068) );
  OR2X2 OR2X2_927 ( .A(_abc_17692_n3066), .B(_abc_17692_n3063), .Y(_abc_17692_n3069) );
  OR2X2 OR2X2_928 ( .A(_abc_17692_n2853), .B(_abc_17692_n2849_1), .Y(_abc_17692_n3072) );
  OR2X2 OR2X2_929 ( .A(sum_7_), .B(\key_in[71] ), .Y(_abc_17692_n3075) );
  OR2X2 OR2X2_93 ( .A(_abc_17692_n727_bF_buf6), .B(workunit2_25_), .Y(_abc_17692_n803) );
  OR2X2 OR2X2_930 ( .A(_abc_17692_n3072), .B(_abc_17692_n3077), .Y(_abc_17692_n3078) );
  OR2X2 OR2X2_931 ( .A(_abc_17692_n3083), .B(_abc_17692_n3084), .Y(_abc_17692_n3085) );
  OR2X2 OR2X2_932 ( .A(_abc_17692_n3086), .B(_abc_17692_n3060), .Y(_abc_17692_n3087) );
  OR2X2 OR2X2_933 ( .A(_abc_17692_n3085), .B(workunit2_7_), .Y(_abc_17692_n3088) );
  OR2X2 OR2X2_934 ( .A(_abc_17692_n2869), .B(_abc_17692_n3091), .Y(_abc_17692_n3092) );
  OR2X2 OR2X2_935 ( .A(_abc_17692_n3093), .B(_abc_17692_n3090), .Y(_abc_17692_n3094) );
  OR2X2 OR2X2_936 ( .A(_abc_17692_n3092), .B(_abc_17692_n3089), .Y(_abc_17692_n3095) );
  OR2X2 OR2X2_937 ( .A(_abc_17692_n2920), .B(_abc_17692_n2921), .Y(_abc_17692_n3098) );
  OR2X2 OR2X2_938 ( .A(sum_7_), .B(\key_in[39] ), .Y(_abc_17692_n3102) );
  OR2X2 OR2X2_939 ( .A(_abc_17692_n2916_1), .B(_abc_17692_n2912), .Y(_abc_17692_n3105) );
  OR2X2 OR2X2_94 ( .A(_abc_17692_n725_bF_buf4), .B(_auto_iopadmap_cc_313_execute_30065_26_), .Y(_abc_17692_n805) );
  OR2X2 OR2X2_940 ( .A(_abc_17692_n3104), .B(_abc_17692_n3107), .Y(_abc_17692_n3108) );
  OR2X2 OR2X2_941 ( .A(_abc_17692_n3055), .B(_abc_17692_n3108), .Y(_abc_17692_n3109) );
  OR2X2 OR2X2_942 ( .A(_abc_17692_n3105), .B(_abc_17692_n3106), .Y(_abc_17692_n3110) );
  OR2X2 OR2X2_943 ( .A(_abc_17692_n3099), .B(_abc_17692_n3103), .Y(_abc_17692_n3111) );
  OR2X2 OR2X2_944 ( .A(_abc_17692_n3041), .B(_abc_17692_n3112), .Y(_abc_17692_n3113) );
  OR2X2 OR2X2_945 ( .A(_abc_17692_n3055), .B(_abc_17692_n3112), .Y(_abc_17692_n3116) );
  OR2X2 OR2X2_946 ( .A(_abc_17692_n3041), .B(_abc_17692_n3108), .Y(_abc_17692_n3117) );
  OR2X2 OR2X2_947 ( .A(_abc_17692_n3115), .B(_abc_17692_n3119), .Y(_abc_17692_n3120) );
  OR2X2 OR2X2_948 ( .A(_abc_17692_n3125), .B(_abc_17692_n3121), .Y(_abc_17692_n3126) );
  OR2X2 OR2X2_949 ( .A(_abc_17692_n3124), .B(_abc_17692_n3120), .Y(_abc_17692_n3127) );
  OR2X2 OR2X2_95 ( .A(_abc_17692_n727_bF_buf5), .B(workunit2_26_), .Y(_abc_17692_n806) );
  OR2X2 OR2X2_950 ( .A(_abc_17692_n3097), .B(_abc_17692_n3129), .Y(_abc_17692_n3130) );
  OR2X2 OR2X2_951 ( .A(_abc_17692_n3130), .B(_abc_17692_n3071), .Y(_abc_17692_n3131) );
  OR2X2 OR2X2_952 ( .A(_abc_17692_n2959), .B(_abc_17692_n2955), .Y(_abc_17692_n3132) );
  OR2X2 OR2X2_953 ( .A(sum_7_), .B(\key_in[103] ), .Y(_abc_17692_n3135) );
  OR2X2 OR2X2_954 ( .A(_abc_17692_n3132), .B(_abc_17692_n3137), .Y(_abc_17692_n3138) );
  OR2X2 OR2X2_955 ( .A(_abc_17692_n3143), .B(_abc_17692_n3144_1), .Y(_abc_17692_n3145) );
  OR2X2 OR2X2_956 ( .A(_abc_17692_n3146), .B(_abc_17692_n3060), .Y(_abc_17692_n3147) );
  OR2X2 OR2X2_957 ( .A(_abc_17692_n3145), .B(workunit2_7_), .Y(_abc_17692_n3148) );
  OR2X2 OR2X2_958 ( .A(_abc_17692_n3151), .B(_abc_17692_n3149), .Y(_abc_17692_n3152) );
  OR2X2 OR2X2_959 ( .A(_abc_17692_n3150), .B(_abc_17692_n3153_1), .Y(_abc_17692_n3154) );
  OR2X2 OR2X2_96 ( .A(_abc_17692_n725_bF_buf3), .B(_auto_iopadmap_cc_313_execute_30065_27_), .Y(_abc_17692_n808) );
  OR2X2 OR2X2_960 ( .A(_abc_17692_n3131), .B(_abc_17692_n3156), .Y(_abc_17692_n3157) );
  OR2X2 OR2X2_961 ( .A(_abc_17692_n3159), .B(_abc_17692_n3064), .Y(_abc_17692_n3160) );
  OR2X2 OR2X2_962 ( .A(_abc_17692_n3161), .B(_abc_17692_n3063), .Y(_abc_17692_n3162) );
  OR2X2 OR2X2_963 ( .A(_abc_17692_n3166_1), .B(_abc_17692_n3120), .Y(_abc_17692_n3167) );
  OR2X2 OR2X2_964 ( .A(_abc_17692_n3165), .B(_abc_17692_n3121), .Y(_abc_17692_n3168) );
  OR2X2 OR2X2_965 ( .A(_abc_17692_n3164), .B(_abc_17692_n3170), .Y(_abc_17692_n3171) );
  OR2X2 OR2X2_966 ( .A(_abc_17692_n2968), .B(_abc_17692_n2862), .Y(_abc_17692_n3172) );
  OR2X2 OR2X2_967 ( .A(_abc_17692_n3174), .B(_abc_17692_n3173), .Y(_abc_17692_n3175) );
  OR2X2 OR2X2_968 ( .A(_abc_17692_n3175), .B(_abc_17692_n3153_1), .Y(_abc_17692_n3176) );
  OR2X2 OR2X2_969 ( .A(_abc_17692_n3177), .B(_abc_17692_n3149), .Y(_abc_17692_n3178_1) );
  OR2X2 OR2X2_97 ( .A(_abc_17692_n727_bF_buf4), .B(workunit2_27_), .Y(_abc_17692_n809) );
  OR2X2 OR2X2_970 ( .A(_abc_17692_n3090), .B(_abc_17692_n2861), .Y(_abc_17692_n3182) );
  OR2X2 OR2X2_971 ( .A(_abc_17692_n3181), .B(_abc_17692_n3182), .Y(_abc_17692_n3183) );
  OR2X2 OR2X2_972 ( .A(_abc_17692_n3089), .B(_abc_17692_n3184), .Y(_abc_17692_n3185) );
  OR2X2 OR2X2_973 ( .A(_abc_17692_n3007), .B(_abc_17692_n3089), .Y(_abc_17692_n3187) );
  OR2X2 OR2X2_974 ( .A(_abc_17692_n3180), .B(_abc_17692_n3189_1), .Y(_abc_17692_n3190) );
  OR2X2 OR2X2_975 ( .A(_abc_17692_n3171), .B(_abc_17692_n3190), .Y(_abc_17692_n3191) );
  OR2X2 OR2X2_976 ( .A(_abc_17692_n3193), .B(_abc_17692_n3194), .Y(_abc_17692_n3195) );
  OR2X2 OR2X2_977 ( .A(_abc_17692_n3192), .B(_abc_17692_n3195), .Y(_abc_17692_n3196) );
  OR2X2 OR2X2_978 ( .A(_abc_17692_n3196), .B(_abc_17692_n3158), .Y(workunit2_7__FF_INPUT) );
  OR2X2 OR2X2_979 ( .A(_abc_17692_n3203), .B(_abc_17692_n3038), .Y(_abc_17692_n3204) );
  OR2X2 OR2X2_98 ( .A(_abc_17692_n725_bF_buf2), .B(_auto_iopadmap_cc_313_execute_30065_28_), .Y(_abc_17692_n811) );
  OR2X2 OR2X2_980 ( .A(_abc_17692_n3202), .B(_abc_17692_n3205), .Y(_abc_17692_n3206) );
  OR2X2 OR2X2_981 ( .A(_abc_17692_n3206), .B(_abc_17692_n3201), .Y(_abc_17692_n3207) );
  OR2X2 OR2X2_982 ( .A(_abc_17692_n3209), .B(_abc_17692_n3210), .Y(_abc_17692_n3211) );
  OR2X2 OR2X2_983 ( .A(_abc_17692_n2433), .B(workunit1_13_bF_buf0), .Y(_abc_17692_n3213) );
  OR2X2 OR2X2_984 ( .A(_abc_17692_n3208), .B(workunit1_4_), .Y(_abc_17692_n3214) );
  OR2X2 OR2X2_985 ( .A(_abc_17692_n3212), .B(_abc_17692_n3216), .Y(_abc_17692_n3217) );
  OR2X2 OR2X2_986 ( .A(_abc_17692_n2452), .B(_abc_17692_n2651), .Y(_abc_17692_n3220) );
  OR2X2 OR2X2_987 ( .A(_abc_17692_n2839), .B(_abc_17692_n3039), .Y(_abc_17692_n3221) );
  OR2X2 OR2X2_988 ( .A(_abc_17692_n3220), .B(_abc_17692_n3221), .Y(_abc_17692_n3222) );
  OR2X2 OR2X2_989 ( .A(_abc_17692_n3222), .B(_abc_17692_n2456), .Y(_abc_17692_n3223) );
  OR2X2 OR2X2_99 ( .A(_abc_17692_n727_bF_buf3), .B(workunit2_28_), .Y(_abc_17692_n812) );
  OR2X2 OR2X2_990 ( .A(_abc_17692_n3221), .B(_abc_17692_n2835), .Y(_abc_17692_n3224_1) );
  OR2X2 OR2X2_991 ( .A(_abc_17692_n3227_1), .B(_abc_17692_n3219), .Y(_abc_17692_n3228) );
  OR2X2 OR2X2_992 ( .A(_abc_17692_n3233), .B(_abc_17692_n3073), .Y(_abc_17692_n3234) );
  OR2X2 OR2X2_993 ( .A(_abc_17692_n3232), .B(_abc_17692_n3234), .Y(_abc_17692_n3235) );
  OR2X2 OR2X2_994 ( .A(_abc_17692_n3235), .B(_abc_17692_n3231), .Y(_abc_17692_n3236) );
  OR2X2 OR2X2_995 ( .A(sum_8_), .B(\key_in[72] ), .Y(_abc_17692_n3239) );
  OR2X2 OR2X2_996 ( .A(_abc_17692_n3244), .B(_abc_17692_n3241), .Y(_abc_17692_n3245) );
  OR2X2 OR2X2_997 ( .A(_abc_17692_n3246), .B(_abc_17692_n3228), .Y(_abc_17692_n3247) );
  OR2X2 OR2X2_998 ( .A(_abc_17692_n3248), .B(_abc_17692_n3245), .Y(_abc_17692_n3249) );
  OR2X2 OR2X2_999 ( .A(_abc_17692_n3252), .B(_abc_17692_n3253), .Y(_abc_17692_n3254) );
endmodule
