module b14_reset(clock, RESET_G, nRESET_G, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, ADDR_REG_19_, ADDR_REG_18_, ADDR_REG_17_, ADDR_REG_16_, ADDR_REG_15_, ADDR_REG_14_, ADDR_REG_13_, ADDR_REG_12_, ADDR_REG_11_, ADDR_REG_10_, ADDR_REG_9_, ADDR_REG_8_, ADDR_REG_7_, ADDR_REG_6_, ADDR_REG_5_, ADDR_REG_4_, ADDR_REG_3_, ADDR_REG_2_, ADDR_REG_1_, ADDR_REG_0_, DATAO_REG_31_, DATAO_REG_30_, DATAO_REG_29_, DATAO_REG_28_, DATAO_REG_27_, DATAO_REG_26_, DATAO_REG_25_, DATAO_REG_24_, DATAO_REG_23_, DATAO_REG_22_, DATAO_REG_21_, DATAO_REG_20_, DATAO_REG_19_, DATAO_REG_18_, DATAO_REG_17_, DATAO_REG_16_, DATAO_REG_15_, DATAO_REG_14_, DATAO_REG_13_, DATAO_REG_12_, DATAO_REG_11_, DATAO_REG_10_, DATAO_REG_9_, DATAO_REG_8_, DATAO_REG_7_, DATAO_REG_6_, DATAO_REG_5_, DATAO_REG_4_, DATAO_REG_3_, DATAO_REG_2_, DATAO_REG_1_, DATAO_REG_0_, RD_REG, WR_REG);

output ADDR_REG_0_;
output ADDR_REG_10_;
output ADDR_REG_11_;
output ADDR_REG_12_;
output ADDR_REG_13_;
output ADDR_REG_14_;
output ADDR_REG_15_;
output ADDR_REG_16_;
output ADDR_REG_17_;
output ADDR_REG_18_;
output ADDR_REG_19_;
output ADDR_REG_1_;
output ADDR_REG_2_;
output ADDR_REG_3_;
output ADDR_REG_4_;
output ADDR_REG_5_;
output ADDR_REG_6_;
output ADDR_REG_7_;
output ADDR_REG_8_;
output ADDR_REG_9_;
wire B_REG; 
input DATAI_0_;
input DATAI_10_;
input DATAI_11_;
input DATAI_12_;
input DATAI_13_;
input DATAI_14_;
input DATAI_15_;
input DATAI_16_;
input DATAI_17_;
input DATAI_18_;
input DATAI_19_;
input DATAI_1_;
input DATAI_20_;
input DATAI_21_;
input DATAI_22_;
input DATAI_23_;
input DATAI_24_;
input DATAI_25_;
input DATAI_26_;
input DATAI_27_;
input DATAI_28_;
input DATAI_29_;
input DATAI_2_;
input DATAI_30_;
input DATAI_31_;
input DATAI_3_;
input DATAI_4_;
input DATAI_5_;
input DATAI_6_;
input DATAI_7_;
input DATAI_8_;
input DATAI_9_;
output DATAO_REG_0_;
output DATAO_REG_10_;
output DATAO_REG_11_;
output DATAO_REG_12_;
output DATAO_REG_13_;
output DATAO_REG_14_;
output DATAO_REG_15_;
output DATAO_REG_16_;
output DATAO_REG_17_;
output DATAO_REG_18_;
output DATAO_REG_19_;
output DATAO_REG_1_;
output DATAO_REG_20_;
output DATAO_REG_21_;
output DATAO_REG_22_;
output DATAO_REG_23_;
output DATAO_REG_24_;
output DATAO_REG_25_;
output DATAO_REG_26_;
output DATAO_REG_27_;
output DATAO_REG_28_;
output DATAO_REG_29_;
output DATAO_REG_2_;
output DATAO_REG_30_;
output DATAO_REG_31_;
output DATAO_REG_3_;
output DATAO_REG_4_;
output DATAO_REG_5_;
output DATAO_REG_6_;
output DATAO_REG_7_;
output DATAO_REG_8_;
output DATAO_REG_9_;
wire D_REG_0_; 
wire D_REG_10_; 
wire D_REG_11_; 
wire D_REG_12_; 
wire D_REG_13_; 
wire D_REG_14_; 
wire D_REG_15_; 
wire D_REG_16_; 
wire D_REG_17_; 
wire D_REG_18_; 
wire D_REG_19_; 
wire D_REG_1_; 
wire D_REG_20_; 
wire D_REG_21_; 
wire D_REG_22_; 
wire D_REG_23_; 
wire D_REG_24_; 
wire D_REG_25_; 
wire D_REG_26_; 
wire D_REG_27_; 
wire D_REG_28_; 
wire D_REG_29_; 
wire D_REG_2_; 
wire D_REG_30_; 
wire D_REG_31_; 
wire D_REG_3_; 
wire D_REG_4_; 
wire D_REG_5_; 
wire D_REG_6_; 
wire D_REG_7_; 
wire D_REG_8_; 
wire D_REG_9_; 
wire IR_REG_0_; 
wire IR_REG_10_; 
wire IR_REG_11_; 
wire IR_REG_12_; 
wire IR_REG_13_; 
wire IR_REG_14_; 
wire IR_REG_15_; 
wire IR_REG_16_; 
wire IR_REG_17_; 
wire IR_REG_18_; 
wire IR_REG_19_; 
wire IR_REG_1_; 
wire IR_REG_20_; 
wire IR_REG_21_; 
wire IR_REG_22_; 
wire IR_REG_23_; 
wire IR_REG_24_; 
wire IR_REG_25_; 
wire IR_REG_26_; 
wire IR_REG_27_; 
wire IR_REG_28_; 
wire IR_REG_29_; 
wire IR_REG_2_; 
wire IR_REG_30_; 
wire IR_REG_31_; 
wire IR_REG_3_; 
wire IR_REG_4_; 
wire IR_REG_5_; 
wire IR_REG_6_; 
wire IR_REG_7_; 
wire IR_REG_8_; 
wire IR_REG_9_; 
output RD_REG;
wire REG0_REG_0_; 
wire REG0_REG_10_; 
wire REG0_REG_11_; 
wire REG0_REG_12_; 
wire REG0_REG_13_; 
wire REG0_REG_14_; 
wire REG0_REG_15_; 
wire REG0_REG_16_; 
wire REG0_REG_17_; 
wire REG0_REG_18_; 
wire REG0_REG_19_; 
wire REG0_REG_1_; 
wire REG0_REG_20_; 
wire REG0_REG_21_; 
wire REG0_REG_22_; 
wire REG0_REG_23_; 
wire REG0_REG_24_; 
wire REG0_REG_25_; 
wire REG0_REG_26_; 
wire REG0_REG_27_; 
wire REG0_REG_28_; 
wire REG0_REG_29_; 
wire REG0_REG_2_; 
wire REG0_REG_30_; 
wire REG0_REG_31_; 
wire REG0_REG_3_; 
wire REG0_REG_4_; 
wire REG0_REG_5_; 
wire REG0_REG_6_; 
wire REG0_REG_7_; 
wire REG0_REG_8_; 
wire REG0_REG_9_; 
wire REG1_REG_0_; 
wire REG1_REG_10_; 
wire REG1_REG_11_; 
wire REG1_REG_12_; 
wire REG1_REG_13_; 
wire REG1_REG_14_; 
wire REG1_REG_15_; 
wire REG1_REG_16_; 
wire REG1_REG_17_; 
wire REG1_REG_18_; 
wire REG1_REG_19_; 
wire REG1_REG_1_; 
wire REG1_REG_20_; 
wire REG1_REG_21_; 
wire REG1_REG_22_; 
wire REG1_REG_23_; 
wire REG1_REG_24_; 
wire REG1_REG_25_; 
wire REG1_REG_26_; 
wire REG1_REG_27_; 
wire REG1_REG_28_; 
wire REG1_REG_29_; 
wire REG1_REG_2_; 
wire REG1_REG_30_; 
wire REG1_REG_31_; 
wire REG1_REG_3_; 
wire REG1_REG_4_; 
wire REG1_REG_5_; 
wire REG1_REG_6_; 
wire REG1_REG_7_; 
wire REG1_REG_8_; 
wire REG1_REG_9_; 
wire REG2_REG_0_; 
wire REG2_REG_10_; 
wire REG2_REG_11_; 
wire REG2_REG_12_; 
wire REG2_REG_13_; 
wire REG2_REG_14_; 
wire REG2_REG_15_; 
wire REG2_REG_16_; 
wire REG2_REG_17_; 
wire REG2_REG_18_; 
wire REG2_REG_19_; 
wire REG2_REG_1_; 
wire REG2_REG_20_; 
wire REG2_REG_21_; 
wire REG2_REG_22_; 
wire REG2_REG_23_; 
wire REG2_REG_24_; 
wire REG2_REG_25_; 
wire REG2_REG_26_; 
wire REG2_REG_27_; 
wire REG2_REG_28_; 
wire REG2_REG_29_; 
wire REG2_REG_2_; 
wire REG2_REG_30_; 
wire REG2_REG_31_; 
wire REG2_REG_3_; 
wire REG2_REG_4_; 
wire REG2_REG_5_; 
wire REG2_REG_6_; 
wire REG2_REG_7_; 
wire REG2_REG_8_; 
wire REG2_REG_9_; 
wire REG3_REG_0_; 
wire REG3_REG_10_; 
wire REG3_REG_11_; 
wire REG3_REG_12_; 
wire REG3_REG_13_; 
wire REG3_REG_14_; 
wire REG3_REG_15_; 
wire REG3_REG_16_; 
wire REG3_REG_17_; 
wire REG3_REG_18_; 
wire REG3_REG_19_; 
wire REG3_REG_1_; 
wire REG3_REG_20_; 
wire REG3_REG_21_; 
wire REG3_REG_22_; 
wire REG3_REG_23_; 
wire REG3_REG_24_; 
wire REG3_REG_25_; 
wire REG3_REG_26_; 
wire REG3_REG_27_; 
wire REG3_REG_28_; 
wire REG3_REG_2_; 
wire REG3_REG_3_; 
wire REG3_REG_4_; 
wire REG3_REG_5_; 
wire REG3_REG_6_; 
wire REG3_REG_7_; 
wire REG3_REG_8_; 
wire REG3_REG_9_; 
input RESET_G;
wire STATE_REG; 
output WR_REG;
wire _abc_40319_new_n1000_; 
wire _abc_40319_new_n1001_; 
wire _abc_40319_new_n1002_; 
wire _abc_40319_new_n1003_; 
wire _abc_40319_new_n1004_; 
wire _abc_40319_new_n1005_; 
wire _abc_40319_new_n1006_; 
wire _abc_40319_new_n1007_; 
wire _abc_40319_new_n1008_; 
wire _abc_40319_new_n1009_; 
wire _abc_40319_new_n1010_; 
wire _abc_40319_new_n1011_; 
wire _abc_40319_new_n1012_; 
wire _abc_40319_new_n1013_; 
wire _abc_40319_new_n1014_; 
wire _abc_40319_new_n1015_; 
wire _abc_40319_new_n1016_; 
wire _abc_40319_new_n1017_; 
wire _abc_40319_new_n1018_; 
wire _abc_40319_new_n1019_; 
wire _abc_40319_new_n1020_; 
wire _abc_40319_new_n1021_; 
wire _abc_40319_new_n1022_; 
wire _abc_40319_new_n1023_; 
wire _abc_40319_new_n1024_; 
wire _abc_40319_new_n1025_; 
wire _abc_40319_new_n1026_; 
wire _abc_40319_new_n1027_; 
wire _abc_40319_new_n1028_; 
wire _abc_40319_new_n1029_; 
wire _abc_40319_new_n1030_; 
wire _abc_40319_new_n1031_; 
wire _abc_40319_new_n1032_; 
wire _abc_40319_new_n1033_; 
wire _abc_40319_new_n1034_; 
wire _abc_40319_new_n1035_; 
wire _abc_40319_new_n1036_; 
wire _abc_40319_new_n1037_; 
wire _abc_40319_new_n1038_; 
wire _abc_40319_new_n1039_; 
wire _abc_40319_new_n1040_; 
wire _abc_40319_new_n1041_; 
wire _abc_40319_new_n1042_; 
wire _abc_40319_new_n1043_; 
wire _abc_40319_new_n1044_; 
wire _abc_40319_new_n1045_; 
wire _abc_40319_new_n1046_; 
wire _abc_40319_new_n1047_; 
wire _abc_40319_new_n1048_; 
wire _abc_40319_new_n1049_; 
wire _abc_40319_new_n1050_; 
wire _abc_40319_new_n1051_; 
wire _abc_40319_new_n1052_; 
wire _abc_40319_new_n1053_; 
wire _abc_40319_new_n1054_; 
wire _abc_40319_new_n1055_; 
wire _abc_40319_new_n1056_; 
wire _abc_40319_new_n1057_; 
wire _abc_40319_new_n1058_; 
wire _abc_40319_new_n1059_; 
wire _abc_40319_new_n1060_; 
wire _abc_40319_new_n1061_; 
wire _abc_40319_new_n1062_; 
wire _abc_40319_new_n1063_; 
wire _abc_40319_new_n1064_; 
wire _abc_40319_new_n1065_; 
wire _abc_40319_new_n1066_; 
wire _abc_40319_new_n1067_; 
wire _abc_40319_new_n1068_; 
wire _abc_40319_new_n1069_; 
wire _abc_40319_new_n1070_; 
wire _abc_40319_new_n1071_; 
wire _abc_40319_new_n1072_; 
wire _abc_40319_new_n1073_; 
wire _abc_40319_new_n1074_; 
wire _abc_40319_new_n1075_; 
wire _abc_40319_new_n1076_; 
wire _abc_40319_new_n1077_; 
wire _abc_40319_new_n1078_; 
wire _abc_40319_new_n1079_; 
wire _abc_40319_new_n1080_; 
wire _abc_40319_new_n1081_; 
wire _abc_40319_new_n1082_; 
wire _abc_40319_new_n1083_; 
wire _abc_40319_new_n1084_; 
wire _abc_40319_new_n1085_; 
wire _abc_40319_new_n1086_; 
wire _abc_40319_new_n1087_; 
wire _abc_40319_new_n1088_; 
wire _abc_40319_new_n1089_; 
wire _abc_40319_new_n1090_; 
wire _abc_40319_new_n1091_; 
wire _abc_40319_new_n1092_; 
wire _abc_40319_new_n1093_; 
wire _abc_40319_new_n1094_; 
wire _abc_40319_new_n1095_; 
wire _abc_40319_new_n1096_; 
wire _abc_40319_new_n1097_; 
wire _abc_40319_new_n1098_; 
wire _abc_40319_new_n1099_; 
wire _abc_40319_new_n1100_; 
wire _abc_40319_new_n1101_; 
wire _abc_40319_new_n1102_; 
wire _abc_40319_new_n1103_; 
wire _abc_40319_new_n1104_; 
wire _abc_40319_new_n1105_; 
wire _abc_40319_new_n1106_; 
wire _abc_40319_new_n1107_; 
wire _abc_40319_new_n1108_; 
wire _abc_40319_new_n1109_; 
wire _abc_40319_new_n1110_; 
wire _abc_40319_new_n1111_; 
wire _abc_40319_new_n1112_; 
wire _abc_40319_new_n1113_; 
wire _abc_40319_new_n1114_; 
wire _abc_40319_new_n1115_; 
wire _abc_40319_new_n1116_; 
wire _abc_40319_new_n1117_; 
wire _abc_40319_new_n1118_; 
wire _abc_40319_new_n1119_; 
wire _abc_40319_new_n1120_; 
wire _abc_40319_new_n1121_; 
wire _abc_40319_new_n1122_; 
wire _abc_40319_new_n1123_; 
wire _abc_40319_new_n1124_; 
wire _abc_40319_new_n1125_; 
wire _abc_40319_new_n1126_; 
wire _abc_40319_new_n1127_; 
wire _abc_40319_new_n1128_; 
wire _abc_40319_new_n1129_; 
wire _abc_40319_new_n1130_; 
wire _abc_40319_new_n1131_; 
wire _abc_40319_new_n1132_; 
wire _abc_40319_new_n1133_; 
wire _abc_40319_new_n1134_; 
wire _abc_40319_new_n1135_; 
wire _abc_40319_new_n1136_; 
wire _abc_40319_new_n1137_; 
wire _abc_40319_new_n1138_; 
wire _abc_40319_new_n1139_; 
wire _abc_40319_new_n1140_; 
wire _abc_40319_new_n1141_; 
wire _abc_40319_new_n1142_; 
wire _abc_40319_new_n1143_; 
wire _abc_40319_new_n1144_; 
wire _abc_40319_new_n1145_; 
wire _abc_40319_new_n1146_; 
wire _abc_40319_new_n1147_; 
wire _abc_40319_new_n1148_; 
wire _abc_40319_new_n1149_; 
wire _abc_40319_new_n1150_; 
wire _abc_40319_new_n1151_; 
wire _abc_40319_new_n1152_; 
wire _abc_40319_new_n1153_; 
wire _abc_40319_new_n1154_; 
wire _abc_40319_new_n1155_; 
wire _abc_40319_new_n1156_; 
wire _abc_40319_new_n1157_; 
wire _abc_40319_new_n1158_; 
wire _abc_40319_new_n1159_; 
wire _abc_40319_new_n1160_; 
wire _abc_40319_new_n1161_; 
wire _abc_40319_new_n1162_; 
wire _abc_40319_new_n1163_; 
wire _abc_40319_new_n1164_; 
wire _abc_40319_new_n1165_; 
wire _abc_40319_new_n1166_; 
wire _abc_40319_new_n1167_; 
wire _abc_40319_new_n1168_; 
wire _abc_40319_new_n1169_; 
wire _abc_40319_new_n1170_; 
wire _abc_40319_new_n1171_; 
wire _abc_40319_new_n1172_; 
wire _abc_40319_new_n1173_; 
wire _abc_40319_new_n1174_; 
wire _abc_40319_new_n1175_; 
wire _abc_40319_new_n1176_; 
wire _abc_40319_new_n1177_; 
wire _abc_40319_new_n1178_; 
wire _abc_40319_new_n1180_; 
wire _abc_40319_new_n1181_; 
wire _abc_40319_new_n1182_; 
wire _abc_40319_new_n1183_; 
wire _abc_40319_new_n1184_; 
wire _abc_40319_new_n1185_; 
wire _abc_40319_new_n1186_; 
wire _abc_40319_new_n1187_; 
wire _abc_40319_new_n1188_; 
wire _abc_40319_new_n1189_; 
wire _abc_40319_new_n1190_; 
wire _abc_40319_new_n1191_; 
wire _abc_40319_new_n1192_; 
wire _abc_40319_new_n1193_; 
wire _abc_40319_new_n1194_; 
wire _abc_40319_new_n1195_; 
wire _abc_40319_new_n1196_; 
wire _abc_40319_new_n1197_; 
wire _abc_40319_new_n1198_; 
wire _abc_40319_new_n1199_; 
wire _abc_40319_new_n1200_; 
wire _abc_40319_new_n1201_; 
wire _abc_40319_new_n1202_; 
wire _abc_40319_new_n1203_; 
wire _abc_40319_new_n1204_; 
wire _abc_40319_new_n1205_; 
wire _abc_40319_new_n1206_; 
wire _abc_40319_new_n1207_; 
wire _abc_40319_new_n1208_; 
wire _abc_40319_new_n1209_; 
wire _abc_40319_new_n1210_; 
wire _abc_40319_new_n1211_; 
wire _abc_40319_new_n1212_; 
wire _abc_40319_new_n1213_; 
wire _abc_40319_new_n1214_; 
wire _abc_40319_new_n1215_; 
wire _abc_40319_new_n1216_; 
wire _abc_40319_new_n1217_; 
wire _abc_40319_new_n1218_; 
wire _abc_40319_new_n1219_; 
wire _abc_40319_new_n1220_; 
wire _abc_40319_new_n1221_; 
wire _abc_40319_new_n1222_; 
wire _abc_40319_new_n1223_; 
wire _abc_40319_new_n1224_; 
wire _abc_40319_new_n1225_; 
wire _abc_40319_new_n1226_; 
wire _abc_40319_new_n1227_; 
wire _abc_40319_new_n1228_; 
wire _abc_40319_new_n1229_; 
wire _abc_40319_new_n1230_; 
wire _abc_40319_new_n1231_; 
wire _abc_40319_new_n1232_; 
wire _abc_40319_new_n1233_; 
wire _abc_40319_new_n1234_; 
wire _abc_40319_new_n1235_; 
wire _abc_40319_new_n1236_; 
wire _abc_40319_new_n1237_; 
wire _abc_40319_new_n1238_; 
wire _abc_40319_new_n1239_; 
wire _abc_40319_new_n1240_; 
wire _abc_40319_new_n1241_; 
wire _abc_40319_new_n1242_; 
wire _abc_40319_new_n1243_; 
wire _abc_40319_new_n1244_; 
wire _abc_40319_new_n1245_; 
wire _abc_40319_new_n1246_; 
wire _abc_40319_new_n1247_; 
wire _abc_40319_new_n1248_; 
wire _abc_40319_new_n1249_; 
wire _abc_40319_new_n1250_; 
wire _abc_40319_new_n1251_; 
wire _abc_40319_new_n1252_; 
wire _abc_40319_new_n1253_; 
wire _abc_40319_new_n1254_; 
wire _abc_40319_new_n1255_; 
wire _abc_40319_new_n1256_; 
wire _abc_40319_new_n1257_; 
wire _abc_40319_new_n1258_; 
wire _abc_40319_new_n1259_; 
wire _abc_40319_new_n1260_; 
wire _abc_40319_new_n1261_; 
wire _abc_40319_new_n1262_; 
wire _abc_40319_new_n1263_; 
wire _abc_40319_new_n1264_; 
wire _abc_40319_new_n1265_; 
wire _abc_40319_new_n1266_; 
wire _abc_40319_new_n1267_; 
wire _abc_40319_new_n1268_; 
wire _abc_40319_new_n1269_; 
wire _abc_40319_new_n1270_; 
wire _abc_40319_new_n1271_; 
wire _abc_40319_new_n1272_; 
wire _abc_40319_new_n1273_; 
wire _abc_40319_new_n1274_; 
wire _abc_40319_new_n1275_; 
wire _abc_40319_new_n1276_; 
wire _abc_40319_new_n1277_; 
wire _abc_40319_new_n1278_; 
wire _abc_40319_new_n1279_; 
wire _abc_40319_new_n1280_; 
wire _abc_40319_new_n1281_; 
wire _abc_40319_new_n1282_; 
wire _abc_40319_new_n1283_; 
wire _abc_40319_new_n1284_; 
wire _abc_40319_new_n1285_; 
wire _abc_40319_new_n1286_; 
wire _abc_40319_new_n1287_; 
wire _abc_40319_new_n1288_; 
wire _abc_40319_new_n1289_; 
wire _abc_40319_new_n1290_; 
wire _abc_40319_new_n1291_; 
wire _abc_40319_new_n1292_; 
wire _abc_40319_new_n1293_; 
wire _abc_40319_new_n1294_; 
wire _abc_40319_new_n1295_; 
wire _abc_40319_new_n1296_; 
wire _abc_40319_new_n1297_; 
wire _abc_40319_new_n1298_; 
wire _abc_40319_new_n1299_; 
wire _abc_40319_new_n1300_; 
wire _abc_40319_new_n1301_; 
wire _abc_40319_new_n1302_; 
wire _abc_40319_new_n1303_; 
wire _abc_40319_new_n1304_; 
wire _abc_40319_new_n1305_; 
wire _abc_40319_new_n1306_; 
wire _abc_40319_new_n1307_; 
wire _abc_40319_new_n1308_; 
wire _abc_40319_new_n1309_; 
wire _abc_40319_new_n1310_; 
wire _abc_40319_new_n1311_; 
wire _abc_40319_new_n1312_; 
wire _abc_40319_new_n1313_; 
wire _abc_40319_new_n1314_; 
wire _abc_40319_new_n1315_; 
wire _abc_40319_new_n1316_; 
wire _abc_40319_new_n1317_; 
wire _abc_40319_new_n1318_; 
wire _abc_40319_new_n1319_; 
wire _abc_40319_new_n1320_; 
wire _abc_40319_new_n1321_; 
wire _abc_40319_new_n1322_; 
wire _abc_40319_new_n1323_; 
wire _abc_40319_new_n1324_; 
wire _abc_40319_new_n1325_; 
wire _abc_40319_new_n1326_; 
wire _abc_40319_new_n1327_; 
wire _abc_40319_new_n1328_; 
wire _abc_40319_new_n1329_; 
wire _abc_40319_new_n1330_; 
wire _abc_40319_new_n1331_; 
wire _abc_40319_new_n1332_; 
wire _abc_40319_new_n1333_; 
wire _abc_40319_new_n1334_; 
wire _abc_40319_new_n1335_; 
wire _abc_40319_new_n1336_; 
wire _abc_40319_new_n1337_; 
wire _abc_40319_new_n1338_; 
wire _abc_40319_new_n1339_; 
wire _abc_40319_new_n1340_; 
wire _abc_40319_new_n1341_; 
wire _abc_40319_new_n1342_; 
wire _abc_40319_new_n1343_; 
wire _abc_40319_new_n1344_; 
wire _abc_40319_new_n1345_; 
wire _abc_40319_new_n1346_; 
wire _abc_40319_new_n1347_; 
wire _abc_40319_new_n1348_; 
wire _abc_40319_new_n1349_; 
wire _abc_40319_new_n1350_; 
wire _abc_40319_new_n1351_; 
wire _abc_40319_new_n1352_; 
wire _abc_40319_new_n1353_; 
wire _abc_40319_new_n1354_; 
wire _abc_40319_new_n1355_; 
wire _abc_40319_new_n1356_; 
wire _abc_40319_new_n1357_; 
wire _abc_40319_new_n1358_; 
wire _abc_40319_new_n1359_; 
wire _abc_40319_new_n1360_; 
wire _abc_40319_new_n1361_; 
wire _abc_40319_new_n1362_; 
wire _abc_40319_new_n1363_; 
wire _abc_40319_new_n1364_; 
wire _abc_40319_new_n1365_; 
wire _abc_40319_new_n1366_; 
wire _abc_40319_new_n1367_; 
wire _abc_40319_new_n1368_; 
wire _abc_40319_new_n1369_; 
wire _abc_40319_new_n1370_; 
wire _abc_40319_new_n1371_; 
wire _abc_40319_new_n1372_; 
wire _abc_40319_new_n1373_; 
wire _abc_40319_new_n1374_; 
wire _abc_40319_new_n1375_; 
wire _abc_40319_new_n1376_; 
wire _abc_40319_new_n1377_; 
wire _abc_40319_new_n1378_; 
wire _abc_40319_new_n1379_; 
wire _abc_40319_new_n1380_; 
wire _abc_40319_new_n1381_; 
wire _abc_40319_new_n1382_; 
wire _abc_40319_new_n1383_; 
wire _abc_40319_new_n1384_; 
wire _abc_40319_new_n1385_; 
wire _abc_40319_new_n1386_; 
wire _abc_40319_new_n1387_; 
wire _abc_40319_new_n1388_; 
wire _abc_40319_new_n1389_; 
wire _abc_40319_new_n1390_; 
wire _abc_40319_new_n1391_; 
wire _abc_40319_new_n1392_; 
wire _abc_40319_new_n1393_; 
wire _abc_40319_new_n1394_; 
wire _abc_40319_new_n1395_; 
wire _abc_40319_new_n1396_; 
wire _abc_40319_new_n1397_; 
wire _abc_40319_new_n1398_; 
wire _abc_40319_new_n1399_; 
wire _abc_40319_new_n1400_; 
wire _abc_40319_new_n1401_; 
wire _abc_40319_new_n1402_; 
wire _abc_40319_new_n1403_; 
wire _abc_40319_new_n1404_; 
wire _abc_40319_new_n1405_; 
wire _abc_40319_new_n1406_; 
wire _abc_40319_new_n1407_; 
wire _abc_40319_new_n1408_; 
wire _abc_40319_new_n1409_; 
wire _abc_40319_new_n1410_; 
wire _abc_40319_new_n1411_; 
wire _abc_40319_new_n1412_; 
wire _abc_40319_new_n1413_; 
wire _abc_40319_new_n1414_; 
wire _abc_40319_new_n1415_; 
wire _abc_40319_new_n1416_; 
wire _abc_40319_new_n1417_; 
wire _abc_40319_new_n1418_; 
wire _abc_40319_new_n1419_; 
wire _abc_40319_new_n1420_; 
wire _abc_40319_new_n1421_; 
wire _abc_40319_new_n1422_; 
wire _abc_40319_new_n1423_; 
wire _abc_40319_new_n1424_; 
wire _abc_40319_new_n1425_; 
wire _abc_40319_new_n1426_; 
wire _abc_40319_new_n1427_; 
wire _abc_40319_new_n1428_; 
wire _abc_40319_new_n1429_; 
wire _abc_40319_new_n1430_; 
wire _abc_40319_new_n1431_; 
wire _abc_40319_new_n1432_; 
wire _abc_40319_new_n1433_; 
wire _abc_40319_new_n1434_; 
wire _abc_40319_new_n1435_; 
wire _abc_40319_new_n1436_; 
wire _abc_40319_new_n1437_; 
wire _abc_40319_new_n1438_; 
wire _abc_40319_new_n1439_; 
wire _abc_40319_new_n1440_; 
wire _abc_40319_new_n1441_; 
wire _abc_40319_new_n1442_; 
wire _abc_40319_new_n1443_; 
wire _abc_40319_new_n1444_; 
wire _abc_40319_new_n1445_; 
wire _abc_40319_new_n1446_; 
wire _abc_40319_new_n1447_; 
wire _abc_40319_new_n1448_; 
wire _abc_40319_new_n1449_; 
wire _abc_40319_new_n1450_; 
wire _abc_40319_new_n1451_; 
wire _abc_40319_new_n1452_; 
wire _abc_40319_new_n1453_; 
wire _abc_40319_new_n1454_; 
wire _abc_40319_new_n1455_; 
wire _abc_40319_new_n1456_; 
wire _abc_40319_new_n1457_; 
wire _abc_40319_new_n1458_; 
wire _abc_40319_new_n1459_; 
wire _abc_40319_new_n1460_; 
wire _abc_40319_new_n1461_; 
wire _abc_40319_new_n1462_; 
wire _abc_40319_new_n1463_; 
wire _abc_40319_new_n1464_; 
wire _abc_40319_new_n1465_; 
wire _abc_40319_new_n1466_; 
wire _abc_40319_new_n1467_; 
wire _abc_40319_new_n1468_; 
wire _abc_40319_new_n1469_; 
wire _abc_40319_new_n1470_; 
wire _abc_40319_new_n1471_; 
wire _abc_40319_new_n1472_; 
wire _abc_40319_new_n1473_; 
wire _abc_40319_new_n1474_; 
wire _abc_40319_new_n1475_; 
wire _abc_40319_new_n1476_; 
wire _abc_40319_new_n1477_; 
wire _abc_40319_new_n1478_; 
wire _abc_40319_new_n1479_; 
wire _abc_40319_new_n1480_; 
wire _abc_40319_new_n1481_; 
wire _abc_40319_new_n1482_; 
wire _abc_40319_new_n1483_; 
wire _abc_40319_new_n1484_; 
wire _abc_40319_new_n1485_; 
wire _abc_40319_new_n1486_; 
wire _abc_40319_new_n1487_; 
wire _abc_40319_new_n1488_; 
wire _abc_40319_new_n1489_; 
wire _abc_40319_new_n1490_; 
wire _abc_40319_new_n1491_; 
wire _abc_40319_new_n1492_; 
wire _abc_40319_new_n1493_; 
wire _abc_40319_new_n1494_; 
wire _abc_40319_new_n1495_; 
wire _abc_40319_new_n1496_; 
wire _abc_40319_new_n1497_; 
wire _abc_40319_new_n1498_; 
wire _abc_40319_new_n1499_; 
wire _abc_40319_new_n1500_; 
wire _abc_40319_new_n1501_; 
wire _abc_40319_new_n1502_; 
wire _abc_40319_new_n1503_; 
wire _abc_40319_new_n1504_; 
wire _abc_40319_new_n1505_; 
wire _abc_40319_new_n1506_; 
wire _abc_40319_new_n1507_; 
wire _abc_40319_new_n1508_; 
wire _abc_40319_new_n1509_; 
wire _abc_40319_new_n1510_; 
wire _abc_40319_new_n1511_; 
wire _abc_40319_new_n1512_; 
wire _abc_40319_new_n1513_; 
wire _abc_40319_new_n1514_; 
wire _abc_40319_new_n1515_; 
wire _abc_40319_new_n1516_; 
wire _abc_40319_new_n1517_; 
wire _abc_40319_new_n1518_; 
wire _abc_40319_new_n1519_; 
wire _abc_40319_new_n1520_; 
wire _abc_40319_new_n1521_; 
wire _abc_40319_new_n1522_; 
wire _abc_40319_new_n1523_; 
wire _abc_40319_new_n1524_; 
wire _abc_40319_new_n1525_; 
wire _abc_40319_new_n1526_; 
wire _abc_40319_new_n1527_; 
wire _abc_40319_new_n1528_; 
wire _abc_40319_new_n1529_; 
wire _abc_40319_new_n1530_; 
wire _abc_40319_new_n1531_; 
wire _abc_40319_new_n1532_; 
wire _abc_40319_new_n1533_; 
wire _abc_40319_new_n1534_; 
wire _abc_40319_new_n1535_; 
wire _abc_40319_new_n1536_; 
wire _abc_40319_new_n1537_; 
wire _abc_40319_new_n1538_; 
wire _abc_40319_new_n1539_; 
wire _abc_40319_new_n1540_; 
wire _abc_40319_new_n1541_; 
wire _abc_40319_new_n1542_; 
wire _abc_40319_new_n1543_; 
wire _abc_40319_new_n1544_; 
wire _abc_40319_new_n1545_; 
wire _abc_40319_new_n1546_; 
wire _abc_40319_new_n1547_; 
wire _abc_40319_new_n1548_; 
wire _abc_40319_new_n1549_; 
wire _abc_40319_new_n1550_; 
wire _abc_40319_new_n1551_; 
wire _abc_40319_new_n1552_; 
wire _abc_40319_new_n1553_; 
wire _abc_40319_new_n1554_; 
wire _abc_40319_new_n1555_; 
wire _abc_40319_new_n1556_; 
wire _abc_40319_new_n1557_; 
wire _abc_40319_new_n1558_; 
wire _abc_40319_new_n1559_; 
wire _abc_40319_new_n1560_; 
wire _abc_40319_new_n1561_; 
wire _abc_40319_new_n1562_; 
wire _abc_40319_new_n1563_; 
wire _abc_40319_new_n1564_; 
wire _abc_40319_new_n1565_; 
wire _abc_40319_new_n1566_; 
wire _abc_40319_new_n1567_; 
wire _abc_40319_new_n1568_; 
wire _abc_40319_new_n1569_; 
wire _abc_40319_new_n1570_; 
wire _abc_40319_new_n1571_; 
wire _abc_40319_new_n1572_; 
wire _abc_40319_new_n1573_; 
wire _abc_40319_new_n1574_; 
wire _abc_40319_new_n1575_; 
wire _abc_40319_new_n1576_; 
wire _abc_40319_new_n1577_; 
wire _abc_40319_new_n1578_; 
wire _abc_40319_new_n1579_; 
wire _abc_40319_new_n1580_; 
wire _abc_40319_new_n1581_; 
wire _abc_40319_new_n1582_; 
wire _abc_40319_new_n1583_; 
wire _abc_40319_new_n1584_; 
wire _abc_40319_new_n1585_; 
wire _abc_40319_new_n1586_; 
wire _abc_40319_new_n1587_; 
wire _abc_40319_new_n1588_; 
wire _abc_40319_new_n1589_; 
wire _abc_40319_new_n1590_; 
wire _abc_40319_new_n1591_; 
wire _abc_40319_new_n1592_; 
wire _abc_40319_new_n1593_; 
wire _abc_40319_new_n1594_; 
wire _abc_40319_new_n1595_; 
wire _abc_40319_new_n1596_; 
wire _abc_40319_new_n1597_; 
wire _abc_40319_new_n1598_; 
wire _abc_40319_new_n1599_; 
wire _abc_40319_new_n1600_; 
wire _abc_40319_new_n1601_; 
wire _abc_40319_new_n1602_; 
wire _abc_40319_new_n1603_; 
wire _abc_40319_new_n1604_; 
wire _abc_40319_new_n1605_; 
wire _abc_40319_new_n1606_; 
wire _abc_40319_new_n1607_; 
wire _abc_40319_new_n1608_; 
wire _abc_40319_new_n1609_; 
wire _abc_40319_new_n1610_; 
wire _abc_40319_new_n1611_; 
wire _abc_40319_new_n1612_; 
wire _abc_40319_new_n1613_; 
wire _abc_40319_new_n1614_; 
wire _abc_40319_new_n1615_; 
wire _abc_40319_new_n1616_; 
wire _abc_40319_new_n1617_; 
wire _abc_40319_new_n1618_; 
wire _abc_40319_new_n1619_; 
wire _abc_40319_new_n1620_; 
wire _abc_40319_new_n1621_; 
wire _abc_40319_new_n1622_; 
wire _abc_40319_new_n1623_; 
wire _abc_40319_new_n1624_; 
wire _abc_40319_new_n1625_; 
wire _abc_40319_new_n1626_; 
wire _abc_40319_new_n1627_; 
wire _abc_40319_new_n1628_; 
wire _abc_40319_new_n1629_; 
wire _abc_40319_new_n1630_; 
wire _abc_40319_new_n1631_; 
wire _abc_40319_new_n1632_; 
wire _abc_40319_new_n1633_; 
wire _abc_40319_new_n1634_; 
wire _abc_40319_new_n1635_; 
wire _abc_40319_new_n1636_; 
wire _abc_40319_new_n1637_; 
wire _abc_40319_new_n1638_; 
wire _abc_40319_new_n1639_; 
wire _abc_40319_new_n1640_; 
wire _abc_40319_new_n1641_; 
wire _abc_40319_new_n1642_; 
wire _abc_40319_new_n1643_; 
wire _abc_40319_new_n1644_; 
wire _abc_40319_new_n1645_; 
wire _abc_40319_new_n1646_; 
wire _abc_40319_new_n1647_; 
wire _abc_40319_new_n1648_; 
wire _abc_40319_new_n1649_; 
wire _abc_40319_new_n1650_; 
wire _abc_40319_new_n1651_; 
wire _abc_40319_new_n1652_; 
wire _abc_40319_new_n1653_; 
wire _abc_40319_new_n1654_; 
wire _abc_40319_new_n1655_; 
wire _abc_40319_new_n1656_; 
wire _abc_40319_new_n1657_; 
wire _abc_40319_new_n1658_; 
wire _abc_40319_new_n1659_; 
wire _abc_40319_new_n1660_; 
wire _abc_40319_new_n1661_; 
wire _abc_40319_new_n1662_; 
wire _abc_40319_new_n1663_; 
wire _abc_40319_new_n1664_; 
wire _abc_40319_new_n1665_; 
wire _abc_40319_new_n1666_; 
wire _abc_40319_new_n1667_; 
wire _abc_40319_new_n1668_; 
wire _abc_40319_new_n1669_; 
wire _abc_40319_new_n1670_; 
wire _abc_40319_new_n1671_; 
wire _abc_40319_new_n1672_; 
wire _abc_40319_new_n1673_; 
wire _abc_40319_new_n1674_; 
wire _abc_40319_new_n1675_; 
wire _abc_40319_new_n1676_; 
wire _abc_40319_new_n1677_; 
wire _abc_40319_new_n1678_; 
wire _abc_40319_new_n1679_; 
wire _abc_40319_new_n1680_; 
wire _abc_40319_new_n1681_; 
wire _abc_40319_new_n1682_; 
wire _abc_40319_new_n1683_; 
wire _abc_40319_new_n1684_; 
wire _abc_40319_new_n1685_; 
wire _abc_40319_new_n1686_; 
wire _abc_40319_new_n1687_; 
wire _abc_40319_new_n1688_; 
wire _abc_40319_new_n1689_; 
wire _abc_40319_new_n1690_; 
wire _abc_40319_new_n1691_; 
wire _abc_40319_new_n1692_; 
wire _abc_40319_new_n1693_; 
wire _abc_40319_new_n1694_; 
wire _abc_40319_new_n1695_; 
wire _abc_40319_new_n1696_; 
wire _abc_40319_new_n1697_; 
wire _abc_40319_new_n1698_; 
wire _abc_40319_new_n1699_; 
wire _abc_40319_new_n1700_; 
wire _abc_40319_new_n1701_; 
wire _abc_40319_new_n1702_; 
wire _abc_40319_new_n1703_; 
wire _abc_40319_new_n1704_; 
wire _abc_40319_new_n1705_; 
wire _abc_40319_new_n1706_; 
wire _abc_40319_new_n1707_; 
wire _abc_40319_new_n1708_; 
wire _abc_40319_new_n1709_; 
wire _abc_40319_new_n1710_; 
wire _abc_40319_new_n1711_; 
wire _abc_40319_new_n1712_; 
wire _abc_40319_new_n1713_; 
wire _abc_40319_new_n1714_; 
wire _abc_40319_new_n1715_; 
wire _abc_40319_new_n1716_; 
wire _abc_40319_new_n1717_; 
wire _abc_40319_new_n1718_; 
wire _abc_40319_new_n1719_; 
wire _abc_40319_new_n1720_; 
wire _abc_40319_new_n1721_; 
wire _abc_40319_new_n1722_; 
wire _abc_40319_new_n1723_; 
wire _abc_40319_new_n1724_; 
wire _abc_40319_new_n1725_; 
wire _abc_40319_new_n1726_; 
wire _abc_40319_new_n1727_; 
wire _abc_40319_new_n1728_; 
wire _abc_40319_new_n1729_; 
wire _abc_40319_new_n1730_; 
wire _abc_40319_new_n1731_; 
wire _abc_40319_new_n1732_; 
wire _abc_40319_new_n1733_; 
wire _abc_40319_new_n1734_; 
wire _abc_40319_new_n1735_; 
wire _abc_40319_new_n1736_; 
wire _abc_40319_new_n1737_; 
wire _abc_40319_new_n1738_; 
wire _abc_40319_new_n1739_; 
wire _abc_40319_new_n1740_; 
wire _abc_40319_new_n1741_; 
wire _abc_40319_new_n1742_; 
wire _abc_40319_new_n1743_; 
wire _abc_40319_new_n1744_; 
wire _abc_40319_new_n1745_; 
wire _abc_40319_new_n1746_; 
wire _abc_40319_new_n1747_; 
wire _abc_40319_new_n1748_; 
wire _abc_40319_new_n1749_; 
wire _abc_40319_new_n1750_; 
wire _abc_40319_new_n1751_; 
wire _abc_40319_new_n1752_; 
wire _abc_40319_new_n1753_; 
wire _abc_40319_new_n1754_; 
wire _abc_40319_new_n1755_; 
wire _abc_40319_new_n1756_; 
wire _abc_40319_new_n1757_; 
wire _abc_40319_new_n1758_; 
wire _abc_40319_new_n1759_; 
wire _abc_40319_new_n1760_; 
wire _abc_40319_new_n1761_; 
wire _abc_40319_new_n1762_; 
wire _abc_40319_new_n1763_; 
wire _abc_40319_new_n1764_; 
wire _abc_40319_new_n1765_; 
wire _abc_40319_new_n1766_; 
wire _abc_40319_new_n1767_; 
wire _abc_40319_new_n1768_; 
wire _abc_40319_new_n1769_; 
wire _abc_40319_new_n1770_; 
wire _abc_40319_new_n1771_; 
wire _abc_40319_new_n1772_; 
wire _abc_40319_new_n1773_; 
wire _abc_40319_new_n1774_; 
wire _abc_40319_new_n1775_; 
wire _abc_40319_new_n1776_; 
wire _abc_40319_new_n1777_; 
wire _abc_40319_new_n1778_; 
wire _abc_40319_new_n1779_; 
wire _abc_40319_new_n1780_; 
wire _abc_40319_new_n1781_; 
wire _abc_40319_new_n1782_; 
wire _abc_40319_new_n1783_; 
wire _abc_40319_new_n1784_; 
wire _abc_40319_new_n1785_; 
wire _abc_40319_new_n1786_; 
wire _abc_40319_new_n1787_; 
wire _abc_40319_new_n1788_; 
wire _abc_40319_new_n1789_; 
wire _abc_40319_new_n1790_; 
wire _abc_40319_new_n1791_; 
wire _abc_40319_new_n1792_; 
wire _abc_40319_new_n1793_; 
wire _abc_40319_new_n1794_; 
wire _abc_40319_new_n1795_; 
wire _abc_40319_new_n1796_; 
wire _abc_40319_new_n1797_; 
wire _abc_40319_new_n1798_; 
wire _abc_40319_new_n1799_; 
wire _abc_40319_new_n1800_; 
wire _abc_40319_new_n1801_; 
wire _abc_40319_new_n1802_; 
wire _abc_40319_new_n1803_; 
wire _abc_40319_new_n1804_; 
wire _abc_40319_new_n1805_; 
wire _abc_40319_new_n1806_; 
wire _abc_40319_new_n1807_; 
wire _abc_40319_new_n1808_; 
wire _abc_40319_new_n1809_; 
wire _abc_40319_new_n1810_; 
wire _abc_40319_new_n1811_; 
wire _abc_40319_new_n1812_; 
wire _abc_40319_new_n1813_; 
wire _abc_40319_new_n1814_; 
wire _abc_40319_new_n1815_; 
wire _abc_40319_new_n1816_; 
wire _abc_40319_new_n1817_; 
wire _abc_40319_new_n1818_; 
wire _abc_40319_new_n1819_; 
wire _abc_40319_new_n1820_; 
wire _abc_40319_new_n1821_; 
wire _abc_40319_new_n1822_; 
wire _abc_40319_new_n1823_; 
wire _abc_40319_new_n1824_; 
wire _abc_40319_new_n1825_; 
wire _abc_40319_new_n1826_; 
wire _abc_40319_new_n1827_; 
wire _abc_40319_new_n1828_; 
wire _abc_40319_new_n1829_; 
wire _abc_40319_new_n1830_; 
wire _abc_40319_new_n1831_; 
wire _abc_40319_new_n1832_; 
wire _abc_40319_new_n1833_; 
wire _abc_40319_new_n1834_; 
wire _abc_40319_new_n1835_; 
wire _abc_40319_new_n1836_; 
wire _abc_40319_new_n1837_; 
wire _abc_40319_new_n1838_; 
wire _abc_40319_new_n1839_; 
wire _abc_40319_new_n1840_; 
wire _abc_40319_new_n1841_; 
wire _abc_40319_new_n1842_; 
wire _abc_40319_new_n1843_; 
wire _abc_40319_new_n1844_; 
wire _abc_40319_new_n1845_; 
wire _abc_40319_new_n1846_; 
wire _abc_40319_new_n1847_; 
wire _abc_40319_new_n1848_; 
wire _abc_40319_new_n1849_; 
wire _abc_40319_new_n1850_; 
wire _abc_40319_new_n1851_; 
wire _abc_40319_new_n1852_; 
wire _abc_40319_new_n1853_; 
wire _abc_40319_new_n1854_; 
wire _abc_40319_new_n1855_; 
wire _abc_40319_new_n1856_; 
wire _abc_40319_new_n1857_; 
wire _abc_40319_new_n1858_; 
wire _abc_40319_new_n1859_; 
wire _abc_40319_new_n1860_; 
wire _abc_40319_new_n1861_; 
wire _abc_40319_new_n1862_; 
wire _abc_40319_new_n1863_; 
wire _abc_40319_new_n1864_; 
wire _abc_40319_new_n1865_; 
wire _abc_40319_new_n1866_; 
wire _abc_40319_new_n1867_; 
wire _abc_40319_new_n1868_; 
wire _abc_40319_new_n1869_; 
wire _abc_40319_new_n1870_; 
wire _abc_40319_new_n1871_; 
wire _abc_40319_new_n1872_; 
wire _abc_40319_new_n1873_; 
wire _abc_40319_new_n1874_; 
wire _abc_40319_new_n1875_; 
wire _abc_40319_new_n1876_; 
wire _abc_40319_new_n1877_; 
wire _abc_40319_new_n1878_; 
wire _abc_40319_new_n1879_; 
wire _abc_40319_new_n1880_; 
wire _abc_40319_new_n1881_; 
wire _abc_40319_new_n1882_; 
wire _abc_40319_new_n1883_; 
wire _abc_40319_new_n1884_; 
wire _abc_40319_new_n1885_; 
wire _abc_40319_new_n1886_; 
wire _abc_40319_new_n1887_; 
wire _abc_40319_new_n1888_; 
wire _abc_40319_new_n1889_; 
wire _abc_40319_new_n1890_; 
wire _abc_40319_new_n1891_; 
wire _abc_40319_new_n1892_; 
wire _abc_40319_new_n1893_; 
wire _abc_40319_new_n1894_; 
wire _abc_40319_new_n1895_; 
wire _abc_40319_new_n1896_; 
wire _abc_40319_new_n1897_; 
wire _abc_40319_new_n1898_; 
wire _abc_40319_new_n1899_; 
wire _abc_40319_new_n1900_; 
wire _abc_40319_new_n1901_; 
wire _abc_40319_new_n1902_; 
wire _abc_40319_new_n1903_; 
wire _abc_40319_new_n1904_; 
wire _abc_40319_new_n1905_; 
wire _abc_40319_new_n1906_; 
wire _abc_40319_new_n1907_; 
wire _abc_40319_new_n1908_; 
wire _abc_40319_new_n1909_; 
wire _abc_40319_new_n1910_; 
wire _abc_40319_new_n1911_; 
wire _abc_40319_new_n1912_; 
wire _abc_40319_new_n1913_; 
wire _abc_40319_new_n1914_; 
wire _abc_40319_new_n1915_; 
wire _abc_40319_new_n1916_; 
wire _abc_40319_new_n1917_; 
wire _abc_40319_new_n1918_; 
wire _abc_40319_new_n1919_; 
wire _abc_40319_new_n1920_; 
wire _abc_40319_new_n1921_; 
wire _abc_40319_new_n1922_; 
wire _abc_40319_new_n1923_; 
wire _abc_40319_new_n1924_; 
wire _abc_40319_new_n1925_; 
wire _abc_40319_new_n1926_; 
wire _abc_40319_new_n1927_; 
wire _abc_40319_new_n1928_; 
wire _abc_40319_new_n1929_; 
wire _abc_40319_new_n1930_; 
wire _abc_40319_new_n1931_; 
wire _abc_40319_new_n1932_; 
wire _abc_40319_new_n1933_; 
wire _abc_40319_new_n1934_; 
wire _abc_40319_new_n1935_; 
wire _abc_40319_new_n1936_; 
wire _abc_40319_new_n1937_; 
wire _abc_40319_new_n1938_; 
wire _abc_40319_new_n1939_; 
wire _abc_40319_new_n1940_; 
wire _abc_40319_new_n1941_; 
wire _abc_40319_new_n1942_; 
wire _abc_40319_new_n1943_; 
wire _abc_40319_new_n1944_; 
wire _abc_40319_new_n1945_; 
wire _abc_40319_new_n1946_; 
wire _abc_40319_new_n1947_; 
wire _abc_40319_new_n1948_; 
wire _abc_40319_new_n1949_; 
wire _abc_40319_new_n1950_; 
wire _abc_40319_new_n1951_; 
wire _abc_40319_new_n1952_; 
wire _abc_40319_new_n1953_; 
wire _abc_40319_new_n1954_; 
wire _abc_40319_new_n1955_; 
wire _abc_40319_new_n1956_; 
wire _abc_40319_new_n1957_; 
wire _abc_40319_new_n1958_; 
wire _abc_40319_new_n1959_; 
wire _abc_40319_new_n1960_; 
wire _abc_40319_new_n1961_; 
wire _abc_40319_new_n1962_; 
wire _abc_40319_new_n1963_; 
wire _abc_40319_new_n1964_; 
wire _abc_40319_new_n1965_; 
wire _abc_40319_new_n1966_; 
wire _abc_40319_new_n1967_; 
wire _abc_40319_new_n1968_; 
wire _abc_40319_new_n1969_; 
wire _abc_40319_new_n1970_; 
wire _abc_40319_new_n1971_; 
wire _abc_40319_new_n1972_; 
wire _abc_40319_new_n1973_; 
wire _abc_40319_new_n1974_; 
wire _abc_40319_new_n1975_; 
wire _abc_40319_new_n1976_; 
wire _abc_40319_new_n1977_; 
wire _abc_40319_new_n1978_; 
wire _abc_40319_new_n1979_; 
wire _abc_40319_new_n1980_; 
wire _abc_40319_new_n1981_; 
wire _abc_40319_new_n1982_; 
wire _abc_40319_new_n1983_; 
wire _abc_40319_new_n1984_; 
wire _abc_40319_new_n1985_; 
wire _abc_40319_new_n1986_; 
wire _abc_40319_new_n1987_; 
wire _abc_40319_new_n1988_; 
wire _abc_40319_new_n1989_; 
wire _abc_40319_new_n1990_; 
wire _abc_40319_new_n1992_; 
wire _abc_40319_new_n1993_; 
wire _abc_40319_new_n1994_; 
wire _abc_40319_new_n1995_; 
wire _abc_40319_new_n1996_; 
wire _abc_40319_new_n1997_; 
wire _abc_40319_new_n1998_; 
wire _abc_40319_new_n1999_; 
wire _abc_40319_new_n2000_; 
wire _abc_40319_new_n2001_; 
wire _abc_40319_new_n2002_; 
wire _abc_40319_new_n2003_; 
wire _abc_40319_new_n2004_; 
wire _abc_40319_new_n2005_; 
wire _abc_40319_new_n2006_; 
wire _abc_40319_new_n2007_; 
wire _abc_40319_new_n2008_; 
wire _abc_40319_new_n2010_; 
wire _abc_40319_new_n2011_; 
wire _abc_40319_new_n2012_; 
wire _abc_40319_new_n2013_; 
wire _abc_40319_new_n2014_; 
wire _abc_40319_new_n2015_; 
wire _abc_40319_new_n2016_; 
wire _abc_40319_new_n2017_; 
wire _abc_40319_new_n2018_; 
wire _abc_40319_new_n2019_; 
wire _abc_40319_new_n2020_; 
wire _abc_40319_new_n2021_; 
wire _abc_40319_new_n2022_; 
wire _abc_40319_new_n2023_; 
wire _abc_40319_new_n2024_; 
wire _abc_40319_new_n2025_; 
wire _abc_40319_new_n2026_; 
wire _abc_40319_new_n2028_; 
wire _abc_40319_new_n2029_; 
wire _abc_40319_new_n2030_; 
wire _abc_40319_new_n2031_; 
wire _abc_40319_new_n2032_; 
wire _abc_40319_new_n2033_; 
wire _abc_40319_new_n2034_; 
wire _abc_40319_new_n2035_; 
wire _abc_40319_new_n2036_; 
wire _abc_40319_new_n2037_; 
wire _abc_40319_new_n2038_; 
wire _abc_40319_new_n2039_; 
wire _abc_40319_new_n2040_; 
wire _abc_40319_new_n2041_; 
wire _abc_40319_new_n2042_; 
wire _abc_40319_new_n2043_; 
wire _abc_40319_new_n2044_; 
wire _abc_40319_new_n2045_; 
wire _abc_40319_new_n2047_; 
wire _abc_40319_new_n2048_; 
wire _abc_40319_new_n2049_; 
wire _abc_40319_new_n2050_; 
wire _abc_40319_new_n2051_; 
wire _abc_40319_new_n2052_; 
wire _abc_40319_new_n2053_; 
wire _abc_40319_new_n2054_; 
wire _abc_40319_new_n2055_; 
wire _abc_40319_new_n2056_; 
wire _abc_40319_new_n2057_; 
wire _abc_40319_new_n2058_; 
wire _abc_40319_new_n2059_; 
wire _abc_40319_new_n2060_; 
wire _abc_40319_new_n2061_; 
wire _abc_40319_new_n2062_; 
wire _abc_40319_new_n2063_; 
wire _abc_40319_new_n2064_; 
wire _abc_40319_new_n2065_; 
wire _abc_40319_new_n2066_; 
wire _abc_40319_new_n2067_; 
wire _abc_40319_new_n2068_; 
wire _abc_40319_new_n2070_; 
wire _abc_40319_new_n2071_; 
wire _abc_40319_new_n2072_; 
wire _abc_40319_new_n2073_; 
wire _abc_40319_new_n2074_; 
wire _abc_40319_new_n2075_; 
wire _abc_40319_new_n2076_; 
wire _abc_40319_new_n2077_; 
wire _abc_40319_new_n2078_; 
wire _abc_40319_new_n2079_; 
wire _abc_40319_new_n2080_; 
wire _abc_40319_new_n2081_; 
wire _abc_40319_new_n2082_; 
wire _abc_40319_new_n2083_; 
wire _abc_40319_new_n2084_; 
wire _abc_40319_new_n2085_; 
wire _abc_40319_new_n2086_; 
wire _abc_40319_new_n2088_; 
wire _abc_40319_new_n2089_; 
wire _abc_40319_new_n2090_; 
wire _abc_40319_new_n2091_; 
wire _abc_40319_new_n2092_; 
wire _abc_40319_new_n2093_; 
wire _abc_40319_new_n2094_; 
wire _abc_40319_new_n2095_; 
wire _abc_40319_new_n2096_; 
wire _abc_40319_new_n2097_; 
wire _abc_40319_new_n2098_; 
wire _abc_40319_new_n2099_; 
wire _abc_40319_new_n2100_; 
wire _abc_40319_new_n2101_; 
wire _abc_40319_new_n2102_; 
wire _abc_40319_new_n2103_; 
wire _abc_40319_new_n2104_; 
wire _abc_40319_new_n2105_; 
wire _abc_40319_new_n2106_; 
wire _abc_40319_new_n2107_; 
wire _abc_40319_new_n2108_; 
wire _abc_40319_new_n2109_; 
wire _abc_40319_new_n2110_; 
wire _abc_40319_new_n2111_; 
wire _abc_40319_new_n2112_; 
wire _abc_40319_new_n2113_; 
wire _abc_40319_new_n2114_; 
wire _abc_40319_new_n2115_; 
wire _abc_40319_new_n2116_; 
wire _abc_40319_new_n2117_; 
wire _abc_40319_new_n2118_; 
wire _abc_40319_new_n2119_; 
wire _abc_40319_new_n2120_; 
wire _abc_40319_new_n2121_; 
wire _abc_40319_new_n2122_; 
wire _abc_40319_new_n2123_; 
wire _abc_40319_new_n2124_; 
wire _abc_40319_new_n2125_; 
wire _abc_40319_new_n2126_; 
wire _abc_40319_new_n2127_; 
wire _abc_40319_new_n2128_; 
wire _abc_40319_new_n2129_; 
wire _abc_40319_new_n2130_; 
wire _abc_40319_new_n2131_; 
wire _abc_40319_new_n2132_; 
wire _abc_40319_new_n2133_; 
wire _abc_40319_new_n2135_; 
wire _abc_40319_new_n2136_; 
wire _abc_40319_new_n2137_; 
wire _abc_40319_new_n2138_; 
wire _abc_40319_new_n2139_; 
wire _abc_40319_new_n2140_; 
wire _abc_40319_new_n2141_; 
wire _abc_40319_new_n2142_; 
wire _abc_40319_new_n2143_; 
wire _abc_40319_new_n2144_; 
wire _abc_40319_new_n2145_; 
wire _abc_40319_new_n2146_; 
wire _abc_40319_new_n2147_; 
wire _abc_40319_new_n2148_; 
wire _abc_40319_new_n2149_; 
wire _abc_40319_new_n2150_; 
wire _abc_40319_new_n2151_; 
wire _abc_40319_new_n2152_; 
wire _abc_40319_new_n2153_; 
wire _abc_40319_new_n2154_; 
wire _abc_40319_new_n2155_; 
wire _abc_40319_new_n2157_; 
wire _abc_40319_new_n2158_; 
wire _abc_40319_new_n2159_; 
wire _abc_40319_new_n2160_; 
wire _abc_40319_new_n2161_; 
wire _abc_40319_new_n2162_; 
wire _abc_40319_new_n2163_; 
wire _abc_40319_new_n2164_; 
wire _abc_40319_new_n2165_; 
wire _abc_40319_new_n2166_; 
wire _abc_40319_new_n2167_; 
wire _abc_40319_new_n2168_; 
wire _abc_40319_new_n2169_; 
wire _abc_40319_new_n2170_; 
wire _abc_40319_new_n2171_; 
wire _abc_40319_new_n2172_; 
wire _abc_40319_new_n2174_; 
wire _abc_40319_new_n2175_; 
wire _abc_40319_new_n2176_; 
wire _abc_40319_new_n2177_; 
wire _abc_40319_new_n2178_; 
wire _abc_40319_new_n2179_; 
wire _abc_40319_new_n2180_; 
wire _abc_40319_new_n2181_; 
wire _abc_40319_new_n2182_; 
wire _abc_40319_new_n2183_; 
wire _abc_40319_new_n2184_; 
wire _abc_40319_new_n2185_; 
wire _abc_40319_new_n2186_; 
wire _abc_40319_new_n2187_; 
wire _abc_40319_new_n2188_; 
wire _abc_40319_new_n2189_; 
wire _abc_40319_new_n2190_; 
wire _abc_40319_new_n2191_; 
wire _abc_40319_new_n2192_; 
wire _abc_40319_new_n2193_; 
wire _abc_40319_new_n2194_; 
wire _abc_40319_new_n2195_; 
wire _abc_40319_new_n2196_; 
wire _abc_40319_new_n2197_; 
wire _abc_40319_new_n2198_; 
wire _abc_40319_new_n2199_; 
wire _abc_40319_new_n2200_; 
wire _abc_40319_new_n2202_; 
wire _abc_40319_new_n2203_; 
wire _abc_40319_new_n2204_; 
wire _abc_40319_new_n2205_; 
wire _abc_40319_new_n2206_; 
wire _abc_40319_new_n2207_; 
wire _abc_40319_new_n2208_; 
wire _abc_40319_new_n2209_; 
wire _abc_40319_new_n2210_; 
wire _abc_40319_new_n2211_; 
wire _abc_40319_new_n2212_; 
wire _abc_40319_new_n2213_; 
wire _abc_40319_new_n2214_; 
wire _abc_40319_new_n2215_; 
wire _abc_40319_new_n2216_; 
wire _abc_40319_new_n2217_; 
wire _abc_40319_new_n2218_; 
wire _abc_40319_new_n2219_; 
wire _abc_40319_new_n2220_; 
wire _abc_40319_new_n2221_; 
wire _abc_40319_new_n2222_; 
wire _abc_40319_new_n2223_; 
wire _abc_40319_new_n2225_; 
wire _abc_40319_new_n2226_; 
wire _abc_40319_new_n2227_; 
wire _abc_40319_new_n2228_; 
wire _abc_40319_new_n2229_; 
wire _abc_40319_new_n2230_; 
wire _abc_40319_new_n2231_; 
wire _abc_40319_new_n2232_; 
wire _abc_40319_new_n2233_; 
wire _abc_40319_new_n2234_; 
wire _abc_40319_new_n2235_; 
wire _abc_40319_new_n2236_; 
wire _abc_40319_new_n2237_; 
wire _abc_40319_new_n2238_; 
wire _abc_40319_new_n2239_; 
wire _abc_40319_new_n2240_; 
wire _abc_40319_new_n2241_; 
wire _abc_40319_new_n2242_; 
wire _abc_40319_new_n2243_; 
wire _abc_40319_new_n2244_; 
wire _abc_40319_new_n2246_; 
wire _abc_40319_new_n2247_; 
wire _abc_40319_new_n2248_; 
wire _abc_40319_new_n2249_; 
wire _abc_40319_new_n2250_; 
wire _abc_40319_new_n2251_; 
wire _abc_40319_new_n2252_; 
wire _abc_40319_new_n2253_; 
wire _abc_40319_new_n2254_; 
wire _abc_40319_new_n2255_; 
wire _abc_40319_new_n2256_; 
wire _abc_40319_new_n2257_; 
wire _abc_40319_new_n2258_; 
wire _abc_40319_new_n2259_; 
wire _abc_40319_new_n2260_; 
wire _abc_40319_new_n2261_; 
wire _abc_40319_new_n2262_; 
wire _abc_40319_new_n2264_; 
wire _abc_40319_new_n2265_; 
wire _abc_40319_new_n2266_; 
wire _abc_40319_new_n2267_; 
wire _abc_40319_new_n2268_; 
wire _abc_40319_new_n2269_; 
wire _abc_40319_new_n2270_; 
wire _abc_40319_new_n2271_; 
wire _abc_40319_new_n2272_; 
wire _abc_40319_new_n2273_; 
wire _abc_40319_new_n2274_; 
wire _abc_40319_new_n2275_; 
wire _abc_40319_new_n2276_; 
wire _abc_40319_new_n2277_; 
wire _abc_40319_new_n2278_; 
wire _abc_40319_new_n2279_; 
wire _abc_40319_new_n2280_; 
wire _abc_40319_new_n2282_; 
wire _abc_40319_new_n2283_; 
wire _abc_40319_new_n2284_; 
wire _abc_40319_new_n2285_; 
wire _abc_40319_new_n2286_; 
wire _abc_40319_new_n2287_; 
wire _abc_40319_new_n2288_; 
wire _abc_40319_new_n2289_; 
wire _abc_40319_new_n2290_; 
wire _abc_40319_new_n2291_; 
wire _abc_40319_new_n2292_; 
wire _abc_40319_new_n2293_; 
wire _abc_40319_new_n2294_; 
wire _abc_40319_new_n2295_; 
wire _abc_40319_new_n2296_; 
wire _abc_40319_new_n2297_; 
wire _abc_40319_new_n2298_; 
wire _abc_40319_new_n2299_; 
wire _abc_40319_new_n2300_; 
wire _abc_40319_new_n2301_; 
wire _abc_40319_new_n2303_; 
wire _abc_40319_new_n2304_; 
wire _abc_40319_new_n2305_; 
wire _abc_40319_new_n2306_; 
wire _abc_40319_new_n2307_; 
wire _abc_40319_new_n2308_; 
wire _abc_40319_new_n2309_; 
wire _abc_40319_new_n2310_; 
wire _abc_40319_new_n2311_; 
wire _abc_40319_new_n2312_; 
wire _abc_40319_new_n2313_; 
wire _abc_40319_new_n2314_; 
wire _abc_40319_new_n2315_; 
wire _abc_40319_new_n2316_; 
wire _abc_40319_new_n2317_; 
wire _abc_40319_new_n2318_; 
wire _abc_40319_new_n2319_; 
wire _abc_40319_new_n2320_; 
wire _abc_40319_new_n2322_; 
wire _abc_40319_new_n2323_; 
wire _abc_40319_new_n2324_; 
wire _abc_40319_new_n2325_; 
wire _abc_40319_new_n2326_; 
wire _abc_40319_new_n2327_; 
wire _abc_40319_new_n2328_; 
wire _abc_40319_new_n2329_; 
wire _abc_40319_new_n2330_; 
wire _abc_40319_new_n2331_; 
wire _abc_40319_new_n2332_; 
wire _abc_40319_new_n2333_; 
wire _abc_40319_new_n2334_; 
wire _abc_40319_new_n2335_; 
wire _abc_40319_new_n2336_; 
wire _abc_40319_new_n2337_; 
wire _abc_40319_new_n2338_; 
wire _abc_40319_new_n2340_; 
wire _abc_40319_new_n2341_; 
wire _abc_40319_new_n2342_; 
wire _abc_40319_new_n2343_; 
wire _abc_40319_new_n2344_; 
wire _abc_40319_new_n2345_; 
wire _abc_40319_new_n2346_; 
wire _abc_40319_new_n2347_; 
wire _abc_40319_new_n2348_; 
wire _abc_40319_new_n2349_; 
wire _abc_40319_new_n2350_; 
wire _abc_40319_new_n2351_; 
wire _abc_40319_new_n2352_; 
wire _abc_40319_new_n2353_; 
wire _abc_40319_new_n2354_; 
wire _abc_40319_new_n2355_; 
wire _abc_40319_new_n2357_; 
wire _abc_40319_new_n2358_; 
wire _abc_40319_new_n2359_; 
wire _abc_40319_new_n2360_; 
wire _abc_40319_new_n2361_; 
wire _abc_40319_new_n2362_; 
wire _abc_40319_new_n2363_; 
wire _abc_40319_new_n2364_; 
wire _abc_40319_new_n2365_; 
wire _abc_40319_new_n2366_; 
wire _abc_40319_new_n2367_; 
wire _abc_40319_new_n2368_; 
wire _abc_40319_new_n2369_; 
wire _abc_40319_new_n2370_; 
wire _abc_40319_new_n2371_; 
wire _abc_40319_new_n2373_; 
wire _abc_40319_new_n2374_; 
wire _abc_40319_new_n2375_; 
wire _abc_40319_new_n2376_; 
wire _abc_40319_new_n2377_; 
wire _abc_40319_new_n2378_; 
wire _abc_40319_new_n2379_; 
wire _abc_40319_new_n2380_; 
wire _abc_40319_new_n2381_; 
wire _abc_40319_new_n2382_; 
wire _abc_40319_new_n2383_; 
wire _abc_40319_new_n2384_; 
wire _abc_40319_new_n2385_; 
wire _abc_40319_new_n2386_; 
wire _abc_40319_new_n2387_; 
wire _abc_40319_new_n2388_; 
wire _abc_40319_new_n2389_; 
wire _abc_40319_new_n2391_; 
wire _abc_40319_new_n2392_; 
wire _abc_40319_new_n2393_; 
wire _abc_40319_new_n2394_; 
wire _abc_40319_new_n2395_; 
wire _abc_40319_new_n2396_; 
wire _abc_40319_new_n2397_; 
wire _abc_40319_new_n2398_; 
wire _abc_40319_new_n2399_; 
wire _abc_40319_new_n2400_; 
wire _abc_40319_new_n2401_; 
wire _abc_40319_new_n2402_; 
wire _abc_40319_new_n2403_; 
wire _abc_40319_new_n2404_; 
wire _abc_40319_new_n2405_; 
wire _abc_40319_new_n2406_; 
wire _abc_40319_new_n2407_; 
wire _abc_40319_new_n2408_; 
wire _abc_40319_new_n2409_; 
wire _abc_40319_new_n2410_; 
wire _abc_40319_new_n2411_; 
wire _abc_40319_new_n2412_; 
wire _abc_40319_new_n2413_; 
wire _abc_40319_new_n2414_; 
wire _abc_40319_new_n2415_; 
wire _abc_40319_new_n2417_; 
wire _abc_40319_new_n2418_; 
wire _abc_40319_new_n2419_; 
wire _abc_40319_new_n2420_; 
wire _abc_40319_new_n2421_; 
wire _abc_40319_new_n2422_; 
wire _abc_40319_new_n2423_; 
wire _abc_40319_new_n2424_; 
wire _abc_40319_new_n2425_; 
wire _abc_40319_new_n2426_; 
wire _abc_40319_new_n2427_; 
wire _abc_40319_new_n2428_; 
wire _abc_40319_new_n2429_; 
wire _abc_40319_new_n2430_; 
wire _abc_40319_new_n2431_; 
wire _abc_40319_new_n2432_; 
wire _abc_40319_new_n2433_; 
wire _abc_40319_new_n2435_; 
wire _abc_40319_new_n2436_; 
wire _abc_40319_new_n2437_; 
wire _abc_40319_new_n2438_; 
wire _abc_40319_new_n2439_; 
wire _abc_40319_new_n2440_; 
wire _abc_40319_new_n2441_; 
wire _abc_40319_new_n2442_; 
wire _abc_40319_new_n2443_; 
wire _abc_40319_new_n2444_; 
wire _abc_40319_new_n2445_; 
wire _abc_40319_new_n2446_; 
wire _abc_40319_new_n2447_; 
wire _abc_40319_new_n2448_; 
wire _abc_40319_new_n2449_; 
wire _abc_40319_new_n2450_; 
wire _abc_40319_new_n2451_; 
wire _abc_40319_new_n2452_; 
wire _abc_40319_new_n2454_; 
wire _abc_40319_new_n2455_; 
wire _abc_40319_new_n2456_; 
wire _abc_40319_new_n2457_; 
wire _abc_40319_new_n2458_; 
wire _abc_40319_new_n2459_; 
wire _abc_40319_new_n2460_; 
wire _abc_40319_new_n2461_; 
wire _abc_40319_new_n2462_; 
wire _abc_40319_new_n2463_; 
wire _abc_40319_new_n2464_; 
wire _abc_40319_new_n2465_; 
wire _abc_40319_new_n2466_; 
wire _abc_40319_new_n2467_; 
wire _abc_40319_new_n2468_; 
wire _abc_40319_new_n2469_; 
wire _abc_40319_new_n2470_; 
wire _abc_40319_new_n2472_; 
wire _abc_40319_new_n2473_; 
wire _abc_40319_new_n2474_; 
wire _abc_40319_new_n2475_; 
wire _abc_40319_new_n2476_; 
wire _abc_40319_new_n2477_; 
wire _abc_40319_new_n2478_; 
wire _abc_40319_new_n2479_; 
wire _abc_40319_new_n2480_; 
wire _abc_40319_new_n2481_; 
wire _abc_40319_new_n2482_; 
wire _abc_40319_new_n2483_; 
wire _abc_40319_new_n2484_; 
wire _abc_40319_new_n2485_; 
wire _abc_40319_new_n2486_; 
wire _abc_40319_new_n2487_; 
wire _abc_40319_new_n2488_; 
wire _abc_40319_new_n2490_; 
wire _abc_40319_new_n2491_; 
wire _abc_40319_new_n2492_; 
wire _abc_40319_new_n2493_; 
wire _abc_40319_new_n2494_; 
wire _abc_40319_new_n2495_; 
wire _abc_40319_new_n2496_; 
wire _abc_40319_new_n2497_; 
wire _abc_40319_new_n2498_; 
wire _abc_40319_new_n2499_; 
wire _abc_40319_new_n2500_; 
wire _abc_40319_new_n2501_; 
wire _abc_40319_new_n2502_; 
wire _abc_40319_new_n2503_; 
wire _abc_40319_new_n2504_; 
wire _abc_40319_new_n2505_; 
wire _abc_40319_new_n2506_; 
wire _abc_40319_new_n2508_; 
wire _abc_40319_new_n2509_; 
wire _abc_40319_new_n2510_; 
wire _abc_40319_new_n2511_; 
wire _abc_40319_new_n2512_; 
wire _abc_40319_new_n2513_; 
wire _abc_40319_new_n2514_; 
wire _abc_40319_new_n2515_; 
wire _abc_40319_new_n2516_; 
wire _abc_40319_new_n2517_; 
wire _abc_40319_new_n2518_; 
wire _abc_40319_new_n2519_; 
wire _abc_40319_new_n2520_; 
wire _abc_40319_new_n2521_; 
wire _abc_40319_new_n2522_; 
wire _abc_40319_new_n2523_; 
wire _abc_40319_new_n2524_; 
wire _abc_40319_new_n2525_; 
wire _abc_40319_new_n2526_; 
wire _abc_40319_new_n2527_; 
wire _abc_40319_new_n2528_; 
wire _abc_40319_new_n2529_; 
wire _abc_40319_new_n2531_; 
wire _abc_40319_new_n2532_; 
wire _abc_40319_new_n2533_; 
wire _abc_40319_new_n2534_; 
wire _abc_40319_new_n2535_; 
wire _abc_40319_new_n2536_; 
wire _abc_40319_new_n2537_; 
wire _abc_40319_new_n2538_; 
wire _abc_40319_new_n2539_; 
wire _abc_40319_new_n2540_; 
wire _abc_40319_new_n2541_; 
wire _abc_40319_new_n2542_; 
wire _abc_40319_new_n2543_; 
wire _abc_40319_new_n2544_; 
wire _abc_40319_new_n2545_; 
wire _abc_40319_new_n2546_; 
wire _abc_40319_new_n2547_; 
wire _abc_40319_new_n2549_; 
wire _abc_40319_new_n2550_; 
wire _abc_40319_new_n2551_; 
wire _abc_40319_new_n2552_; 
wire _abc_40319_new_n2553_; 
wire _abc_40319_new_n2554_; 
wire _abc_40319_new_n2555_; 
wire _abc_40319_new_n2556_; 
wire _abc_40319_new_n2557_; 
wire _abc_40319_new_n2558_; 
wire _abc_40319_new_n2559_; 
wire _abc_40319_new_n2560_; 
wire _abc_40319_new_n2561_; 
wire _abc_40319_new_n2562_; 
wire _abc_40319_new_n2563_; 
wire _abc_40319_new_n2564_; 
wire _abc_40319_new_n2565_; 
wire _abc_40319_new_n2566_; 
wire _abc_40319_new_n2567_; 
wire _abc_40319_new_n2568_; 
wire _abc_40319_new_n2569_; 
wire _abc_40319_new_n2570_; 
wire _abc_40319_new_n2571_; 
wire _abc_40319_new_n2572_; 
wire _abc_40319_new_n2573_; 
wire _abc_40319_new_n2574_; 
wire _abc_40319_new_n2575_; 
wire _abc_40319_new_n2576_; 
wire _abc_40319_new_n2577_; 
wire _abc_40319_new_n2578_; 
wire _abc_40319_new_n2579_; 
wire _abc_40319_new_n2580_; 
wire _abc_40319_new_n2581_; 
wire _abc_40319_new_n2582_; 
wire _abc_40319_new_n2583_; 
wire _abc_40319_new_n2584_; 
wire _abc_40319_new_n2585_; 
wire _abc_40319_new_n2586_; 
wire _abc_40319_new_n2587_; 
wire _abc_40319_new_n2588_; 
wire _abc_40319_new_n2589_; 
wire _abc_40319_new_n2590_; 
wire _abc_40319_new_n2591_; 
wire _abc_40319_new_n2592_; 
wire _abc_40319_new_n2593_; 
wire _abc_40319_new_n2594_; 
wire _abc_40319_new_n2595_; 
wire _abc_40319_new_n2596_; 
wire _abc_40319_new_n2597_; 
wire _abc_40319_new_n2598_; 
wire _abc_40319_new_n2599_; 
wire _abc_40319_new_n2600_; 
wire _abc_40319_new_n2601_; 
wire _abc_40319_new_n2602_; 
wire _abc_40319_new_n2603_; 
wire _abc_40319_new_n2604_; 
wire _abc_40319_new_n2605_; 
wire _abc_40319_new_n2606_; 
wire _abc_40319_new_n2607_; 
wire _abc_40319_new_n2608_; 
wire _abc_40319_new_n2609_; 
wire _abc_40319_new_n2610_; 
wire _abc_40319_new_n2611_; 
wire _abc_40319_new_n2612_; 
wire _abc_40319_new_n2613_; 
wire _abc_40319_new_n2614_; 
wire _abc_40319_new_n2615_; 
wire _abc_40319_new_n2616_; 
wire _abc_40319_new_n2617_; 
wire _abc_40319_new_n2618_; 
wire _abc_40319_new_n2619_; 
wire _abc_40319_new_n2620_; 
wire _abc_40319_new_n2621_; 
wire _abc_40319_new_n2622_; 
wire _abc_40319_new_n2623_; 
wire _abc_40319_new_n2624_; 
wire _abc_40319_new_n2625_; 
wire _abc_40319_new_n2626_; 
wire _abc_40319_new_n2627_; 
wire _abc_40319_new_n2628_; 
wire _abc_40319_new_n2629_; 
wire _abc_40319_new_n2630_; 
wire _abc_40319_new_n2631_; 
wire _abc_40319_new_n2632_; 
wire _abc_40319_new_n2633_; 
wire _abc_40319_new_n2634_; 
wire _abc_40319_new_n2635_; 
wire _abc_40319_new_n2636_; 
wire _abc_40319_new_n2637_; 
wire _abc_40319_new_n2638_; 
wire _abc_40319_new_n2639_; 
wire _abc_40319_new_n2640_; 
wire _abc_40319_new_n2641_; 
wire _abc_40319_new_n2642_; 
wire _abc_40319_new_n2643_; 
wire _abc_40319_new_n2644_; 
wire _abc_40319_new_n2645_; 
wire _abc_40319_new_n2646_; 
wire _abc_40319_new_n2647_; 
wire _abc_40319_new_n2648_; 
wire _abc_40319_new_n2649_; 
wire _abc_40319_new_n2650_; 
wire _abc_40319_new_n2651_; 
wire _abc_40319_new_n2652_; 
wire _abc_40319_new_n2653_; 
wire _abc_40319_new_n2654_; 
wire _abc_40319_new_n2655_; 
wire _abc_40319_new_n2656_; 
wire _abc_40319_new_n2657_; 
wire _abc_40319_new_n2658_; 
wire _abc_40319_new_n2659_; 
wire _abc_40319_new_n2660_; 
wire _abc_40319_new_n2661_; 
wire _abc_40319_new_n2662_; 
wire _abc_40319_new_n2663_; 
wire _abc_40319_new_n2664_; 
wire _abc_40319_new_n2665_; 
wire _abc_40319_new_n2666_; 
wire _abc_40319_new_n2667_; 
wire _abc_40319_new_n2668_; 
wire _abc_40319_new_n2669_; 
wire _abc_40319_new_n2670_; 
wire _abc_40319_new_n2671_; 
wire _abc_40319_new_n2672_; 
wire _abc_40319_new_n2673_; 
wire _abc_40319_new_n2674_; 
wire _abc_40319_new_n2675_; 
wire _abc_40319_new_n2676_; 
wire _abc_40319_new_n2677_; 
wire _abc_40319_new_n2678_; 
wire _abc_40319_new_n2679_; 
wire _abc_40319_new_n2680_; 
wire _abc_40319_new_n2681_; 
wire _abc_40319_new_n2682_; 
wire _abc_40319_new_n2683_; 
wire _abc_40319_new_n2684_; 
wire _abc_40319_new_n2685_; 
wire _abc_40319_new_n2686_; 
wire _abc_40319_new_n2687_; 
wire _abc_40319_new_n2688_; 
wire _abc_40319_new_n2689_; 
wire _abc_40319_new_n2690_; 
wire _abc_40319_new_n2691_; 
wire _abc_40319_new_n2692_; 
wire _abc_40319_new_n2693_; 
wire _abc_40319_new_n2694_; 
wire _abc_40319_new_n2695_; 
wire _abc_40319_new_n2696_; 
wire _abc_40319_new_n2697_; 
wire _abc_40319_new_n2698_; 
wire _abc_40319_new_n2699_; 
wire _abc_40319_new_n2700_; 
wire _abc_40319_new_n2701_; 
wire _abc_40319_new_n2702_; 
wire _abc_40319_new_n2703_; 
wire _abc_40319_new_n2704_; 
wire _abc_40319_new_n2705_; 
wire _abc_40319_new_n2706_; 
wire _abc_40319_new_n2707_; 
wire _abc_40319_new_n2708_; 
wire _abc_40319_new_n2709_; 
wire _abc_40319_new_n2710_; 
wire _abc_40319_new_n2711_; 
wire _abc_40319_new_n2712_; 
wire _abc_40319_new_n2713_; 
wire _abc_40319_new_n2714_; 
wire _abc_40319_new_n2715_; 
wire _abc_40319_new_n2716_; 
wire _abc_40319_new_n2717_; 
wire _abc_40319_new_n2718_; 
wire _abc_40319_new_n2719_; 
wire _abc_40319_new_n2720_; 
wire _abc_40319_new_n2721_; 
wire _abc_40319_new_n2722_; 
wire _abc_40319_new_n2723_; 
wire _abc_40319_new_n2724_; 
wire _abc_40319_new_n2725_; 
wire _abc_40319_new_n2726_; 
wire _abc_40319_new_n2727_; 
wire _abc_40319_new_n2728_; 
wire _abc_40319_new_n2729_; 
wire _abc_40319_new_n2730_; 
wire _abc_40319_new_n2731_; 
wire _abc_40319_new_n2732_; 
wire _abc_40319_new_n2733_; 
wire _abc_40319_new_n2734_; 
wire _abc_40319_new_n2735_; 
wire _abc_40319_new_n2736_; 
wire _abc_40319_new_n2737_; 
wire _abc_40319_new_n2738_; 
wire _abc_40319_new_n2739_; 
wire _abc_40319_new_n2740_; 
wire _abc_40319_new_n2741_; 
wire _abc_40319_new_n2742_; 
wire _abc_40319_new_n2743_; 
wire _abc_40319_new_n2744_; 
wire _abc_40319_new_n2745_; 
wire _abc_40319_new_n2746_; 
wire _abc_40319_new_n2747_; 
wire _abc_40319_new_n2748_; 
wire _abc_40319_new_n2749_; 
wire _abc_40319_new_n2750_; 
wire _abc_40319_new_n2751_; 
wire _abc_40319_new_n2752_; 
wire _abc_40319_new_n2753_; 
wire _abc_40319_new_n2754_; 
wire _abc_40319_new_n2755_; 
wire _abc_40319_new_n2756_; 
wire _abc_40319_new_n2757_; 
wire _abc_40319_new_n2758_; 
wire _abc_40319_new_n2759_; 
wire _abc_40319_new_n2760_; 
wire _abc_40319_new_n2761_; 
wire _abc_40319_new_n2762_; 
wire _abc_40319_new_n2763_; 
wire _abc_40319_new_n2764_; 
wire _abc_40319_new_n2765_; 
wire _abc_40319_new_n2766_; 
wire _abc_40319_new_n2767_; 
wire _abc_40319_new_n2768_; 
wire _abc_40319_new_n2769_; 
wire _abc_40319_new_n2770_; 
wire _abc_40319_new_n2771_; 
wire _abc_40319_new_n2772_; 
wire _abc_40319_new_n2773_; 
wire _abc_40319_new_n2774_; 
wire _abc_40319_new_n2775_; 
wire _abc_40319_new_n2776_; 
wire _abc_40319_new_n2777_; 
wire _abc_40319_new_n2778_; 
wire _abc_40319_new_n2779_; 
wire _abc_40319_new_n2780_; 
wire _abc_40319_new_n2781_; 
wire _abc_40319_new_n2782_; 
wire _abc_40319_new_n2783_; 
wire _abc_40319_new_n2784_; 
wire _abc_40319_new_n2785_; 
wire _abc_40319_new_n2786_; 
wire _abc_40319_new_n2787_; 
wire _abc_40319_new_n2788_; 
wire _abc_40319_new_n2789_; 
wire _abc_40319_new_n2790_; 
wire _abc_40319_new_n2791_; 
wire _abc_40319_new_n2792_; 
wire _abc_40319_new_n2793_; 
wire _abc_40319_new_n2794_; 
wire _abc_40319_new_n2795_; 
wire _abc_40319_new_n2796_; 
wire _abc_40319_new_n2797_; 
wire _abc_40319_new_n2798_; 
wire _abc_40319_new_n2799_; 
wire _abc_40319_new_n2800_; 
wire _abc_40319_new_n2801_; 
wire _abc_40319_new_n2802_; 
wire _abc_40319_new_n2803_; 
wire _abc_40319_new_n2804_; 
wire _abc_40319_new_n2805_; 
wire _abc_40319_new_n2806_; 
wire _abc_40319_new_n2807_; 
wire _abc_40319_new_n2808_; 
wire _abc_40319_new_n2809_; 
wire _abc_40319_new_n2810_; 
wire _abc_40319_new_n2811_; 
wire _abc_40319_new_n2812_; 
wire _abc_40319_new_n2813_; 
wire _abc_40319_new_n2814_; 
wire _abc_40319_new_n2815_; 
wire _abc_40319_new_n2816_; 
wire _abc_40319_new_n2817_; 
wire _abc_40319_new_n2818_; 
wire _abc_40319_new_n2819_; 
wire _abc_40319_new_n2820_; 
wire _abc_40319_new_n2821_; 
wire _abc_40319_new_n2822_; 
wire _abc_40319_new_n2823_; 
wire _abc_40319_new_n2824_; 
wire _abc_40319_new_n2825_; 
wire _abc_40319_new_n2826_; 
wire _abc_40319_new_n2827_; 
wire _abc_40319_new_n2828_; 
wire _abc_40319_new_n2829_; 
wire _abc_40319_new_n2830_; 
wire _abc_40319_new_n2831_; 
wire _abc_40319_new_n2832_; 
wire _abc_40319_new_n2833_; 
wire _abc_40319_new_n2834_; 
wire _abc_40319_new_n2835_; 
wire _abc_40319_new_n2836_; 
wire _abc_40319_new_n2837_; 
wire _abc_40319_new_n2838_; 
wire _abc_40319_new_n2839_; 
wire _abc_40319_new_n2840_; 
wire _abc_40319_new_n2841_; 
wire _abc_40319_new_n2842_; 
wire _abc_40319_new_n2843_; 
wire _abc_40319_new_n2844_; 
wire _abc_40319_new_n2845_; 
wire _abc_40319_new_n2846_; 
wire _abc_40319_new_n2847_; 
wire _abc_40319_new_n2848_; 
wire _abc_40319_new_n2849_; 
wire _abc_40319_new_n2850_; 
wire _abc_40319_new_n2851_; 
wire _abc_40319_new_n2852_; 
wire _abc_40319_new_n2853_; 
wire _abc_40319_new_n2854_; 
wire _abc_40319_new_n2855_; 
wire _abc_40319_new_n2856_; 
wire _abc_40319_new_n2857_; 
wire _abc_40319_new_n2858_; 
wire _abc_40319_new_n2859_; 
wire _abc_40319_new_n2860_; 
wire _abc_40319_new_n2861_; 
wire _abc_40319_new_n2862_; 
wire _abc_40319_new_n2863_; 
wire _abc_40319_new_n2864_; 
wire _abc_40319_new_n2865_; 
wire _abc_40319_new_n2866_; 
wire _abc_40319_new_n2867_; 
wire _abc_40319_new_n2868_; 
wire _abc_40319_new_n2869_; 
wire _abc_40319_new_n2870_; 
wire _abc_40319_new_n2871_; 
wire _abc_40319_new_n2872_; 
wire _abc_40319_new_n2873_; 
wire _abc_40319_new_n2874_; 
wire _abc_40319_new_n2875_; 
wire _abc_40319_new_n2876_; 
wire _abc_40319_new_n2877_; 
wire _abc_40319_new_n2878_; 
wire _abc_40319_new_n2879_; 
wire _abc_40319_new_n2880_; 
wire _abc_40319_new_n2881_; 
wire _abc_40319_new_n2882_; 
wire _abc_40319_new_n2883_; 
wire _abc_40319_new_n2884_; 
wire _abc_40319_new_n2885_; 
wire _abc_40319_new_n2886_; 
wire _abc_40319_new_n2887_; 
wire _abc_40319_new_n2888_; 
wire _abc_40319_new_n2889_; 
wire _abc_40319_new_n2890_; 
wire _abc_40319_new_n2891_; 
wire _abc_40319_new_n2892_; 
wire _abc_40319_new_n2893_; 
wire _abc_40319_new_n2894_; 
wire _abc_40319_new_n2895_; 
wire _abc_40319_new_n2896_; 
wire _abc_40319_new_n2897_; 
wire _abc_40319_new_n2898_; 
wire _abc_40319_new_n2899_; 
wire _abc_40319_new_n2900_; 
wire _abc_40319_new_n2901_; 
wire _abc_40319_new_n2902_; 
wire _abc_40319_new_n2903_; 
wire _abc_40319_new_n2904_; 
wire _abc_40319_new_n2905_; 
wire _abc_40319_new_n2906_; 
wire _abc_40319_new_n2907_; 
wire _abc_40319_new_n2908_; 
wire _abc_40319_new_n2909_; 
wire _abc_40319_new_n2910_; 
wire _abc_40319_new_n2911_; 
wire _abc_40319_new_n2912_; 
wire _abc_40319_new_n2913_; 
wire _abc_40319_new_n2914_; 
wire _abc_40319_new_n2915_; 
wire _abc_40319_new_n2916_; 
wire _abc_40319_new_n2917_; 
wire _abc_40319_new_n2918_; 
wire _abc_40319_new_n2919_; 
wire _abc_40319_new_n2920_; 
wire _abc_40319_new_n2921_; 
wire _abc_40319_new_n2922_; 
wire _abc_40319_new_n2923_; 
wire _abc_40319_new_n2924_; 
wire _abc_40319_new_n2925_; 
wire _abc_40319_new_n2926_; 
wire _abc_40319_new_n2927_; 
wire _abc_40319_new_n2928_; 
wire _abc_40319_new_n2929_; 
wire _abc_40319_new_n2930_; 
wire _abc_40319_new_n2931_; 
wire _abc_40319_new_n2932_; 
wire _abc_40319_new_n2933_; 
wire _abc_40319_new_n2934_; 
wire _abc_40319_new_n2935_; 
wire _abc_40319_new_n2936_; 
wire _abc_40319_new_n2937_; 
wire _abc_40319_new_n2938_; 
wire _abc_40319_new_n2939_; 
wire _abc_40319_new_n2940_; 
wire _abc_40319_new_n2941_; 
wire _abc_40319_new_n2942_; 
wire _abc_40319_new_n2943_; 
wire _abc_40319_new_n2944_; 
wire _abc_40319_new_n2945_; 
wire _abc_40319_new_n2946_; 
wire _abc_40319_new_n2947_; 
wire _abc_40319_new_n2948_; 
wire _abc_40319_new_n2949_; 
wire _abc_40319_new_n2950_; 
wire _abc_40319_new_n2951_; 
wire _abc_40319_new_n2952_; 
wire _abc_40319_new_n2953_; 
wire _abc_40319_new_n2954_; 
wire _abc_40319_new_n2955_; 
wire _abc_40319_new_n2956_; 
wire _abc_40319_new_n2957_; 
wire _abc_40319_new_n2958_; 
wire _abc_40319_new_n2959_; 
wire _abc_40319_new_n2960_; 
wire _abc_40319_new_n2961_; 
wire _abc_40319_new_n2962_; 
wire _abc_40319_new_n2963_; 
wire _abc_40319_new_n2964_; 
wire _abc_40319_new_n2965_; 
wire _abc_40319_new_n2966_; 
wire _abc_40319_new_n2967_; 
wire _abc_40319_new_n2968_; 
wire _abc_40319_new_n2969_; 
wire _abc_40319_new_n2970_; 
wire _abc_40319_new_n2971_; 
wire _abc_40319_new_n2972_; 
wire _abc_40319_new_n2973_; 
wire _abc_40319_new_n2974_; 
wire _abc_40319_new_n2975_; 
wire _abc_40319_new_n2976_; 
wire _abc_40319_new_n2977_; 
wire _abc_40319_new_n2978_; 
wire _abc_40319_new_n2979_; 
wire _abc_40319_new_n2980_; 
wire _abc_40319_new_n2981_; 
wire _abc_40319_new_n2982_; 
wire _abc_40319_new_n2983_; 
wire _abc_40319_new_n2984_; 
wire _abc_40319_new_n2985_; 
wire _abc_40319_new_n2986_; 
wire _abc_40319_new_n2987_; 
wire _abc_40319_new_n2988_; 
wire _abc_40319_new_n2989_; 
wire _abc_40319_new_n2990_; 
wire _abc_40319_new_n2991_; 
wire _abc_40319_new_n2992_; 
wire _abc_40319_new_n2993_; 
wire _abc_40319_new_n2994_; 
wire _abc_40319_new_n2995_; 
wire _abc_40319_new_n2996_; 
wire _abc_40319_new_n2997_; 
wire _abc_40319_new_n2998_; 
wire _abc_40319_new_n2999_; 
wire _abc_40319_new_n3000_; 
wire _abc_40319_new_n3001_; 
wire _abc_40319_new_n3002_; 
wire _abc_40319_new_n3003_; 
wire _abc_40319_new_n3004_; 
wire _abc_40319_new_n3005_; 
wire _abc_40319_new_n3006_; 
wire _abc_40319_new_n3007_; 
wire _abc_40319_new_n3008_; 
wire _abc_40319_new_n3009_; 
wire _abc_40319_new_n3010_; 
wire _abc_40319_new_n3011_; 
wire _abc_40319_new_n3012_; 
wire _abc_40319_new_n3013_; 
wire _abc_40319_new_n3014_; 
wire _abc_40319_new_n3015_; 
wire _abc_40319_new_n3016_; 
wire _abc_40319_new_n3017_; 
wire _abc_40319_new_n3018_; 
wire _abc_40319_new_n3019_; 
wire _abc_40319_new_n3020_; 
wire _abc_40319_new_n3021_; 
wire _abc_40319_new_n3022_; 
wire _abc_40319_new_n3023_; 
wire _abc_40319_new_n3024_; 
wire _abc_40319_new_n3025_; 
wire _abc_40319_new_n3026_; 
wire _abc_40319_new_n3027_; 
wire _abc_40319_new_n3028_; 
wire _abc_40319_new_n3029_; 
wire _abc_40319_new_n3030_; 
wire _abc_40319_new_n3031_; 
wire _abc_40319_new_n3032_; 
wire _abc_40319_new_n3033_; 
wire _abc_40319_new_n3034_; 
wire _abc_40319_new_n3035_; 
wire _abc_40319_new_n3036_; 
wire _abc_40319_new_n3037_; 
wire _abc_40319_new_n3038_; 
wire _abc_40319_new_n3039_; 
wire _abc_40319_new_n3040_; 
wire _abc_40319_new_n3041_; 
wire _abc_40319_new_n3042_; 
wire _abc_40319_new_n3043_; 
wire _abc_40319_new_n3044_; 
wire _abc_40319_new_n3045_; 
wire _abc_40319_new_n3046_; 
wire _abc_40319_new_n3047_; 
wire _abc_40319_new_n3048_; 
wire _abc_40319_new_n3049_; 
wire _abc_40319_new_n3050_; 
wire _abc_40319_new_n3051_; 
wire _abc_40319_new_n3052_; 
wire _abc_40319_new_n3053_; 
wire _abc_40319_new_n3054_; 
wire _abc_40319_new_n3055_; 
wire _abc_40319_new_n3056_; 
wire _abc_40319_new_n3057_; 
wire _abc_40319_new_n3058_; 
wire _abc_40319_new_n3059_; 
wire _abc_40319_new_n3060_; 
wire _abc_40319_new_n3061_; 
wire _abc_40319_new_n3062_; 
wire _abc_40319_new_n3063_; 
wire _abc_40319_new_n3064_; 
wire _abc_40319_new_n3065_; 
wire _abc_40319_new_n3066_; 
wire _abc_40319_new_n3067_; 
wire _abc_40319_new_n3068_; 
wire _abc_40319_new_n3069_; 
wire _abc_40319_new_n3070_; 
wire _abc_40319_new_n3071_; 
wire _abc_40319_new_n3072_; 
wire _abc_40319_new_n3073_; 
wire _abc_40319_new_n3074_; 
wire _abc_40319_new_n3075_; 
wire _abc_40319_new_n3076_; 
wire _abc_40319_new_n3077_; 
wire _abc_40319_new_n3078_; 
wire _abc_40319_new_n3079_; 
wire _abc_40319_new_n3080_; 
wire _abc_40319_new_n3081_; 
wire _abc_40319_new_n3082_; 
wire _abc_40319_new_n3083_; 
wire _abc_40319_new_n3084_; 
wire _abc_40319_new_n3085_; 
wire _abc_40319_new_n3086_; 
wire _abc_40319_new_n3087_; 
wire _abc_40319_new_n3088_; 
wire _abc_40319_new_n3089_; 
wire _abc_40319_new_n3090_; 
wire _abc_40319_new_n3091_; 
wire _abc_40319_new_n3092_; 
wire _abc_40319_new_n3093_; 
wire _abc_40319_new_n3094_; 
wire _abc_40319_new_n3095_; 
wire _abc_40319_new_n3096_; 
wire _abc_40319_new_n3097_; 
wire _abc_40319_new_n3098_; 
wire _abc_40319_new_n3099_; 
wire _abc_40319_new_n3100_; 
wire _abc_40319_new_n3101_; 
wire _abc_40319_new_n3102_; 
wire _abc_40319_new_n3103_; 
wire _abc_40319_new_n3104_; 
wire _abc_40319_new_n3105_; 
wire _abc_40319_new_n3106_; 
wire _abc_40319_new_n3107_; 
wire _abc_40319_new_n3108_; 
wire _abc_40319_new_n3109_; 
wire _abc_40319_new_n3110_; 
wire _abc_40319_new_n3111_; 
wire _abc_40319_new_n3112_; 
wire _abc_40319_new_n3113_; 
wire _abc_40319_new_n3114_; 
wire _abc_40319_new_n3115_; 
wire _abc_40319_new_n3116_; 
wire _abc_40319_new_n3117_; 
wire _abc_40319_new_n3118_; 
wire _abc_40319_new_n3119_; 
wire _abc_40319_new_n3120_; 
wire _abc_40319_new_n3121_; 
wire _abc_40319_new_n3122_; 
wire _abc_40319_new_n3123_; 
wire _abc_40319_new_n3124_; 
wire _abc_40319_new_n3125_; 
wire _abc_40319_new_n3126_; 
wire _abc_40319_new_n3127_; 
wire _abc_40319_new_n3128_; 
wire _abc_40319_new_n3129_; 
wire _abc_40319_new_n3130_; 
wire _abc_40319_new_n3131_; 
wire _abc_40319_new_n3132_; 
wire _abc_40319_new_n3133_; 
wire _abc_40319_new_n3134_; 
wire _abc_40319_new_n3135_; 
wire _abc_40319_new_n3136_; 
wire _abc_40319_new_n3137_; 
wire _abc_40319_new_n3138_; 
wire _abc_40319_new_n3139_; 
wire _abc_40319_new_n3140_; 
wire _abc_40319_new_n3141_; 
wire _abc_40319_new_n3142_; 
wire _abc_40319_new_n3143_; 
wire _abc_40319_new_n3144_; 
wire _abc_40319_new_n3145_; 
wire _abc_40319_new_n3146_; 
wire _abc_40319_new_n3147_; 
wire _abc_40319_new_n3148_; 
wire _abc_40319_new_n3149_; 
wire _abc_40319_new_n3150_; 
wire _abc_40319_new_n3151_; 
wire _abc_40319_new_n3152_; 
wire _abc_40319_new_n3153_; 
wire _abc_40319_new_n3154_; 
wire _abc_40319_new_n3155_; 
wire _abc_40319_new_n3156_; 
wire _abc_40319_new_n3157_; 
wire _abc_40319_new_n3158_; 
wire _abc_40319_new_n3159_; 
wire _abc_40319_new_n3160_; 
wire _abc_40319_new_n3161_; 
wire _abc_40319_new_n3162_; 
wire _abc_40319_new_n3163_; 
wire _abc_40319_new_n3164_; 
wire _abc_40319_new_n3165_; 
wire _abc_40319_new_n3166_; 
wire _abc_40319_new_n3167_; 
wire _abc_40319_new_n3168_; 
wire _abc_40319_new_n3169_; 
wire _abc_40319_new_n3170_; 
wire _abc_40319_new_n3171_; 
wire _abc_40319_new_n3172_; 
wire _abc_40319_new_n3173_; 
wire _abc_40319_new_n3174_; 
wire _abc_40319_new_n3175_; 
wire _abc_40319_new_n3176_; 
wire _abc_40319_new_n3177_; 
wire _abc_40319_new_n3178_; 
wire _abc_40319_new_n3179_; 
wire _abc_40319_new_n3180_; 
wire _abc_40319_new_n3181_; 
wire _abc_40319_new_n3182_; 
wire _abc_40319_new_n3183_; 
wire _abc_40319_new_n3184_; 
wire _abc_40319_new_n3185_; 
wire _abc_40319_new_n3186_; 
wire _abc_40319_new_n3187_; 
wire _abc_40319_new_n3188_; 
wire _abc_40319_new_n3189_; 
wire _abc_40319_new_n3190_; 
wire _abc_40319_new_n3191_; 
wire _abc_40319_new_n3192_; 
wire _abc_40319_new_n3193_; 
wire _abc_40319_new_n3194_; 
wire _abc_40319_new_n3195_; 
wire _abc_40319_new_n3196_; 
wire _abc_40319_new_n3197_; 
wire _abc_40319_new_n3198_; 
wire _abc_40319_new_n3199_; 
wire _abc_40319_new_n3200_; 
wire _abc_40319_new_n3201_; 
wire _abc_40319_new_n3202_; 
wire _abc_40319_new_n3203_; 
wire _abc_40319_new_n3204_; 
wire _abc_40319_new_n3205_; 
wire _abc_40319_new_n3206_; 
wire _abc_40319_new_n3207_; 
wire _abc_40319_new_n3208_; 
wire _abc_40319_new_n3209_; 
wire _abc_40319_new_n3210_; 
wire _abc_40319_new_n3211_; 
wire _abc_40319_new_n3212_; 
wire _abc_40319_new_n3213_; 
wire _abc_40319_new_n3214_; 
wire _abc_40319_new_n3215_; 
wire _abc_40319_new_n3216_; 
wire _abc_40319_new_n3217_; 
wire _abc_40319_new_n3218_; 
wire _abc_40319_new_n3219_; 
wire _abc_40319_new_n3220_; 
wire _abc_40319_new_n3221_; 
wire _abc_40319_new_n3222_; 
wire _abc_40319_new_n3223_; 
wire _abc_40319_new_n3224_; 
wire _abc_40319_new_n3225_; 
wire _abc_40319_new_n3226_; 
wire _abc_40319_new_n3227_; 
wire _abc_40319_new_n3228_; 
wire _abc_40319_new_n3229_; 
wire _abc_40319_new_n3230_; 
wire _abc_40319_new_n3231_; 
wire _abc_40319_new_n3232_; 
wire _abc_40319_new_n3233_; 
wire _abc_40319_new_n3234_; 
wire _abc_40319_new_n3235_; 
wire _abc_40319_new_n3236_; 
wire _abc_40319_new_n3237_; 
wire _abc_40319_new_n3238_; 
wire _abc_40319_new_n3239_; 
wire _abc_40319_new_n3240_; 
wire _abc_40319_new_n3241_; 
wire _abc_40319_new_n3242_; 
wire _abc_40319_new_n3243_; 
wire _abc_40319_new_n3244_; 
wire _abc_40319_new_n3245_; 
wire _abc_40319_new_n3246_; 
wire _abc_40319_new_n3247_; 
wire _abc_40319_new_n3248_; 
wire _abc_40319_new_n3249_; 
wire _abc_40319_new_n3250_; 
wire _abc_40319_new_n3251_; 
wire _abc_40319_new_n3252_; 
wire _abc_40319_new_n3253_; 
wire _abc_40319_new_n3254_; 
wire _abc_40319_new_n3255_; 
wire _abc_40319_new_n3256_; 
wire _abc_40319_new_n3257_; 
wire _abc_40319_new_n3258_; 
wire _abc_40319_new_n3259_; 
wire _abc_40319_new_n3260_; 
wire _abc_40319_new_n3261_; 
wire _abc_40319_new_n3262_; 
wire _abc_40319_new_n3263_; 
wire _abc_40319_new_n3264_; 
wire _abc_40319_new_n3265_; 
wire _abc_40319_new_n3266_; 
wire _abc_40319_new_n3267_; 
wire _abc_40319_new_n3268_; 
wire _abc_40319_new_n3269_; 
wire _abc_40319_new_n3270_; 
wire _abc_40319_new_n3271_; 
wire _abc_40319_new_n3272_; 
wire _abc_40319_new_n3273_; 
wire _abc_40319_new_n3274_; 
wire _abc_40319_new_n3275_; 
wire _abc_40319_new_n3276_; 
wire _abc_40319_new_n3277_; 
wire _abc_40319_new_n3278_; 
wire _abc_40319_new_n3279_; 
wire _abc_40319_new_n3280_; 
wire _abc_40319_new_n3281_; 
wire _abc_40319_new_n3282_; 
wire _abc_40319_new_n3283_; 
wire _abc_40319_new_n3284_; 
wire _abc_40319_new_n3285_; 
wire _abc_40319_new_n3286_; 
wire _abc_40319_new_n3287_; 
wire _abc_40319_new_n3288_; 
wire _abc_40319_new_n3289_; 
wire _abc_40319_new_n3290_; 
wire _abc_40319_new_n3291_; 
wire _abc_40319_new_n3292_; 
wire _abc_40319_new_n3293_; 
wire _abc_40319_new_n3294_; 
wire _abc_40319_new_n3295_; 
wire _abc_40319_new_n3296_; 
wire _abc_40319_new_n3297_; 
wire _abc_40319_new_n3298_; 
wire _abc_40319_new_n3299_; 
wire _abc_40319_new_n3300_; 
wire _abc_40319_new_n3301_; 
wire _abc_40319_new_n3302_; 
wire _abc_40319_new_n3303_; 
wire _abc_40319_new_n3304_; 
wire _abc_40319_new_n3305_; 
wire _abc_40319_new_n3306_; 
wire _abc_40319_new_n3307_; 
wire _abc_40319_new_n3308_; 
wire _abc_40319_new_n3309_; 
wire _abc_40319_new_n3310_; 
wire _abc_40319_new_n3311_; 
wire _abc_40319_new_n3312_; 
wire _abc_40319_new_n3313_; 
wire _abc_40319_new_n3314_; 
wire _abc_40319_new_n3315_; 
wire _abc_40319_new_n3316_; 
wire _abc_40319_new_n3317_; 
wire _abc_40319_new_n3318_; 
wire _abc_40319_new_n3319_; 
wire _abc_40319_new_n3320_; 
wire _abc_40319_new_n3321_; 
wire _abc_40319_new_n3322_; 
wire _abc_40319_new_n3323_; 
wire _abc_40319_new_n3324_; 
wire _abc_40319_new_n3325_; 
wire _abc_40319_new_n3326_; 
wire _abc_40319_new_n3327_; 
wire _abc_40319_new_n3328_; 
wire _abc_40319_new_n3329_; 
wire _abc_40319_new_n3330_; 
wire _abc_40319_new_n3331_; 
wire _abc_40319_new_n3332_; 
wire _abc_40319_new_n3333_; 
wire _abc_40319_new_n3334_; 
wire _abc_40319_new_n3335_; 
wire _abc_40319_new_n3336_; 
wire _abc_40319_new_n3337_; 
wire _abc_40319_new_n3338_; 
wire _abc_40319_new_n3339_; 
wire _abc_40319_new_n3340_; 
wire _abc_40319_new_n3341_; 
wire _abc_40319_new_n3342_; 
wire _abc_40319_new_n3343_; 
wire _abc_40319_new_n3344_; 
wire _abc_40319_new_n3345_; 
wire _abc_40319_new_n3346_; 
wire _abc_40319_new_n3347_; 
wire _abc_40319_new_n3348_; 
wire _abc_40319_new_n3349_; 
wire _abc_40319_new_n3350_; 
wire _abc_40319_new_n3351_; 
wire _abc_40319_new_n3352_; 
wire _abc_40319_new_n3353_; 
wire _abc_40319_new_n3354_; 
wire _abc_40319_new_n3355_; 
wire _abc_40319_new_n3356_; 
wire _abc_40319_new_n3357_; 
wire _abc_40319_new_n3358_; 
wire _abc_40319_new_n3359_; 
wire _abc_40319_new_n3360_; 
wire _abc_40319_new_n3361_; 
wire _abc_40319_new_n3362_; 
wire _abc_40319_new_n3363_; 
wire _abc_40319_new_n3364_; 
wire _abc_40319_new_n3365_; 
wire _abc_40319_new_n3366_; 
wire _abc_40319_new_n3367_; 
wire _abc_40319_new_n3368_; 
wire _abc_40319_new_n3369_; 
wire _abc_40319_new_n3370_; 
wire _abc_40319_new_n3371_; 
wire _abc_40319_new_n3372_; 
wire _abc_40319_new_n3373_; 
wire _abc_40319_new_n3374_; 
wire _abc_40319_new_n3375_; 
wire _abc_40319_new_n3376_; 
wire _abc_40319_new_n3377_; 
wire _abc_40319_new_n3378_; 
wire _abc_40319_new_n3379_; 
wire _abc_40319_new_n3380_; 
wire _abc_40319_new_n3381_; 
wire _abc_40319_new_n3382_; 
wire _abc_40319_new_n3383_; 
wire _abc_40319_new_n3384_; 
wire _abc_40319_new_n3385_; 
wire _abc_40319_new_n3386_; 
wire _abc_40319_new_n3387_; 
wire _abc_40319_new_n3388_; 
wire _abc_40319_new_n3389_; 
wire _abc_40319_new_n3390_; 
wire _abc_40319_new_n3391_; 
wire _abc_40319_new_n3392_; 
wire _abc_40319_new_n3393_; 
wire _abc_40319_new_n3394_; 
wire _abc_40319_new_n3395_; 
wire _abc_40319_new_n3396_; 
wire _abc_40319_new_n3397_; 
wire _abc_40319_new_n3398_; 
wire _abc_40319_new_n3399_; 
wire _abc_40319_new_n3400_; 
wire _abc_40319_new_n3401_; 
wire _abc_40319_new_n3402_; 
wire _abc_40319_new_n3403_; 
wire _abc_40319_new_n3404_; 
wire _abc_40319_new_n3405_; 
wire _abc_40319_new_n3406_; 
wire _abc_40319_new_n3407_; 
wire _abc_40319_new_n3408_; 
wire _abc_40319_new_n3409_; 
wire _abc_40319_new_n3410_; 
wire _abc_40319_new_n3411_; 
wire _abc_40319_new_n3412_; 
wire _abc_40319_new_n3413_; 
wire _abc_40319_new_n3414_; 
wire _abc_40319_new_n3415_; 
wire _abc_40319_new_n3416_; 
wire _abc_40319_new_n3417_; 
wire _abc_40319_new_n3418_; 
wire _abc_40319_new_n3419_; 
wire _abc_40319_new_n3420_; 
wire _abc_40319_new_n3421_; 
wire _abc_40319_new_n3422_; 
wire _abc_40319_new_n3423_; 
wire _abc_40319_new_n3424_; 
wire _abc_40319_new_n3425_; 
wire _abc_40319_new_n3426_; 
wire _abc_40319_new_n3427_; 
wire _abc_40319_new_n3428_; 
wire _abc_40319_new_n3429_; 
wire _abc_40319_new_n3430_; 
wire _abc_40319_new_n3431_; 
wire _abc_40319_new_n3432_; 
wire _abc_40319_new_n3433_; 
wire _abc_40319_new_n3434_; 
wire _abc_40319_new_n3435_; 
wire _abc_40319_new_n3436_; 
wire _abc_40319_new_n3437_; 
wire _abc_40319_new_n3438_; 
wire _abc_40319_new_n3439_; 
wire _abc_40319_new_n3440_; 
wire _abc_40319_new_n3441_; 
wire _abc_40319_new_n3442_; 
wire _abc_40319_new_n3443_; 
wire _abc_40319_new_n3444_; 
wire _abc_40319_new_n3445_; 
wire _abc_40319_new_n3446_; 
wire _abc_40319_new_n3447_; 
wire _abc_40319_new_n3448_; 
wire _abc_40319_new_n3449_; 
wire _abc_40319_new_n3450_; 
wire _abc_40319_new_n3451_; 
wire _abc_40319_new_n3452_; 
wire _abc_40319_new_n3453_; 
wire _abc_40319_new_n3454_; 
wire _abc_40319_new_n3455_; 
wire _abc_40319_new_n3456_; 
wire _abc_40319_new_n3457_; 
wire _abc_40319_new_n3458_; 
wire _abc_40319_new_n3459_; 
wire _abc_40319_new_n3460_; 
wire _abc_40319_new_n3461_; 
wire _abc_40319_new_n3462_; 
wire _abc_40319_new_n3463_; 
wire _abc_40319_new_n3464_; 
wire _abc_40319_new_n3465_; 
wire _abc_40319_new_n3466_; 
wire _abc_40319_new_n3467_; 
wire _abc_40319_new_n3468_; 
wire _abc_40319_new_n3469_; 
wire _abc_40319_new_n3470_; 
wire _abc_40319_new_n3471_; 
wire _abc_40319_new_n3472_; 
wire _abc_40319_new_n3473_; 
wire _abc_40319_new_n3474_; 
wire _abc_40319_new_n3475_; 
wire _abc_40319_new_n3476_; 
wire _abc_40319_new_n3477_; 
wire _abc_40319_new_n3478_; 
wire _abc_40319_new_n3479_; 
wire _abc_40319_new_n3480_; 
wire _abc_40319_new_n3481_; 
wire _abc_40319_new_n3482_; 
wire _abc_40319_new_n3483_; 
wire _abc_40319_new_n3484_; 
wire _abc_40319_new_n3485_; 
wire _abc_40319_new_n3486_; 
wire _abc_40319_new_n3487_; 
wire _abc_40319_new_n3488_; 
wire _abc_40319_new_n3489_; 
wire _abc_40319_new_n3490_; 
wire _abc_40319_new_n3491_; 
wire _abc_40319_new_n3492_; 
wire _abc_40319_new_n3493_; 
wire _abc_40319_new_n3494_; 
wire _abc_40319_new_n3495_; 
wire _abc_40319_new_n3496_; 
wire _abc_40319_new_n3497_; 
wire _abc_40319_new_n3498_; 
wire _abc_40319_new_n3499_; 
wire _abc_40319_new_n3500_; 
wire _abc_40319_new_n3501_; 
wire _abc_40319_new_n3502_; 
wire _abc_40319_new_n3503_; 
wire _abc_40319_new_n3504_; 
wire _abc_40319_new_n3505_; 
wire _abc_40319_new_n3506_; 
wire _abc_40319_new_n3507_; 
wire _abc_40319_new_n3508_; 
wire _abc_40319_new_n3509_; 
wire _abc_40319_new_n3510_; 
wire _abc_40319_new_n3511_; 
wire _abc_40319_new_n3512_; 
wire _abc_40319_new_n3513_; 
wire _abc_40319_new_n3514_; 
wire _abc_40319_new_n3515_; 
wire _abc_40319_new_n3516_; 
wire _abc_40319_new_n3517_; 
wire _abc_40319_new_n3518_; 
wire _abc_40319_new_n3519_; 
wire _abc_40319_new_n3520_; 
wire _abc_40319_new_n3521_; 
wire _abc_40319_new_n3522_; 
wire _abc_40319_new_n3523_; 
wire _abc_40319_new_n3524_; 
wire _abc_40319_new_n3525_; 
wire _abc_40319_new_n3526_; 
wire _abc_40319_new_n3527_; 
wire _abc_40319_new_n3528_; 
wire _abc_40319_new_n3529_; 
wire _abc_40319_new_n3530_; 
wire _abc_40319_new_n3531_; 
wire _abc_40319_new_n3532_; 
wire _abc_40319_new_n3533_; 
wire _abc_40319_new_n3534_; 
wire _abc_40319_new_n3535_; 
wire _abc_40319_new_n3536_; 
wire _abc_40319_new_n3537_; 
wire _abc_40319_new_n3538_; 
wire _abc_40319_new_n3539_; 
wire _abc_40319_new_n3540_; 
wire _abc_40319_new_n3541_; 
wire _abc_40319_new_n3542_; 
wire _abc_40319_new_n3543_; 
wire _abc_40319_new_n3544_; 
wire _abc_40319_new_n3545_; 
wire _abc_40319_new_n3546_; 
wire _abc_40319_new_n3547_; 
wire _abc_40319_new_n3548_; 
wire _abc_40319_new_n3549_; 
wire _abc_40319_new_n3550_; 
wire _abc_40319_new_n3551_; 
wire _abc_40319_new_n3552_; 
wire _abc_40319_new_n3553_; 
wire _abc_40319_new_n3554_; 
wire _abc_40319_new_n3555_; 
wire _abc_40319_new_n3556_; 
wire _abc_40319_new_n3557_; 
wire _abc_40319_new_n3558_; 
wire _abc_40319_new_n3559_; 
wire _abc_40319_new_n3560_; 
wire _abc_40319_new_n3561_; 
wire _abc_40319_new_n3562_; 
wire _abc_40319_new_n3563_; 
wire _abc_40319_new_n3564_; 
wire _abc_40319_new_n3566_; 
wire _abc_40319_new_n3567_; 
wire _abc_40319_new_n3568_; 
wire _abc_40319_new_n3569_; 
wire _abc_40319_new_n3570_; 
wire _abc_40319_new_n3571_; 
wire _abc_40319_new_n3572_; 
wire _abc_40319_new_n3573_; 
wire _abc_40319_new_n3574_; 
wire _abc_40319_new_n3575_; 
wire _abc_40319_new_n3576_; 
wire _abc_40319_new_n3577_; 
wire _abc_40319_new_n3578_; 
wire _abc_40319_new_n3579_; 
wire _abc_40319_new_n3580_; 
wire _abc_40319_new_n3581_; 
wire _abc_40319_new_n3582_; 
wire _abc_40319_new_n3583_; 
wire _abc_40319_new_n3584_; 
wire _abc_40319_new_n3585_; 
wire _abc_40319_new_n3586_; 
wire _abc_40319_new_n3587_; 
wire _abc_40319_new_n3589_; 
wire _abc_40319_new_n3590_; 
wire _abc_40319_new_n3591_; 
wire _abc_40319_new_n3592_; 
wire _abc_40319_new_n3593_; 
wire _abc_40319_new_n3594_; 
wire _abc_40319_new_n3595_; 
wire _abc_40319_new_n3596_; 
wire _abc_40319_new_n3597_; 
wire _abc_40319_new_n3598_; 
wire _abc_40319_new_n3599_; 
wire _abc_40319_new_n3600_; 
wire _abc_40319_new_n3601_; 
wire _abc_40319_new_n3602_; 
wire _abc_40319_new_n3603_; 
wire _abc_40319_new_n3604_; 
wire _abc_40319_new_n3605_; 
wire _abc_40319_new_n3606_; 
wire _abc_40319_new_n3607_; 
wire _abc_40319_new_n3608_; 
wire _abc_40319_new_n3609_; 
wire _abc_40319_new_n3610_; 
wire _abc_40319_new_n3611_; 
wire _abc_40319_new_n3612_; 
wire _abc_40319_new_n3613_; 
wire _abc_40319_new_n3614_; 
wire _abc_40319_new_n3615_; 
wire _abc_40319_new_n3616_; 
wire _abc_40319_new_n3617_; 
wire _abc_40319_new_n3619_; 
wire _abc_40319_new_n3620_; 
wire _abc_40319_new_n3621_; 
wire _abc_40319_new_n3622_; 
wire _abc_40319_new_n3623_; 
wire _abc_40319_new_n3624_; 
wire _abc_40319_new_n3625_; 
wire _abc_40319_new_n3626_; 
wire _abc_40319_new_n3627_; 
wire _abc_40319_new_n3628_; 
wire _abc_40319_new_n3629_; 
wire _abc_40319_new_n3630_; 
wire _abc_40319_new_n3631_; 
wire _abc_40319_new_n3632_; 
wire _abc_40319_new_n3633_; 
wire _abc_40319_new_n3634_; 
wire _abc_40319_new_n3635_; 
wire _abc_40319_new_n3636_; 
wire _abc_40319_new_n3637_; 
wire _abc_40319_new_n3638_; 
wire _abc_40319_new_n3639_; 
wire _abc_40319_new_n3640_; 
wire _abc_40319_new_n3641_; 
wire _abc_40319_new_n3642_; 
wire _abc_40319_new_n3643_; 
wire _abc_40319_new_n3644_; 
wire _abc_40319_new_n3645_; 
wire _abc_40319_new_n3646_; 
wire _abc_40319_new_n3647_; 
wire _abc_40319_new_n3648_; 
wire _abc_40319_new_n3649_; 
wire _abc_40319_new_n3650_; 
wire _abc_40319_new_n3651_; 
wire _abc_40319_new_n3652_; 
wire _abc_40319_new_n3653_; 
wire _abc_40319_new_n3654_; 
wire _abc_40319_new_n3655_; 
wire _abc_40319_new_n3656_; 
wire _abc_40319_new_n3657_; 
wire _abc_40319_new_n3658_; 
wire _abc_40319_new_n3660_; 
wire _abc_40319_new_n3661_; 
wire _abc_40319_new_n3662_; 
wire _abc_40319_new_n3663_; 
wire _abc_40319_new_n3664_; 
wire _abc_40319_new_n3665_; 
wire _abc_40319_new_n3666_; 
wire _abc_40319_new_n3667_; 
wire _abc_40319_new_n3668_; 
wire _abc_40319_new_n3669_; 
wire _abc_40319_new_n3670_; 
wire _abc_40319_new_n3671_; 
wire _abc_40319_new_n3672_; 
wire _abc_40319_new_n3673_; 
wire _abc_40319_new_n3674_; 
wire _abc_40319_new_n3675_; 
wire _abc_40319_new_n3676_; 
wire _abc_40319_new_n3677_; 
wire _abc_40319_new_n3678_; 
wire _abc_40319_new_n3679_; 
wire _abc_40319_new_n3680_; 
wire _abc_40319_new_n3681_; 
wire _abc_40319_new_n3682_; 
wire _abc_40319_new_n3683_; 
wire _abc_40319_new_n3684_; 
wire _abc_40319_new_n3685_; 
wire _abc_40319_new_n3686_; 
wire _abc_40319_new_n3687_; 
wire _abc_40319_new_n3688_; 
wire _abc_40319_new_n3689_; 
wire _abc_40319_new_n3690_; 
wire _abc_40319_new_n3691_; 
wire _abc_40319_new_n3692_; 
wire _abc_40319_new_n3693_; 
wire _abc_40319_new_n3695_; 
wire _abc_40319_new_n3696_; 
wire _abc_40319_new_n3697_; 
wire _abc_40319_new_n3698_; 
wire _abc_40319_new_n3699_; 
wire _abc_40319_new_n3700_; 
wire _abc_40319_new_n3701_; 
wire _abc_40319_new_n3702_; 
wire _abc_40319_new_n3703_; 
wire _abc_40319_new_n3704_; 
wire _abc_40319_new_n3705_; 
wire _abc_40319_new_n3706_; 
wire _abc_40319_new_n3707_; 
wire _abc_40319_new_n3708_; 
wire _abc_40319_new_n3709_; 
wire _abc_40319_new_n3710_; 
wire _abc_40319_new_n3711_; 
wire _abc_40319_new_n3712_; 
wire _abc_40319_new_n3713_; 
wire _abc_40319_new_n3714_; 
wire _abc_40319_new_n3715_; 
wire _abc_40319_new_n3716_; 
wire _abc_40319_new_n3717_; 
wire _abc_40319_new_n3718_; 
wire _abc_40319_new_n3719_; 
wire _abc_40319_new_n3720_; 
wire _abc_40319_new_n3721_; 
wire _abc_40319_new_n3722_; 
wire _abc_40319_new_n3723_; 
wire _abc_40319_new_n3724_; 
wire _abc_40319_new_n3725_; 
wire _abc_40319_new_n3726_; 
wire _abc_40319_new_n3727_; 
wire _abc_40319_new_n3728_; 
wire _abc_40319_new_n3729_; 
wire _abc_40319_new_n3730_; 
wire _abc_40319_new_n3731_; 
wire _abc_40319_new_n3733_; 
wire _abc_40319_new_n3734_; 
wire _abc_40319_new_n3735_; 
wire _abc_40319_new_n3736_; 
wire _abc_40319_new_n3737_; 
wire _abc_40319_new_n3738_; 
wire _abc_40319_new_n3739_; 
wire _abc_40319_new_n3740_; 
wire _abc_40319_new_n3741_; 
wire _abc_40319_new_n3742_; 
wire _abc_40319_new_n3743_; 
wire _abc_40319_new_n3744_; 
wire _abc_40319_new_n3745_; 
wire _abc_40319_new_n3746_; 
wire _abc_40319_new_n3747_; 
wire _abc_40319_new_n3748_; 
wire _abc_40319_new_n3749_; 
wire _abc_40319_new_n3750_; 
wire _abc_40319_new_n3751_; 
wire _abc_40319_new_n3752_; 
wire _abc_40319_new_n3753_; 
wire _abc_40319_new_n3754_; 
wire _abc_40319_new_n3755_; 
wire _abc_40319_new_n3756_; 
wire _abc_40319_new_n3757_; 
wire _abc_40319_new_n3758_; 
wire _abc_40319_new_n3759_; 
wire _abc_40319_new_n3760_; 
wire _abc_40319_new_n3761_; 
wire _abc_40319_new_n3762_; 
wire _abc_40319_new_n3763_; 
wire _abc_40319_new_n3764_; 
wire _abc_40319_new_n3766_; 
wire _abc_40319_new_n3767_; 
wire _abc_40319_new_n3768_; 
wire _abc_40319_new_n3769_; 
wire _abc_40319_new_n3770_; 
wire _abc_40319_new_n3771_; 
wire _abc_40319_new_n3772_; 
wire _abc_40319_new_n3773_; 
wire _abc_40319_new_n3774_; 
wire _abc_40319_new_n3775_; 
wire _abc_40319_new_n3776_; 
wire _abc_40319_new_n3777_; 
wire _abc_40319_new_n3778_; 
wire _abc_40319_new_n3779_; 
wire _abc_40319_new_n3780_; 
wire _abc_40319_new_n3781_; 
wire _abc_40319_new_n3782_; 
wire _abc_40319_new_n3783_; 
wire _abc_40319_new_n3784_; 
wire _abc_40319_new_n3785_; 
wire _abc_40319_new_n3786_; 
wire _abc_40319_new_n3787_; 
wire _abc_40319_new_n3788_; 
wire _abc_40319_new_n3789_; 
wire _abc_40319_new_n3790_; 
wire _abc_40319_new_n3791_; 
wire _abc_40319_new_n3792_; 
wire _abc_40319_new_n3793_; 
wire _abc_40319_new_n3794_; 
wire _abc_40319_new_n3795_; 
wire _abc_40319_new_n3796_; 
wire _abc_40319_new_n3797_; 
wire _abc_40319_new_n3799_; 
wire _abc_40319_new_n3800_; 
wire _abc_40319_new_n3801_; 
wire _abc_40319_new_n3802_; 
wire _abc_40319_new_n3803_; 
wire _abc_40319_new_n3804_; 
wire _abc_40319_new_n3805_; 
wire _abc_40319_new_n3806_; 
wire _abc_40319_new_n3807_; 
wire _abc_40319_new_n3808_; 
wire _abc_40319_new_n3809_; 
wire _abc_40319_new_n3810_; 
wire _abc_40319_new_n3811_; 
wire _abc_40319_new_n3812_; 
wire _abc_40319_new_n3813_; 
wire _abc_40319_new_n3814_; 
wire _abc_40319_new_n3815_; 
wire _abc_40319_new_n3816_; 
wire _abc_40319_new_n3817_; 
wire _abc_40319_new_n3818_; 
wire _abc_40319_new_n3819_; 
wire _abc_40319_new_n3820_; 
wire _abc_40319_new_n3821_; 
wire _abc_40319_new_n3822_; 
wire _abc_40319_new_n3823_; 
wire _abc_40319_new_n3824_; 
wire _abc_40319_new_n3825_; 
wire _abc_40319_new_n3826_; 
wire _abc_40319_new_n3827_; 
wire _abc_40319_new_n3828_; 
wire _abc_40319_new_n3830_; 
wire _abc_40319_new_n3831_; 
wire _abc_40319_new_n3832_; 
wire _abc_40319_new_n3833_; 
wire _abc_40319_new_n3834_; 
wire _abc_40319_new_n3835_; 
wire _abc_40319_new_n3836_; 
wire _abc_40319_new_n3837_; 
wire _abc_40319_new_n3838_; 
wire _abc_40319_new_n3839_; 
wire _abc_40319_new_n3840_; 
wire _abc_40319_new_n3841_; 
wire _abc_40319_new_n3842_; 
wire _abc_40319_new_n3843_; 
wire _abc_40319_new_n3844_; 
wire _abc_40319_new_n3845_; 
wire _abc_40319_new_n3846_; 
wire _abc_40319_new_n3847_; 
wire _abc_40319_new_n3848_; 
wire _abc_40319_new_n3849_; 
wire _abc_40319_new_n3850_; 
wire _abc_40319_new_n3851_; 
wire _abc_40319_new_n3852_; 
wire _abc_40319_new_n3853_; 
wire _abc_40319_new_n3854_; 
wire _abc_40319_new_n3855_; 
wire _abc_40319_new_n3856_; 
wire _abc_40319_new_n3857_; 
wire _abc_40319_new_n3858_; 
wire _abc_40319_new_n3859_; 
wire _abc_40319_new_n3860_; 
wire _abc_40319_new_n3861_; 
wire _abc_40319_new_n3862_; 
wire _abc_40319_new_n3863_; 
wire _abc_40319_new_n3865_; 
wire _abc_40319_new_n3866_; 
wire _abc_40319_new_n3867_; 
wire _abc_40319_new_n3868_; 
wire _abc_40319_new_n3869_; 
wire _abc_40319_new_n3870_; 
wire _abc_40319_new_n3871_; 
wire _abc_40319_new_n3872_; 
wire _abc_40319_new_n3873_; 
wire _abc_40319_new_n3874_; 
wire _abc_40319_new_n3875_; 
wire _abc_40319_new_n3876_; 
wire _abc_40319_new_n3877_; 
wire _abc_40319_new_n3878_; 
wire _abc_40319_new_n3879_; 
wire _abc_40319_new_n3880_; 
wire _abc_40319_new_n3881_; 
wire _abc_40319_new_n3882_; 
wire _abc_40319_new_n3883_; 
wire _abc_40319_new_n3884_; 
wire _abc_40319_new_n3885_; 
wire _abc_40319_new_n3886_; 
wire _abc_40319_new_n3887_; 
wire _abc_40319_new_n3888_; 
wire _abc_40319_new_n3889_; 
wire _abc_40319_new_n3890_; 
wire _abc_40319_new_n3891_; 
wire _abc_40319_new_n3892_; 
wire _abc_40319_new_n3893_; 
wire _abc_40319_new_n3894_; 
wire _abc_40319_new_n3895_; 
wire _abc_40319_new_n3897_; 
wire _abc_40319_new_n3898_; 
wire _abc_40319_new_n3899_; 
wire _abc_40319_new_n3900_; 
wire _abc_40319_new_n3901_; 
wire _abc_40319_new_n3902_; 
wire _abc_40319_new_n3903_; 
wire _abc_40319_new_n3904_; 
wire _abc_40319_new_n3905_; 
wire _abc_40319_new_n3906_; 
wire _abc_40319_new_n3907_; 
wire _abc_40319_new_n3908_; 
wire _abc_40319_new_n3909_; 
wire _abc_40319_new_n3910_; 
wire _abc_40319_new_n3911_; 
wire _abc_40319_new_n3912_; 
wire _abc_40319_new_n3913_; 
wire _abc_40319_new_n3914_; 
wire _abc_40319_new_n3915_; 
wire _abc_40319_new_n3916_; 
wire _abc_40319_new_n3917_; 
wire _abc_40319_new_n3918_; 
wire _abc_40319_new_n3919_; 
wire _abc_40319_new_n3920_; 
wire _abc_40319_new_n3921_; 
wire _abc_40319_new_n3922_; 
wire _abc_40319_new_n3923_; 
wire _abc_40319_new_n3924_; 
wire _abc_40319_new_n3925_; 
wire _abc_40319_new_n3926_; 
wire _abc_40319_new_n3927_; 
wire _abc_40319_new_n3928_; 
wire _abc_40319_new_n3929_; 
wire _abc_40319_new_n3930_; 
wire _abc_40319_new_n3931_; 
wire _abc_40319_new_n3932_; 
wire _abc_40319_new_n3933_; 
wire _abc_40319_new_n3934_; 
wire _abc_40319_new_n3935_; 
wire _abc_40319_new_n3936_; 
wire _abc_40319_new_n3937_; 
wire _abc_40319_new_n3938_; 
wire _abc_40319_new_n3940_; 
wire _abc_40319_new_n3941_; 
wire _abc_40319_new_n3942_; 
wire _abc_40319_new_n3943_; 
wire _abc_40319_new_n3944_; 
wire _abc_40319_new_n3945_; 
wire _abc_40319_new_n3946_; 
wire _abc_40319_new_n3947_; 
wire _abc_40319_new_n3948_; 
wire _abc_40319_new_n3949_; 
wire _abc_40319_new_n3950_; 
wire _abc_40319_new_n3951_; 
wire _abc_40319_new_n3952_; 
wire _abc_40319_new_n3953_; 
wire _abc_40319_new_n3954_; 
wire _abc_40319_new_n3955_; 
wire _abc_40319_new_n3956_; 
wire _abc_40319_new_n3957_; 
wire _abc_40319_new_n3958_; 
wire _abc_40319_new_n3959_; 
wire _abc_40319_new_n3960_; 
wire _abc_40319_new_n3961_; 
wire _abc_40319_new_n3962_; 
wire _abc_40319_new_n3963_; 
wire _abc_40319_new_n3964_; 
wire _abc_40319_new_n3965_; 
wire _abc_40319_new_n3966_; 
wire _abc_40319_new_n3967_; 
wire _abc_40319_new_n3968_; 
wire _abc_40319_new_n3969_; 
wire _abc_40319_new_n3970_; 
wire _abc_40319_new_n3971_; 
wire _abc_40319_new_n3972_; 
wire _abc_40319_new_n3973_; 
wire _abc_40319_new_n3974_; 
wire _abc_40319_new_n3976_; 
wire _abc_40319_new_n3977_; 
wire _abc_40319_new_n3978_; 
wire _abc_40319_new_n3979_; 
wire _abc_40319_new_n3980_; 
wire _abc_40319_new_n3981_; 
wire _abc_40319_new_n3982_; 
wire _abc_40319_new_n3983_; 
wire _abc_40319_new_n3984_; 
wire _abc_40319_new_n3985_; 
wire _abc_40319_new_n3986_; 
wire _abc_40319_new_n3987_; 
wire _abc_40319_new_n3988_; 
wire _abc_40319_new_n3989_; 
wire _abc_40319_new_n3990_; 
wire _abc_40319_new_n3991_; 
wire _abc_40319_new_n3992_; 
wire _abc_40319_new_n3993_; 
wire _abc_40319_new_n3994_; 
wire _abc_40319_new_n3995_; 
wire _abc_40319_new_n3996_; 
wire _abc_40319_new_n3997_; 
wire _abc_40319_new_n3998_; 
wire _abc_40319_new_n3999_; 
wire _abc_40319_new_n4000_; 
wire _abc_40319_new_n4001_; 
wire _abc_40319_new_n4002_; 
wire _abc_40319_new_n4003_; 
wire _abc_40319_new_n4004_; 
wire _abc_40319_new_n4005_; 
wire _abc_40319_new_n4006_; 
wire _abc_40319_new_n4007_; 
wire _abc_40319_new_n4008_; 
wire _abc_40319_new_n4009_; 
wire _abc_40319_new_n4011_; 
wire _abc_40319_new_n4012_; 
wire _abc_40319_new_n4013_; 
wire _abc_40319_new_n4014_; 
wire _abc_40319_new_n4015_; 
wire _abc_40319_new_n4016_; 
wire _abc_40319_new_n4017_; 
wire _abc_40319_new_n4018_; 
wire _abc_40319_new_n4019_; 
wire _abc_40319_new_n4020_; 
wire _abc_40319_new_n4021_; 
wire _abc_40319_new_n4022_; 
wire _abc_40319_new_n4023_; 
wire _abc_40319_new_n4024_; 
wire _abc_40319_new_n4025_; 
wire _abc_40319_new_n4026_; 
wire _abc_40319_new_n4027_; 
wire _abc_40319_new_n4028_; 
wire _abc_40319_new_n4029_; 
wire _abc_40319_new_n4030_; 
wire _abc_40319_new_n4031_; 
wire _abc_40319_new_n4032_; 
wire _abc_40319_new_n4033_; 
wire _abc_40319_new_n4034_; 
wire _abc_40319_new_n4035_; 
wire _abc_40319_new_n4036_; 
wire _abc_40319_new_n4037_; 
wire _abc_40319_new_n4038_; 
wire _abc_40319_new_n4039_; 
wire _abc_40319_new_n4040_; 
wire _abc_40319_new_n4041_; 
wire _abc_40319_new_n4042_; 
wire _abc_40319_new_n4043_; 
wire _abc_40319_new_n4044_; 
wire _abc_40319_new_n4045_; 
wire _abc_40319_new_n4046_; 
wire _abc_40319_new_n4048_; 
wire _abc_40319_new_n4049_; 
wire _abc_40319_new_n4050_; 
wire _abc_40319_new_n4051_; 
wire _abc_40319_new_n4052_; 
wire _abc_40319_new_n4053_; 
wire _abc_40319_new_n4054_; 
wire _abc_40319_new_n4055_; 
wire _abc_40319_new_n4056_; 
wire _abc_40319_new_n4057_; 
wire _abc_40319_new_n4058_; 
wire _abc_40319_new_n4059_; 
wire _abc_40319_new_n4060_; 
wire _abc_40319_new_n4061_; 
wire _abc_40319_new_n4062_; 
wire _abc_40319_new_n4063_; 
wire _abc_40319_new_n4064_; 
wire _abc_40319_new_n4065_; 
wire _abc_40319_new_n4066_; 
wire _abc_40319_new_n4067_; 
wire _abc_40319_new_n4068_; 
wire _abc_40319_new_n4069_; 
wire _abc_40319_new_n4070_; 
wire _abc_40319_new_n4071_; 
wire _abc_40319_new_n4072_; 
wire _abc_40319_new_n4073_; 
wire _abc_40319_new_n4074_; 
wire _abc_40319_new_n4075_; 
wire _abc_40319_new_n4076_; 
wire _abc_40319_new_n4077_; 
wire _abc_40319_new_n4078_; 
wire _abc_40319_new_n4079_; 
wire _abc_40319_new_n4080_; 
wire _abc_40319_new_n4081_; 
wire _abc_40319_new_n4082_; 
wire _abc_40319_new_n4084_; 
wire _abc_40319_new_n4085_; 
wire _abc_40319_new_n4086_; 
wire _abc_40319_new_n4087_; 
wire _abc_40319_new_n4088_; 
wire _abc_40319_new_n4089_; 
wire _abc_40319_new_n4090_; 
wire _abc_40319_new_n4091_; 
wire _abc_40319_new_n4092_; 
wire _abc_40319_new_n4093_; 
wire _abc_40319_new_n4094_; 
wire _abc_40319_new_n4095_; 
wire _abc_40319_new_n4096_; 
wire _abc_40319_new_n4097_; 
wire _abc_40319_new_n4098_; 
wire _abc_40319_new_n4099_; 
wire _abc_40319_new_n4100_; 
wire _abc_40319_new_n4101_; 
wire _abc_40319_new_n4102_; 
wire _abc_40319_new_n4103_; 
wire _abc_40319_new_n4104_; 
wire _abc_40319_new_n4105_; 
wire _abc_40319_new_n4106_; 
wire _abc_40319_new_n4107_; 
wire _abc_40319_new_n4108_; 
wire _abc_40319_new_n4109_; 
wire _abc_40319_new_n4110_; 
wire _abc_40319_new_n4111_; 
wire _abc_40319_new_n4112_; 
wire _abc_40319_new_n4113_; 
wire _abc_40319_new_n4114_; 
wire _abc_40319_new_n4115_; 
wire _abc_40319_new_n4116_; 
wire _abc_40319_new_n4117_; 
wire _abc_40319_new_n4118_; 
wire _abc_40319_new_n4120_; 
wire _abc_40319_new_n4121_; 
wire _abc_40319_new_n4122_; 
wire _abc_40319_new_n4123_; 
wire _abc_40319_new_n4124_; 
wire _abc_40319_new_n4125_; 
wire _abc_40319_new_n4126_; 
wire _abc_40319_new_n4127_; 
wire _abc_40319_new_n4128_; 
wire _abc_40319_new_n4129_; 
wire _abc_40319_new_n4130_; 
wire _abc_40319_new_n4131_; 
wire _abc_40319_new_n4132_; 
wire _abc_40319_new_n4133_; 
wire _abc_40319_new_n4134_; 
wire _abc_40319_new_n4135_; 
wire _abc_40319_new_n4136_; 
wire _abc_40319_new_n4137_; 
wire _abc_40319_new_n4138_; 
wire _abc_40319_new_n4139_; 
wire _abc_40319_new_n4140_; 
wire _abc_40319_new_n4141_; 
wire _abc_40319_new_n4142_; 
wire _abc_40319_new_n4143_; 
wire _abc_40319_new_n4144_; 
wire _abc_40319_new_n4145_; 
wire _abc_40319_new_n4146_; 
wire _abc_40319_new_n4147_; 
wire _abc_40319_new_n4148_; 
wire _abc_40319_new_n4149_; 
wire _abc_40319_new_n4150_; 
wire _abc_40319_new_n4151_; 
wire _abc_40319_new_n4152_; 
wire _abc_40319_new_n4153_; 
wire _abc_40319_new_n4154_; 
wire _abc_40319_new_n4156_; 
wire _abc_40319_new_n4157_; 
wire _abc_40319_new_n4158_; 
wire _abc_40319_new_n4159_; 
wire _abc_40319_new_n4160_; 
wire _abc_40319_new_n4161_; 
wire _abc_40319_new_n4162_; 
wire _abc_40319_new_n4163_; 
wire _abc_40319_new_n4164_; 
wire _abc_40319_new_n4165_; 
wire _abc_40319_new_n4166_; 
wire _abc_40319_new_n4167_; 
wire _abc_40319_new_n4168_; 
wire _abc_40319_new_n4169_; 
wire _abc_40319_new_n4170_; 
wire _abc_40319_new_n4171_; 
wire _abc_40319_new_n4172_; 
wire _abc_40319_new_n4173_; 
wire _abc_40319_new_n4174_; 
wire _abc_40319_new_n4175_; 
wire _abc_40319_new_n4176_; 
wire _abc_40319_new_n4177_; 
wire _abc_40319_new_n4178_; 
wire _abc_40319_new_n4179_; 
wire _abc_40319_new_n4180_; 
wire _abc_40319_new_n4181_; 
wire _abc_40319_new_n4182_; 
wire _abc_40319_new_n4183_; 
wire _abc_40319_new_n4184_; 
wire _abc_40319_new_n4185_; 
wire _abc_40319_new_n4186_; 
wire _abc_40319_new_n4187_; 
wire _abc_40319_new_n4188_; 
wire _abc_40319_new_n4189_; 
wire _abc_40319_new_n4191_; 
wire _abc_40319_new_n4192_; 
wire _abc_40319_new_n4193_; 
wire _abc_40319_new_n4194_; 
wire _abc_40319_new_n4195_; 
wire _abc_40319_new_n4196_; 
wire _abc_40319_new_n4197_; 
wire _abc_40319_new_n4198_; 
wire _abc_40319_new_n4199_; 
wire _abc_40319_new_n4200_; 
wire _abc_40319_new_n4201_; 
wire _abc_40319_new_n4202_; 
wire _abc_40319_new_n4203_; 
wire _abc_40319_new_n4204_; 
wire _abc_40319_new_n4205_; 
wire _abc_40319_new_n4206_; 
wire _abc_40319_new_n4207_; 
wire _abc_40319_new_n4208_; 
wire _abc_40319_new_n4209_; 
wire _abc_40319_new_n4210_; 
wire _abc_40319_new_n4211_; 
wire _abc_40319_new_n4212_; 
wire _abc_40319_new_n4213_; 
wire _abc_40319_new_n4214_; 
wire _abc_40319_new_n4215_; 
wire _abc_40319_new_n4216_; 
wire _abc_40319_new_n4217_; 
wire _abc_40319_new_n4218_; 
wire _abc_40319_new_n4219_; 
wire _abc_40319_new_n4220_; 
wire _abc_40319_new_n4221_; 
wire _abc_40319_new_n4222_; 
wire _abc_40319_new_n4223_; 
wire _abc_40319_new_n4224_; 
wire _abc_40319_new_n4225_; 
wire _abc_40319_new_n4226_; 
wire _abc_40319_new_n4227_; 
wire _abc_40319_new_n4229_; 
wire _abc_40319_new_n4230_; 
wire _abc_40319_new_n4231_; 
wire _abc_40319_new_n4232_; 
wire _abc_40319_new_n4233_; 
wire _abc_40319_new_n4234_; 
wire _abc_40319_new_n4235_; 
wire _abc_40319_new_n4236_; 
wire _abc_40319_new_n4237_; 
wire _abc_40319_new_n4238_; 
wire _abc_40319_new_n4239_; 
wire _abc_40319_new_n4240_; 
wire _abc_40319_new_n4241_; 
wire _abc_40319_new_n4242_; 
wire _abc_40319_new_n4243_; 
wire _abc_40319_new_n4244_; 
wire _abc_40319_new_n4245_; 
wire _abc_40319_new_n4246_; 
wire _abc_40319_new_n4247_; 
wire _abc_40319_new_n4248_; 
wire _abc_40319_new_n4249_; 
wire _abc_40319_new_n4250_; 
wire _abc_40319_new_n4251_; 
wire _abc_40319_new_n4252_; 
wire _abc_40319_new_n4253_; 
wire _abc_40319_new_n4254_; 
wire _abc_40319_new_n4255_; 
wire _abc_40319_new_n4256_; 
wire _abc_40319_new_n4257_; 
wire _abc_40319_new_n4258_; 
wire _abc_40319_new_n4259_; 
wire _abc_40319_new_n4260_; 
wire _abc_40319_new_n4261_; 
wire _abc_40319_new_n4262_; 
wire _abc_40319_new_n4264_; 
wire _abc_40319_new_n4265_; 
wire _abc_40319_new_n4266_; 
wire _abc_40319_new_n4267_; 
wire _abc_40319_new_n4268_; 
wire _abc_40319_new_n4269_; 
wire _abc_40319_new_n4270_; 
wire _abc_40319_new_n4271_; 
wire _abc_40319_new_n4272_; 
wire _abc_40319_new_n4273_; 
wire _abc_40319_new_n4274_; 
wire _abc_40319_new_n4275_; 
wire _abc_40319_new_n4276_; 
wire _abc_40319_new_n4277_; 
wire _abc_40319_new_n4278_; 
wire _abc_40319_new_n4279_; 
wire _abc_40319_new_n4280_; 
wire _abc_40319_new_n4281_; 
wire _abc_40319_new_n4282_; 
wire _abc_40319_new_n4283_; 
wire _abc_40319_new_n4284_; 
wire _abc_40319_new_n4285_; 
wire _abc_40319_new_n4286_; 
wire _abc_40319_new_n4287_; 
wire _abc_40319_new_n4288_; 
wire _abc_40319_new_n4289_; 
wire _abc_40319_new_n4290_; 
wire _abc_40319_new_n4291_; 
wire _abc_40319_new_n4292_; 
wire _abc_40319_new_n4293_; 
wire _abc_40319_new_n4294_; 
wire _abc_40319_new_n4295_; 
wire _abc_40319_new_n4296_; 
wire _abc_40319_new_n4297_; 
wire _abc_40319_new_n4298_; 
wire _abc_40319_new_n4299_; 
wire _abc_40319_new_n4300_; 
wire _abc_40319_new_n4301_; 
wire _abc_40319_new_n4302_; 
wire _abc_40319_new_n4303_; 
wire _abc_40319_new_n4304_; 
wire _abc_40319_new_n4305_; 
wire _abc_40319_new_n4306_; 
wire _abc_40319_new_n4307_; 
wire _abc_40319_new_n4308_; 
wire _abc_40319_new_n4309_; 
wire _abc_40319_new_n4310_; 
wire _abc_40319_new_n4311_; 
wire _abc_40319_new_n4312_; 
wire _abc_40319_new_n4313_; 
wire _abc_40319_new_n4314_; 
wire _abc_40319_new_n4315_; 
wire _abc_40319_new_n4316_; 
wire _abc_40319_new_n4317_; 
wire _abc_40319_new_n4318_; 
wire _abc_40319_new_n4319_; 
wire _abc_40319_new_n4320_; 
wire _abc_40319_new_n4322_; 
wire _abc_40319_new_n4323_; 
wire _abc_40319_new_n4324_; 
wire _abc_40319_new_n4325_; 
wire _abc_40319_new_n4326_; 
wire _abc_40319_new_n4327_; 
wire _abc_40319_new_n4328_; 
wire _abc_40319_new_n4329_; 
wire _abc_40319_new_n4331_; 
wire _abc_40319_new_n4332_; 
wire _abc_40319_new_n4333_; 
wire _abc_40319_new_n4334_; 
wire _abc_40319_new_n4335_; 
wire _abc_40319_new_n4336_; 
wire _abc_40319_new_n4337_; 
wire _abc_40319_new_n4338_; 
wire _abc_40319_new_n4339_; 
wire _abc_40319_new_n4340_; 
wire _abc_40319_new_n4341_; 
wire _abc_40319_new_n4342_; 
wire _abc_40319_new_n4343_; 
wire _abc_40319_new_n4344_; 
wire _abc_40319_new_n4345_; 
wire _abc_40319_new_n4346_; 
wire _abc_40319_new_n4347_; 
wire _abc_40319_new_n4348_; 
wire _abc_40319_new_n4349_; 
wire _abc_40319_new_n4350_; 
wire _abc_40319_new_n4351_; 
wire _abc_40319_new_n4352_; 
wire _abc_40319_new_n4353_; 
wire _abc_40319_new_n4354_; 
wire _abc_40319_new_n4355_; 
wire _abc_40319_new_n4356_; 
wire _abc_40319_new_n4357_; 
wire _abc_40319_new_n4358_; 
wire _abc_40319_new_n4359_; 
wire _abc_40319_new_n4360_; 
wire _abc_40319_new_n4361_; 
wire _abc_40319_new_n4362_; 
wire _abc_40319_new_n4363_; 
wire _abc_40319_new_n4364_; 
wire _abc_40319_new_n4365_; 
wire _abc_40319_new_n4366_; 
wire _abc_40319_new_n4367_; 
wire _abc_40319_new_n4368_; 
wire _abc_40319_new_n4369_; 
wire _abc_40319_new_n4370_; 
wire _abc_40319_new_n4371_; 
wire _abc_40319_new_n4372_; 
wire _abc_40319_new_n4373_; 
wire _abc_40319_new_n4374_; 
wire _abc_40319_new_n4375_; 
wire _abc_40319_new_n4376_; 
wire _abc_40319_new_n4377_; 
wire _abc_40319_new_n4378_; 
wire _abc_40319_new_n4379_; 
wire _abc_40319_new_n4380_; 
wire _abc_40319_new_n4381_; 
wire _abc_40319_new_n4382_; 
wire _abc_40319_new_n4383_; 
wire _abc_40319_new_n4384_; 
wire _abc_40319_new_n4385_; 
wire _abc_40319_new_n4386_; 
wire _abc_40319_new_n4387_; 
wire _abc_40319_new_n4388_; 
wire _abc_40319_new_n4389_; 
wire _abc_40319_new_n4390_; 
wire _abc_40319_new_n4391_; 
wire _abc_40319_new_n4392_; 
wire _abc_40319_new_n4393_; 
wire _abc_40319_new_n4394_; 
wire _abc_40319_new_n4395_; 
wire _abc_40319_new_n4396_; 
wire _abc_40319_new_n4397_; 
wire _abc_40319_new_n4398_; 
wire _abc_40319_new_n4399_; 
wire _abc_40319_new_n4400_; 
wire _abc_40319_new_n4401_; 
wire _abc_40319_new_n4402_; 
wire _abc_40319_new_n4403_; 
wire _abc_40319_new_n4404_; 
wire _abc_40319_new_n4405_; 
wire _abc_40319_new_n4406_; 
wire _abc_40319_new_n4407_; 
wire _abc_40319_new_n4408_; 
wire _abc_40319_new_n4409_; 
wire _abc_40319_new_n4410_; 
wire _abc_40319_new_n4411_; 
wire _abc_40319_new_n4412_; 
wire _abc_40319_new_n4413_; 
wire _abc_40319_new_n4414_; 
wire _abc_40319_new_n4415_; 
wire _abc_40319_new_n4416_; 
wire _abc_40319_new_n4417_; 
wire _abc_40319_new_n4418_; 
wire _abc_40319_new_n4419_; 
wire _abc_40319_new_n4420_; 
wire _abc_40319_new_n4421_; 
wire _abc_40319_new_n4422_; 
wire _abc_40319_new_n4423_; 
wire _abc_40319_new_n4424_; 
wire _abc_40319_new_n4425_; 
wire _abc_40319_new_n4426_; 
wire _abc_40319_new_n4427_; 
wire _abc_40319_new_n4428_; 
wire _abc_40319_new_n4429_; 
wire _abc_40319_new_n4430_; 
wire _abc_40319_new_n4431_; 
wire _abc_40319_new_n4432_; 
wire _abc_40319_new_n4433_; 
wire _abc_40319_new_n4434_; 
wire _abc_40319_new_n4435_; 
wire _abc_40319_new_n4436_; 
wire _abc_40319_new_n4437_; 
wire _abc_40319_new_n4438_; 
wire _abc_40319_new_n4439_; 
wire _abc_40319_new_n4440_; 
wire _abc_40319_new_n4441_; 
wire _abc_40319_new_n4442_; 
wire _abc_40319_new_n4443_; 
wire _abc_40319_new_n4444_; 
wire _abc_40319_new_n4445_; 
wire _abc_40319_new_n4446_; 
wire _abc_40319_new_n4447_; 
wire _abc_40319_new_n4448_; 
wire _abc_40319_new_n4449_; 
wire _abc_40319_new_n4450_; 
wire _abc_40319_new_n4451_; 
wire _abc_40319_new_n4452_; 
wire _abc_40319_new_n4453_; 
wire _abc_40319_new_n4454_; 
wire _abc_40319_new_n4455_; 
wire _abc_40319_new_n4456_; 
wire _abc_40319_new_n4457_; 
wire _abc_40319_new_n4458_; 
wire _abc_40319_new_n4459_; 
wire _abc_40319_new_n4460_; 
wire _abc_40319_new_n4461_; 
wire _abc_40319_new_n4462_; 
wire _abc_40319_new_n4463_; 
wire _abc_40319_new_n4464_; 
wire _abc_40319_new_n4465_; 
wire _abc_40319_new_n4466_; 
wire _abc_40319_new_n4467_; 
wire _abc_40319_new_n4468_; 
wire _abc_40319_new_n4469_; 
wire _abc_40319_new_n4470_; 
wire _abc_40319_new_n4471_; 
wire _abc_40319_new_n4472_; 
wire _abc_40319_new_n4473_; 
wire _abc_40319_new_n4474_; 
wire _abc_40319_new_n4475_; 
wire _abc_40319_new_n4476_; 
wire _abc_40319_new_n4477_; 
wire _abc_40319_new_n4478_; 
wire _abc_40319_new_n4479_; 
wire _abc_40319_new_n4480_; 
wire _abc_40319_new_n4481_; 
wire _abc_40319_new_n4482_; 
wire _abc_40319_new_n4483_; 
wire _abc_40319_new_n4484_; 
wire _abc_40319_new_n4485_; 
wire _abc_40319_new_n4486_; 
wire _abc_40319_new_n4487_; 
wire _abc_40319_new_n4488_; 
wire _abc_40319_new_n4489_; 
wire _abc_40319_new_n4490_; 
wire _abc_40319_new_n4491_; 
wire _abc_40319_new_n4492_; 
wire _abc_40319_new_n4493_; 
wire _abc_40319_new_n4494_; 
wire _abc_40319_new_n4495_; 
wire _abc_40319_new_n4496_; 
wire _abc_40319_new_n4497_; 
wire _abc_40319_new_n4498_; 
wire _abc_40319_new_n4499_; 
wire _abc_40319_new_n4500_; 
wire _abc_40319_new_n4501_; 
wire _abc_40319_new_n4502_; 
wire _abc_40319_new_n4503_; 
wire _abc_40319_new_n4504_; 
wire _abc_40319_new_n4505_; 
wire _abc_40319_new_n4506_; 
wire _abc_40319_new_n4507_; 
wire _abc_40319_new_n4508_; 
wire _abc_40319_new_n4509_; 
wire _abc_40319_new_n4510_; 
wire _abc_40319_new_n4511_; 
wire _abc_40319_new_n4512_; 
wire _abc_40319_new_n4513_; 
wire _abc_40319_new_n4514_; 
wire _abc_40319_new_n4515_; 
wire _abc_40319_new_n4516_; 
wire _abc_40319_new_n4517_; 
wire _abc_40319_new_n4518_; 
wire _abc_40319_new_n4519_; 
wire _abc_40319_new_n4520_; 
wire _abc_40319_new_n4521_; 
wire _abc_40319_new_n4522_; 
wire _abc_40319_new_n4523_; 
wire _abc_40319_new_n4524_; 
wire _abc_40319_new_n4525_; 
wire _abc_40319_new_n4526_; 
wire _abc_40319_new_n4527_; 
wire _abc_40319_new_n4528_; 
wire _abc_40319_new_n4529_; 
wire _abc_40319_new_n4531_; 
wire _abc_40319_new_n4532_; 
wire _abc_40319_new_n4533_; 
wire _abc_40319_new_n4534_; 
wire _abc_40319_new_n4535_; 
wire _abc_40319_new_n4536_; 
wire _abc_40319_new_n4537_; 
wire _abc_40319_new_n4538_; 
wire _abc_40319_new_n4539_; 
wire _abc_40319_new_n4540_; 
wire _abc_40319_new_n4541_; 
wire _abc_40319_new_n4542_; 
wire _abc_40319_new_n4543_; 
wire _abc_40319_new_n4544_; 
wire _abc_40319_new_n4545_; 
wire _abc_40319_new_n4546_; 
wire _abc_40319_new_n4547_; 
wire _abc_40319_new_n4548_; 
wire _abc_40319_new_n4549_; 
wire _abc_40319_new_n4550_; 
wire _abc_40319_new_n4551_; 
wire _abc_40319_new_n4552_; 
wire _abc_40319_new_n4553_; 
wire _abc_40319_new_n4554_; 
wire _abc_40319_new_n4555_; 
wire _abc_40319_new_n4556_; 
wire _abc_40319_new_n4557_; 
wire _abc_40319_new_n4558_; 
wire _abc_40319_new_n4559_; 
wire _abc_40319_new_n4560_; 
wire _abc_40319_new_n4561_; 
wire _abc_40319_new_n4562_; 
wire _abc_40319_new_n4563_; 
wire _abc_40319_new_n4564_; 
wire _abc_40319_new_n4565_; 
wire _abc_40319_new_n4567_; 
wire _abc_40319_new_n4568_; 
wire _abc_40319_new_n4569_; 
wire _abc_40319_new_n4570_; 
wire _abc_40319_new_n4571_; 
wire _abc_40319_new_n4572_; 
wire _abc_40319_new_n4573_; 
wire _abc_40319_new_n4574_; 
wire _abc_40319_new_n4575_; 
wire _abc_40319_new_n4576_; 
wire _abc_40319_new_n4577_; 
wire _abc_40319_new_n4578_; 
wire _abc_40319_new_n4579_; 
wire _abc_40319_new_n4580_; 
wire _abc_40319_new_n4581_; 
wire _abc_40319_new_n4582_; 
wire _abc_40319_new_n4583_; 
wire _abc_40319_new_n4584_; 
wire _abc_40319_new_n4585_; 
wire _abc_40319_new_n4586_; 
wire _abc_40319_new_n4587_; 
wire _abc_40319_new_n4588_; 
wire _abc_40319_new_n4589_; 
wire _abc_40319_new_n4590_; 
wire _abc_40319_new_n4591_; 
wire _abc_40319_new_n4592_; 
wire _abc_40319_new_n4593_; 
wire _abc_40319_new_n4594_; 
wire _abc_40319_new_n4595_; 
wire _abc_40319_new_n4596_; 
wire _abc_40319_new_n4597_; 
wire _abc_40319_new_n4598_; 
wire _abc_40319_new_n4599_; 
wire _abc_40319_new_n4600_; 
wire _abc_40319_new_n4601_; 
wire _abc_40319_new_n4602_; 
wire _abc_40319_new_n4603_; 
wire _abc_40319_new_n4604_; 
wire _abc_40319_new_n4606_; 
wire _abc_40319_new_n4607_; 
wire _abc_40319_new_n4608_; 
wire _abc_40319_new_n4609_; 
wire _abc_40319_new_n4610_; 
wire _abc_40319_new_n4611_; 
wire _abc_40319_new_n4612_; 
wire _abc_40319_new_n4613_; 
wire _abc_40319_new_n4614_; 
wire _abc_40319_new_n4615_; 
wire _abc_40319_new_n4616_; 
wire _abc_40319_new_n4617_; 
wire _abc_40319_new_n4618_; 
wire _abc_40319_new_n4619_; 
wire _abc_40319_new_n4620_; 
wire _abc_40319_new_n4621_; 
wire _abc_40319_new_n4622_; 
wire _abc_40319_new_n4623_; 
wire _abc_40319_new_n4624_; 
wire _abc_40319_new_n4625_; 
wire _abc_40319_new_n4626_; 
wire _abc_40319_new_n4627_; 
wire _abc_40319_new_n4628_; 
wire _abc_40319_new_n4629_; 
wire _abc_40319_new_n4630_; 
wire _abc_40319_new_n4631_; 
wire _abc_40319_new_n4632_; 
wire _abc_40319_new_n4633_; 
wire _abc_40319_new_n4634_; 
wire _abc_40319_new_n4635_; 
wire _abc_40319_new_n4637_; 
wire _abc_40319_new_n4638_; 
wire _abc_40319_new_n4639_; 
wire _abc_40319_new_n4640_; 
wire _abc_40319_new_n4641_; 
wire _abc_40319_new_n4642_; 
wire _abc_40319_new_n4643_; 
wire _abc_40319_new_n4644_; 
wire _abc_40319_new_n4645_; 
wire _abc_40319_new_n4646_; 
wire _abc_40319_new_n4647_; 
wire _abc_40319_new_n4648_; 
wire _abc_40319_new_n4649_; 
wire _abc_40319_new_n4650_; 
wire _abc_40319_new_n4651_; 
wire _abc_40319_new_n4652_; 
wire _abc_40319_new_n4653_; 
wire _abc_40319_new_n4654_; 
wire _abc_40319_new_n4655_; 
wire _abc_40319_new_n4656_; 
wire _abc_40319_new_n4657_; 
wire _abc_40319_new_n4658_; 
wire _abc_40319_new_n4659_; 
wire _abc_40319_new_n4660_; 
wire _abc_40319_new_n4661_; 
wire _abc_40319_new_n4662_; 
wire _abc_40319_new_n4663_; 
wire _abc_40319_new_n4664_; 
wire _abc_40319_new_n4665_; 
wire _abc_40319_new_n4666_; 
wire _abc_40319_new_n4667_; 
wire _abc_40319_new_n4668_; 
wire _abc_40319_new_n4669_; 
wire _abc_40319_new_n4670_; 
wire _abc_40319_new_n4671_; 
wire _abc_40319_new_n4672_; 
wire _abc_40319_new_n4673_; 
wire _abc_40319_new_n4674_; 
wire _abc_40319_new_n4675_; 
wire _abc_40319_new_n4676_; 
wire _abc_40319_new_n4677_; 
wire _abc_40319_new_n4678_; 
wire _abc_40319_new_n4679_; 
wire _abc_40319_new_n4680_; 
wire _abc_40319_new_n4681_; 
wire _abc_40319_new_n4683_; 
wire _abc_40319_new_n4684_; 
wire _abc_40319_new_n4685_; 
wire _abc_40319_new_n4686_; 
wire _abc_40319_new_n4687_; 
wire _abc_40319_new_n4688_; 
wire _abc_40319_new_n4689_; 
wire _abc_40319_new_n4690_; 
wire _abc_40319_new_n4691_; 
wire _abc_40319_new_n4692_; 
wire _abc_40319_new_n4693_; 
wire _abc_40319_new_n4694_; 
wire _abc_40319_new_n4695_; 
wire _abc_40319_new_n4696_; 
wire _abc_40319_new_n4697_; 
wire _abc_40319_new_n4698_; 
wire _abc_40319_new_n4699_; 
wire _abc_40319_new_n4700_; 
wire _abc_40319_new_n4701_; 
wire _abc_40319_new_n4702_; 
wire _abc_40319_new_n4703_; 
wire _abc_40319_new_n4704_; 
wire _abc_40319_new_n4705_; 
wire _abc_40319_new_n4706_; 
wire _abc_40319_new_n4707_; 
wire _abc_40319_new_n4708_; 
wire _abc_40319_new_n4709_; 
wire _abc_40319_new_n4710_; 
wire _abc_40319_new_n4711_; 
wire _abc_40319_new_n4712_; 
wire _abc_40319_new_n4713_; 
wire _abc_40319_new_n4714_; 
wire _abc_40319_new_n4715_; 
wire _abc_40319_new_n4716_; 
wire _abc_40319_new_n4717_; 
wire _abc_40319_new_n4718_; 
wire _abc_40319_new_n4719_; 
wire _abc_40319_new_n4720_; 
wire _abc_40319_new_n4721_; 
wire _abc_40319_new_n4722_; 
wire _abc_40319_new_n4723_; 
wire _abc_40319_new_n4725_; 
wire _abc_40319_new_n4726_; 
wire _abc_40319_new_n4727_; 
wire _abc_40319_new_n4728_; 
wire _abc_40319_new_n4729_; 
wire _abc_40319_new_n4730_; 
wire _abc_40319_new_n4731_; 
wire _abc_40319_new_n4732_; 
wire _abc_40319_new_n4733_; 
wire _abc_40319_new_n4734_; 
wire _abc_40319_new_n4735_; 
wire _abc_40319_new_n4736_; 
wire _abc_40319_new_n4737_; 
wire _abc_40319_new_n4738_; 
wire _abc_40319_new_n4739_; 
wire _abc_40319_new_n4740_; 
wire _abc_40319_new_n4741_; 
wire _abc_40319_new_n4742_; 
wire _abc_40319_new_n4743_; 
wire _abc_40319_new_n4744_; 
wire _abc_40319_new_n4745_; 
wire _abc_40319_new_n4746_; 
wire _abc_40319_new_n4747_; 
wire _abc_40319_new_n4748_; 
wire _abc_40319_new_n4749_; 
wire _abc_40319_new_n4750_; 
wire _abc_40319_new_n4751_; 
wire _abc_40319_new_n4752_; 
wire _abc_40319_new_n4753_; 
wire _abc_40319_new_n4754_; 
wire _abc_40319_new_n4756_; 
wire _abc_40319_new_n4757_; 
wire _abc_40319_new_n4758_; 
wire _abc_40319_new_n4759_; 
wire _abc_40319_new_n4760_; 
wire _abc_40319_new_n4761_; 
wire _abc_40319_new_n4762_; 
wire _abc_40319_new_n4763_; 
wire _abc_40319_new_n4764_; 
wire _abc_40319_new_n4765_; 
wire _abc_40319_new_n4766_; 
wire _abc_40319_new_n4767_; 
wire _abc_40319_new_n4768_; 
wire _abc_40319_new_n4769_; 
wire _abc_40319_new_n4770_; 
wire _abc_40319_new_n4771_; 
wire _abc_40319_new_n4772_; 
wire _abc_40319_new_n4773_; 
wire _abc_40319_new_n4774_; 
wire _abc_40319_new_n4775_; 
wire _abc_40319_new_n4776_; 
wire _abc_40319_new_n4777_; 
wire _abc_40319_new_n4778_; 
wire _abc_40319_new_n4779_; 
wire _abc_40319_new_n4780_; 
wire _abc_40319_new_n4781_; 
wire _abc_40319_new_n4782_; 
wire _abc_40319_new_n4783_; 
wire _abc_40319_new_n4784_; 
wire _abc_40319_new_n4785_; 
wire _abc_40319_new_n4786_; 
wire _abc_40319_new_n4787_; 
wire _abc_40319_new_n4788_; 
wire _abc_40319_new_n4789_; 
wire _abc_40319_new_n4790_; 
wire _abc_40319_new_n4791_; 
wire _abc_40319_new_n4793_; 
wire _abc_40319_new_n4794_; 
wire _abc_40319_new_n4795_; 
wire _abc_40319_new_n4796_; 
wire _abc_40319_new_n4797_; 
wire _abc_40319_new_n4798_; 
wire _abc_40319_new_n4799_; 
wire _abc_40319_new_n4800_; 
wire _abc_40319_new_n4801_; 
wire _abc_40319_new_n4802_; 
wire _abc_40319_new_n4803_; 
wire _abc_40319_new_n4804_; 
wire _abc_40319_new_n4805_; 
wire _abc_40319_new_n4806_; 
wire _abc_40319_new_n4807_; 
wire _abc_40319_new_n4808_; 
wire _abc_40319_new_n4809_; 
wire _abc_40319_new_n4810_; 
wire _abc_40319_new_n4811_; 
wire _abc_40319_new_n4812_; 
wire _abc_40319_new_n4813_; 
wire _abc_40319_new_n4814_; 
wire _abc_40319_new_n4815_; 
wire _abc_40319_new_n4816_; 
wire _abc_40319_new_n4817_; 
wire _abc_40319_new_n4818_; 
wire _abc_40319_new_n4819_; 
wire _abc_40319_new_n4820_; 
wire _abc_40319_new_n4821_; 
wire _abc_40319_new_n4822_; 
wire _abc_40319_new_n4823_; 
wire _abc_40319_new_n4824_; 
wire _abc_40319_new_n4825_; 
wire _abc_40319_new_n4826_; 
wire _abc_40319_new_n4827_; 
wire _abc_40319_new_n4829_; 
wire _abc_40319_new_n4830_; 
wire _abc_40319_new_n4831_; 
wire _abc_40319_new_n4832_; 
wire _abc_40319_new_n4833_; 
wire _abc_40319_new_n4834_; 
wire _abc_40319_new_n4835_; 
wire _abc_40319_new_n4836_; 
wire _abc_40319_new_n4837_; 
wire _abc_40319_new_n4838_; 
wire _abc_40319_new_n4839_; 
wire _abc_40319_new_n4840_; 
wire _abc_40319_new_n4841_; 
wire _abc_40319_new_n4842_; 
wire _abc_40319_new_n4843_; 
wire _abc_40319_new_n4844_; 
wire _abc_40319_new_n4845_; 
wire _abc_40319_new_n4846_; 
wire _abc_40319_new_n4847_; 
wire _abc_40319_new_n4848_; 
wire _abc_40319_new_n4849_; 
wire _abc_40319_new_n4850_; 
wire _abc_40319_new_n4851_; 
wire _abc_40319_new_n4852_; 
wire _abc_40319_new_n4853_; 
wire _abc_40319_new_n4854_; 
wire _abc_40319_new_n4855_; 
wire _abc_40319_new_n4856_; 
wire _abc_40319_new_n4857_; 
wire _abc_40319_new_n4858_; 
wire _abc_40319_new_n4860_; 
wire _abc_40319_new_n4861_; 
wire _abc_40319_new_n4862_; 
wire _abc_40319_new_n4863_; 
wire _abc_40319_new_n4864_; 
wire _abc_40319_new_n4865_; 
wire _abc_40319_new_n4866_; 
wire _abc_40319_new_n4867_; 
wire _abc_40319_new_n4868_; 
wire _abc_40319_new_n4869_; 
wire _abc_40319_new_n4870_; 
wire _abc_40319_new_n4871_; 
wire _abc_40319_new_n4872_; 
wire _abc_40319_new_n4873_; 
wire _abc_40319_new_n4874_; 
wire _abc_40319_new_n4875_; 
wire _abc_40319_new_n4876_; 
wire _abc_40319_new_n4877_; 
wire _abc_40319_new_n4878_; 
wire _abc_40319_new_n4879_; 
wire _abc_40319_new_n4880_; 
wire _abc_40319_new_n4881_; 
wire _abc_40319_new_n4882_; 
wire _abc_40319_new_n4883_; 
wire _abc_40319_new_n4884_; 
wire _abc_40319_new_n4885_; 
wire _abc_40319_new_n4886_; 
wire _abc_40319_new_n4887_; 
wire _abc_40319_new_n4888_; 
wire _abc_40319_new_n4889_; 
wire _abc_40319_new_n4890_; 
wire _abc_40319_new_n4892_; 
wire _abc_40319_new_n4893_; 
wire _abc_40319_new_n4894_; 
wire _abc_40319_new_n4895_; 
wire _abc_40319_new_n4896_; 
wire _abc_40319_new_n4897_; 
wire _abc_40319_new_n4898_; 
wire _abc_40319_new_n4899_; 
wire _abc_40319_new_n4900_; 
wire _abc_40319_new_n4901_; 
wire _abc_40319_new_n4902_; 
wire _abc_40319_new_n4903_; 
wire _abc_40319_new_n4904_; 
wire _abc_40319_new_n4905_; 
wire _abc_40319_new_n4906_; 
wire _abc_40319_new_n4907_; 
wire _abc_40319_new_n4908_; 
wire _abc_40319_new_n4909_; 
wire _abc_40319_new_n4910_; 
wire _abc_40319_new_n4911_; 
wire _abc_40319_new_n4912_; 
wire _abc_40319_new_n4913_; 
wire _abc_40319_new_n4914_; 
wire _abc_40319_new_n4915_; 
wire _abc_40319_new_n4916_; 
wire _abc_40319_new_n4917_; 
wire _abc_40319_new_n4918_; 
wire _abc_40319_new_n4919_; 
wire _abc_40319_new_n4920_; 
wire _abc_40319_new_n4921_; 
wire _abc_40319_new_n4922_; 
wire _abc_40319_new_n4923_; 
wire _abc_40319_new_n4924_; 
wire _abc_40319_new_n4925_; 
wire _abc_40319_new_n4926_; 
wire _abc_40319_new_n4928_; 
wire _abc_40319_new_n4929_; 
wire _abc_40319_new_n4930_; 
wire _abc_40319_new_n4931_; 
wire _abc_40319_new_n4932_; 
wire _abc_40319_new_n4933_; 
wire _abc_40319_new_n4934_; 
wire _abc_40319_new_n4935_; 
wire _abc_40319_new_n4936_; 
wire _abc_40319_new_n4937_; 
wire _abc_40319_new_n4938_; 
wire _abc_40319_new_n4939_; 
wire _abc_40319_new_n4940_; 
wire _abc_40319_new_n4941_; 
wire _abc_40319_new_n4942_; 
wire _abc_40319_new_n4943_; 
wire _abc_40319_new_n4944_; 
wire _abc_40319_new_n4945_; 
wire _abc_40319_new_n4946_; 
wire _abc_40319_new_n4947_; 
wire _abc_40319_new_n4948_; 
wire _abc_40319_new_n4949_; 
wire _abc_40319_new_n4950_; 
wire _abc_40319_new_n4951_; 
wire _abc_40319_new_n4952_; 
wire _abc_40319_new_n4953_; 
wire _abc_40319_new_n4954_; 
wire _abc_40319_new_n4955_; 
wire _abc_40319_new_n4956_; 
wire _abc_40319_new_n4957_; 
wire _abc_40319_new_n4958_; 
wire _abc_40319_new_n4959_; 
wire _abc_40319_new_n4960_; 
wire _abc_40319_new_n4961_; 
wire _abc_40319_new_n4962_; 
wire _abc_40319_new_n4964_; 
wire _abc_40319_new_n4965_; 
wire _abc_40319_new_n4966_; 
wire _abc_40319_new_n4967_; 
wire _abc_40319_new_n4968_; 
wire _abc_40319_new_n4969_; 
wire _abc_40319_new_n4970_; 
wire _abc_40319_new_n4971_; 
wire _abc_40319_new_n4972_; 
wire _abc_40319_new_n4973_; 
wire _abc_40319_new_n4974_; 
wire _abc_40319_new_n4975_; 
wire _abc_40319_new_n4976_; 
wire _abc_40319_new_n4977_; 
wire _abc_40319_new_n4978_; 
wire _abc_40319_new_n4979_; 
wire _abc_40319_new_n4980_; 
wire _abc_40319_new_n4981_; 
wire _abc_40319_new_n4982_; 
wire _abc_40319_new_n4983_; 
wire _abc_40319_new_n4984_; 
wire _abc_40319_new_n4985_; 
wire _abc_40319_new_n4986_; 
wire _abc_40319_new_n4987_; 
wire _abc_40319_new_n4988_; 
wire _abc_40319_new_n4989_; 
wire _abc_40319_new_n4990_; 
wire _abc_40319_new_n4991_; 
wire _abc_40319_new_n4992_; 
wire _abc_40319_new_n4993_; 
wire _abc_40319_new_n4995_; 
wire _abc_40319_new_n4996_; 
wire _abc_40319_new_n4997_; 
wire _abc_40319_new_n4998_; 
wire _abc_40319_new_n4999_; 
wire _abc_40319_new_n5000_; 
wire _abc_40319_new_n5001_; 
wire _abc_40319_new_n5002_; 
wire _abc_40319_new_n5003_; 
wire _abc_40319_new_n5004_; 
wire _abc_40319_new_n5005_; 
wire _abc_40319_new_n5006_; 
wire _abc_40319_new_n5007_; 
wire _abc_40319_new_n5008_; 
wire _abc_40319_new_n5009_; 
wire _abc_40319_new_n5010_; 
wire _abc_40319_new_n5011_; 
wire _abc_40319_new_n5012_; 
wire _abc_40319_new_n5013_; 
wire _abc_40319_new_n5014_; 
wire _abc_40319_new_n5015_; 
wire _abc_40319_new_n5016_; 
wire _abc_40319_new_n5017_; 
wire _abc_40319_new_n5018_; 
wire _abc_40319_new_n5019_; 
wire _abc_40319_new_n5020_; 
wire _abc_40319_new_n5021_; 
wire _abc_40319_new_n5022_; 
wire _abc_40319_new_n5024_; 
wire _abc_40319_new_n5025_; 
wire _abc_40319_new_n5026_; 
wire _abc_40319_new_n5027_; 
wire _abc_40319_new_n5028_; 
wire _abc_40319_new_n5029_; 
wire _abc_40319_new_n5030_; 
wire _abc_40319_new_n5031_; 
wire _abc_40319_new_n5032_; 
wire _abc_40319_new_n5033_; 
wire _abc_40319_new_n5034_; 
wire _abc_40319_new_n5035_; 
wire _abc_40319_new_n5036_; 
wire _abc_40319_new_n5037_; 
wire _abc_40319_new_n5038_; 
wire _abc_40319_new_n5039_; 
wire _abc_40319_new_n5040_; 
wire _abc_40319_new_n5041_; 
wire _abc_40319_new_n5042_; 
wire _abc_40319_new_n5043_; 
wire _abc_40319_new_n5044_; 
wire _abc_40319_new_n5045_; 
wire _abc_40319_new_n5046_; 
wire _abc_40319_new_n5047_; 
wire _abc_40319_new_n5048_; 
wire _abc_40319_new_n5049_; 
wire _abc_40319_new_n5050_; 
wire _abc_40319_new_n5051_; 
wire _abc_40319_new_n5052_; 
wire _abc_40319_new_n5053_; 
wire _abc_40319_new_n5054_; 
wire _abc_40319_new_n5055_; 
wire _abc_40319_new_n5056_; 
wire _abc_40319_new_n5058_; 
wire _abc_40319_new_n5059_; 
wire _abc_40319_new_n5060_; 
wire _abc_40319_new_n5061_; 
wire _abc_40319_new_n5062_; 
wire _abc_40319_new_n5063_; 
wire _abc_40319_new_n5064_; 
wire _abc_40319_new_n5065_; 
wire _abc_40319_new_n5066_; 
wire _abc_40319_new_n5067_; 
wire _abc_40319_new_n5068_; 
wire _abc_40319_new_n5069_; 
wire _abc_40319_new_n5070_; 
wire _abc_40319_new_n5071_; 
wire _abc_40319_new_n5072_; 
wire _abc_40319_new_n5073_; 
wire _abc_40319_new_n5074_; 
wire _abc_40319_new_n5075_; 
wire _abc_40319_new_n5076_; 
wire _abc_40319_new_n5077_; 
wire _abc_40319_new_n5078_; 
wire _abc_40319_new_n5079_; 
wire _abc_40319_new_n5080_; 
wire _abc_40319_new_n5081_; 
wire _abc_40319_new_n5082_; 
wire _abc_40319_new_n5083_; 
wire _abc_40319_new_n5084_; 
wire _abc_40319_new_n5085_; 
wire _abc_40319_new_n5086_; 
wire _abc_40319_new_n5087_; 
wire _abc_40319_new_n5089_; 
wire _abc_40319_new_n5090_; 
wire _abc_40319_new_n5091_; 
wire _abc_40319_new_n5092_; 
wire _abc_40319_new_n5093_; 
wire _abc_40319_new_n5094_; 
wire _abc_40319_new_n5095_; 
wire _abc_40319_new_n5096_; 
wire _abc_40319_new_n5097_; 
wire _abc_40319_new_n5098_; 
wire _abc_40319_new_n5099_; 
wire _abc_40319_new_n5100_; 
wire _abc_40319_new_n5101_; 
wire _abc_40319_new_n5102_; 
wire _abc_40319_new_n5103_; 
wire _abc_40319_new_n5104_; 
wire _abc_40319_new_n5105_; 
wire _abc_40319_new_n5106_; 
wire _abc_40319_new_n5107_; 
wire _abc_40319_new_n5108_; 
wire _abc_40319_new_n5109_; 
wire _abc_40319_new_n5110_; 
wire _abc_40319_new_n5111_; 
wire _abc_40319_new_n5112_; 
wire _abc_40319_new_n5113_; 
wire _abc_40319_new_n5114_; 
wire _abc_40319_new_n5115_; 
wire _abc_40319_new_n5116_; 
wire _abc_40319_new_n5117_; 
wire _abc_40319_new_n5118_; 
wire _abc_40319_new_n5119_; 
wire _abc_40319_new_n5120_; 
wire _abc_40319_new_n5121_; 
wire _abc_40319_new_n5122_; 
wire _abc_40319_new_n5123_; 
wire _abc_40319_new_n5125_; 
wire _abc_40319_new_n5126_; 
wire _abc_40319_new_n5127_; 
wire _abc_40319_new_n5128_; 
wire _abc_40319_new_n5129_; 
wire _abc_40319_new_n5130_; 
wire _abc_40319_new_n5131_; 
wire _abc_40319_new_n5132_; 
wire _abc_40319_new_n5133_; 
wire _abc_40319_new_n5134_; 
wire _abc_40319_new_n5135_; 
wire _abc_40319_new_n5136_; 
wire _abc_40319_new_n5137_; 
wire _abc_40319_new_n5138_; 
wire _abc_40319_new_n5139_; 
wire _abc_40319_new_n5140_; 
wire _abc_40319_new_n5141_; 
wire _abc_40319_new_n5142_; 
wire _abc_40319_new_n5143_; 
wire _abc_40319_new_n5144_; 
wire _abc_40319_new_n5145_; 
wire _abc_40319_new_n5146_; 
wire _abc_40319_new_n5147_; 
wire _abc_40319_new_n5148_; 
wire _abc_40319_new_n5149_; 
wire _abc_40319_new_n5150_; 
wire _abc_40319_new_n5151_; 
wire _abc_40319_new_n5152_; 
wire _abc_40319_new_n5153_; 
wire _abc_40319_new_n5154_; 
wire _abc_40319_new_n5155_; 
wire _abc_40319_new_n5156_; 
wire _abc_40319_new_n5157_; 
wire _abc_40319_new_n5158_; 
wire _abc_40319_new_n5160_; 
wire _abc_40319_new_n5161_; 
wire _abc_40319_new_n5162_; 
wire _abc_40319_new_n5163_; 
wire _abc_40319_new_n5164_; 
wire _abc_40319_new_n5165_; 
wire _abc_40319_new_n5166_; 
wire _abc_40319_new_n5167_; 
wire _abc_40319_new_n5168_; 
wire _abc_40319_new_n5169_; 
wire _abc_40319_new_n5170_; 
wire _abc_40319_new_n5171_; 
wire _abc_40319_new_n5172_; 
wire _abc_40319_new_n5173_; 
wire _abc_40319_new_n5174_; 
wire _abc_40319_new_n5175_; 
wire _abc_40319_new_n5176_; 
wire _abc_40319_new_n5177_; 
wire _abc_40319_new_n5178_; 
wire _abc_40319_new_n5179_; 
wire _abc_40319_new_n5180_; 
wire _abc_40319_new_n5181_; 
wire _abc_40319_new_n5182_; 
wire _abc_40319_new_n5183_; 
wire _abc_40319_new_n5184_; 
wire _abc_40319_new_n5185_; 
wire _abc_40319_new_n5186_; 
wire _abc_40319_new_n5187_; 
wire _abc_40319_new_n5188_; 
wire _abc_40319_new_n5190_; 
wire _abc_40319_new_n5191_; 
wire _abc_40319_new_n5192_; 
wire _abc_40319_new_n5193_; 
wire _abc_40319_new_n5194_; 
wire _abc_40319_new_n5195_; 
wire _abc_40319_new_n5196_; 
wire _abc_40319_new_n5197_; 
wire _abc_40319_new_n5198_; 
wire _abc_40319_new_n5199_; 
wire _abc_40319_new_n5200_; 
wire _abc_40319_new_n5201_; 
wire _abc_40319_new_n5202_; 
wire _abc_40319_new_n5203_; 
wire _abc_40319_new_n5204_; 
wire _abc_40319_new_n5205_; 
wire _abc_40319_new_n5206_; 
wire _abc_40319_new_n5207_; 
wire _abc_40319_new_n5208_; 
wire _abc_40319_new_n5209_; 
wire _abc_40319_new_n5210_; 
wire _abc_40319_new_n5211_; 
wire _abc_40319_new_n5212_; 
wire _abc_40319_new_n5213_; 
wire _abc_40319_new_n5214_; 
wire _abc_40319_new_n5215_; 
wire _abc_40319_new_n5216_; 
wire _abc_40319_new_n5217_; 
wire _abc_40319_new_n5218_; 
wire _abc_40319_new_n5219_; 
wire _abc_40319_new_n5220_; 
wire _abc_40319_new_n5222_; 
wire _abc_40319_new_n5223_; 
wire _abc_40319_new_n5224_; 
wire _abc_40319_new_n5225_; 
wire _abc_40319_new_n5226_; 
wire _abc_40319_new_n5227_; 
wire _abc_40319_new_n5228_; 
wire _abc_40319_new_n5229_; 
wire _abc_40319_new_n5230_; 
wire _abc_40319_new_n5231_; 
wire _abc_40319_new_n5232_; 
wire _abc_40319_new_n5233_; 
wire _abc_40319_new_n5234_; 
wire _abc_40319_new_n5235_; 
wire _abc_40319_new_n5236_; 
wire _abc_40319_new_n5237_; 
wire _abc_40319_new_n5238_; 
wire _abc_40319_new_n5239_; 
wire _abc_40319_new_n523_; 
wire _abc_40319_new_n5240_; 
wire _abc_40319_new_n5241_; 
wire _abc_40319_new_n5242_; 
wire _abc_40319_new_n5243_; 
wire _abc_40319_new_n5244_; 
wire _abc_40319_new_n5245_; 
wire _abc_40319_new_n5246_; 
wire _abc_40319_new_n5247_; 
wire _abc_40319_new_n5248_; 
wire _abc_40319_new_n5249_; 
wire _abc_40319_new_n524_; 
wire _abc_40319_new_n5250_; 
wire _abc_40319_new_n5251_; 
wire _abc_40319_new_n5253_; 
wire _abc_40319_new_n5254_; 
wire _abc_40319_new_n5255_; 
wire _abc_40319_new_n5256_; 
wire _abc_40319_new_n5257_; 
wire _abc_40319_new_n5258_; 
wire _abc_40319_new_n5259_; 
wire _abc_40319_new_n525_; 
wire _abc_40319_new_n5260_; 
wire _abc_40319_new_n5261_; 
wire _abc_40319_new_n5262_; 
wire _abc_40319_new_n5263_; 
wire _abc_40319_new_n5264_; 
wire _abc_40319_new_n5265_; 
wire _abc_40319_new_n5266_; 
wire _abc_40319_new_n5267_; 
wire _abc_40319_new_n5268_; 
wire _abc_40319_new_n5269_; 
wire _abc_40319_new_n526_; 
wire _abc_40319_new_n5270_; 
wire _abc_40319_new_n5271_; 
wire _abc_40319_new_n5272_; 
wire _abc_40319_new_n5273_; 
wire _abc_40319_new_n5274_; 
wire _abc_40319_new_n5275_; 
wire _abc_40319_new_n5276_; 
wire _abc_40319_new_n5277_; 
wire _abc_40319_new_n5278_; 
wire _abc_40319_new_n5279_; 
wire _abc_40319_new_n527_; 
wire _abc_40319_new_n5280_; 
wire _abc_40319_new_n5281_; 
wire _abc_40319_new_n5282_; 
wire _abc_40319_new_n5283_; 
wire _abc_40319_new_n5284_; 
wire _abc_40319_new_n5285_; 
wire _abc_40319_new_n5286_; 
wire _abc_40319_new_n5287_; 
wire _abc_40319_new_n5288_; 
wire _abc_40319_new_n528_; 
wire _abc_40319_new_n5290_; 
wire _abc_40319_new_n5291_; 
wire _abc_40319_new_n5292_; 
wire _abc_40319_new_n5293_; 
wire _abc_40319_new_n5294_; 
wire _abc_40319_new_n5295_; 
wire _abc_40319_new_n5296_; 
wire _abc_40319_new_n5297_; 
wire _abc_40319_new_n5298_; 
wire _abc_40319_new_n5299_; 
wire _abc_40319_new_n529_; 
wire _abc_40319_new_n5300_; 
wire _abc_40319_new_n5301_; 
wire _abc_40319_new_n5302_; 
wire _abc_40319_new_n5303_; 
wire _abc_40319_new_n5304_; 
wire _abc_40319_new_n5305_; 
wire _abc_40319_new_n5306_; 
wire _abc_40319_new_n5307_; 
wire _abc_40319_new_n5308_; 
wire _abc_40319_new_n5309_; 
wire _abc_40319_new_n530_; 
wire _abc_40319_new_n5310_; 
wire _abc_40319_new_n5311_; 
wire _abc_40319_new_n5312_; 
wire _abc_40319_new_n5313_; 
wire _abc_40319_new_n5314_; 
wire _abc_40319_new_n5315_; 
wire _abc_40319_new_n5316_; 
wire _abc_40319_new_n5317_; 
wire _abc_40319_new_n5318_; 
wire _abc_40319_new_n5319_; 
wire _abc_40319_new_n531_; 
wire _abc_40319_new_n5320_; 
wire _abc_40319_new_n5321_; 
wire _abc_40319_new_n5322_; 
wire _abc_40319_new_n5323_; 
wire _abc_40319_new_n5325_; 
wire _abc_40319_new_n5326_; 
wire _abc_40319_new_n5327_; 
wire _abc_40319_new_n5328_; 
wire _abc_40319_new_n5329_; 
wire _abc_40319_new_n532_; 
wire _abc_40319_new_n5330_; 
wire _abc_40319_new_n5331_; 
wire _abc_40319_new_n5332_; 
wire _abc_40319_new_n5333_; 
wire _abc_40319_new_n5334_; 
wire _abc_40319_new_n5335_; 
wire _abc_40319_new_n5336_; 
wire _abc_40319_new_n5337_; 
wire _abc_40319_new_n5338_; 
wire _abc_40319_new_n5339_; 
wire _abc_40319_new_n533_; 
wire _abc_40319_new_n5340_; 
wire _abc_40319_new_n5341_; 
wire _abc_40319_new_n5342_; 
wire _abc_40319_new_n5343_; 
wire _abc_40319_new_n5344_; 
wire _abc_40319_new_n5345_; 
wire _abc_40319_new_n5346_; 
wire _abc_40319_new_n5347_; 
wire _abc_40319_new_n5348_; 
wire _abc_40319_new_n5349_; 
wire _abc_40319_new_n534_; 
wire _abc_40319_new_n5350_; 
wire _abc_40319_new_n5351_; 
wire _abc_40319_new_n5352_; 
wire _abc_40319_new_n5353_; 
wire _abc_40319_new_n5354_; 
wire _abc_40319_new_n5356_; 
wire _abc_40319_new_n5357_; 
wire _abc_40319_new_n5358_; 
wire _abc_40319_new_n5359_; 
wire _abc_40319_new_n535_; 
wire _abc_40319_new_n5360_; 
wire _abc_40319_new_n5361_; 
wire _abc_40319_new_n5362_; 
wire _abc_40319_new_n5363_; 
wire _abc_40319_new_n5364_; 
wire _abc_40319_new_n5365_; 
wire _abc_40319_new_n5366_; 
wire _abc_40319_new_n5367_; 
wire _abc_40319_new_n5368_; 
wire _abc_40319_new_n5369_; 
wire _abc_40319_new_n536_; 
wire _abc_40319_new_n5370_; 
wire _abc_40319_new_n5371_; 
wire _abc_40319_new_n5372_; 
wire _abc_40319_new_n5373_; 
wire _abc_40319_new_n5374_; 
wire _abc_40319_new_n5375_; 
wire _abc_40319_new_n5376_; 
wire _abc_40319_new_n5377_; 
wire _abc_40319_new_n5378_; 
wire _abc_40319_new_n5379_; 
wire _abc_40319_new_n537_; 
wire _abc_40319_new_n5380_; 
wire _abc_40319_new_n5381_; 
wire _abc_40319_new_n5382_; 
wire _abc_40319_new_n5383_; 
wire _abc_40319_new_n5384_; 
wire _abc_40319_new_n5385_; 
wire _abc_40319_new_n5387_; 
wire _abc_40319_new_n5388_; 
wire _abc_40319_new_n5389_; 
wire _abc_40319_new_n538_; 
wire _abc_40319_new_n5390_; 
wire _abc_40319_new_n5391_; 
wire _abc_40319_new_n5392_; 
wire _abc_40319_new_n5393_; 
wire _abc_40319_new_n5394_; 
wire _abc_40319_new_n5395_; 
wire _abc_40319_new_n5396_; 
wire _abc_40319_new_n5397_; 
wire _abc_40319_new_n5398_; 
wire _abc_40319_new_n5399_; 
wire _abc_40319_new_n539_; 
wire _abc_40319_new_n5400_; 
wire _abc_40319_new_n5401_; 
wire _abc_40319_new_n5402_; 
wire _abc_40319_new_n5403_; 
wire _abc_40319_new_n5404_; 
wire _abc_40319_new_n5405_; 
wire _abc_40319_new_n5406_; 
wire _abc_40319_new_n5407_; 
wire _abc_40319_new_n5408_; 
wire _abc_40319_new_n5409_; 
wire _abc_40319_new_n540_; 
wire _abc_40319_new_n5410_; 
wire _abc_40319_new_n5411_; 
wire _abc_40319_new_n5412_; 
wire _abc_40319_new_n5413_; 
wire _abc_40319_new_n5414_; 
wire _abc_40319_new_n5415_; 
wire _abc_40319_new_n5416_; 
wire _abc_40319_new_n5418_; 
wire _abc_40319_new_n5419_; 
wire _abc_40319_new_n541_; 
wire _abc_40319_new_n5420_; 
wire _abc_40319_new_n5421_; 
wire _abc_40319_new_n5422_; 
wire _abc_40319_new_n5423_; 
wire _abc_40319_new_n5424_; 
wire _abc_40319_new_n5425_; 
wire _abc_40319_new_n5426_; 
wire _abc_40319_new_n5427_; 
wire _abc_40319_new_n5428_; 
wire _abc_40319_new_n5429_; 
wire _abc_40319_new_n542_; 
wire _abc_40319_new_n5430_; 
wire _abc_40319_new_n5431_; 
wire _abc_40319_new_n5432_; 
wire _abc_40319_new_n5433_; 
wire _abc_40319_new_n5434_; 
wire _abc_40319_new_n5435_; 
wire _abc_40319_new_n5436_; 
wire _abc_40319_new_n5437_; 
wire _abc_40319_new_n5438_; 
wire _abc_40319_new_n5439_; 
wire _abc_40319_new_n543_; 
wire _abc_40319_new_n5440_; 
wire _abc_40319_new_n5441_; 
wire _abc_40319_new_n5442_; 
wire _abc_40319_new_n5443_; 
wire _abc_40319_new_n5444_; 
wire _abc_40319_new_n5445_; 
wire _abc_40319_new_n5446_; 
wire _abc_40319_new_n5448_; 
wire _abc_40319_new_n5449_; 
wire _abc_40319_new_n544_; 
wire _abc_40319_new_n5450_; 
wire _abc_40319_new_n5451_; 
wire _abc_40319_new_n5452_; 
wire _abc_40319_new_n5453_; 
wire _abc_40319_new_n5454_; 
wire _abc_40319_new_n5455_; 
wire _abc_40319_new_n5456_; 
wire _abc_40319_new_n5457_; 
wire _abc_40319_new_n5458_; 
wire _abc_40319_new_n5459_; 
wire _abc_40319_new_n545_; 
wire _abc_40319_new_n5460_; 
wire _abc_40319_new_n5461_; 
wire _abc_40319_new_n5463_; 
wire _abc_40319_new_n5464_; 
wire _abc_40319_new_n5465_; 
wire _abc_40319_new_n5466_; 
wire _abc_40319_new_n5468_; 
wire _abc_40319_new_n5469_; 
wire _abc_40319_new_n546_; 
wire _abc_40319_new_n5470_; 
wire _abc_40319_new_n547_; 
wire _abc_40319_new_n548_; 
wire _abc_40319_new_n549_; 
wire _abc_40319_new_n5501_; 
wire _abc_40319_new_n5502_; 
wire _abc_40319_new_n5503_; 
wire _abc_40319_new_n5504_; 
wire _abc_40319_new_n5505_; 
wire _abc_40319_new_n5506_; 
wire _abc_40319_new_n5508_; 
wire _abc_40319_new_n5509_; 
wire _abc_40319_new_n550_; 
wire _abc_40319_new_n5510_; 
wire _abc_40319_new_n5511_; 
wire _abc_40319_new_n5512_; 
wire _abc_40319_new_n5514_; 
wire _abc_40319_new_n5515_; 
wire _abc_40319_new_n5516_; 
wire _abc_40319_new_n5517_; 
wire _abc_40319_new_n5518_; 
wire _abc_40319_new_n551_; 
wire _abc_40319_new_n5520_; 
wire _abc_40319_new_n5521_; 
wire _abc_40319_new_n5522_; 
wire _abc_40319_new_n5523_; 
wire _abc_40319_new_n5524_; 
wire _abc_40319_new_n5526_; 
wire _abc_40319_new_n5527_; 
wire _abc_40319_new_n5528_; 
wire _abc_40319_new_n5529_; 
wire _abc_40319_new_n552_; 
wire _abc_40319_new_n5530_; 
wire _abc_40319_new_n5532_; 
wire _abc_40319_new_n5533_; 
wire _abc_40319_new_n5534_; 
wire _abc_40319_new_n5535_; 
wire _abc_40319_new_n5536_; 
wire _abc_40319_new_n5538_; 
wire _abc_40319_new_n5539_; 
wire _abc_40319_new_n553_; 
wire _abc_40319_new_n5540_; 
wire _abc_40319_new_n5541_; 
wire _abc_40319_new_n5542_; 
wire _abc_40319_new_n5544_; 
wire _abc_40319_new_n5545_; 
wire _abc_40319_new_n5547_; 
wire _abc_40319_new_n5548_; 
wire _abc_40319_new_n5549_; 
wire _abc_40319_new_n554_; 
wire _abc_40319_new_n5550_; 
wire _abc_40319_new_n5551_; 
wire _abc_40319_new_n5552_; 
wire _abc_40319_new_n5554_; 
wire _abc_40319_new_n5555_; 
wire _abc_40319_new_n5556_; 
wire _abc_40319_new_n5557_; 
wire _abc_40319_new_n5558_; 
wire _abc_40319_new_n555_; 
wire _abc_40319_new_n5560_; 
wire _abc_40319_new_n5561_; 
wire _abc_40319_new_n5562_; 
wire _abc_40319_new_n5563_; 
wire _abc_40319_new_n5564_; 
wire _abc_40319_new_n5566_; 
wire _abc_40319_new_n5567_; 
wire _abc_40319_new_n5568_; 
wire _abc_40319_new_n5569_; 
wire _abc_40319_new_n556_; 
wire _abc_40319_new_n5570_; 
wire _abc_40319_new_n5572_; 
wire _abc_40319_new_n5573_; 
wire _abc_40319_new_n5574_; 
wire _abc_40319_new_n5575_; 
wire _abc_40319_new_n5576_; 
wire _abc_40319_new_n5578_; 
wire _abc_40319_new_n5579_; 
wire _abc_40319_new_n557_; 
wire _abc_40319_new_n5580_; 
wire _abc_40319_new_n5581_; 
wire _abc_40319_new_n5582_; 
wire _abc_40319_new_n5584_; 
wire _abc_40319_new_n5585_; 
wire _abc_40319_new_n5586_; 
wire _abc_40319_new_n5587_; 
wire _abc_40319_new_n5588_; 
wire _abc_40319_new_n5589_; 
wire _abc_40319_new_n558_; 
wire _abc_40319_new_n5591_; 
wire _abc_40319_new_n5592_; 
wire _abc_40319_new_n5593_; 
wire _abc_40319_new_n5594_; 
wire _abc_40319_new_n5595_; 
wire _abc_40319_new_n5597_; 
wire _abc_40319_new_n5598_; 
wire _abc_40319_new_n5599_; 
wire _abc_40319_new_n559_; 
wire _abc_40319_new_n5600_; 
wire _abc_40319_new_n5601_; 
wire _abc_40319_new_n5603_; 
wire _abc_40319_new_n5604_; 
wire _abc_40319_new_n5605_; 
wire _abc_40319_new_n5606_; 
wire _abc_40319_new_n5607_; 
wire _abc_40319_new_n5608_; 
wire _abc_40319_new_n560_; 
wire _abc_40319_new_n5610_; 
wire _abc_40319_new_n5611_; 
wire _abc_40319_new_n5612_; 
wire _abc_40319_new_n5613_; 
wire _abc_40319_new_n5614_; 
wire _abc_40319_new_n5615_; 
wire _abc_40319_new_n5617_; 
wire _abc_40319_new_n5618_; 
wire _abc_40319_new_n5619_; 
wire _abc_40319_new_n561_; 
wire _abc_40319_new_n5620_; 
wire _abc_40319_new_n5621_; 
wire _abc_40319_new_n5622_; 
wire _abc_40319_new_n5624_; 
wire _abc_40319_new_n5625_; 
wire _abc_40319_new_n5626_; 
wire _abc_40319_new_n5627_; 
wire _abc_40319_new_n5628_; 
wire _abc_40319_new_n5629_; 
wire _abc_40319_new_n562_; 
wire _abc_40319_new_n5631_; 
wire _abc_40319_new_n5632_; 
wire _abc_40319_new_n5633_; 
wire _abc_40319_new_n5634_; 
wire _abc_40319_new_n5635_; 
wire _abc_40319_new_n5637_; 
wire _abc_40319_new_n5638_; 
wire _abc_40319_new_n5639_; 
wire _abc_40319_new_n563_; 
wire _abc_40319_new_n5640_; 
wire _abc_40319_new_n5641_; 
wire _abc_40319_new_n5643_; 
wire _abc_40319_new_n5644_; 
wire _abc_40319_new_n5645_; 
wire _abc_40319_new_n5646_; 
wire _abc_40319_new_n5647_; 
wire _abc_40319_new_n5649_; 
wire _abc_40319_new_n564_; 
wire _abc_40319_new_n5650_; 
wire _abc_40319_new_n5651_; 
wire _abc_40319_new_n5652_; 
wire _abc_40319_new_n5653_; 
wire _abc_40319_new_n5655_; 
wire _abc_40319_new_n5656_; 
wire _abc_40319_new_n5657_; 
wire _abc_40319_new_n5658_; 
wire _abc_40319_new_n5659_; 
wire _abc_40319_new_n565_; 
wire _abc_40319_new_n5661_; 
wire _abc_40319_new_n5662_; 
wire _abc_40319_new_n5663_; 
wire _abc_40319_new_n5664_; 
wire _abc_40319_new_n5665_; 
wire _abc_40319_new_n5667_; 
wire _abc_40319_new_n5668_; 
wire _abc_40319_new_n5669_; 
wire _abc_40319_new_n566_; 
wire _abc_40319_new_n5670_; 
wire _abc_40319_new_n5671_; 
wire _abc_40319_new_n5673_; 
wire _abc_40319_new_n5674_; 
wire _abc_40319_new_n5675_; 
wire _abc_40319_new_n5676_; 
wire _abc_40319_new_n5677_; 
wire _abc_40319_new_n5678_; 
wire _abc_40319_new_n5679_; 
wire _abc_40319_new_n567_; 
wire _abc_40319_new_n5681_; 
wire _abc_40319_new_n5682_; 
wire _abc_40319_new_n5683_; 
wire _abc_40319_new_n5685_; 
wire _abc_40319_new_n5686_; 
wire _abc_40319_new_n5687_; 
wire _abc_40319_new_n5689_; 
wire _abc_40319_new_n568_; 
wire _abc_40319_new_n5690_; 
wire _abc_40319_new_n5691_; 
wire _abc_40319_new_n5692_; 
wire _abc_40319_new_n5693_; 
wire _abc_40319_new_n5694_; 
wire _abc_40319_new_n5695_; 
wire _abc_40319_new_n5696_; 
wire _abc_40319_new_n5697_; 
wire _abc_40319_new_n5698_; 
wire _abc_40319_new_n5699_; 
wire _abc_40319_new_n569_; 
wire _abc_40319_new_n5700_; 
wire _abc_40319_new_n5701_; 
wire _abc_40319_new_n5702_; 
wire _abc_40319_new_n5703_; 
wire _abc_40319_new_n5704_; 
wire _abc_40319_new_n5705_; 
wire _abc_40319_new_n5706_; 
wire _abc_40319_new_n5707_; 
wire _abc_40319_new_n5708_; 
wire _abc_40319_new_n5709_; 
wire _abc_40319_new_n570_; 
wire _abc_40319_new_n5710_; 
wire _abc_40319_new_n5711_; 
wire _abc_40319_new_n5712_; 
wire _abc_40319_new_n5713_; 
wire _abc_40319_new_n5714_; 
wire _abc_40319_new_n5715_; 
wire _abc_40319_new_n5716_; 
wire _abc_40319_new_n5717_; 
wire _abc_40319_new_n5718_; 
wire _abc_40319_new_n5719_; 
wire _abc_40319_new_n571_; 
wire _abc_40319_new_n5720_; 
wire _abc_40319_new_n5721_; 
wire _abc_40319_new_n5722_; 
wire _abc_40319_new_n5723_; 
wire _abc_40319_new_n5724_; 
wire _abc_40319_new_n5725_; 
wire _abc_40319_new_n5726_; 
wire _abc_40319_new_n5727_; 
wire _abc_40319_new_n5728_; 
wire _abc_40319_new_n572_; 
wire _abc_40319_new_n5730_; 
wire _abc_40319_new_n5731_; 
wire _abc_40319_new_n5732_; 
wire _abc_40319_new_n5733_; 
wire _abc_40319_new_n5734_; 
wire _abc_40319_new_n5736_; 
wire _abc_40319_new_n5737_; 
wire _abc_40319_new_n5738_; 
wire _abc_40319_new_n573_; 
wire _abc_40319_new_n5740_; 
wire _abc_40319_new_n5741_; 
wire _abc_40319_new_n5742_; 
wire _abc_40319_new_n5743_; 
wire _abc_40319_new_n5744_; 
wire _abc_40319_new_n5745_; 
wire _abc_40319_new_n5746_; 
wire _abc_40319_new_n5747_; 
wire _abc_40319_new_n5748_; 
wire _abc_40319_new_n5749_; 
wire _abc_40319_new_n574_; 
wire _abc_40319_new_n5750_; 
wire _abc_40319_new_n5751_; 
wire _abc_40319_new_n5752_; 
wire _abc_40319_new_n5753_; 
wire _abc_40319_new_n5754_; 
wire _abc_40319_new_n5755_; 
wire _abc_40319_new_n5757_; 
wire _abc_40319_new_n5758_; 
wire _abc_40319_new_n5759_; 
wire _abc_40319_new_n575_; 
wire _abc_40319_new_n5760_; 
wire _abc_40319_new_n5761_; 
wire _abc_40319_new_n5762_; 
wire _abc_40319_new_n5763_; 
wire _abc_40319_new_n5765_; 
wire _abc_40319_new_n5766_; 
wire _abc_40319_new_n5767_; 
wire _abc_40319_new_n5768_; 
wire _abc_40319_new_n5769_; 
wire _abc_40319_new_n576_; 
wire _abc_40319_new_n5770_; 
wire _abc_40319_new_n5771_; 
wire _abc_40319_new_n5773_; 
wire _abc_40319_new_n5774_; 
wire _abc_40319_new_n5775_; 
wire _abc_40319_new_n5776_; 
wire _abc_40319_new_n5777_; 
wire _abc_40319_new_n5778_; 
wire _abc_40319_new_n577_; 
wire _abc_40319_new_n5780_; 
wire _abc_40319_new_n5781_; 
wire _abc_40319_new_n5782_; 
wire _abc_40319_new_n5783_; 
wire _abc_40319_new_n5784_; 
wire _abc_40319_new_n5785_; 
wire _abc_40319_new_n5786_; 
wire _abc_40319_new_n5787_; 
wire _abc_40319_new_n5789_; 
wire _abc_40319_new_n578_; 
wire _abc_40319_new_n5790_; 
wire _abc_40319_new_n5791_; 
wire _abc_40319_new_n5792_; 
wire _abc_40319_new_n5793_; 
wire _abc_40319_new_n5794_; 
wire _abc_40319_new_n5795_; 
wire _abc_40319_new_n5796_; 
wire _abc_40319_new_n5798_; 
wire _abc_40319_new_n5799_; 
wire _abc_40319_new_n579_; 
wire _abc_40319_new_n5800_; 
wire _abc_40319_new_n5801_; 
wire _abc_40319_new_n5802_; 
wire _abc_40319_new_n5803_; 
wire _abc_40319_new_n5804_; 
wire _abc_40319_new_n5805_; 
wire _abc_40319_new_n5807_; 
wire _abc_40319_new_n5808_; 
wire _abc_40319_new_n5809_; 
wire _abc_40319_new_n580_; 
wire _abc_40319_new_n5810_; 
wire _abc_40319_new_n5811_; 
wire _abc_40319_new_n5812_; 
wire _abc_40319_new_n5813_; 
wire _abc_40319_new_n5814_; 
wire _abc_40319_new_n5816_; 
wire _abc_40319_new_n5817_; 
wire _abc_40319_new_n5818_; 
wire _abc_40319_new_n5819_; 
wire _abc_40319_new_n581_; 
wire _abc_40319_new_n5820_; 
wire _abc_40319_new_n5821_; 
wire _abc_40319_new_n5822_; 
wire _abc_40319_new_n5823_; 
wire _abc_40319_new_n5825_; 
wire _abc_40319_new_n5826_; 
wire _abc_40319_new_n5827_; 
wire _abc_40319_new_n5828_; 
wire _abc_40319_new_n5829_; 
wire _abc_40319_new_n582_; 
wire _abc_40319_new_n5830_; 
wire _abc_40319_new_n5831_; 
wire _abc_40319_new_n5832_; 
wire _abc_40319_new_n5834_; 
wire _abc_40319_new_n5835_; 
wire _abc_40319_new_n5836_; 
wire _abc_40319_new_n5837_; 
wire _abc_40319_new_n5838_; 
wire _abc_40319_new_n5839_; 
wire _abc_40319_new_n583_; 
wire _abc_40319_new_n5840_; 
wire _abc_40319_new_n5841_; 
wire _abc_40319_new_n5843_; 
wire _abc_40319_new_n5844_; 
wire _abc_40319_new_n5845_; 
wire _abc_40319_new_n5846_; 
wire _abc_40319_new_n5847_; 
wire _abc_40319_new_n5848_; 
wire _abc_40319_new_n5849_; 
wire _abc_40319_new_n584_; 
wire _abc_40319_new_n5850_; 
wire _abc_40319_new_n5851_; 
wire _abc_40319_new_n5853_; 
wire _abc_40319_new_n5854_; 
wire _abc_40319_new_n5855_; 
wire _abc_40319_new_n5856_; 
wire _abc_40319_new_n5857_; 
wire _abc_40319_new_n5858_; 
wire _abc_40319_new_n5859_; 
wire _abc_40319_new_n585_; 
wire _abc_40319_new_n5860_; 
wire _abc_40319_new_n5862_; 
wire _abc_40319_new_n5863_; 
wire _abc_40319_new_n5864_; 
wire _abc_40319_new_n5865_; 
wire _abc_40319_new_n5866_; 
wire _abc_40319_new_n5867_; 
wire _abc_40319_new_n5868_; 
wire _abc_40319_new_n5869_; 
wire _abc_40319_new_n586_; 
wire _abc_40319_new_n5870_; 
wire _abc_40319_new_n5872_; 
wire _abc_40319_new_n5873_; 
wire _abc_40319_new_n5874_; 
wire _abc_40319_new_n5875_; 
wire _abc_40319_new_n5876_; 
wire _abc_40319_new_n5877_; 
wire _abc_40319_new_n5878_; 
wire _abc_40319_new_n5879_; 
wire _abc_40319_new_n587_; 
wire _abc_40319_new_n5880_; 
wire _abc_40319_new_n5882_; 
wire _abc_40319_new_n5883_; 
wire _abc_40319_new_n5884_; 
wire _abc_40319_new_n5885_; 
wire _abc_40319_new_n5886_; 
wire _abc_40319_new_n5887_; 
wire _abc_40319_new_n5888_; 
wire _abc_40319_new_n5889_; 
wire _abc_40319_new_n588_; 
wire _abc_40319_new_n5891_; 
wire _abc_40319_new_n5892_; 
wire _abc_40319_new_n5893_; 
wire _abc_40319_new_n5894_; 
wire _abc_40319_new_n5895_; 
wire _abc_40319_new_n5896_; 
wire _abc_40319_new_n5897_; 
wire _abc_40319_new_n5898_; 
wire _abc_40319_new_n5899_; 
wire _abc_40319_new_n589_; 
wire _abc_40319_new_n5901_; 
wire _abc_40319_new_n5902_; 
wire _abc_40319_new_n5903_; 
wire _abc_40319_new_n5904_; 
wire _abc_40319_new_n5905_; 
wire _abc_40319_new_n5906_; 
wire _abc_40319_new_n5907_; 
wire _abc_40319_new_n5908_; 
wire _abc_40319_new_n5909_; 
wire _abc_40319_new_n590_; 
wire _abc_40319_new_n5911_; 
wire _abc_40319_new_n5912_; 
wire _abc_40319_new_n5913_; 
wire _abc_40319_new_n5914_; 
wire _abc_40319_new_n5915_; 
wire _abc_40319_new_n5916_; 
wire _abc_40319_new_n5917_; 
wire _abc_40319_new_n5918_; 
wire _abc_40319_new_n5919_; 
wire _abc_40319_new_n591_; 
wire _abc_40319_new_n5921_; 
wire _abc_40319_new_n5922_; 
wire _abc_40319_new_n5923_; 
wire _abc_40319_new_n5924_; 
wire _abc_40319_new_n5925_; 
wire _abc_40319_new_n5926_; 
wire _abc_40319_new_n5927_; 
wire _abc_40319_new_n5928_; 
wire _abc_40319_new_n5929_; 
wire _abc_40319_new_n592_; 
wire _abc_40319_new_n5930_; 
wire _abc_40319_new_n5932_; 
wire _abc_40319_new_n5933_; 
wire _abc_40319_new_n5934_; 
wire _abc_40319_new_n5935_; 
wire _abc_40319_new_n5936_; 
wire _abc_40319_new_n5937_; 
wire _abc_40319_new_n5938_; 
wire _abc_40319_new_n5939_; 
wire _abc_40319_new_n593_; 
wire _abc_40319_new_n5940_; 
wire _abc_40319_new_n5941_; 
wire _abc_40319_new_n5943_; 
wire _abc_40319_new_n5944_; 
wire _abc_40319_new_n5945_; 
wire _abc_40319_new_n5946_; 
wire _abc_40319_new_n5947_; 
wire _abc_40319_new_n5948_; 
wire _abc_40319_new_n5949_; 
wire _abc_40319_new_n594_; 
wire _abc_40319_new_n5950_; 
wire _abc_40319_new_n5951_; 
wire _abc_40319_new_n5952_; 
wire _abc_40319_new_n5954_; 
wire _abc_40319_new_n5955_; 
wire _abc_40319_new_n5956_; 
wire _abc_40319_new_n5957_; 
wire _abc_40319_new_n5958_; 
wire _abc_40319_new_n5959_; 
wire _abc_40319_new_n595_; 
wire _abc_40319_new_n5960_; 
wire _abc_40319_new_n5961_; 
wire _abc_40319_new_n5962_; 
wire _abc_40319_new_n5963_; 
wire _abc_40319_new_n5965_; 
wire _abc_40319_new_n5966_; 
wire _abc_40319_new_n5967_; 
wire _abc_40319_new_n5968_; 
wire _abc_40319_new_n5969_; 
wire _abc_40319_new_n596_; 
wire _abc_40319_new_n5970_; 
wire _abc_40319_new_n5971_; 
wire _abc_40319_new_n5972_; 
wire _abc_40319_new_n5973_; 
wire _abc_40319_new_n5974_; 
wire _abc_40319_new_n5976_; 
wire _abc_40319_new_n5977_; 
wire _abc_40319_new_n5978_; 
wire _abc_40319_new_n5979_; 
wire _abc_40319_new_n597_; 
wire _abc_40319_new_n5980_; 
wire _abc_40319_new_n5981_; 
wire _abc_40319_new_n5982_; 
wire _abc_40319_new_n5983_; 
wire _abc_40319_new_n5984_; 
wire _abc_40319_new_n5985_; 
wire _abc_40319_new_n5987_; 
wire _abc_40319_new_n5988_; 
wire _abc_40319_new_n5989_; 
wire _abc_40319_new_n598_; 
wire _abc_40319_new_n5990_; 
wire _abc_40319_new_n5991_; 
wire _abc_40319_new_n5992_; 
wire _abc_40319_new_n5993_; 
wire _abc_40319_new_n5994_; 
wire _abc_40319_new_n5995_; 
wire _abc_40319_new_n5996_; 
wire _abc_40319_new_n5998_; 
wire _abc_40319_new_n5999_; 
wire _abc_40319_new_n599_; 
wire _abc_40319_new_n6000_; 
wire _abc_40319_new_n6001_; 
wire _abc_40319_new_n6002_; 
wire _abc_40319_new_n6003_; 
wire _abc_40319_new_n6004_; 
wire _abc_40319_new_n6005_; 
wire _abc_40319_new_n6006_; 
wire _abc_40319_new_n6007_; 
wire _abc_40319_new_n6009_; 
wire _abc_40319_new_n600_; 
wire _abc_40319_new_n6010_; 
wire _abc_40319_new_n6011_; 
wire _abc_40319_new_n6012_; 
wire _abc_40319_new_n6013_; 
wire _abc_40319_new_n6014_; 
wire _abc_40319_new_n6015_; 
wire _abc_40319_new_n6016_; 
wire _abc_40319_new_n6017_; 
wire _abc_40319_new_n6018_; 
wire _abc_40319_new_n601_; 
wire _abc_40319_new_n6020_; 
wire _abc_40319_new_n6021_; 
wire _abc_40319_new_n6022_; 
wire _abc_40319_new_n6023_; 
wire _abc_40319_new_n6024_; 
wire _abc_40319_new_n6025_; 
wire _abc_40319_new_n6026_; 
wire _abc_40319_new_n6027_; 
wire _abc_40319_new_n6028_; 
wire _abc_40319_new_n6029_; 
wire _abc_40319_new_n602_; 
wire _abc_40319_new_n6031_; 
wire _abc_40319_new_n6032_; 
wire _abc_40319_new_n6033_; 
wire _abc_40319_new_n6034_; 
wire _abc_40319_new_n6035_; 
wire _abc_40319_new_n6036_; 
wire _abc_40319_new_n6037_; 
wire _abc_40319_new_n6038_; 
wire _abc_40319_new_n6039_; 
wire _abc_40319_new_n603_; 
wire _abc_40319_new_n6041_; 
wire _abc_40319_new_n6042_; 
wire _abc_40319_new_n6043_; 
wire _abc_40319_new_n6044_; 
wire _abc_40319_new_n6045_; 
wire _abc_40319_new_n6046_; 
wire _abc_40319_new_n6047_; 
wire _abc_40319_new_n6049_; 
wire _abc_40319_new_n604_; 
wire _abc_40319_new_n6050_; 
wire _abc_40319_new_n6051_; 
wire _abc_40319_new_n6052_; 
wire _abc_40319_new_n6053_; 
wire _abc_40319_new_n6054_; 
wire _abc_40319_new_n6055_; 
wire _abc_40319_new_n6057_; 
wire _abc_40319_new_n6058_; 
wire _abc_40319_new_n6059_; 
wire _abc_40319_new_n605_; 
wire _abc_40319_new_n6060_; 
wire _abc_40319_new_n6061_; 
wire _abc_40319_new_n6063_; 
wire _abc_40319_new_n6064_; 
wire _abc_40319_new_n6065_; 
wire _abc_40319_new_n6067_; 
wire _abc_40319_new_n6068_; 
wire _abc_40319_new_n6069_; 
wire _abc_40319_new_n606_; 
wire _abc_40319_new_n6071_; 
wire _abc_40319_new_n6072_; 
wire _abc_40319_new_n6073_; 
wire _abc_40319_new_n6075_; 
wire _abc_40319_new_n6076_; 
wire _abc_40319_new_n6077_; 
wire _abc_40319_new_n6079_; 
wire _abc_40319_new_n607_; 
wire _abc_40319_new_n6080_; 
wire _abc_40319_new_n6081_; 
wire _abc_40319_new_n6083_; 
wire _abc_40319_new_n6084_; 
wire _abc_40319_new_n6085_; 
wire _abc_40319_new_n6087_; 
wire _abc_40319_new_n6088_; 
wire _abc_40319_new_n6089_; 
wire _abc_40319_new_n608_; 
wire _abc_40319_new_n6091_; 
wire _abc_40319_new_n6092_; 
wire _abc_40319_new_n6093_; 
wire _abc_40319_new_n6095_; 
wire _abc_40319_new_n6096_; 
wire _abc_40319_new_n6097_; 
wire _abc_40319_new_n6099_; 
wire _abc_40319_new_n609_; 
wire _abc_40319_new_n6100_; 
wire _abc_40319_new_n6101_; 
wire _abc_40319_new_n6103_; 
wire _abc_40319_new_n6104_; 
wire _abc_40319_new_n6105_; 
wire _abc_40319_new_n6107_; 
wire _abc_40319_new_n6108_; 
wire _abc_40319_new_n6109_; 
wire _abc_40319_new_n610_; 
wire _abc_40319_new_n6111_; 
wire _abc_40319_new_n6112_; 
wire _abc_40319_new_n6113_; 
wire _abc_40319_new_n6115_; 
wire _abc_40319_new_n6116_; 
wire _abc_40319_new_n6117_; 
wire _abc_40319_new_n6119_; 
wire _abc_40319_new_n611_; 
wire _abc_40319_new_n6120_; 
wire _abc_40319_new_n6121_; 
wire _abc_40319_new_n6123_; 
wire _abc_40319_new_n6124_; 
wire _abc_40319_new_n6125_; 
wire _abc_40319_new_n6127_; 
wire _abc_40319_new_n6128_; 
wire _abc_40319_new_n6129_; 
wire _abc_40319_new_n612_; 
wire _abc_40319_new_n6131_; 
wire _abc_40319_new_n6132_; 
wire _abc_40319_new_n6133_; 
wire _abc_40319_new_n6135_; 
wire _abc_40319_new_n6136_; 
wire _abc_40319_new_n6137_; 
wire _abc_40319_new_n6139_; 
wire _abc_40319_new_n613_; 
wire _abc_40319_new_n6140_; 
wire _abc_40319_new_n6141_; 
wire _abc_40319_new_n6143_; 
wire _abc_40319_new_n6144_; 
wire _abc_40319_new_n6145_; 
wire _abc_40319_new_n6147_; 
wire _abc_40319_new_n6148_; 
wire _abc_40319_new_n6149_; 
wire _abc_40319_new_n614_; 
wire _abc_40319_new_n6151_; 
wire _abc_40319_new_n6152_; 
wire _abc_40319_new_n6153_; 
wire _abc_40319_new_n6155_; 
wire _abc_40319_new_n6156_; 
wire _abc_40319_new_n6157_; 
wire _abc_40319_new_n6159_; 
wire _abc_40319_new_n615_; 
wire _abc_40319_new_n6160_; 
wire _abc_40319_new_n6161_; 
wire _abc_40319_new_n6163_; 
wire _abc_40319_new_n6164_; 
wire _abc_40319_new_n6165_; 
wire _abc_40319_new_n6167_; 
wire _abc_40319_new_n6168_; 
wire _abc_40319_new_n6169_; 
wire _abc_40319_new_n6171_; 
wire _abc_40319_new_n6172_; 
wire _abc_40319_new_n6173_; 
wire _abc_40319_new_n6175_; 
wire _abc_40319_new_n6176_; 
wire _abc_40319_new_n6177_; 
wire _abc_40319_new_n6179_; 
wire _abc_40319_new_n617_; 
wire _abc_40319_new_n6180_; 
wire _abc_40319_new_n6181_; 
wire _abc_40319_new_n6183_; 
wire _abc_40319_new_n6184_; 
wire _abc_40319_new_n6185_; 
wire _abc_40319_new_n6187_; 
wire _abc_40319_new_n6188_; 
wire _abc_40319_new_n6189_; 
wire _abc_40319_new_n6190_; 
wire _abc_40319_new_n6192_; 
wire _abc_40319_new_n6193_; 
wire _abc_40319_new_n6194_; 
wire _abc_40319_new_n6196_; 
wire _abc_40319_new_n6197_; 
wire _abc_40319_new_n6198_; 
wire _abc_40319_new_n619_; 
wire _abc_40319_new_n6200_; 
wire _abc_40319_new_n6201_; 
wire _abc_40319_new_n6202_; 
wire _abc_40319_new_n6204_; 
wire _abc_40319_new_n6205_; 
wire _abc_40319_new_n6206_; 
wire _abc_40319_new_n6208_; 
wire _abc_40319_new_n6209_; 
wire _abc_40319_new_n620_; 
wire _abc_40319_new_n6210_; 
wire _abc_40319_new_n6212_; 
wire _abc_40319_new_n6213_; 
wire _abc_40319_new_n6214_; 
wire _abc_40319_new_n6216_; 
wire _abc_40319_new_n6217_; 
wire _abc_40319_new_n6218_; 
wire _abc_40319_new_n621_; 
wire _abc_40319_new_n6220_; 
wire _abc_40319_new_n6221_; 
wire _abc_40319_new_n6222_; 
wire _abc_40319_new_n6224_; 
wire _abc_40319_new_n6225_; 
wire _abc_40319_new_n6226_; 
wire _abc_40319_new_n6228_; 
wire _abc_40319_new_n6229_; 
wire _abc_40319_new_n622_; 
wire _abc_40319_new_n6230_; 
wire _abc_40319_new_n6232_; 
wire _abc_40319_new_n6233_; 
wire _abc_40319_new_n6234_; 
wire _abc_40319_new_n6236_; 
wire _abc_40319_new_n6237_; 
wire _abc_40319_new_n6238_; 
wire _abc_40319_new_n623_; 
wire _abc_40319_new_n6240_; 
wire _abc_40319_new_n6241_; 
wire _abc_40319_new_n6242_; 
wire _abc_40319_new_n6244_; 
wire _abc_40319_new_n6245_; 
wire _abc_40319_new_n6246_; 
wire _abc_40319_new_n6248_; 
wire _abc_40319_new_n6249_; 
wire _abc_40319_new_n624_; 
wire _abc_40319_new_n6250_; 
wire _abc_40319_new_n6252_; 
wire _abc_40319_new_n6253_; 
wire _abc_40319_new_n6254_; 
wire _abc_40319_new_n6256_; 
wire _abc_40319_new_n6257_; 
wire _abc_40319_new_n6258_; 
wire _abc_40319_new_n625_; 
wire _abc_40319_new_n6260_; 
wire _abc_40319_new_n6261_; 
wire _abc_40319_new_n6262_; 
wire _abc_40319_new_n6264_; 
wire _abc_40319_new_n6265_; 
wire _abc_40319_new_n6266_; 
wire _abc_40319_new_n6268_; 
wire _abc_40319_new_n6269_; 
wire _abc_40319_new_n626_; 
wire _abc_40319_new_n6270_; 
wire _abc_40319_new_n6272_; 
wire _abc_40319_new_n6273_; 
wire _abc_40319_new_n6274_; 
wire _abc_40319_new_n6276_; 
wire _abc_40319_new_n6277_; 
wire _abc_40319_new_n6278_; 
wire _abc_40319_new_n627_; 
wire _abc_40319_new_n6280_; 
wire _abc_40319_new_n6281_; 
wire _abc_40319_new_n6282_; 
wire _abc_40319_new_n6284_; 
wire _abc_40319_new_n6285_; 
wire _abc_40319_new_n6286_; 
wire _abc_40319_new_n6288_; 
wire _abc_40319_new_n6289_; 
wire _abc_40319_new_n628_; 
wire _abc_40319_new_n6290_; 
wire _abc_40319_new_n6292_; 
wire _abc_40319_new_n6293_; 
wire _abc_40319_new_n6294_; 
wire _abc_40319_new_n6296_; 
wire _abc_40319_new_n6297_; 
wire _abc_40319_new_n6298_; 
wire _abc_40319_new_n629_; 
wire _abc_40319_new_n6300_; 
wire _abc_40319_new_n6301_; 
wire _abc_40319_new_n6302_; 
wire _abc_40319_new_n6304_; 
wire _abc_40319_new_n6305_; 
wire _abc_40319_new_n6306_; 
wire _abc_40319_new_n6308_; 
wire _abc_40319_new_n6309_; 
wire _abc_40319_new_n630_; 
wire _abc_40319_new_n6310_; 
wire _abc_40319_new_n6312_; 
wire _abc_40319_new_n6313_; 
wire _abc_40319_new_n6314_; 
wire _abc_40319_new_n631_; 
wire _abc_40319_new_n632_; 
wire _abc_40319_new_n633_; 
wire _abc_40319_new_n634_; 
wire _abc_40319_new_n635_; 
wire _abc_40319_new_n636_; 
wire _abc_40319_new_n637_; 
wire _abc_40319_new_n638_; 
wire _abc_40319_new_n639_; 
wire _abc_40319_new_n640_; 
wire _abc_40319_new_n641_; 
wire _abc_40319_new_n642_; 
wire _abc_40319_new_n643_; 
wire _abc_40319_new_n644_; 
wire _abc_40319_new_n645_; 
wire _abc_40319_new_n646_; 
wire _abc_40319_new_n647_; 
wire _abc_40319_new_n648_; 
wire _abc_40319_new_n649_; 
wire _abc_40319_new_n650_; 
wire _abc_40319_new_n651_; 
wire _abc_40319_new_n652_; 
wire _abc_40319_new_n653_; 
wire _abc_40319_new_n654_; 
wire _abc_40319_new_n655_; 
wire _abc_40319_new_n656_; 
wire _abc_40319_new_n657_; 
wire _abc_40319_new_n658_; 
wire _abc_40319_new_n659_; 
wire _abc_40319_new_n660_; 
wire _abc_40319_new_n661_; 
wire _abc_40319_new_n663_; 
wire _abc_40319_new_n664_; 
wire _abc_40319_new_n665_; 
wire _abc_40319_new_n666_; 
wire _abc_40319_new_n667_; 
wire _abc_40319_new_n668_; 
wire _abc_40319_new_n669_; 
wire _abc_40319_new_n670_; 
wire _abc_40319_new_n671_; 
wire _abc_40319_new_n672_; 
wire _abc_40319_new_n673_; 
wire _abc_40319_new_n674_; 
wire _abc_40319_new_n675_; 
wire _abc_40319_new_n676_; 
wire _abc_40319_new_n677_; 
wire _abc_40319_new_n678_; 
wire _abc_40319_new_n679_; 
wire _abc_40319_new_n680_; 
wire _abc_40319_new_n681_; 
wire _abc_40319_new_n682_; 
wire _abc_40319_new_n683_; 
wire _abc_40319_new_n684_; 
wire _abc_40319_new_n685_; 
wire _abc_40319_new_n686_; 
wire _abc_40319_new_n687_; 
wire _abc_40319_new_n688_; 
wire _abc_40319_new_n689_; 
wire _abc_40319_new_n690_; 
wire _abc_40319_new_n691_; 
wire _abc_40319_new_n692_; 
wire _abc_40319_new_n693_; 
wire _abc_40319_new_n694_; 
wire _abc_40319_new_n695_; 
wire _abc_40319_new_n696_; 
wire _abc_40319_new_n697_; 
wire _abc_40319_new_n698_; 
wire _abc_40319_new_n699_; 
wire _abc_40319_new_n700_; 
wire _abc_40319_new_n701_; 
wire _abc_40319_new_n702_; 
wire _abc_40319_new_n703_; 
wire _abc_40319_new_n704_; 
wire _abc_40319_new_n705_; 
wire _abc_40319_new_n706_; 
wire _abc_40319_new_n707_; 
wire _abc_40319_new_n708_; 
wire _abc_40319_new_n709_; 
wire _abc_40319_new_n710_; 
wire _abc_40319_new_n711_; 
wire _abc_40319_new_n712_; 
wire _abc_40319_new_n713_; 
wire _abc_40319_new_n714_; 
wire _abc_40319_new_n715_; 
wire _abc_40319_new_n716_; 
wire _abc_40319_new_n717_; 
wire _abc_40319_new_n718_; 
wire _abc_40319_new_n719_; 
wire _abc_40319_new_n720_; 
wire _abc_40319_new_n721_; 
wire _abc_40319_new_n722_; 
wire _abc_40319_new_n723_; 
wire _abc_40319_new_n724_; 
wire _abc_40319_new_n725_; 
wire _abc_40319_new_n726_; 
wire _abc_40319_new_n727_; 
wire _abc_40319_new_n728_; 
wire _abc_40319_new_n729_; 
wire _abc_40319_new_n730_; 
wire _abc_40319_new_n731_; 
wire _abc_40319_new_n732_; 
wire _abc_40319_new_n733_; 
wire _abc_40319_new_n734_; 
wire _abc_40319_new_n735_; 
wire _abc_40319_new_n736_; 
wire _abc_40319_new_n737_; 
wire _abc_40319_new_n738_; 
wire _abc_40319_new_n739_; 
wire _abc_40319_new_n740_; 
wire _abc_40319_new_n741_; 
wire _abc_40319_new_n742_; 
wire _abc_40319_new_n743_; 
wire _abc_40319_new_n744_; 
wire _abc_40319_new_n745_; 
wire _abc_40319_new_n746_; 
wire _abc_40319_new_n747_; 
wire _abc_40319_new_n748_; 
wire _abc_40319_new_n749_; 
wire _abc_40319_new_n750_; 
wire _abc_40319_new_n751_; 
wire _abc_40319_new_n752_; 
wire _abc_40319_new_n753_; 
wire _abc_40319_new_n754_; 
wire _abc_40319_new_n755_; 
wire _abc_40319_new_n756_; 
wire _abc_40319_new_n757_; 
wire _abc_40319_new_n758_; 
wire _abc_40319_new_n759_; 
wire _abc_40319_new_n760_; 
wire _abc_40319_new_n761_; 
wire _abc_40319_new_n762_; 
wire _abc_40319_new_n763_; 
wire _abc_40319_new_n764_; 
wire _abc_40319_new_n765_; 
wire _abc_40319_new_n766_; 
wire _abc_40319_new_n767_; 
wire _abc_40319_new_n768_; 
wire _abc_40319_new_n769_; 
wire _abc_40319_new_n770_; 
wire _abc_40319_new_n771_; 
wire _abc_40319_new_n772_; 
wire _abc_40319_new_n773_; 
wire _abc_40319_new_n774_; 
wire _abc_40319_new_n775_; 
wire _abc_40319_new_n776_; 
wire _abc_40319_new_n777_; 
wire _abc_40319_new_n778_; 
wire _abc_40319_new_n779_; 
wire _abc_40319_new_n780_; 
wire _abc_40319_new_n781_; 
wire _abc_40319_new_n782_; 
wire _abc_40319_new_n783_; 
wire _abc_40319_new_n784_; 
wire _abc_40319_new_n785_; 
wire _abc_40319_new_n786_; 
wire _abc_40319_new_n787_; 
wire _abc_40319_new_n788_; 
wire _abc_40319_new_n789_; 
wire _abc_40319_new_n790_; 
wire _abc_40319_new_n791_; 
wire _abc_40319_new_n792_; 
wire _abc_40319_new_n793_; 
wire _abc_40319_new_n794_; 
wire _abc_40319_new_n795_; 
wire _abc_40319_new_n796_; 
wire _abc_40319_new_n797_; 
wire _abc_40319_new_n798_; 
wire _abc_40319_new_n799_; 
wire _abc_40319_new_n800_; 
wire _abc_40319_new_n801_; 
wire _abc_40319_new_n802_; 
wire _abc_40319_new_n803_; 
wire _abc_40319_new_n804_; 
wire _abc_40319_new_n805_; 
wire _abc_40319_new_n806_; 
wire _abc_40319_new_n807_; 
wire _abc_40319_new_n808_; 
wire _abc_40319_new_n809_; 
wire _abc_40319_new_n810_; 
wire _abc_40319_new_n811_; 
wire _abc_40319_new_n812_; 
wire _abc_40319_new_n813_; 
wire _abc_40319_new_n814_; 
wire _abc_40319_new_n815_; 
wire _abc_40319_new_n816_; 
wire _abc_40319_new_n817_; 
wire _abc_40319_new_n818_; 
wire _abc_40319_new_n819_; 
wire _abc_40319_new_n820_; 
wire _abc_40319_new_n821_; 
wire _abc_40319_new_n822_; 
wire _abc_40319_new_n823_; 
wire _abc_40319_new_n824_; 
wire _abc_40319_new_n825_; 
wire _abc_40319_new_n826_; 
wire _abc_40319_new_n827_; 
wire _abc_40319_new_n828_; 
wire _abc_40319_new_n829_; 
wire _abc_40319_new_n830_; 
wire _abc_40319_new_n831_; 
wire _abc_40319_new_n832_; 
wire _abc_40319_new_n833_; 
wire _abc_40319_new_n834_; 
wire _abc_40319_new_n835_; 
wire _abc_40319_new_n836_; 
wire _abc_40319_new_n837_; 
wire _abc_40319_new_n838_; 
wire _abc_40319_new_n839_; 
wire _abc_40319_new_n840_; 
wire _abc_40319_new_n841_; 
wire _abc_40319_new_n842_; 
wire _abc_40319_new_n843_; 
wire _abc_40319_new_n844_; 
wire _abc_40319_new_n845_; 
wire _abc_40319_new_n846_; 
wire _abc_40319_new_n847_; 
wire _abc_40319_new_n848_; 
wire _abc_40319_new_n849_; 
wire _abc_40319_new_n850_; 
wire _abc_40319_new_n851_; 
wire _abc_40319_new_n852_; 
wire _abc_40319_new_n853_; 
wire _abc_40319_new_n854_; 
wire _abc_40319_new_n855_; 
wire _abc_40319_new_n856_; 
wire _abc_40319_new_n857_; 
wire _abc_40319_new_n858_; 
wire _abc_40319_new_n859_; 
wire _abc_40319_new_n860_; 
wire _abc_40319_new_n861_; 
wire _abc_40319_new_n862_; 
wire _abc_40319_new_n863_; 
wire _abc_40319_new_n864_; 
wire _abc_40319_new_n865_; 
wire _abc_40319_new_n866_; 
wire _abc_40319_new_n867_; 
wire _abc_40319_new_n868_; 
wire _abc_40319_new_n869_; 
wire _abc_40319_new_n870_; 
wire _abc_40319_new_n871_; 
wire _abc_40319_new_n872_; 
wire _abc_40319_new_n873_; 
wire _abc_40319_new_n874_; 
wire _abc_40319_new_n875_; 
wire _abc_40319_new_n876_; 
wire _abc_40319_new_n877_; 
wire _abc_40319_new_n878_; 
wire _abc_40319_new_n879_; 
wire _abc_40319_new_n880_; 
wire _abc_40319_new_n881_; 
wire _abc_40319_new_n882_; 
wire _abc_40319_new_n883_; 
wire _abc_40319_new_n884_; 
wire _abc_40319_new_n885_; 
wire _abc_40319_new_n886_; 
wire _abc_40319_new_n887_; 
wire _abc_40319_new_n888_; 
wire _abc_40319_new_n889_; 
wire _abc_40319_new_n890_; 
wire _abc_40319_new_n891_; 
wire _abc_40319_new_n892_; 
wire _abc_40319_new_n893_; 
wire _abc_40319_new_n894_; 
wire _abc_40319_new_n895_; 
wire _abc_40319_new_n896_; 
wire _abc_40319_new_n897_; 
wire _abc_40319_new_n898_; 
wire _abc_40319_new_n899_; 
wire _abc_40319_new_n900_; 
wire _abc_40319_new_n901_; 
wire _abc_40319_new_n902_; 
wire _abc_40319_new_n903_; 
wire _abc_40319_new_n904_; 
wire _abc_40319_new_n905_; 
wire _abc_40319_new_n906_; 
wire _abc_40319_new_n907_; 
wire _abc_40319_new_n908_; 
wire _abc_40319_new_n909_; 
wire _abc_40319_new_n910_; 
wire _abc_40319_new_n911_; 
wire _abc_40319_new_n912_; 
wire _abc_40319_new_n913_; 
wire _abc_40319_new_n914_; 
wire _abc_40319_new_n915_; 
wire _abc_40319_new_n916_; 
wire _abc_40319_new_n917_; 
wire _abc_40319_new_n918_; 
wire _abc_40319_new_n919_; 
wire _abc_40319_new_n920_; 
wire _abc_40319_new_n921_; 
wire _abc_40319_new_n922_; 
wire _abc_40319_new_n923_; 
wire _abc_40319_new_n924_; 
wire _abc_40319_new_n925_; 
wire _abc_40319_new_n926_; 
wire _abc_40319_new_n927_; 
wire _abc_40319_new_n928_; 
wire _abc_40319_new_n929_; 
wire _abc_40319_new_n930_; 
wire _abc_40319_new_n931_; 
wire _abc_40319_new_n932_; 
wire _abc_40319_new_n933_; 
wire _abc_40319_new_n934_; 
wire _abc_40319_new_n935_; 
wire _abc_40319_new_n936_; 
wire _abc_40319_new_n937_; 
wire _abc_40319_new_n938_; 
wire _abc_40319_new_n939_; 
wire _abc_40319_new_n940_; 
wire _abc_40319_new_n941_; 
wire _abc_40319_new_n942_; 
wire _abc_40319_new_n943_; 
wire _abc_40319_new_n944_; 
wire _abc_40319_new_n945_; 
wire _abc_40319_new_n946_; 
wire _abc_40319_new_n947_; 
wire _abc_40319_new_n948_; 
wire _abc_40319_new_n949_; 
wire _abc_40319_new_n950_; 
wire _abc_40319_new_n951_; 
wire _abc_40319_new_n952_; 
wire _abc_40319_new_n953_; 
wire _abc_40319_new_n954_; 
wire _abc_40319_new_n955_; 
wire _abc_40319_new_n956_; 
wire _abc_40319_new_n957_; 
wire _abc_40319_new_n958_; 
wire _abc_40319_new_n959_; 
wire _abc_40319_new_n960_; 
wire _abc_40319_new_n961_; 
wire _abc_40319_new_n962_; 
wire _abc_40319_new_n963_; 
wire _abc_40319_new_n964_; 
wire _abc_40319_new_n965_; 
wire _abc_40319_new_n966_; 
wire _abc_40319_new_n967_; 
wire _abc_40319_new_n968_; 
wire _abc_40319_new_n969_; 
wire _abc_40319_new_n970_; 
wire _abc_40319_new_n971_; 
wire _abc_40319_new_n972_; 
wire _abc_40319_new_n973_; 
wire _abc_40319_new_n974_; 
wire _abc_40319_new_n975_; 
wire _abc_40319_new_n976_; 
wire _abc_40319_new_n977_; 
wire _abc_40319_new_n978_; 
wire _abc_40319_new_n979_; 
wire _abc_40319_new_n980_; 
wire _abc_40319_new_n981_; 
wire _abc_40319_new_n982_; 
wire _abc_40319_new_n983_; 
wire _abc_40319_new_n984_; 
wire _abc_40319_new_n985_; 
wire _abc_40319_new_n986_; 
wire _abc_40319_new_n987_; 
wire _abc_40319_new_n988_; 
wire _abc_40319_new_n989_; 
wire _abc_40319_new_n990_; 
wire _abc_40319_new_n991_; 
wire _abc_40319_new_n992_; 
wire _abc_40319_new_n993_; 
wire _abc_40319_new_n994_; 
wire _abc_40319_new_n995_; 
wire _abc_40319_new_n996_; 
wire _abc_40319_new_n997_; 
wire _abc_40319_new_n998_; 
wire _abc_40319_new_n999_; 
input clock;
wire n1002; 
wire n1006; 
wire n1010; 
wire n1014; 
wire n1018; 
wire n1022; 
wire n1026; 
wire n1030; 
wire n1034; 
wire n1038; 
wire n1042; 
wire n1046; 
wire n1050; 
wire n1054; 
wire n1058; 
wire n1062; 
wire n1066; 
wire n1070; 
wire n1074; 
wire n1078; 
wire n1082; 
wire n1086; 
wire n1090; 
wire n1094; 
wire n1098; 
wire n1102; 
wire n1106; 
wire n1110; 
wire n1114; 
wire n1118; 
wire n1122; 
wire n1126; 
wire n1130; 
wire n1134; 
wire n1138; 
wire n1142; 
wire n1146; 
wire n1150; 
wire n1154; 
wire n1158; 
wire n1162; 
wire n1166; 
wire n1170; 
wire n1174; 
wire n1178; 
wire n1182; 
wire n1186; 
wire n1191; 
wire n1196; 
wire n1201; 
wire n1206; 
wire n1211; 
wire n1216; 
wire n1221; 
wire n1226; 
wire n1231; 
wire n1236; 
wire n1241; 
wire n1246; 
wire n1251; 
wire n1256; 
wire n1261; 
wire n1266; 
wire n1271; 
wire n1276; 
wire n1281; 
wire n1286; 
wire n1291; 
wire n1296; 
wire n1301; 
wire n1306; 
wire n1311; 
wire n1316; 
wire n1321; 
wire n1326; 
wire n1331; 
wire n1336; 
wire n1341; 
wire n1345; 
wire n178; 
wire n183; 
wire n188; 
wire n193; 
wire n198; 
wire n203; 
wire n208; 
wire n213; 
wire n218; 
wire n223; 
wire n228; 
wire n233; 
wire n238; 
wire n243; 
wire n248; 
wire n253; 
wire n258; 
wire n263; 
wire n268; 
wire n273; 
wire n278; 
wire n283; 
wire n288; 
wire n293; 
wire n298; 
wire n303; 
wire n308; 
wire n313; 
wire n318; 
wire n323; 
wire n328; 
wire n333; 
wire n338; 
wire n343; 
wire n348; 
wire n353; 
wire n358; 
wire n363; 
wire n368; 
wire n373; 
wire n378; 
wire n383; 
wire n388; 
wire n393; 
wire n398; 
wire n403; 
wire n408; 
wire n413; 
wire n418; 
wire n423; 
wire n428; 
wire n433; 
wire n438; 
wire n443; 
wire n448; 
wire n453; 
wire n458; 
wire n463; 
wire n468; 
wire n473; 
wire n478; 
wire n483; 
wire n488; 
wire n493; 
wire n498; 
wire n503; 
wire n508; 
wire n513; 
wire n518; 
wire n523; 
wire n528; 
wire n533; 
wire n538; 
wire n543; 
wire n548; 
wire n553; 
wire n558; 
wire n563; 
wire n568; 
wire n573; 
wire n578; 
wire n583; 
wire n588; 
wire n593; 
wire n598; 
wire n603; 
wire n608; 
wire n613; 
wire n618; 
wire n623; 
wire n628; 
wire n633; 
wire n638; 
wire n643; 
wire n648; 
wire n653; 
wire n658; 
wire n663; 
wire n668; 
wire n673; 
wire n678; 
wire n683; 
wire n688; 
wire n693; 
wire n698; 
wire n703; 
wire n708; 
wire n713; 
wire n718; 
wire n723; 
wire n728; 
wire n733; 
wire n738; 
wire n743; 
wire n748; 
wire n753; 
wire n758; 
wire n763; 
wire n768; 
wire n773; 
wire n778; 
wire n783; 
wire n788; 
wire n793; 
wire n798; 
wire n803; 
wire n808; 
wire n813; 
wire n818; 
wire n823; 
wire n828; 
wire n833; 
wire n838; 
wire n843; 
wire n848; 
wire n853; 
wire n858; 
wire n863; 
wire n868; 
wire n873; 
wire n878; 
wire n883; 
wire n888; 
wire n893; 
wire n898; 
wire n903; 
wire n908; 
wire n913; 
wire n918; 
wire n923; 
wire n928; 
wire n933; 
wire n938; 
wire n943; 
wire n948; 
wire n953; 
wire n958; 
wire n963; 
wire n968; 
wire n973; 
wire n978; 
wire n982; 
wire n986; 
wire n990; 
wire n994; 
wire n998; 
input nRESET_G;
AND2X2 AND2X2_1 ( .A(_abc_40319_new_n524_), .B(_abc_40319_new_n525_), .Y(_abc_40319_new_n526_));
AND2X2 AND2X2_10 ( .A(_abc_40319_new_n548_), .B(_abc_40319_new_n549_), .Y(_abc_40319_new_n550_));
AND2X2 AND2X2_100 ( .A(_abc_40319_new_n730_), .B(_abc_40319_new_n731_), .Y(_abc_40319_new_n732_));
AND2X2 AND2X2_1000 ( .A(_abc_40319_new_n2560_), .B(_abc_40319_new_n2555_), .Y(_abc_40319_new_n2561_));
AND2X2 AND2X2_1001 ( .A(_abc_40319_new_n2553_), .B(_abc_40319_new_n2555_), .Y(_abc_40319_new_n2563_));
AND2X2 AND2X2_1002 ( .A(_abc_40319_new_n2560_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2564_));
AND2X2 AND2X2_1003 ( .A(_abc_40319_new_n2566_), .B(_abc_40319_new_n2562_), .Y(_abc_40319_new_n2567_));
AND2X2 AND2X2_1004 ( .A(_abc_40319_new_n1046_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2569_));
AND2X2 AND2X2_1005 ( .A(_abc_40319_new_n1034_), .B(_abc_40319_new_n2555_), .Y(_abc_40319_new_n2570_));
AND2X2 AND2X2_1006 ( .A(_abc_40319_new_n1010_), .B(_abc_40319_new_n613_), .Y(_abc_40319_new_n2571_));
AND2X2 AND2X2_1007 ( .A(_abc_40319_new_n2555_), .B(_abc_40319_new_n2549_), .Y(_abc_40319_new_n2576_));
AND2X2 AND2X2_1008 ( .A(_abc_40319_new_n2575_), .B(_abc_40319_new_n2576_), .Y(_abc_40319_new_n2577_));
AND2X2 AND2X2_1009 ( .A(_abc_40319_new_n2578_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2579_));
AND2X2 AND2X2_101 ( .A(_abc_40319_new_n729_), .B(_abc_40319_new_n732_), .Y(_abc_40319_new_n733_));
AND2X2 AND2X2_1010 ( .A(_abc_40319_new_n2574_), .B(_abc_40319_new_n2581_), .Y(_abc_40319_new_n2582_));
AND2X2 AND2X2_1011 ( .A(_abc_40319_new_n2583_), .B(_abc_40319_new_n2576_), .Y(_abc_40319_new_n2584_));
AND2X2 AND2X2_1012 ( .A(_abc_40319_new_n2585_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2586_));
AND2X2 AND2X2_1013 ( .A(_abc_40319_new_n998_), .B(_abc_40319_new_n2555_), .Y(_abc_40319_new_n2589_));
AND2X2 AND2X2_1014 ( .A(_abc_40319_new_n1010_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2590_));
AND2X2 AND2X2_1015 ( .A(_abc_40319_new_n746_), .B(_abc_40319_new_n613_), .Y(_abc_40319_new_n2591_));
AND2X2 AND2X2_1016 ( .A(_abc_40319_new_n2594_), .B(_abc_40319_new_n2588_), .Y(_abc_40319_new_n2595_));
AND2X2 AND2X2_1017 ( .A(_abc_40319_new_n689_), .B(_abc_40319_new_n2555_), .Y(_abc_40319_new_n2598_));
AND2X2 AND2X2_1018 ( .A(_abc_40319_new_n746_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2599_));
AND2X2 AND2X2_1019 ( .A(_abc_40319_new_n795_), .B(_abc_40319_new_n613_), .Y(_abc_40319_new_n2600_));
AND2X2 AND2X2_102 ( .A(_abc_40319_new_n733_), .B(REG2_REG_5_), .Y(_abc_40319_new_n734_));
AND2X2 AND2X2_1020 ( .A(_abc_40319_new_n2603_), .B(_abc_40319_new_n2576_), .Y(_abc_40319_new_n2604_));
AND2X2 AND2X2_1021 ( .A(_abc_40319_new_n2605_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2606_));
AND2X2 AND2X2_1022 ( .A(_abc_40319_new_n2597_), .B(_abc_40319_new_n2608_), .Y(_abc_40319_new_n2609_));
AND2X2 AND2X2_1023 ( .A(_abc_40319_new_n848_), .B(_abc_40319_new_n2555_), .Y(_abc_40319_new_n2613_));
AND2X2 AND2X2_1024 ( .A(_abc_40319_new_n2614_), .B(_abc_40319_new_n2615_), .Y(_abc_40319_new_n2616_));
AND2X2 AND2X2_1025 ( .A(_abc_40319_new_n2616_), .B(_abc_40319_new_n2612_), .Y(_abc_40319_new_n2617_));
AND2X2 AND2X2_1026 ( .A(_abc_40319_new_n864_), .B(_abc_40319_new_n2576_), .Y(_abc_40319_new_n2619_));
AND2X2 AND2X2_1027 ( .A(_abc_40319_new_n847_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2620_));
AND2X2 AND2X2_1028 ( .A(_abc_40319_new_n2618_), .B(_abc_40319_new_n2621_), .Y(_abc_40319_new_n2622_));
AND2X2 AND2X2_1029 ( .A(_abc_40319_new_n904_), .B(_abc_40319_new_n645_), .Y(_abc_40319_new_n2624_));
AND2X2 AND2X2_103 ( .A(_abc_40319_new_n716_), .B(_abc_40319_new_n732_), .Y(_abc_40319_new_n736_));
AND2X2 AND2X2_1030 ( .A(_abc_40319_new_n891_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2626_));
AND2X2 AND2X2_1031 ( .A(_abc_40319_new_n904_), .B(_abc_40319_new_n670_), .Y(_abc_40319_new_n2628_));
AND2X2 AND2X2_1032 ( .A(_abc_40319_new_n904_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2630_));
AND2X2 AND2X2_1033 ( .A(_abc_40319_new_n924_), .B(_abc_40319_new_n613_), .Y(_abc_40319_new_n2631_));
AND2X2 AND2X2_1034 ( .A(_abc_40319_new_n891_), .B(_abc_40319_new_n2555_), .Y(_abc_40319_new_n2633_));
AND2X2 AND2X2_1035 ( .A(_abc_40319_new_n924_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2636_));
AND2X2 AND2X2_1036 ( .A(_abc_40319_new_n930_), .B(_abc_40319_new_n2555_), .Y(_abc_40319_new_n2637_));
AND2X2 AND2X2_1037 ( .A(_abc_40319_new_n924_), .B(_abc_40319_new_n645_), .Y(_abc_40319_new_n2640_));
AND2X2 AND2X2_1038 ( .A(_abc_40319_new_n930_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2642_));
AND2X2 AND2X2_1039 ( .A(_abc_40319_new_n924_), .B(_abc_40319_new_n670_), .Y(_abc_40319_new_n2644_));
AND2X2 AND2X2_104 ( .A(_abc_40319_new_n736_), .B(REG0_REG_5_), .Y(_abc_40319_new_n737_));
AND2X2 AND2X2_1040 ( .A(_abc_40319_new_n2646_), .B(_abc_40319_new_n2635_), .Y(_abc_40319_new_n2647_));
AND2X2 AND2X2_1041 ( .A(_abc_40319_new_n2648_), .B(_abc_40319_new_n2623_), .Y(_abc_40319_new_n2649_));
AND2X2 AND2X2_1042 ( .A(_abc_40319_new_n2652_), .B(_abc_40319_new_n2653_), .Y(_abc_40319_new_n2654_));
AND2X2 AND2X2_1043 ( .A(_abc_40319_new_n2654_), .B(_abc_40319_new_n2651_), .Y(_abc_40319_new_n2655_));
AND2X2 AND2X2_1044 ( .A(_abc_40319_new_n2658_), .B(_abc_40319_new_n2657_), .Y(_abc_40319_new_n2659_));
AND2X2 AND2X2_1045 ( .A(_abc_40319_new_n784_), .B(_abc_40319_new_n2551_), .Y(_abc_40319_new_n2661_));
AND2X2 AND2X2_1046 ( .A(_abc_40319_new_n795_), .B(_abc_40319_new_n2555_), .Y(_abc_40319_new_n2662_));
AND2X2 AND2X2_1047 ( .A(_abc_40319_new_n784_), .B(_abc_40319_new_n2555_), .Y(_abc_40319_new_n2665_));
AND2X2 AND2X2_1048 ( .A(_abc_40319_new_n795_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2667_));
AND2X2 AND2X2_1049 ( .A(_abc_40319_new_n2669_), .B(_abc_40319_new_n2668_), .Y(_abc_40319_new_n2670_));
AND2X2 AND2X2_105 ( .A(_abc_40319_new_n729_), .B(_abc_40319_new_n721_), .Y(_abc_40319_new_n738_));
AND2X2 AND2X2_1050 ( .A(_abc_40319_new_n2670_), .B(_abc_40319_new_n2666_), .Y(_abc_40319_new_n2671_));
AND2X2 AND2X2_1051 ( .A(_abc_40319_new_n2673_), .B(_abc_40319_new_n2549_), .Y(_abc_40319_new_n2674_));
AND2X2 AND2X2_1052 ( .A(_abc_40319_new_n2674_), .B(_abc_40319_new_n2675_), .Y(_abc_40319_new_n2676_));
AND2X2 AND2X2_1053 ( .A(_abc_40319_new_n2676_), .B(_abc_40319_new_n2677_), .Y(_abc_40319_new_n2678_));
AND2X2 AND2X2_1054 ( .A(_abc_40319_new_n2678_), .B(_abc_40319_new_n2638_), .Y(_abc_40319_new_n2679_));
AND2X2 AND2X2_1055 ( .A(_abc_40319_new_n2679_), .B(_abc_40319_new_n2634_), .Y(_abc_40319_new_n2680_));
AND2X2 AND2X2_1056 ( .A(_abc_40319_new_n2681_), .B(_abc_40319_new_n2672_), .Y(_abc_40319_new_n2682_));
AND2X2 AND2X2_1057 ( .A(_abc_40319_new_n2682_), .B(_abc_40319_new_n2660_), .Y(_abc_40319_new_n2683_));
AND2X2 AND2X2_1058 ( .A(_abc_40319_new_n2649_), .B(_abc_40319_new_n2683_), .Y(_abc_40319_new_n2684_));
AND2X2 AND2X2_1059 ( .A(_abc_40319_new_n2655_), .B(_abc_40319_new_n2659_), .Y(_abc_40319_new_n2685_));
AND2X2 AND2X2_106 ( .A(REG3_REG_3_), .B(REG3_REG_4_), .Y(_abc_40319_new_n739_));
AND2X2 AND2X2_1060 ( .A(_abc_40319_new_n2672_), .B(_abc_40319_new_n2685_), .Y(_abc_40319_new_n2686_));
AND2X2 AND2X2_1061 ( .A(_abc_40319_new_n2671_), .B(_abc_40319_new_n2664_), .Y(_abc_40319_new_n2687_));
AND2X2 AND2X2_1062 ( .A(_abc_40319_new_n2660_), .B(_abc_40319_new_n2617_), .Y(_abc_40319_new_n2689_));
AND2X2 AND2X2_1063 ( .A(_abc_40319_new_n2689_), .B(_abc_40319_new_n2688_), .Y(_abc_40319_new_n2690_));
AND2X2 AND2X2_1064 ( .A(_abc_40319_new_n2690_), .B(_abc_40319_new_n2672_), .Y(_abc_40319_new_n2691_));
AND2X2 AND2X2_1065 ( .A(_abc_40319_new_n1758_), .B(_abc_40319_new_n2555_), .Y(_abc_40319_new_n2696_));
AND2X2 AND2X2_1066 ( .A(_abc_40319_new_n1769_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2697_));
AND2X2 AND2X2_1067 ( .A(_abc_40319_new_n1625_), .B(_abc_40319_new_n613_), .Y(_abc_40319_new_n2698_));
AND2X2 AND2X2_1068 ( .A(_abc_40319_new_n2701_), .B(_abc_40319_new_n2576_), .Y(_abc_40319_new_n2702_));
AND2X2 AND2X2_1069 ( .A(_abc_40319_new_n2703_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2704_));
AND2X2 AND2X2_107 ( .A(_abc_40319_new_n739_), .B(REG3_REG_5_), .Y(_abc_40319_new_n740_));
AND2X2 AND2X2_1070 ( .A(_abc_40319_new_n2700_), .B(_abc_40319_new_n2705_), .Y(_abc_40319_new_n2706_));
AND2X2 AND2X2_1071 ( .A(_abc_40319_new_n1614_), .B(_abc_40319_new_n2555_), .Y(_abc_40319_new_n2707_));
AND2X2 AND2X2_1072 ( .A(_abc_40319_new_n1625_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2708_));
AND2X2 AND2X2_1073 ( .A(_abc_40319_new_n1146_), .B(_abc_40319_new_n613_), .Y(_abc_40319_new_n2709_));
AND2X2 AND2X2_1074 ( .A(_abc_40319_new_n2712_), .B(_abc_40319_new_n2576_), .Y(_abc_40319_new_n2713_));
AND2X2 AND2X2_1075 ( .A(_abc_40319_new_n2714_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2715_));
AND2X2 AND2X2_1076 ( .A(_abc_40319_new_n2711_), .B(_abc_40319_new_n2716_), .Y(_abc_40319_new_n2717_));
AND2X2 AND2X2_1077 ( .A(_abc_40319_new_n2573_), .B(_abc_40319_new_n2580_), .Y(_abc_40319_new_n2722_));
AND2X2 AND2X2_1078 ( .A(_abc_40319_new_n1572_), .B(_abc_40319_new_n2555_), .Y(_abc_40319_new_n2723_));
AND2X2 AND2X2_1079 ( .A(_abc_40319_new_n1146_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2724_));
AND2X2 AND2X2_108 ( .A(_abc_40319_new_n741_), .B(_abc_40319_new_n742_), .Y(_abc_40319_new_n743_));
AND2X2 AND2X2_1080 ( .A(_abc_40319_new_n1046_), .B(_abc_40319_new_n613_), .Y(_abc_40319_new_n2725_));
AND2X2 AND2X2_1081 ( .A(_abc_40319_new_n2728_), .B(_abc_40319_new_n2576_), .Y(_abc_40319_new_n2729_));
AND2X2 AND2X2_1082 ( .A(_abc_40319_new_n2730_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2731_));
AND2X2 AND2X2_1083 ( .A(_abc_40319_new_n2727_), .B(_abc_40319_new_n2732_), .Y(_abc_40319_new_n2733_));
AND2X2 AND2X2_1084 ( .A(_abc_40319_new_n2721_), .B(_abc_40319_new_n2735_), .Y(_abc_40319_new_n2736_));
AND2X2 AND2X2_1085 ( .A(_abc_40319_new_n2736_), .B(_abc_40319_new_n2719_), .Y(_abc_40319_new_n2737_));
AND2X2 AND2X2_1086 ( .A(_abc_40319_new_n2602_), .B(_abc_40319_new_n2607_), .Y(_abc_40319_new_n2738_));
AND2X2 AND2X2_1087 ( .A(_abc_40319_new_n2597_), .B(_abc_40319_new_n2738_), .Y(_abc_40319_new_n2739_));
AND2X2 AND2X2_1088 ( .A(_abc_40319_new_n2740_), .B(_abc_40319_new_n2737_), .Y(_abc_40319_new_n2741_));
AND2X2 AND2X2_1089 ( .A(_abc_40319_new_n2695_), .B(_abc_40319_new_n2741_), .Y(_abc_40319_new_n2742_));
AND2X2 AND2X2_109 ( .A(_abc_40319_new_n738_), .B(_abc_40319_new_n743_), .Y(_abc_40319_new_n744_));
AND2X2 AND2X2_1090 ( .A(_abc_40319_new_n1667_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2747_));
AND2X2 AND2X2_1091 ( .A(_abc_40319_new_n1655_), .B(_abc_40319_new_n2555_), .Y(_abc_40319_new_n2748_));
AND2X2 AND2X2_1092 ( .A(_abc_40319_new_n1701_), .B(_abc_40319_new_n613_), .Y(_abc_40319_new_n2749_));
AND2X2 AND2X2_1093 ( .A(_abc_40319_new_n2753_), .B(_abc_40319_new_n2576_), .Y(_abc_40319_new_n2754_));
AND2X2 AND2X2_1094 ( .A(_abc_40319_new_n2755_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2756_));
AND2X2 AND2X2_1095 ( .A(_abc_40319_new_n2752_), .B(_abc_40319_new_n2758_), .Y(_abc_40319_new_n2759_));
AND2X2 AND2X2_1096 ( .A(_abc_40319_new_n2760_), .B(_abc_40319_new_n2576_), .Y(_abc_40319_new_n2761_));
AND2X2 AND2X2_1097 ( .A(_abc_40319_new_n2762_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2763_));
AND2X2 AND2X2_1098 ( .A(_abc_40319_new_n1701_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2766_));
AND2X2 AND2X2_1099 ( .A(_abc_40319_new_n1690_), .B(_abc_40319_new_n2555_), .Y(_abc_40319_new_n2767_));
AND2X2 AND2X2_11 ( .A(_abc_40319_new_n547_), .B(_abc_40319_new_n550_), .Y(_abc_40319_new_n551_));
AND2X2 AND2X2_110 ( .A(_abc_40319_new_n705_), .B(_abc_40319_new_n746_), .Y(_abc_40319_new_n747_));
AND2X2 AND2X2_1100 ( .A(_abc_40319_new_n1735_), .B(_abc_40319_new_n613_), .Y(_abc_40319_new_n2768_));
AND2X2 AND2X2_1101 ( .A(_abc_40319_new_n2771_), .B(_abc_40319_new_n2765_), .Y(_abc_40319_new_n2772_));
AND2X2 AND2X2_1102 ( .A(_abc_40319_new_n1735_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2776_));
AND2X2 AND2X2_1103 ( .A(_abc_40319_new_n1724_), .B(_abc_40319_new_n2555_), .Y(_abc_40319_new_n2777_));
AND2X2 AND2X2_1104 ( .A(_abc_40319_new_n1769_), .B(_abc_40319_new_n613_), .Y(_abc_40319_new_n2778_));
AND2X2 AND2X2_1105 ( .A(_abc_40319_new_n2782_), .B(_abc_40319_new_n2576_), .Y(_abc_40319_new_n2783_));
AND2X2 AND2X2_1106 ( .A(_abc_40319_new_n2784_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2785_));
AND2X2 AND2X2_1107 ( .A(_abc_40319_new_n2781_), .B(_abc_40319_new_n2787_), .Y(_abc_40319_new_n2788_));
AND2X2 AND2X2_1108 ( .A(_abc_40319_new_n2789_), .B(_abc_40319_new_n2775_), .Y(_abc_40319_new_n2790_));
AND2X2 AND2X2_1109 ( .A(_abc_40319_new_n2774_), .B(_abc_40319_new_n2790_), .Y(_abc_40319_new_n2791_));
AND2X2 AND2X2_111 ( .A(_abc_40319_new_n749_), .B(_abc_40319_new_n750_), .Y(_abc_40319_new_n751_));
AND2X2 AND2X2_1110 ( .A(_abc_40319_new_n2791_), .B(_abc_40319_new_n2746_), .Y(_abc_40319_new_n2792_));
AND2X2 AND2X2_1111 ( .A(_abc_40319_new_n2792_), .B(_abc_40319_new_n2744_), .Y(_abc_40319_new_n2793_));
AND2X2 AND2X2_1112 ( .A(_abc_40319_new_n2780_), .B(_abc_40319_new_n2786_), .Y(_abc_40319_new_n2796_));
AND2X2 AND2X2_1113 ( .A(_abc_40319_new_n2774_), .B(_abc_40319_new_n2796_), .Y(_abc_40319_new_n2797_));
AND2X2 AND2X2_1114 ( .A(_abc_40319_new_n2770_), .B(_abc_40319_new_n2764_), .Y(_abc_40319_new_n2799_));
AND2X2 AND2X2_1115 ( .A(_abc_40319_new_n2798_), .B(_abc_40319_new_n2799_), .Y(_abc_40319_new_n2800_));
AND2X2 AND2X2_1116 ( .A(_abc_40319_new_n2751_), .B(_abc_40319_new_n2757_), .Y(_abc_40319_new_n2801_));
AND2X2 AND2X2_1117 ( .A(_abc_40319_new_n1506_), .B(_abc_40319_new_n2555_), .Y(_abc_40319_new_n2802_));
AND2X2 AND2X2_1118 ( .A(_abc_40319_new_n1517_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2803_));
AND2X2 AND2X2_1119 ( .A(_abc_40319_new_n1667_), .B(_abc_40319_new_n613_), .Y(_abc_40319_new_n2804_));
AND2X2 AND2X2_112 ( .A(_abc_40319_new_n751_), .B(_abc_40319_new_n645_), .Y(_abc_40319_new_n752_));
AND2X2 AND2X2_1120 ( .A(_abc_40319_new_n2807_), .B(_abc_40319_new_n2576_), .Y(_abc_40319_new_n2808_));
AND2X2 AND2X2_1121 ( .A(_abc_40319_new_n2809_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2810_));
AND2X2 AND2X2_1122 ( .A(_abc_40319_new_n2806_), .B(_abc_40319_new_n2811_), .Y(_abc_40319_new_n2812_));
AND2X2 AND2X2_1123 ( .A(_abc_40319_new_n2795_), .B(_abc_40319_new_n2816_), .Y(_abc_40319_new_n2817_));
AND2X2 AND2X2_1124 ( .A(_abc_40319_new_n1483_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2819_));
AND2X2 AND2X2_1125 ( .A(_abc_40319_new_n1471_), .B(_abc_40319_new_n2555_), .Y(_abc_40319_new_n2820_));
AND2X2 AND2X2_1126 ( .A(_abc_40319_new_n1517_), .B(_abc_40319_new_n613_), .Y(_abc_40319_new_n2821_));
AND2X2 AND2X2_1127 ( .A(_abc_40319_new_n2825_), .B(_abc_40319_new_n2576_), .Y(_abc_40319_new_n2826_));
AND2X2 AND2X2_1128 ( .A(_abc_40319_new_n2827_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2828_));
AND2X2 AND2X2_1129 ( .A(_abc_40319_new_n2824_), .B(_abc_40319_new_n2830_), .Y(_abc_40319_new_n2831_));
AND2X2 AND2X2_113 ( .A(_abc_40319_new_n751_), .B(_abc_40319_new_n697_), .Y(_abc_40319_new_n753_));
AND2X2 AND2X2_1130 ( .A(_abc_40319_new_n2832_), .B(_abc_40319_new_n2818_), .Y(_abc_40319_new_n2833_));
AND2X2 AND2X2_1131 ( .A(_abc_40319_new_n2823_), .B(_abc_40319_new_n2829_), .Y(_abc_40319_new_n2836_));
AND2X2 AND2X2_1132 ( .A(_abc_40319_new_n1398_), .B(_abc_40319_new_n2555_), .Y(_abc_40319_new_n2837_));
AND2X2 AND2X2_1133 ( .A(_abc_40319_new_n1483_), .B(_abc_40319_new_n613_), .Y(_abc_40319_new_n2838_));
AND2X2 AND2X2_1134 ( .A(_abc_40319_new_n1410_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2839_));
AND2X2 AND2X2_1135 ( .A(_abc_40319_new_n2842_), .B(_abc_40319_new_n2576_), .Y(_abc_40319_new_n2843_));
AND2X2 AND2X2_1136 ( .A(_abc_40319_new_n2844_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2845_));
AND2X2 AND2X2_1137 ( .A(_abc_40319_new_n2841_), .B(_abc_40319_new_n2846_), .Y(_abc_40319_new_n2847_));
AND2X2 AND2X2_1138 ( .A(_abc_40319_new_n2835_), .B(_abc_40319_new_n2849_), .Y(_abc_40319_new_n2850_));
AND2X2 AND2X2_1139 ( .A(_abc_40319_new_n1444_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2852_));
AND2X2 AND2X2_114 ( .A(_abc_40319_new_n655_), .B(_abc_40319_new_n670_), .Y(_abc_40319_new_n754_));
AND2X2 AND2X2_1140 ( .A(_abc_40319_new_n1433_), .B(_abc_40319_new_n2555_), .Y(_abc_40319_new_n2853_));
AND2X2 AND2X2_1141 ( .A(_abc_40319_new_n1410_), .B(_abc_40319_new_n613_), .Y(_abc_40319_new_n2854_));
AND2X2 AND2X2_1142 ( .A(_abc_40319_new_n2858_), .B(_abc_40319_new_n2576_), .Y(_abc_40319_new_n2859_));
AND2X2 AND2X2_1143 ( .A(_abc_40319_new_n2860_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2861_));
AND2X2 AND2X2_1144 ( .A(_abc_40319_new_n2857_), .B(_abc_40319_new_n2863_), .Y(_abc_40319_new_n2864_));
AND2X2 AND2X2_1145 ( .A(_abc_40319_new_n2865_), .B(_abc_40319_new_n2851_), .Y(_abc_40319_new_n2866_));
AND2X2 AND2X2_1146 ( .A(_abc_40319_new_n2856_), .B(_abc_40319_new_n2862_), .Y(_abc_40319_new_n2869_));
AND2X2 AND2X2_1147 ( .A(_abc_40319_new_n1374_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2870_));
AND2X2 AND2X2_1148 ( .A(_abc_40319_new_n1363_), .B(_abc_40319_new_n2555_), .Y(_abc_40319_new_n2871_));
AND2X2 AND2X2_1149 ( .A(_abc_40319_new_n1444_), .B(_abc_40319_new_n613_), .Y(_abc_40319_new_n2872_));
AND2X2 AND2X2_115 ( .A(_abc_40319_new_n756_), .B(_abc_40319_new_n663_), .Y(_abc_40319_new_n757_));
AND2X2 AND2X2_1150 ( .A(_abc_40319_new_n2875_), .B(_abc_40319_new_n2576_), .Y(_abc_40319_new_n2876_));
AND2X2 AND2X2_1151 ( .A(_abc_40319_new_n2877_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2878_));
AND2X2 AND2X2_1152 ( .A(_abc_40319_new_n2879_), .B(_abc_40319_new_n2874_), .Y(_abc_40319_new_n2880_));
AND2X2 AND2X2_1153 ( .A(_abc_40319_new_n2868_), .B(_abc_40319_new_n2882_), .Y(_abc_40319_new_n2883_));
AND2X2 AND2X2_1154 ( .A(_abc_40319_new_n1374_), .B(_abc_40319_new_n613_), .Y(_abc_40319_new_n2885_));
AND2X2 AND2X2_1155 ( .A(_abc_40319_new_n1817_), .B(_abc_40319_new_n2555_), .Y(_abc_40319_new_n2886_));
AND2X2 AND2X2_1156 ( .A(_abc_40319_new_n1828_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2887_));
AND2X2 AND2X2_1157 ( .A(_abc_40319_new_n2891_), .B(_abc_40319_new_n2576_), .Y(_abc_40319_new_n2892_));
AND2X2 AND2X2_1158 ( .A(_abc_40319_new_n2893_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2894_));
AND2X2 AND2X2_1159 ( .A(_abc_40319_new_n2890_), .B(_abc_40319_new_n2896_), .Y(_abc_40319_new_n2897_));
AND2X2 AND2X2_116 ( .A(_abc_40319_new_n700_), .B(_abc_40319_new_n663_), .Y(_abc_40319_new_n758_));
AND2X2 AND2X2_1160 ( .A(_abc_40319_new_n2898_), .B(_abc_40319_new_n2884_), .Y(_abc_40319_new_n2899_));
AND2X2 AND2X2_1161 ( .A(_abc_40319_new_n2889_), .B(_abc_40319_new_n2895_), .Y(_abc_40319_new_n2902_));
AND2X2 AND2X2_1162 ( .A(_abc_40319_new_n1852_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2903_));
AND2X2 AND2X2_1163 ( .A(_abc_40319_new_n1841_), .B(_abc_40319_new_n2555_), .Y(_abc_40319_new_n2904_));
AND2X2 AND2X2_1164 ( .A(_abc_40319_new_n1828_), .B(_abc_40319_new_n613_), .Y(_abc_40319_new_n2905_));
AND2X2 AND2X2_1165 ( .A(_abc_40319_new_n2908_), .B(_abc_40319_new_n2576_), .Y(_abc_40319_new_n2909_));
AND2X2 AND2X2_1166 ( .A(_abc_40319_new_n2910_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2911_));
AND2X2 AND2X2_1167 ( .A(_abc_40319_new_n2907_), .B(_abc_40319_new_n2912_), .Y(_abc_40319_new_n2913_));
AND2X2 AND2X2_1168 ( .A(_abc_40319_new_n2901_), .B(_abc_40319_new_n2915_), .Y(_abc_40319_new_n2916_));
AND2X2 AND2X2_1169 ( .A(_abc_40319_new_n1876_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2918_));
AND2X2 AND2X2_117 ( .A(_abc_40319_new_n759_), .B(_abc_40319_new_n702_), .Y(_abc_40319_new_n760_));
AND2X2 AND2X2_1170 ( .A(_abc_40319_new_n1865_), .B(_abc_40319_new_n2555_), .Y(_abc_40319_new_n2919_));
AND2X2 AND2X2_1171 ( .A(_abc_40319_new_n1852_), .B(_abc_40319_new_n613_), .Y(_abc_40319_new_n2920_));
AND2X2 AND2X2_1172 ( .A(_abc_40319_new_n2924_), .B(_abc_40319_new_n2576_), .Y(_abc_40319_new_n2925_));
AND2X2 AND2X2_1173 ( .A(_abc_40319_new_n2926_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2927_));
AND2X2 AND2X2_1174 ( .A(_abc_40319_new_n2923_), .B(_abc_40319_new_n2929_), .Y(_abc_40319_new_n2930_));
AND2X2 AND2X2_1175 ( .A(_abc_40319_new_n2931_), .B(_abc_40319_new_n2917_), .Y(_abc_40319_new_n2932_));
AND2X2 AND2X2_1176 ( .A(_abc_40319_new_n2922_), .B(_abc_40319_new_n2928_), .Y(_abc_40319_new_n2935_));
AND2X2 AND2X2_1177 ( .A(_abc_40319_new_n1340_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2936_));
AND2X2 AND2X2_1178 ( .A(_abc_40319_new_n1329_), .B(_abc_40319_new_n2555_), .Y(_abc_40319_new_n2937_));
AND2X2 AND2X2_1179 ( .A(_abc_40319_new_n1876_), .B(_abc_40319_new_n613_), .Y(_abc_40319_new_n2938_));
AND2X2 AND2X2_118 ( .A(_abc_40319_new_n761_), .B(_abc_40319_new_n663_), .Y(_abc_40319_new_n762_));
AND2X2 AND2X2_1180 ( .A(_abc_40319_new_n2941_), .B(_abc_40319_new_n2576_), .Y(_abc_40319_new_n2942_));
AND2X2 AND2X2_1181 ( .A(_abc_40319_new_n2943_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2944_));
AND2X2 AND2X2_1182 ( .A(_abc_40319_new_n2945_), .B(_abc_40319_new_n2940_), .Y(_abc_40319_new_n2946_));
AND2X2 AND2X2_1183 ( .A(_abc_40319_new_n2934_), .B(_abc_40319_new_n2948_), .Y(_abc_40319_new_n2949_));
AND2X2 AND2X2_1184 ( .A(_abc_40319_new_n1317_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2951_));
AND2X2 AND2X2_1185 ( .A(_abc_40319_new_n1306_), .B(_abc_40319_new_n2555_), .Y(_abc_40319_new_n2952_));
AND2X2 AND2X2_1186 ( .A(_abc_40319_new_n1340_), .B(_abc_40319_new_n613_), .Y(_abc_40319_new_n2953_));
AND2X2 AND2X2_1187 ( .A(_abc_40319_new_n2957_), .B(_abc_40319_new_n2576_), .Y(_abc_40319_new_n2958_));
AND2X2 AND2X2_1188 ( .A(_abc_40319_new_n2959_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2960_));
AND2X2 AND2X2_1189 ( .A(_abc_40319_new_n2962_), .B(_abc_40319_new_n2956_), .Y(_abc_40319_new_n2963_));
AND2X2 AND2X2_119 ( .A(_abc_40319_new_n689_), .B(_abc_40319_new_n763_), .Y(_abc_40319_new_n764_));
AND2X2 AND2X2_1190 ( .A(_abc_40319_new_n2964_), .B(_abc_40319_new_n2950_), .Y(_abc_40319_new_n2965_));
AND2X2 AND2X2_1191 ( .A(_abc_40319_new_n2961_), .B(_abc_40319_new_n2955_), .Y(_abc_40319_new_n2968_));
AND2X2 AND2X2_1192 ( .A(_abc_40319_new_n1285_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2969_));
AND2X2 AND2X2_1193 ( .A(_abc_40319_new_n1274_), .B(_abc_40319_new_n2555_), .Y(_abc_40319_new_n2970_));
AND2X2 AND2X2_1194 ( .A(_abc_40319_new_n1317_), .B(_abc_40319_new_n613_), .Y(_abc_40319_new_n2971_));
AND2X2 AND2X2_1195 ( .A(_abc_40319_new_n2974_), .B(_abc_40319_new_n2576_), .Y(_abc_40319_new_n2975_));
AND2X2 AND2X2_1196 ( .A(_abc_40319_new_n2976_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2977_));
AND2X2 AND2X2_1197 ( .A(_abc_40319_new_n2978_), .B(_abc_40319_new_n2973_), .Y(_abc_40319_new_n2979_));
AND2X2 AND2X2_1198 ( .A(_abc_40319_new_n2967_), .B(_abc_40319_new_n2981_), .Y(_abc_40319_new_n2982_));
AND2X2 AND2X2_1199 ( .A(_abc_40319_new_n1260_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2984_));
AND2X2 AND2X2_12 ( .A(_abc_40319_new_n544_), .B(_abc_40319_new_n551_), .Y(_abc_40319_new_n552_));
AND2X2 AND2X2_120 ( .A(_abc_40319_new_n746_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n765_));
AND2X2 AND2X2_1200 ( .A(_abc_40319_new_n1249_), .B(_abc_40319_new_n2555_), .Y(_abc_40319_new_n2985_));
AND2X2 AND2X2_1201 ( .A(_abc_40319_new_n1285_), .B(_abc_40319_new_n613_), .Y(_abc_40319_new_n2986_));
AND2X2 AND2X2_1202 ( .A(_abc_40319_new_n2990_), .B(_abc_40319_new_n2576_), .Y(_abc_40319_new_n2991_));
AND2X2 AND2X2_1203 ( .A(_abc_40319_new_n2992_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2993_));
AND2X2 AND2X2_1204 ( .A(_abc_40319_new_n2995_), .B(_abc_40319_new_n2989_), .Y(_abc_40319_new_n2996_));
AND2X2 AND2X2_1205 ( .A(_abc_40319_new_n2997_), .B(_abc_40319_new_n2983_), .Y(_abc_40319_new_n2998_));
AND2X2 AND2X2_1206 ( .A(_abc_40319_new_n2994_), .B(_abc_40319_new_n2988_), .Y(_abc_40319_new_n3001_));
AND2X2 AND2X2_1207 ( .A(_abc_40319_new_n1235_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n3002_));
AND2X2 AND2X2_1208 ( .A(_abc_40319_new_n1224_), .B(_abc_40319_new_n2555_), .Y(_abc_40319_new_n3003_));
AND2X2 AND2X2_1209 ( .A(_abc_40319_new_n1260_), .B(_abc_40319_new_n613_), .Y(_abc_40319_new_n3004_));
AND2X2 AND2X2_121 ( .A(_abc_40319_new_n770_), .B(_abc_40319_new_n767_), .Y(_abc_40319_new_n771_));
AND2X2 AND2X2_1210 ( .A(_abc_40319_new_n3007_), .B(_abc_40319_new_n2576_), .Y(_abc_40319_new_n3008_));
AND2X2 AND2X2_1211 ( .A(_abc_40319_new_n3009_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n3010_));
AND2X2 AND2X2_1212 ( .A(_abc_40319_new_n3011_), .B(_abc_40319_new_n3006_), .Y(_abc_40319_new_n3012_));
AND2X2 AND2X2_1213 ( .A(_abc_40319_new_n3000_), .B(_abc_40319_new_n3014_), .Y(_abc_40319_new_n3015_));
AND2X2 AND2X2_1214 ( .A(_abc_40319_new_n1210_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n3017_));
AND2X2 AND2X2_1215 ( .A(_abc_40319_new_n1180_), .B(_abc_40319_new_n2555_), .Y(_abc_40319_new_n3018_));
AND2X2 AND2X2_1216 ( .A(_abc_40319_new_n1235_), .B(_abc_40319_new_n613_), .Y(_abc_40319_new_n3019_));
AND2X2 AND2X2_1217 ( .A(_abc_40319_new_n3023_), .B(_abc_40319_new_n2576_), .Y(_abc_40319_new_n3024_));
AND2X2 AND2X2_1218 ( .A(_abc_40319_new_n3025_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n3026_));
AND2X2 AND2X2_1219 ( .A(_abc_40319_new_n3028_), .B(_abc_40319_new_n3022_), .Y(_abc_40319_new_n3029_));
AND2X2 AND2X2_122 ( .A(_abc_40319_new_n771_), .B(_abc_40319_new_n748_), .Y(_abc_40319_new_n772_));
AND2X2 AND2X2_1220 ( .A(_abc_40319_new_n3030_), .B(_abc_40319_new_n3016_), .Y(_abc_40319_new_n3031_));
AND2X2 AND2X2_1221 ( .A(_abc_40319_new_n3027_), .B(_abc_40319_new_n3021_), .Y(_abc_40319_new_n3034_));
AND2X2 AND2X2_1222 ( .A(_abc_40319_new_n1980_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n3035_));
AND2X2 AND2X2_1223 ( .A(_abc_40319_new_n2089_), .B(_abc_40319_new_n2555_), .Y(_abc_40319_new_n3036_));
AND2X2 AND2X2_1224 ( .A(_abc_40319_new_n1210_), .B(_abc_40319_new_n613_), .Y(_abc_40319_new_n3037_));
AND2X2 AND2X2_1225 ( .A(_abc_40319_new_n3040_), .B(_abc_40319_new_n2576_), .Y(_abc_40319_new_n3041_));
AND2X2 AND2X2_1226 ( .A(_abc_40319_new_n3042_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n3043_));
AND2X2 AND2X2_1227 ( .A(_abc_40319_new_n3044_), .B(_abc_40319_new_n3039_), .Y(_abc_40319_new_n3045_));
AND2X2 AND2X2_1228 ( .A(_abc_40319_new_n3033_), .B(_abc_40319_new_n3047_), .Y(_abc_40319_new_n3048_));
AND2X2 AND2X2_1229 ( .A(_abc_40319_new_n1980_), .B(_abc_40319_new_n613_), .Y(_abc_40319_new_n3050_));
AND2X2 AND2X2_123 ( .A(_abc_40319_new_n675_), .B(IR_REG_4_), .Y(_abc_40319_new_n774_));
AND2X2 AND2X2_1230 ( .A(_abc_40319_new_n817_), .B(DATAI_29_), .Y(_abc_40319_new_n3051_));
AND2X2 AND2X2_1231 ( .A(_abc_40319_new_n3051_), .B(_abc_40319_new_n2555_), .Y(_abc_40319_new_n3052_));
AND2X2 AND2X2_1232 ( .A(_abc_40319_new_n2123_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n3053_));
AND2X2 AND2X2_1233 ( .A(_abc_40319_new_n3057_), .B(_abc_40319_new_n2576_), .Y(_abc_40319_new_n3058_));
AND2X2 AND2X2_1234 ( .A(_abc_40319_new_n3059_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n3060_));
AND2X2 AND2X2_1235 ( .A(_abc_40319_new_n3056_), .B(_abc_40319_new_n3062_), .Y(_abc_40319_new_n3063_));
AND2X2 AND2X2_1236 ( .A(_abc_40319_new_n3064_), .B(_abc_40319_new_n3049_), .Y(_abc_40319_new_n3065_));
AND2X2 AND2X2_1237 ( .A(_abc_40319_new_n3055_), .B(_abc_40319_new_n3061_), .Y(_abc_40319_new_n3068_));
AND2X2 AND2X2_1238 ( .A(_abc_40319_new_n817_), .B(DATAI_30_), .Y(_abc_40319_new_n3069_));
AND2X2 AND2X2_1239 ( .A(_abc_40319_new_n3069_), .B(_abc_40319_new_n2555_), .Y(_abc_40319_new_n3070_));
AND2X2 AND2X2_124 ( .A(_abc_40319_new_n776_), .B(IR_REG_31_), .Y(_abc_40319_new_n777_));
AND2X2 AND2X2_1240 ( .A(_abc_40319_new_n736_), .B(REG0_REG_30_), .Y(_abc_40319_new_n3071_));
AND2X2 AND2X2_1241 ( .A(_abc_40319_new_n733_), .B(REG2_REG_30_), .Y(_abc_40319_new_n3072_));
AND2X2 AND2X2_1242 ( .A(_abc_40319_new_n722_), .B(REG1_REG_30_), .Y(_abc_40319_new_n3073_));
AND2X2 AND2X2_1243 ( .A(_abc_40319_new_n3075_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n3076_));
AND2X2 AND2X2_1244 ( .A(_abc_40319_new_n2560_), .B(_abc_40319_new_n3075_), .Y(_abc_40319_new_n3078_));
AND2X2 AND2X2_1245 ( .A(_abc_40319_new_n3078_), .B(_abc_40319_new_n670_), .Y(_abc_40319_new_n3079_));
AND2X2 AND2X2_1246 ( .A(_abc_40319_new_n3075_), .B(_abc_40319_new_n645_), .Y(_abc_40319_new_n3080_));
AND2X2 AND2X2_1247 ( .A(_abc_40319_new_n3069_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n3081_));
AND2X2 AND2X2_1248 ( .A(_abc_40319_new_n3084_), .B(_abc_40319_new_n3077_), .Y(_abc_40319_new_n3085_));
AND2X2 AND2X2_1249 ( .A(_abc_40319_new_n3067_), .B(_abc_40319_new_n3087_), .Y(_abc_40319_new_n3088_));
AND2X2 AND2X2_125 ( .A(_abc_40319_new_n524_), .B(IR_REG_4_), .Y(_abc_40319_new_n778_));
AND2X2 AND2X2_1250 ( .A(_abc_40319_new_n3089_), .B(_abc_40319_new_n3090_), .Y(_abc_40319_new_n3091_));
AND2X2 AND2X2_1251 ( .A(_abc_40319_new_n3093_), .B(_abc_40319_new_n2568_), .Y(_abc_40319_new_n3094_));
AND2X2 AND2X2_1252 ( .A(_abc_40319_new_n3096_), .B(_abc_40319_new_n670_), .Y(_abc_40319_new_n3097_));
AND2X2 AND2X2_1253 ( .A(_abc_40319_new_n751_), .B(_abc_40319_new_n670_), .Y(_abc_40319_new_n3098_));
AND2X2 AND2X2_1254 ( .A(_abc_40319_new_n2123_), .B(_abc_40319_new_n3059_), .Y(_abc_40319_new_n3099_));
AND2X2 AND2X2_1255 ( .A(_abc_40319_new_n3057_), .B(_abc_40319_new_n3051_), .Y(_abc_40319_new_n3101_));
AND2X2 AND2X2_1256 ( .A(_abc_40319_new_n3102_), .B(_abc_40319_new_n3100_), .Y(_abc_40319_new_n3103_));
AND2X2 AND2X2_1257 ( .A(_abc_40319_new_n1235_), .B(_abc_40319_new_n3009_), .Y(_abc_40319_new_n3104_));
AND2X2 AND2X2_1258 ( .A(_abc_40319_new_n3007_), .B(_abc_40319_new_n1224_), .Y(_abc_40319_new_n3105_));
AND2X2 AND2X2_1259 ( .A(_abc_40319_new_n2908_), .B(_abc_40319_new_n2910_), .Y(_abc_40319_new_n3108_));
AND2X2 AND2X2_126 ( .A(_abc_40319_new_n640_), .B(_abc_40319_new_n780_), .Y(_abc_40319_new_n781_));
AND2X2 AND2X2_1260 ( .A(_abc_40319_new_n1852_), .B(_abc_40319_new_n1841_), .Y(_abc_40319_new_n3109_));
AND2X2 AND2X2_1261 ( .A(_abc_40319_new_n2827_), .B(_abc_40319_new_n1483_), .Y(_abc_40319_new_n3111_));
AND2X2 AND2X2_1262 ( .A(_abc_40319_new_n2825_), .B(_abc_40319_new_n1471_), .Y(_abc_40319_new_n3112_));
AND2X2 AND2X2_1263 ( .A(_abc_40319_new_n903_), .B(_abc_40319_new_n891_), .Y(_abc_40319_new_n3117_));
AND2X2 AND2X2_1264 ( .A(_abc_40319_new_n3114_), .B(_abc_40319_new_n3119_), .Y(_abc_40319_new_n3120_));
AND2X2 AND2X2_1265 ( .A(_abc_40319_new_n2605_), .B(_abc_40319_new_n746_), .Y(_abc_40319_new_n3121_));
AND2X2 AND2X2_1266 ( .A(_abc_40319_new_n2603_), .B(_abc_40319_new_n689_), .Y(_abc_40319_new_n3122_));
AND2X2 AND2X2_1267 ( .A(_abc_40319_new_n865_), .B(_abc_40319_new_n847_), .Y(_abc_40319_new_n3125_));
AND2X2 AND2X2_1268 ( .A(_abc_40319_new_n848_), .B(_abc_40319_new_n864_), .Y(_abc_40319_new_n3126_));
AND2X2 AND2X2_1269 ( .A(_abc_40319_new_n3124_), .B(_abc_40319_new_n3128_), .Y(_abc_40319_new_n3129_));
AND2X2 AND2X2_127 ( .A(_abc_40319_new_n782_), .B(_abc_40319_new_n783_), .Y(_abc_40319_new_n784_));
AND2X2 AND2X2_1270 ( .A(_abc_40319_new_n3120_), .B(_abc_40319_new_n3129_), .Y(_abc_40319_new_n3130_));
AND2X2 AND2X2_1271 ( .A(_abc_40319_new_n2650_), .B(_abc_40319_new_n820_), .Y(_abc_40319_new_n3131_));
AND2X2 AND2X2_1272 ( .A(_abc_40319_new_n829_), .B(_abc_40319_new_n819_), .Y(_abc_40319_new_n3132_));
AND2X2 AND2X2_1273 ( .A(_abc_40319_new_n924_), .B(_abc_40319_new_n942_), .Y(_abc_40319_new_n3135_));
AND2X2 AND2X2_1274 ( .A(_abc_40319_new_n930_), .B(_abc_40319_new_n954_), .Y(_abc_40319_new_n3136_));
AND2X2 AND2X2_1275 ( .A(_abc_40319_new_n3134_), .B(_abc_40319_new_n3138_), .Y(_abc_40319_new_n3139_));
AND2X2 AND2X2_1276 ( .A(_abc_40319_new_n2755_), .B(_abc_40319_new_n1667_), .Y(_abc_40319_new_n3140_));
AND2X2 AND2X2_1277 ( .A(_abc_40319_new_n2753_), .B(_abc_40319_new_n1655_), .Y(_abc_40319_new_n3141_));
AND2X2 AND2X2_1278 ( .A(_abc_40319_new_n2809_), .B(_abc_40319_new_n1517_), .Y(_abc_40319_new_n3144_));
AND2X2 AND2X2_1279 ( .A(_abc_40319_new_n2807_), .B(_abc_40319_new_n1506_), .Y(_abc_40319_new_n3145_));
AND2X2 AND2X2_128 ( .A(_abc_40319_new_n784_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n785_));
AND2X2 AND2X2_1280 ( .A(_abc_40319_new_n3143_), .B(_abc_40319_new_n3147_), .Y(_abc_40319_new_n3148_));
AND2X2 AND2X2_1281 ( .A(_abc_40319_new_n3148_), .B(_abc_40319_new_n3139_), .Y(_abc_40319_new_n3149_));
AND2X2 AND2X2_1282 ( .A(_abc_40319_new_n3149_), .B(_abc_40319_new_n3130_), .Y(_abc_40319_new_n3150_));
AND2X2 AND2X2_1283 ( .A(_abc_40319_new_n1374_), .B(_abc_40319_new_n2877_), .Y(_abc_40319_new_n3151_));
AND2X2 AND2X2_1284 ( .A(_abc_40319_new_n2875_), .B(_abc_40319_new_n1363_), .Y(_abc_40319_new_n3152_));
AND2X2 AND2X2_1285 ( .A(_abc_40319_new_n2714_), .B(_abc_40319_new_n1625_), .Y(_abc_40319_new_n3155_));
AND2X2 AND2X2_1286 ( .A(_abc_40319_new_n2712_), .B(_abc_40319_new_n1614_), .Y(_abc_40319_new_n3156_));
AND2X2 AND2X2_1287 ( .A(_abc_40319_new_n3159_), .B(_abc_40319_new_n2553_), .Y(_abc_40319_new_n3160_));
AND2X2 AND2X2_1288 ( .A(_abc_40319_new_n2560_), .B(_abc_40319_new_n3162_), .Y(_abc_40319_new_n3163_));
AND2X2 AND2X2_1289 ( .A(_abc_40319_new_n3161_), .B(_abc_40319_new_n3164_), .Y(_abc_40319_new_n3165_));
AND2X2 AND2X2_129 ( .A(_abc_40319_new_n722_), .B(REG1_REG_4_), .Y(_abc_40319_new_n786_));
AND2X2 AND2X2_1290 ( .A(_abc_40319_new_n3166_), .B(_abc_40319_new_n3069_), .Y(_abc_40319_new_n3167_));
AND2X2 AND2X2_1291 ( .A(_abc_40319_new_n3075_), .B(_abc_40319_new_n3169_), .Y(_abc_40319_new_n3170_));
AND2X2 AND2X2_1292 ( .A(_abc_40319_new_n3168_), .B(_abc_40319_new_n3171_), .Y(_abc_40319_new_n3172_));
AND2X2 AND2X2_1293 ( .A(_abc_40319_new_n3165_), .B(_abc_40319_new_n3172_), .Y(_abc_40319_new_n3173_));
AND2X2 AND2X2_1294 ( .A(_abc_40319_new_n2730_), .B(_abc_40319_new_n1146_), .Y(_abc_40319_new_n3174_));
AND2X2 AND2X2_1295 ( .A(_abc_40319_new_n2728_), .B(_abc_40319_new_n1572_), .Y(_abc_40319_new_n3175_));
AND2X2 AND2X2_1296 ( .A(_abc_40319_new_n3173_), .B(_abc_40319_new_n3177_), .Y(_abc_40319_new_n3178_));
AND2X2 AND2X2_1297 ( .A(_abc_40319_new_n3178_), .B(_abc_40319_new_n3158_), .Y(_abc_40319_new_n3179_));
AND2X2 AND2X2_1298 ( .A(_abc_40319_new_n3179_), .B(_abc_40319_new_n3154_), .Y(_abc_40319_new_n3180_));
AND2X2 AND2X2_1299 ( .A(_abc_40319_new_n3180_), .B(_abc_40319_new_n3150_), .Y(_abc_40319_new_n3181_));
AND2X2 AND2X2_13 ( .A(_abc_40319_new_n537_), .B(_abc_40319_new_n552_), .Y(_abc_40319_new_n553_));
AND2X2 AND2X2_130 ( .A(_abc_40319_new_n733_), .B(REG2_REG_4_), .Y(_abc_40319_new_n787_));
AND2X2 AND2X2_1300 ( .A(_abc_40319_new_n3181_), .B(_abc_40319_new_n3110_), .Y(_abc_40319_new_n3182_));
AND2X2 AND2X2_1301 ( .A(_abc_40319_new_n2860_), .B(_abc_40319_new_n1444_), .Y(_abc_40319_new_n3183_));
AND2X2 AND2X2_1302 ( .A(_abc_40319_new_n2858_), .B(_abc_40319_new_n1433_), .Y(_abc_40319_new_n3184_));
AND2X2 AND2X2_1303 ( .A(_abc_40319_new_n1828_), .B(_abc_40319_new_n2893_), .Y(_abc_40319_new_n3187_));
AND2X2 AND2X2_1304 ( .A(_abc_40319_new_n2891_), .B(_abc_40319_new_n1817_), .Y(_abc_40319_new_n3188_));
AND2X2 AND2X2_1305 ( .A(_abc_40319_new_n3190_), .B(_abc_40319_new_n3186_), .Y(_abc_40319_new_n3191_));
AND2X2 AND2X2_1306 ( .A(_abc_40319_new_n3182_), .B(_abc_40319_new_n3191_), .Y(_abc_40319_new_n3192_));
AND2X2 AND2X2_1307 ( .A(_abc_40319_new_n2974_), .B(_abc_40319_new_n1274_), .Y(_abc_40319_new_n3193_));
AND2X2 AND2X2_1308 ( .A(_abc_40319_new_n1285_), .B(_abc_40319_new_n2976_), .Y(_abc_40319_new_n3194_));
AND2X2 AND2X2_1309 ( .A(_abc_40319_new_n1340_), .B(_abc_40319_new_n2943_), .Y(_abc_40319_new_n3197_));
AND2X2 AND2X2_131 ( .A(_abc_40319_new_n736_), .B(REG0_REG_4_), .Y(_abc_40319_new_n789_));
AND2X2 AND2X2_1310 ( .A(_abc_40319_new_n2941_), .B(_abc_40319_new_n1329_), .Y(_abc_40319_new_n3198_));
AND2X2 AND2X2_1311 ( .A(_abc_40319_new_n1876_), .B(_abc_40319_new_n2926_), .Y(_abc_40319_new_n3201_));
AND2X2 AND2X2_1312 ( .A(_abc_40319_new_n2924_), .B(_abc_40319_new_n1865_), .Y(_abc_40319_new_n3202_));
AND2X2 AND2X2_1313 ( .A(_abc_40319_new_n2703_), .B(_abc_40319_new_n1769_), .Y(_abc_40319_new_n3205_));
AND2X2 AND2X2_1314 ( .A(_abc_40319_new_n2701_), .B(_abc_40319_new_n1758_), .Y(_abc_40319_new_n3206_));
AND2X2 AND2X2_1315 ( .A(_abc_40319_new_n2578_), .B(_abc_40319_new_n1046_), .Y(_abc_40319_new_n3209_));
AND2X2 AND2X2_1316 ( .A(_abc_40319_new_n2575_), .B(_abc_40319_new_n1034_), .Y(_abc_40319_new_n3210_));
AND2X2 AND2X2_1317 ( .A(_abc_40319_new_n2585_), .B(_abc_40319_new_n1010_), .Y(_abc_40319_new_n3213_));
AND2X2 AND2X2_1318 ( .A(_abc_40319_new_n2583_), .B(_abc_40319_new_n998_), .Y(_abc_40319_new_n3214_));
AND2X2 AND2X2_1319 ( .A(_abc_40319_new_n3212_), .B(_abc_40319_new_n3216_), .Y(_abc_40319_new_n3217_));
AND2X2 AND2X2_132 ( .A(_abc_40319_new_n790_), .B(_abc_40319_new_n791_), .Y(_abc_40319_new_n792_));
AND2X2 AND2X2_1320 ( .A(_abc_40319_new_n3218_), .B(_abc_40319_new_n795_), .Y(_abc_40319_new_n3219_));
AND2X2 AND2X2_1321 ( .A(_abc_40319_new_n3220_), .B(_abc_40319_new_n784_), .Y(_abc_40319_new_n3221_));
AND2X2 AND2X2_1322 ( .A(_abc_40319_new_n2784_), .B(_abc_40319_new_n1735_), .Y(_abc_40319_new_n3224_));
AND2X2 AND2X2_1323 ( .A(_abc_40319_new_n2782_), .B(_abc_40319_new_n1724_), .Y(_abc_40319_new_n3225_));
AND2X2 AND2X2_1324 ( .A(_abc_40319_new_n3227_), .B(_abc_40319_new_n3223_), .Y(_abc_40319_new_n3228_));
AND2X2 AND2X2_1325 ( .A(_abc_40319_new_n2844_), .B(_abc_40319_new_n1410_), .Y(_abc_40319_new_n3229_));
AND2X2 AND2X2_1326 ( .A(_abc_40319_new_n2842_), .B(_abc_40319_new_n1398_), .Y(_abc_40319_new_n3230_));
AND2X2 AND2X2_1327 ( .A(_abc_40319_new_n2762_), .B(_abc_40319_new_n1701_), .Y(_abc_40319_new_n3233_));
AND2X2 AND2X2_1328 ( .A(_abc_40319_new_n2760_), .B(_abc_40319_new_n1690_), .Y(_abc_40319_new_n3234_));
AND2X2 AND2X2_1329 ( .A(_abc_40319_new_n3232_), .B(_abc_40319_new_n3236_), .Y(_abc_40319_new_n3237_));
AND2X2 AND2X2_133 ( .A(_abc_40319_new_n738_), .B(_abc_40319_new_n792_), .Y(_abc_40319_new_n793_));
AND2X2 AND2X2_1330 ( .A(_abc_40319_new_n3237_), .B(_abc_40319_new_n3228_), .Y(_abc_40319_new_n3238_));
AND2X2 AND2X2_1331 ( .A(_abc_40319_new_n3238_), .B(_abc_40319_new_n3217_), .Y(_abc_40319_new_n3239_));
AND2X2 AND2X2_1332 ( .A(_abc_40319_new_n3239_), .B(_abc_40319_new_n3208_), .Y(_abc_40319_new_n3240_));
AND2X2 AND2X2_1333 ( .A(_abc_40319_new_n3240_), .B(_abc_40319_new_n3204_), .Y(_abc_40319_new_n3241_));
AND2X2 AND2X2_1334 ( .A(_abc_40319_new_n3241_), .B(_abc_40319_new_n3200_), .Y(_abc_40319_new_n3242_));
AND2X2 AND2X2_1335 ( .A(_abc_40319_new_n3242_), .B(_abc_40319_new_n3196_), .Y(_abc_40319_new_n3243_));
AND2X2 AND2X2_1336 ( .A(_abc_40319_new_n3243_), .B(_abc_40319_new_n3192_), .Y(_abc_40319_new_n3244_));
AND2X2 AND2X2_1337 ( .A(_abc_40319_new_n3244_), .B(_abc_40319_new_n3107_), .Y(_abc_40319_new_n3245_));
AND2X2 AND2X2_1338 ( .A(_abc_40319_new_n3245_), .B(_abc_40319_new_n3103_), .Y(_abc_40319_new_n3246_));
AND2X2 AND2X2_1339 ( .A(_abc_40319_new_n1980_), .B(_abc_40319_new_n3042_), .Y(_abc_40319_new_n3247_));
AND2X2 AND2X2_134 ( .A(_abc_40319_new_n705_), .B(_abc_40319_new_n795_), .Y(_abc_40319_new_n796_));
AND2X2 AND2X2_1340 ( .A(_abc_40319_new_n3040_), .B(_abc_40319_new_n2089_), .Y(_abc_40319_new_n3248_));
AND2X2 AND2X2_1341 ( .A(_abc_40319_new_n1210_), .B(_abc_40319_new_n3025_), .Y(_abc_40319_new_n3251_));
AND2X2 AND2X2_1342 ( .A(_abc_40319_new_n3023_), .B(_abc_40319_new_n1180_), .Y(_abc_40319_new_n3252_));
AND2X2 AND2X2_1343 ( .A(_abc_40319_new_n1260_), .B(_abc_40319_new_n2992_), .Y(_abc_40319_new_n3255_));
AND2X2 AND2X2_1344 ( .A(_abc_40319_new_n2990_), .B(_abc_40319_new_n1249_), .Y(_abc_40319_new_n3256_));
AND2X2 AND2X2_1345 ( .A(_abc_40319_new_n2957_), .B(_abc_40319_new_n1306_), .Y(_abc_40319_new_n3259_));
AND2X2 AND2X2_1346 ( .A(_abc_40319_new_n1317_), .B(_abc_40319_new_n2959_), .Y(_abc_40319_new_n3260_));
AND2X2 AND2X2_1347 ( .A(_abc_40319_new_n3258_), .B(_abc_40319_new_n3262_), .Y(_abc_40319_new_n3263_));
AND2X2 AND2X2_1348 ( .A(_abc_40319_new_n3254_), .B(_abc_40319_new_n3263_), .Y(_abc_40319_new_n3264_));
AND2X2 AND2X2_1349 ( .A(_abc_40319_new_n3250_), .B(_abc_40319_new_n3264_), .Y(_abc_40319_new_n3265_));
AND2X2 AND2X2_135 ( .A(_abc_40319_new_n784_), .B(_abc_40319_new_n763_), .Y(_abc_40319_new_n798_));
AND2X2 AND2X2_1350 ( .A(_abc_40319_new_n3265_), .B(_abc_40319_new_n3246_), .Y(_abc_40319_new_n3266_));
AND2X2 AND2X2_1351 ( .A(_abc_40319_new_n3266_), .B(_abc_40319_new_n3098_), .Y(_abc_40319_new_n3267_));
AND2X2 AND2X2_1352 ( .A(_abc_40319_new_n3100_), .B(_abc_40319_new_n3171_), .Y(_abc_40319_new_n3269_));
AND2X2 AND2X2_1353 ( .A(_abc_40319_new_n3270_), .B(_abc_40319_new_n3161_), .Y(_abc_40319_new_n3271_));
AND2X2 AND2X2_1354 ( .A(_abc_40319_new_n3269_), .B(_abc_40319_new_n3271_), .Y(_abc_40319_new_n3272_));
AND2X2 AND2X2_1355 ( .A(_abc_40319_new_n3268_), .B(_abc_40319_new_n3272_), .Y(_abc_40319_new_n3273_));
AND2X2 AND2X2_1356 ( .A(_abc_40319_new_n3275_), .B(_abc_40319_new_n3276_), .Y(_abc_40319_new_n3277_));
AND2X2 AND2X2_1357 ( .A(_abc_40319_new_n3277_), .B(_abc_40319_new_n3197_), .Y(_abc_40319_new_n3278_));
AND2X2 AND2X2_1358 ( .A(_abc_40319_new_n3275_), .B(_abc_40319_new_n3260_), .Y(_abc_40319_new_n3280_));
AND2X2 AND2X2_1359 ( .A(_abc_40319_new_n3284_), .B(_abc_40319_new_n3279_), .Y(_abc_40319_new_n3285_));
AND2X2 AND2X2_136 ( .A(_abc_40319_new_n795_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n799_));
AND2X2 AND2X2_1360 ( .A(_abc_40319_new_n1852_), .B(_abc_40319_new_n2910_), .Y(_abc_40319_new_n3287_));
AND2X2 AND2X2_1361 ( .A(_abc_40319_new_n3288_), .B(_abc_40319_new_n3286_), .Y(_abc_40319_new_n3289_));
AND2X2 AND2X2_1362 ( .A(_abc_40319_new_n3291_), .B(_abc_40319_new_n3292_), .Y(_abc_40319_new_n3293_));
AND2X2 AND2X2_1363 ( .A(_abc_40319_new_n3295_), .B(_abc_40319_new_n3183_), .Y(_abc_40319_new_n3296_));
AND2X2 AND2X2_1364 ( .A(_abc_40319_new_n3298_), .B(_abc_40319_new_n3290_), .Y(_abc_40319_new_n3299_));
AND2X2 AND2X2_1365 ( .A(_abc_40319_new_n3299_), .B(_abc_40319_new_n3112_), .Y(_abc_40319_new_n3300_));
AND2X2 AND2X2_1366 ( .A(_abc_40319_new_n3301_), .B(_abc_40319_new_n3289_), .Y(_abc_40319_new_n3302_));
AND2X2 AND2X2_1367 ( .A(_abc_40319_new_n3303_), .B(_abc_40319_new_n3304_), .Y(_abc_40319_new_n3305_));
AND2X2 AND2X2_1368 ( .A(_abc_40319_new_n3299_), .B(_abc_40319_new_n3289_), .Y(_abc_40319_new_n3306_));
AND2X2 AND2X2_1369 ( .A(_abc_40319_new_n3307_), .B(_abc_40319_new_n3308_), .Y(_abc_40319_new_n3309_));
AND2X2 AND2X2_137 ( .A(_abc_40319_new_n803_), .B(_abc_40319_new_n801_), .Y(_abc_40319_new_n804_));
AND2X2 AND2X2_1370 ( .A(_abc_40319_new_n3306_), .B(_abc_40319_new_n3309_), .Y(_abc_40319_new_n3310_));
AND2X2 AND2X2_1371 ( .A(_abc_40319_new_n3310_), .B(_abc_40319_new_n3305_), .Y(_abc_40319_new_n3311_));
AND2X2 AND2X2_1372 ( .A(_abc_40319_new_n3314_), .B(_abc_40319_new_n3312_), .Y(_abc_40319_new_n3315_));
AND2X2 AND2X2_1373 ( .A(_abc_40319_new_n3317_), .B(_abc_40319_new_n3318_), .Y(_abc_40319_new_n3319_));
AND2X2 AND2X2_1374 ( .A(_abc_40319_new_n3319_), .B(_abc_40319_new_n3316_), .Y(_abc_40319_new_n3320_));
AND2X2 AND2X2_1375 ( .A(_abc_40319_new_n3315_), .B(_abc_40319_new_n3320_), .Y(_abc_40319_new_n3321_));
AND2X2 AND2X2_1376 ( .A(_abc_40319_new_n3311_), .B(_abc_40319_new_n3321_), .Y(_abc_40319_new_n3322_));
AND2X2 AND2X2_1377 ( .A(_abc_40319_new_n3322_), .B(_abc_40319_new_n3214_), .Y(_abc_40319_new_n3323_));
AND2X2 AND2X2_1378 ( .A(_abc_40319_new_n3324_), .B(_abc_40319_new_n3285_), .Y(_abc_40319_new_n3325_));
AND2X2 AND2X2_1379 ( .A(_abc_40319_new_n3311_), .B(_abc_40319_new_n3279_), .Y(_abc_40319_new_n3327_));
AND2X2 AND2X2_138 ( .A(_abc_40319_new_n805_), .B(_abc_40319_new_n797_), .Y(_abc_40319_new_n806_));
AND2X2 AND2X2_1380 ( .A(_abc_40319_new_n3321_), .B(_abc_40319_new_n3328_), .Y(_abc_40319_new_n3329_));
AND2X2 AND2X2_1381 ( .A(_abc_40319_new_n3284_), .B(_abc_40319_new_n3329_), .Y(_abc_40319_new_n3330_));
AND2X2 AND2X2_1382 ( .A(_abc_40319_new_n3327_), .B(_abc_40319_new_n3330_), .Y(_abc_40319_new_n3331_));
AND2X2 AND2X2_1383 ( .A(_abc_40319_new_n3331_), .B(_abc_40319_new_n3333_), .Y(_abc_40319_new_n3334_));
AND2X2 AND2X2_1384 ( .A(_abc_40319_new_n3337_), .B(_abc_40319_new_n3336_), .Y(_abc_40319_new_n3338_));
AND2X2 AND2X2_1385 ( .A(_abc_40319_new_n3338_), .B(_abc_40319_new_n3335_), .Y(_abc_40319_new_n3339_));
AND2X2 AND2X2_1386 ( .A(_abc_40319_new_n3339_), .B(_abc_40319_new_n3117_), .Y(_abc_40319_new_n3340_));
AND2X2 AND2X2_1387 ( .A(_abc_40319_new_n3334_), .B(_abc_40319_new_n3340_), .Y(_abc_40319_new_n3341_));
AND2X2 AND2X2_1388 ( .A(_abc_40319_new_n3333_), .B(_abc_40319_new_n3345_), .Y(_abc_40319_new_n3346_));
AND2X2 AND2X2_1389 ( .A(_abc_40319_new_n3346_), .B(_abc_40319_new_n3343_), .Y(_abc_40319_new_n3347_));
AND2X2 AND2X2_139 ( .A(_abc_40319_new_n674_), .B(IR_REG_3_), .Y(_abc_40319_new_n808_));
AND2X2 AND2X2_1390 ( .A(_abc_40319_new_n3347_), .B(_abc_40319_new_n3339_), .Y(_abc_40319_new_n3348_));
AND2X2 AND2X2_1391 ( .A(_abc_40319_new_n3311_), .B(_abc_40319_new_n3349_), .Y(_abc_40319_new_n3350_));
AND2X2 AND2X2_1392 ( .A(_abc_40319_new_n3350_), .B(_abc_40319_new_n3348_), .Y(_abc_40319_new_n3351_));
AND2X2 AND2X2_1393 ( .A(_abc_40319_new_n3351_), .B(_abc_40319_new_n3330_), .Y(_abc_40319_new_n3352_));
AND2X2 AND2X2_1394 ( .A(_abc_40319_new_n3304_), .B(_abc_40319_new_n3234_), .Y(_abc_40319_new_n3355_));
AND2X2 AND2X2_1395 ( .A(_abc_40319_new_n3285_), .B(_abc_40319_new_n3355_), .Y(_abc_40319_new_n3356_));
AND2X2 AND2X2_1396 ( .A(_abc_40319_new_n3356_), .B(_abc_40319_new_n3310_), .Y(_abc_40319_new_n3357_));
AND2X2 AND2X2_1397 ( .A(_abc_40319_new_n3284_), .B(_abc_40319_new_n3315_), .Y(_abc_40319_new_n3358_));
AND2X2 AND2X2_1398 ( .A(_abc_40319_new_n3327_), .B(_abc_40319_new_n3358_), .Y(_abc_40319_new_n3359_));
AND2X2 AND2X2_1399 ( .A(_abc_40319_new_n3359_), .B(_abc_40319_new_n3156_), .Y(_abc_40319_new_n3360_));
AND2X2 AND2X2_14 ( .A(_abc_40319_new_n557_), .B(_abc_40319_new_n558_), .Y(_abc_40319_new_n559_));
AND2X2 AND2X2_140 ( .A(_abc_40319_new_n810_), .B(IR_REG_31_), .Y(_abc_40319_new_n811_));
AND2X2 AND2X2_1400 ( .A(_abc_40319_new_n3310_), .B(_abc_40319_new_n3141_), .Y(_abc_40319_new_n3361_));
AND2X2 AND2X2_1401 ( .A(_abc_40319_new_n3285_), .B(_abc_40319_new_n3361_), .Y(_abc_40319_new_n3362_));
AND2X2 AND2X2_1402 ( .A(_abc_40319_new_n2908_), .B(_abc_40319_new_n1841_), .Y(_abc_40319_new_n3366_));
AND2X2 AND2X2_1403 ( .A(_abc_40319_new_n3298_), .B(_abc_40319_new_n3230_), .Y(_abc_40319_new_n3367_));
AND2X2 AND2X2_1404 ( .A(_abc_40319_new_n3368_), .B(_abc_40319_new_n3289_), .Y(_abc_40319_new_n3369_));
AND2X2 AND2X2_1405 ( .A(_abc_40319_new_n3307_), .B(_abc_40319_new_n3145_), .Y(_abc_40319_new_n3370_));
AND2X2 AND2X2_1406 ( .A(_abc_40319_new_n3306_), .B(_abc_40319_new_n3370_), .Y(_abc_40319_new_n3371_));
AND2X2 AND2X2_1407 ( .A(_abc_40319_new_n3285_), .B(_abc_40319_new_n3372_), .Y(_abc_40319_new_n3373_));
AND2X2 AND2X2_1408 ( .A(_abc_40319_new_n3319_), .B(_abc_40319_new_n3210_), .Y(_abc_40319_new_n3375_));
AND2X2 AND2X2_1409 ( .A(_abc_40319_new_n3359_), .B(_abc_40319_new_n3375_), .Y(_abc_40319_new_n3376_));
AND2X2 AND2X2_141 ( .A(_abc_40319_new_n524_), .B(IR_REG_3_), .Y(_abc_40319_new_n812_));
AND2X2 AND2X2_1410 ( .A(_abc_40319_new_n3378_), .B(_abc_40319_new_n3379_), .Y(_abc_40319_new_n3380_));
AND2X2 AND2X2_1411 ( .A(_abc_40319_new_n3314_), .B(_abc_40319_new_n3206_), .Y(_abc_40319_new_n3382_));
AND2X2 AND2X2_1412 ( .A(_abc_40319_new_n3327_), .B(_abc_40319_new_n3382_), .Y(_abc_40319_new_n3383_));
AND2X2 AND2X2_1413 ( .A(_abc_40319_new_n3383_), .B(_abc_40319_new_n3284_), .Y(_abc_40319_new_n3384_));
AND2X2 AND2X2_1414 ( .A(_abc_40319_new_n3385_), .B(_abc_40319_new_n3381_), .Y(_abc_40319_new_n3386_));
AND2X2 AND2X2_1415 ( .A(_abc_40319_new_n3327_), .B(_abc_40319_new_n3225_), .Y(_abc_40319_new_n3387_));
AND2X2 AND2X2_1416 ( .A(_abc_40319_new_n3387_), .B(_abc_40319_new_n3284_), .Y(_abc_40319_new_n3388_));
AND2X2 AND2X2_1417 ( .A(_abc_40319_new_n3386_), .B(_abc_40319_new_n3389_), .Y(_abc_40319_new_n3390_));
AND2X2 AND2X2_1418 ( .A(_abc_40319_new_n3390_), .B(_abc_40319_new_n3377_), .Y(_abc_40319_new_n3391_));
AND2X2 AND2X2_1419 ( .A(_abc_40319_new_n3391_), .B(_abc_40319_new_n3374_), .Y(_abc_40319_new_n3392_));
AND2X2 AND2X2_142 ( .A(_abc_40319_new_n640_), .B(_abc_40319_new_n814_), .Y(_abc_40319_new_n815_));
AND2X2 AND2X2_1420 ( .A(_abc_40319_new_n3392_), .B(_abc_40319_new_n3365_), .Y(_abc_40319_new_n3393_));
AND2X2 AND2X2_1421 ( .A(_abc_40319_new_n3393_), .B(_abc_40319_new_n3354_), .Y(_abc_40319_new_n3394_));
AND2X2 AND2X2_1422 ( .A(_abc_40319_new_n3394_), .B(_abc_40319_new_n3326_), .Y(_abc_40319_new_n3395_));
AND2X2 AND2X2_1423 ( .A(_abc_40319_new_n3399_), .B(_abc_40319_new_n3398_), .Y(_abc_40319_new_n3400_));
AND2X2 AND2X2_1424 ( .A(_abc_40319_new_n3295_), .B(_abc_40319_new_n3402_), .Y(_abc_40319_new_n3403_));
AND2X2 AND2X2_1425 ( .A(_abc_40319_new_n3405_), .B(_abc_40319_new_n3400_), .Y(_abc_40319_new_n3406_));
AND2X2 AND2X2_1426 ( .A(_abc_40319_new_n3406_), .B(_abc_40319_new_n3277_), .Y(_abc_40319_new_n3407_));
AND2X2 AND2X2_1427 ( .A(_abc_40319_new_n3408_), .B(_abc_40319_new_n3270_), .Y(_abc_40319_new_n3409_));
AND2X2 AND2X2_1428 ( .A(_abc_40319_new_n3285_), .B(_abc_40319_new_n3409_), .Y(_abc_40319_new_n3410_));
AND2X2 AND2X2_1429 ( .A(_abc_40319_new_n3411_), .B(_abc_40319_new_n3268_), .Y(_abc_40319_new_n3412_));
AND2X2 AND2X2_143 ( .A(_abc_40319_new_n817_), .B(_abc_40319_new_n816_), .Y(_abc_40319_new_n818_));
AND2X2 AND2X2_1430 ( .A(_abc_40319_new_n3413_), .B(_abc_40319_new_n3269_), .Y(_abc_40319_new_n3414_));
AND2X2 AND2X2_1431 ( .A(_abc_40319_new_n3415_), .B(_abc_40319_new_n3161_), .Y(_abc_40319_new_n3416_));
AND2X2 AND2X2_1432 ( .A(_abc_40319_new_n3273_), .B(_abc_40319_new_n3221_), .Y(_abc_40319_new_n3417_));
AND2X2 AND2X2_1433 ( .A(_abc_40319_new_n3268_), .B(_abc_40319_new_n3335_), .Y(_abc_40319_new_n3418_));
AND2X2 AND2X2_1434 ( .A(_abc_40319_new_n3272_), .B(_abc_40319_new_n3336_), .Y(_abc_40319_new_n3419_));
AND2X2 AND2X2_1435 ( .A(_abc_40319_new_n3419_), .B(_abc_40319_new_n3126_), .Y(_abc_40319_new_n3420_));
AND2X2 AND2X2_1436 ( .A(_abc_40319_new_n3418_), .B(_abc_40319_new_n3420_), .Y(_abc_40319_new_n3421_));
AND2X2 AND2X2_1437 ( .A(_abc_40319_new_n3422_), .B(_abc_40319_new_n3334_), .Y(_abc_40319_new_n3423_));
AND2X2 AND2X2_1438 ( .A(_abc_40319_new_n3418_), .B(_abc_40319_new_n3131_), .Y(_abc_40319_new_n3424_));
AND2X2 AND2X2_1439 ( .A(_abc_40319_new_n3424_), .B(_abc_40319_new_n3272_), .Y(_abc_40319_new_n3425_));
AND2X2 AND2X2_144 ( .A(_abc_40319_new_n820_), .B(_abc_40319_new_n763_), .Y(_abc_40319_new_n821_));
AND2X2 AND2X2_1440 ( .A(_abc_40319_new_n3425_), .B(_abc_40319_new_n3334_), .Y(_abc_40319_new_n3426_));
AND2X2 AND2X2_1441 ( .A(_abc_40319_new_n3268_), .B(_abc_40319_new_n3317_), .Y(_abc_40319_new_n3428_));
AND2X2 AND2X2_1442 ( .A(_abc_40319_new_n3428_), .B(_abc_40319_new_n3272_), .Y(_abc_40319_new_n3429_));
AND2X2 AND2X2_1443 ( .A(_abc_40319_new_n3429_), .B(_abc_40319_new_n3359_), .Y(_abc_40319_new_n3430_));
AND2X2 AND2X2_1444 ( .A(_abc_40319_new_n3430_), .B(_abc_40319_new_n3175_), .Y(_abc_40319_new_n3431_));
AND2X2 AND2X2_1445 ( .A(_abc_40319_new_n3329_), .B(_abc_40319_new_n3122_), .Y(_abc_40319_new_n3432_));
AND2X2 AND2X2_1446 ( .A(_abc_40319_new_n3327_), .B(_abc_40319_new_n3432_), .Y(_abc_40319_new_n3433_));
AND2X2 AND2X2_1447 ( .A(_abc_40319_new_n3433_), .B(_abc_40319_new_n3284_), .Y(_abc_40319_new_n3434_));
AND2X2 AND2X2_1448 ( .A(_abc_40319_new_n3273_), .B(_abc_40319_new_n3434_), .Y(_abc_40319_new_n3435_));
AND2X2 AND2X2_1449 ( .A(_abc_40319_new_n3396_), .B(_abc_40319_new_n3440_), .Y(_abc_40319_new_n3441_));
AND2X2 AND2X2_145 ( .A(_abc_40319_new_n722_), .B(REG1_REG_3_), .Y(_abc_40319_new_n822_));
AND2X2 AND2X2_1450 ( .A(_abc_40319_new_n3443_), .B(_abc_40319_new_n671_), .Y(_abc_40319_new_n3444_));
AND2X2 AND2X2_1451 ( .A(_abc_40319_new_n3095_), .B(_abc_40319_new_n3444_), .Y(_abc_40319_new_n3445_));
AND2X2 AND2X2_1452 ( .A(_abc_40319_new_n3447_), .B(_abc_40319_new_n698_), .Y(_abc_40319_new_n3448_));
AND2X2 AND2X2_1453 ( .A(_abc_40319_new_n3094_), .B(_abc_40319_new_n1168_), .Y(_abc_40319_new_n3449_));
AND2X2 AND2X2_1454 ( .A(_abc_40319_new_n655_), .B(_abc_40319_new_n697_), .Y(_abc_40319_new_n3450_));
AND2X2 AND2X2_1455 ( .A(_abc_40319_new_n3450_), .B(_abc_40319_new_n671_), .Y(_abc_40319_new_n3451_));
AND2X2 AND2X2_1456 ( .A(_abc_40319_new_n646_), .B(_abc_40319_new_n697_), .Y(_abc_40319_new_n3452_));
AND2X2 AND2X2_1457 ( .A(_abc_40319_new_n3452_), .B(_abc_40319_new_n671_), .Y(_abc_40319_new_n3453_));
AND2X2 AND2X2_1458 ( .A(_abc_40319_new_n3441_), .B(_abc_40319_new_n3454_), .Y(_abc_40319_new_n3455_));
AND2X2 AND2X2_1459 ( .A(_abc_40319_new_n754_), .B(_abc_40319_new_n698_), .Y(_abc_40319_new_n3456_));
AND2X2 AND2X2_146 ( .A(_abc_40319_new_n733_), .B(REG2_REG_3_), .Y(_abc_40319_new_n823_));
AND2X2 AND2X2_1460 ( .A(_abc_40319_new_n3456_), .B(_abc_40319_new_n645_), .Y(_abc_40319_new_n3457_));
AND2X2 AND2X2_1461 ( .A(_abc_40319_new_n3458_), .B(_abc_40319_new_n3164_), .Y(_abc_40319_new_n3459_));
AND2X2 AND2X2_1462 ( .A(_abc_40319_new_n3099_), .B(_abc_40319_new_n3459_), .Y(_abc_40319_new_n3460_));
AND2X2 AND2X2_1463 ( .A(_abc_40319_new_n3170_), .B(_abc_40319_new_n2553_), .Y(_abc_40319_new_n3461_));
AND2X2 AND2X2_1464 ( .A(_abc_40319_new_n3102_), .B(_abc_40319_new_n3459_), .Y(_abc_40319_new_n3464_));
AND2X2 AND2X2_1465 ( .A(_abc_40319_new_n3270_), .B(_abc_40319_new_n3466_), .Y(_abc_40319_new_n3467_));
AND2X2 AND2X2_1466 ( .A(_abc_40319_new_n3277_), .B(_abc_40319_new_n3469_), .Y(_abc_40319_new_n3470_));
AND2X2 AND2X2_1467 ( .A(_abc_40319_new_n3473_), .B(_abc_40319_new_n3472_), .Y(_abc_40319_new_n3474_));
AND2X2 AND2X2_1468 ( .A(_abc_40319_new_n3477_), .B(_abc_40319_new_n3478_), .Y(_abc_40319_new_n3479_));
AND2X2 AND2X2_1469 ( .A(_abc_40319_new_n3479_), .B(_abc_40319_new_n3476_), .Y(_abc_40319_new_n3480_));
AND2X2 AND2X2_147 ( .A(_abc_40319_new_n736_), .B(REG0_REG_3_), .Y(_abc_40319_new_n825_));
AND2X2 AND2X2_1470 ( .A(_abc_40319_new_n3313_), .B(_abc_40319_new_n3312_), .Y(_abc_40319_new_n3482_));
AND2X2 AND2X2_1471 ( .A(_abc_40319_new_n3483_), .B(_abc_40319_new_n3484_), .Y(_abc_40319_new_n3485_));
AND2X2 AND2X2_1472 ( .A(_abc_40319_new_n3485_), .B(_abc_40319_new_n3155_), .Y(_abc_40319_new_n3486_));
AND2X2 AND2X2_1473 ( .A(_abc_40319_new_n3487_), .B(_abc_40319_new_n3482_), .Y(_abc_40319_new_n3488_));
AND2X2 AND2X2_1474 ( .A(_abc_40319_new_n3490_), .B(_abc_40319_new_n3115_), .Y(_abc_40319_new_n3491_));
AND2X2 AND2X2_1475 ( .A(_abc_40319_new_n3492_), .B(_abc_40319_new_n3337_), .Y(_abc_40319_new_n3493_));
AND2X2 AND2X2_1476 ( .A(_abc_40319_new_n3493_), .B(_abc_40319_new_n3336_), .Y(_abc_40319_new_n3494_));
AND2X2 AND2X2_1477 ( .A(_abc_40319_new_n3498_), .B(_abc_40319_new_n3496_), .Y(_abc_40319_new_n3499_));
AND2X2 AND2X2_1478 ( .A(_abc_40319_new_n3335_), .B(_abc_40319_new_n3332_), .Y(_abc_40319_new_n3502_));
AND2X2 AND2X2_1479 ( .A(_abc_40319_new_n3503_), .B(_abc_40319_new_n3328_), .Y(_abc_40319_new_n3504_));
AND2X2 AND2X2_148 ( .A(_abc_40319_new_n738_), .B(_abc_40319_new_n826_), .Y(_abc_40319_new_n827_));
AND2X2 AND2X2_1480 ( .A(_abc_40319_new_n3501_), .B(_abc_40319_new_n3504_), .Y(_abc_40319_new_n3505_));
AND2X2 AND2X2_1481 ( .A(_abc_40319_new_n3316_), .B(_abc_40319_new_n3318_), .Y(_abc_40319_new_n3507_));
AND2X2 AND2X2_1482 ( .A(_abc_40319_new_n3506_), .B(_abc_40319_new_n3507_), .Y(_abc_40319_new_n3508_));
AND2X2 AND2X2_1483 ( .A(_abc_40319_new_n3485_), .B(_abc_40319_new_n3510_), .Y(_abc_40319_new_n3511_));
AND2X2 AND2X2_1484 ( .A(_abc_40319_new_n3513_), .B(_abc_40319_new_n3489_), .Y(_abc_40319_new_n3514_));
AND2X2 AND2X2_1485 ( .A(_abc_40319_new_n3515_), .B(_abc_40319_new_n3303_), .Y(_abc_40319_new_n3516_));
AND2X2 AND2X2_1486 ( .A(_abc_40319_new_n3517_), .B(_abc_40319_new_n3304_), .Y(_abc_40319_new_n3518_));
AND2X2 AND2X2_1487 ( .A(_abc_40319_new_n3479_), .B(_abc_40319_new_n3144_), .Y(_abc_40319_new_n3520_));
AND2X2 AND2X2_1488 ( .A(_abc_40319_new_n3522_), .B(_abc_40319_new_n3290_), .Y(_abc_40319_new_n3523_));
AND2X2 AND2X2_1489 ( .A(_abc_40319_new_n3521_), .B(_abc_40319_new_n3523_), .Y(_abc_40319_new_n3524_));
AND2X2 AND2X2_149 ( .A(_abc_40319_new_n829_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n830_));
AND2X2 AND2X2_1490 ( .A(_abc_40319_new_n3527_), .B(_abc_40319_new_n3293_), .Y(_abc_40319_new_n3528_));
AND2X2 AND2X2_1491 ( .A(_abc_40319_new_n3519_), .B(_abc_40319_new_n3528_), .Y(_abc_40319_new_n3529_));
AND2X2 AND2X2_1492 ( .A(_abc_40319_new_n3530_), .B(_abc_40319_new_n3289_), .Y(_abc_40319_new_n3531_));
AND2X2 AND2X2_1493 ( .A(_abc_40319_new_n3532_), .B(_abc_40319_new_n3471_), .Y(_abc_40319_new_n3533_));
AND2X2 AND2X2_1494 ( .A(_abc_40319_new_n3535_), .B(_abc_40319_new_n3380_), .Y(_abc_40319_new_n3536_));
AND2X2 AND2X2_1495 ( .A(_abc_40319_new_n3537_), .B(_abc_40319_new_n3465_), .Y(_abc_40319_new_n3538_));
AND2X2 AND2X2_1496 ( .A(_abc_40319_new_n3539_), .B(_abc_40319_new_n3464_), .Y(_abc_40319_new_n3540_));
AND2X2 AND2X2_1497 ( .A(_abc_40319_new_n3542_), .B(_abc_40319_new_n3457_), .Y(_abc_40319_new_n3543_));
AND2X2 AND2X2_1498 ( .A(_abc_40319_new_n3098_), .B(_abc_40319_new_n697_), .Y(_abc_40319_new_n3545_));
AND2X2 AND2X2_1499 ( .A(_abc_40319_new_n3544_), .B(_abc_40319_new_n3545_), .Y(_abc_40319_new_n3546_));
AND2X2 AND2X2_15 ( .A(_abc_40319_new_n559_), .B(_abc_40319_new_n556_), .Y(_abc_40319_new_n560_));
AND2X2 AND2X2_150 ( .A(_abc_40319_new_n832_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n833_));
AND2X2 AND2X2_1500 ( .A(_abc_40319_new_n754_), .B(_abc_40319_new_n697_), .Y(_abc_40319_new_n3547_));
AND2X2 AND2X2_1501 ( .A(_abc_40319_new_n3541_), .B(_abc_40319_new_n3547_), .Y(_abc_40319_new_n3548_));
AND2X2 AND2X2_1502 ( .A(_abc_40319_new_n3553_), .B(_abc_40319_new_n2550_), .Y(_abc_40319_new_n3554_));
AND2X2 AND2X2_1503 ( .A(_abc_40319_new_n628_), .B(_abc_40319_new_n638_), .Y(_abc_40319_new_n3555_));
AND2X2 AND2X2_1504 ( .A(_abc_40319_new_n1132_), .B(_abc_40319_new_n3555_), .Y(_abc_40319_new_n3556_));
AND2X2 AND2X2_1505 ( .A(_abc_40319_new_n3557_), .B(_abc_40319_new_n613_), .Y(_abc_40319_new_n3558_));
AND2X2 AND2X2_1506 ( .A(_abc_40319_new_n2549_), .B(_abc_40319_new_n646_), .Y(_abc_40319_new_n3559_));
AND2X2 AND2X2_1507 ( .A(_abc_40319_new_n3562_), .B(B_REG), .Y(_abc_40319_new_n3563_));
AND2X2 AND2X2_1508 ( .A(IR_REG_0_), .B(REG1_REG_0_), .Y(_abc_40319_new_n3567_));
AND2X2 AND2X2_1509 ( .A(_abc_40319_new_n3568_), .B(_abc_40319_new_n3566_), .Y(_abc_40319_new_n3569_));
AND2X2 AND2X2_151 ( .A(_abc_40319_new_n831_), .B(_abc_40319_new_n768_), .Y(_abc_40319_new_n834_));
AND2X2 AND2X2_1510 ( .A(_abc_40319_new_n629_), .B(_abc_40319_new_n3569_), .Y(_abc_40319_new_n3570_));
AND2X2 AND2X2_1511 ( .A(_abc_40319_new_n639_), .B(IR_REG_0_), .Y(_abc_40319_new_n3571_));
AND2X2 AND2X2_1512 ( .A(IR_REG_0_), .B(REG2_REG_0_), .Y(_abc_40319_new_n3573_));
AND2X2 AND2X2_1513 ( .A(_abc_40319_new_n3574_), .B(_abc_40319_new_n3572_), .Y(_abc_40319_new_n3575_));
AND2X2 AND2X2_1514 ( .A(_abc_40319_new_n3555_), .B(_abc_40319_new_n3575_), .Y(_abc_40319_new_n3576_));
AND2X2 AND2X2_1515 ( .A(n1341), .B(_abc_40319_new_n2550_), .Y(_abc_40319_new_n3579_));
AND2X2 AND2X2_1516 ( .A(n1341), .B(_abc_40319_new_n1120_), .Y(_abc_40319_new_n3580_));
AND2X2 AND2X2_1517 ( .A(_abc_40319_new_n3581_), .B(_abc_40319_new_n3578_), .Y(_abc_40319_new_n3582_));
AND2X2 AND2X2_1518 ( .A(_abc_40319_new_n3585_), .B(ADDR_REG_0_), .Y(_abc_40319_new_n3586_));
AND2X2 AND2X2_1519 ( .A(_abc_40319_new_n3574_), .B(_abc_40319_new_n3589_), .Y(_abc_40319_new_n3590_));
AND2X2 AND2X2_152 ( .A(_abc_40319_new_n820_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n836_));
AND2X2 AND2X2_1520 ( .A(_abc_40319_new_n3573_), .B(REG2_REG_1_), .Y(_abc_40319_new_n3592_));
AND2X2 AND2X2_1521 ( .A(_abc_40319_new_n3591_), .B(_abc_40319_new_n3593_), .Y(_abc_40319_new_n3594_));
AND2X2 AND2X2_1522 ( .A(_abc_40319_new_n3598_), .B(_abc_40319_new_n3595_), .Y(_abc_40319_new_n3599_));
AND2X2 AND2X2_1523 ( .A(_abc_40319_new_n3555_), .B(_abc_40319_new_n3599_), .Y(_abc_40319_new_n3600_));
AND2X2 AND2X2_1524 ( .A(_abc_40319_new_n3567_), .B(REG1_REG_1_), .Y(_abc_40319_new_n3601_));
AND2X2 AND2X2_1525 ( .A(_abc_40319_new_n3568_), .B(_abc_40319_new_n3603_), .Y(_abc_40319_new_n3604_));
AND2X2 AND2X2_1526 ( .A(_abc_40319_new_n3605_), .B(_abc_40319_new_n3602_), .Y(_abc_40319_new_n3606_));
AND2X2 AND2X2_1527 ( .A(_abc_40319_new_n3609_), .B(_abc_40319_new_n3607_), .Y(_abc_40319_new_n3610_));
AND2X2 AND2X2_1528 ( .A(_abc_40319_new_n629_), .B(_abc_40319_new_n3610_), .Y(_abc_40319_new_n3611_));
AND2X2 AND2X2_1529 ( .A(_abc_40319_new_n639_), .B(_abc_40319_new_n886_), .Y(_abc_40319_new_n3612_));
AND2X2 AND2X2_153 ( .A(_abc_40319_new_n705_), .B(_abc_40319_new_n829_), .Y(_abc_40319_new_n837_));
AND2X2 AND2X2_1530 ( .A(_abc_40319_new_n3581_), .B(_abc_40319_new_n3614_), .Y(_abc_40319_new_n3615_));
AND2X2 AND2X2_1531 ( .A(_abc_40319_new_n3585_), .B(ADDR_REG_1_), .Y(_abc_40319_new_n3616_));
AND2X2 AND2X2_1532 ( .A(_abc_40319_new_n629_), .B(_abc_40319_new_n638_), .Y(_abc_40319_new_n3619_));
AND2X2 AND2X2_1533 ( .A(_abc_40319_new_n2361_), .B(_abc_40319_new_n3619_), .Y(_abc_40319_new_n3620_));
AND2X2 AND2X2_1534 ( .A(_abc_40319_new_n3621_), .B(n1345), .Y(_abc_40319_new_n3622_));
AND2X2 AND2X2_1535 ( .A(_abc_40319_new_n3585_), .B(ADDR_REG_2_), .Y(_abc_40319_new_n3623_));
AND2X2 AND2X2_1536 ( .A(_abc_40319_new_n3625_), .B(REG2_REG_2_), .Y(_abc_40319_new_n3626_));
AND2X2 AND2X2_1537 ( .A(_abc_40319_new_n843_), .B(_abc_40319_new_n860_), .Y(_abc_40319_new_n3628_));
AND2X2 AND2X2_1538 ( .A(_abc_40319_new_n3627_), .B(_abc_40319_new_n3629_), .Y(_abc_40319_new_n3630_));
AND2X2 AND2X2_1539 ( .A(_abc_40319_new_n3596_), .B(_abc_40319_new_n3593_), .Y(_abc_40319_new_n3632_));
AND2X2 AND2X2_154 ( .A(_abc_40319_new_n529_), .B(IR_REG_31_), .Y(_abc_40319_new_n839_));
AND2X2 AND2X2_1540 ( .A(_abc_40319_new_n3634_), .B(_abc_40319_new_n3636_), .Y(_abc_40319_new_n3637_));
AND2X2 AND2X2_1541 ( .A(_abc_40319_new_n3555_), .B(_abc_40319_new_n3637_), .Y(_abc_40319_new_n3638_));
AND2X2 AND2X2_1542 ( .A(_abc_40319_new_n843_), .B(_abc_40319_new_n853_), .Y(_abc_40319_new_n3639_));
AND2X2 AND2X2_1543 ( .A(_abc_40319_new_n3625_), .B(REG1_REG_2_), .Y(_abc_40319_new_n3641_));
AND2X2 AND2X2_1544 ( .A(_abc_40319_new_n3642_), .B(_abc_40319_new_n3640_), .Y(_abc_40319_new_n3643_));
AND2X2 AND2X2_1545 ( .A(_abc_40319_new_n886_), .B(_abc_40319_new_n3605_), .Y(_abc_40319_new_n3645_));
AND2X2 AND2X2_1546 ( .A(_abc_40319_new_n3648_), .B(_abc_40319_new_n3649_), .Y(_abc_40319_new_n3650_));
AND2X2 AND2X2_1547 ( .A(_abc_40319_new_n629_), .B(_abc_40319_new_n3650_), .Y(_abc_40319_new_n3651_));
AND2X2 AND2X2_1548 ( .A(_abc_40319_new_n639_), .B(_abc_40319_new_n3625_), .Y(_abc_40319_new_n3652_));
AND2X2 AND2X2_1549 ( .A(_abc_40319_new_n3580_), .B(_abc_40319_new_n3654_), .Y(_abc_40319_new_n3655_));
AND2X2 AND2X2_155 ( .A(_abc_40319_new_n839_), .B(_abc_40319_new_n528_), .Y(_abc_40319_new_n841_));
AND2X2 AND2X2_1550 ( .A(_abc_40319_new_n3579_), .B(_abc_40319_new_n3654_), .Y(_abc_40319_new_n3656_));
AND2X2 AND2X2_1551 ( .A(_abc_40319_new_n813_), .B(REG2_REG_3_), .Y(_abc_40319_new_n3660_));
AND2X2 AND2X2_1552 ( .A(_abc_40319_new_n3635_), .B(_abc_40319_new_n3629_), .Y(_abc_40319_new_n3661_));
AND2X2 AND2X2_1553 ( .A(_abc_40319_new_n814_), .B(_abc_40319_new_n3663_), .Y(_abc_40319_new_n3664_));
AND2X2 AND2X2_1554 ( .A(_abc_40319_new_n3665_), .B(_abc_40319_new_n3662_), .Y(_abc_40319_new_n3666_));
AND2X2 AND2X2_1555 ( .A(_abc_40319_new_n3665_), .B(_abc_40319_new_n3669_), .Y(_abc_40319_new_n3670_));
AND2X2 AND2X2_1556 ( .A(_abc_40319_new_n3668_), .B(_abc_40319_new_n3671_), .Y(_abc_40319_new_n3672_));
AND2X2 AND2X2_1557 ( .A(_abc_40319_new_n3555_), .B(_abc_40319_new_n3672_), .Y(_abc_40319_new_n3673_));
AND2X2 AND2X2_1558 ( .A(_abc_40319_new_n3646_), .B(_abc_40319_new_n3640_), .Y(_abc_40319_new_n3675_));
AND2X2 AND2X2_1559 ( .A(_abc_40319_new_n3677_), .B(_abc_40319_new_n3674_), .Y(_abc_40319_new_n3678_));
AND2X2 AND2X2_156 ( .A(_abc_40319_new_n842_), .B(_abc_40319_new_n840_), .Y(_abc_40319_new_n843_));
AND2X2 AND2X2_1560 ( .A(_abc_40319_new_n3676_), .B(REG1_REG_3_), .Y(_abc_40319_new_n3680_));
AND2X2 AND2X2_1561 ( .A(_abc_40319_new_n3679_), .B(_abc_40319_new_n3681_), .Y(_abc_40319_new_n3682_));
AND2X2 AND2X2_1562 ( .A(_abc_40319_new_n3683_), .B(_abc_40319_new_n813_), .Y(_abc_40319_new_n3684_));
AND2X2 AND2X2_1563 ( .A(_abc_40319_new_n3682_), .B(_abc_40319_new_n814_), .Y(_abc_40319_new_n3685_));
AND2X2 AND2X2_1564 ( .A(_abc_40319_new_n629_), .B(_abc_40319_new_n3686_), .Y(_abc_40319_new_n3687_));
AND2X2 AND2X2_1565 ( .A(_abc_40319_new_n639_), .B(_abc_40319_new_n813_), .Y(_abc_40319_new_n3688_));
AND2X2 AND2X2_1566 ( .A(_abc_40319_new_n3581_), .B(_abc_40319_new_n3690_), .Y(_abc_40319_new_n3691_));
AND2X2 AND2X2_1567 ( .A(_abc_40319_new_n3585_), .B(ADDR_REG_3_), .Y(_abc_40319_new_n3692_));
AND2X2 AND2X2_1568 ( .A(_abc_40319_new_n3585_), .B(ADDR_REG_4_), .Y(_abc_40319_new_n3695_));
AND2X2 AND2X2_1569 ( .A(_abc_40319_new_n779_), .B(REG2_REG_4_), .Y(_abc_40319_new_n3696_));
AND2X2 AND2X2_157 ( .A(_abc_40319_new_n640_), .B(_abc_40319_new_n843_), .Y(_abc_40319_new_n844_));
AND2X2 AND2X2_1570 ( .A(_abc_40319_new_n780_), .B(_abc_40319_new_n3698_), .Y(_abc_40319_new_n3699_));
AND2X2 AND2X2_1571 ( .A(_abc_40319_new_n3700_), .B(_abc_40319_new_n3697_), .Y(_abc_40319_new_n3701_));
AND2X2 AND2X2_1572 ( .A(_abc_40319_new_n3667_), .B(_abc_40319_new_n3669_), .Y(_abc_40319_new_n3702_));
AND2X2 AND2X2_1573 ( .A(_abc_40319_new_n3703_), .B(_abc_40319_new_n3700_), .Y(_abc_40319_new_n3705_));
AND2X2 AND2X2_1574 ( .A(_abc_40319_new_n3707_), .B(_abc_40319_new_n3704_), .Y(_abc_40319_new_n3708_));
AND2X2 AND2X2_1575 ( .A(_abc_40319_new_n3708_), .B(_abc_40319_new_n3555_), .Y(_abc_40319_new_n3709_));
AND2X2 AND2X2_1576 ( .A(_abc_40319_new_n779_), .B(REG1_REG_4_), .Y(_abc_40319_new_n3710_));
AND2X2 AND2X2_1577 ( .A(_abc_40319_new_n3711_), .B(_abc_40319_new_n3681_), .Y(_abc_40319_new_n3712_));
AND2X2 AND2X2_1578 ( .A(_abc_40319_new_n780_), .B(_abc_40319_new_n3713_), .Y(_abc_40319_new_n3714_));
AND2X2 AND2X2_1579 ( .A(_abc_40319_new_n3719_), .B(_abc_40319_new_n3718_), .Y(_abc_40319_new_n3720_));
AND2X2 AND2X2_158 ( .A(_abc_40319_new_n817_), .B(_abc_40319_new_n845_), .Y(_abc_40319_new_n846_));
AND2X2 AND2X2_1580 ( .A(_abc_40319_new_n3716_), .B(_abc_40319_new_n3721_), .Y(_abc_40319_new_n3722_));
AND2X2 AND2X2_1581 ( .A(_abc_40319_new_n3722_), .B(_abc_40319_new_n629_), .Y(_abc_40319_new_n3723_));
AND2X2 AND2X2_1582 ( .A(_abc_40319_new_n639_), .B(_abc_40319_new_n779_), .Y(_abc_40319_new_n3724_));
AND2X2 AND2X2_1583 ( .A(_abc_40319_new_n3726_), .B(_abc_40319_new_n3580_), .Y(_abc_40319_new_n3727_));
AND2X2 AND2X2_1584 ( .A(_abc_40319_new_n3726_), .B(_abc_40319_new_n3579_), .Y(_abc_40319_new_n3729_));
AND2X2 AND2X2_1585 ( .A(_abc_40319_new_n3715_), .B(_abc_40319_new_n3718_), .Y(_abc_40319_new_n3733_));
AND2X2 AND2X2_1586 ( .A(_abc_40319_new_n3734_), .B(REG1_REG_5_), .Y(_abc_40319_new_n3735_));
AND2X2 AND2X2_1587 ( .A(_abc_40319_new_n3733_), .B(_abc_40319_new_n3737_), .Y(_abc_40319_new_n3738_));
AND2X2 AND2X2_1588 ( .A(_abc_40319_new_n3736_), .B(_abc_40319_new_n3739_), .Y(_abc_40319_new_n3740_));
AND2X2 AND2X2_1589 ( .A(_abc_40319_new_n3743_), .B(_abc_40319_new_n629_), .Y(_abc_40319_new_n3744_));
AND2X2 AND2X2_159 ( .A(_abc_40319_new_n848_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n849_));
AND2X2 AND2X2_1590 ( .A(_abc_40319_new_n3744_), .B(_abc_40319_new_n3742_), .Y(_abc_40319_new_n3745_));
AND2X2 AND2X2_1591 ( .A(_abc_40319_new_n3706_), .B(_abc_40319_new_n3697_), .Y(_abc_40319_new_n3746_));
AND2X2 AND2X2_1592 ( .A(_abc_40319_new_n685_), .B(_abc_40319_new_n3747_), .Y(_abc_40319_new_n3748_));
AND2X2 AND2X2_1593 ( .A(_abc_40319_new_n684_), .B(REG2_REG_5_), .Y(_abc_40319_new_n3750_));
AND2X2 AND2X2_1594 ( .A(_abc_40319_new_n3749_), .B(_abc_40319_new_n3751_), .Y(_abc_40319_new_n3752_));
AND2X2 AND2X2_1595 ( .A(_abc_40319_new_n3746_), .B(_abc_40319_new_n3752_), .Y(_abc_40319_new_n3753_));
AND2X2 AND2X2_1596 ( .A(_abc_40319_new_n3754_), .B(_abc_40319_new_n3755_), .Y(_abc_40319_new_n3756_));
AND2X2 AND2X2_1597 ( .A(_abc_40319_new_n3757_), .B(_abc_40319_new_n3555_), .Y(_abc_40319_new_n3758_));
AND2X2 AND2X2_1598 ( .A(_abc_40319_new_n639_), .B(_abc_40319_new_n684_), .Y(_abc_40319_new_n3759_));
AND2X2 AND2X2_1599 ( .A(_abc_40319_new_n3761_), .B(_abc_40319_new_n3581_), .Y(_abc_40319_new_n3762_));
AND2X2 AND2X2_16 ( .A(_abc_40319_new_n560_), .B(_abc_40319_new_n555_), .Y(_abc_40319_new_n561_));
AND2X2 AND2X2_160 ( .A(_abc_40319_new_n852_), .B(_abc_40319_new_n855_), .Y(_abc_40319_new_n856_));
AND2X2 AND2X2_1600 ( .A(_abc_40319_new_n3585_), .B(ADDR_REG_5_), .Y(_abc_40319_new_n3763_));
AND2X2 AND2X2_1601 ( .A(_abc_40319_new_n993_), .B(REG2_REG_6_), .Y(_abc_40319_new_n3766_));
AND2X2 AND2X2_1602 ( .A(_abc_40319_new_n3746_), .B(_abc_40319_new_n3751_), .Y(_abc_40319_new_n3767_));
AND2X2 AND2X2_1603 ( .A(_abc_40319_new_n3769_), .B(_abc_40319_new_n3770_), .Y(_abc_40319_new_n3771_));
AND2X2 AND2X2_1604 ( .A(_abc_40319_new_n3774_), .B(_abc_40319_new_n3770_), .Y(_abc_40319_new_n3775_));
AND2X2 AND2X2_1605 ( .A(_abc_40319_new_n3776_), .B(_abc_40319_new_n3555_), .Y(_abc_40319_new_n3777_));
AND2X2 AND2X2_1606 ( .A(_abc_40319_new_n3773_), .B(_abc_40319_new_n3777_), .Y(_abc_40319_new_n3778_));
AND2X2 AND2X2_1607 ( .A(_abc_40319_new_n993_), .B(REG1_REG_6_), .Y(_abc_40319_new_n3779_));
AND2X2 AND2X2_1608 ( .A(_abc_40319_new_n3736_), .B(_abc_40319_new_n3780_), .Y(_abc_40319_new_n3781_));
AND2X2 AND2X2_1609 ( .A(_abc_40319_new_n3787_), .B(_abc_40319_new_n3782_), .Y(_abc_40319_new_n3788_));
AND2X2 AND2X2_161 ( .A(_abc_40319_new_n862_), .B(_abc_40319_new_n859_), .Y(_abc_40319_new_n863_));
AND2X2 AND2X2_1610 ( .A(_abc_40319_new_n3789_), .B(_abc_40319_new_n629_), .Y(_abc_40319_new_n3790_));
AND2X2 AND2X2_1611 ( .A(_abc_40319_new_n3790_), .B(_abc_40319_new_n3785_), .Y(_abc_40319_new_n3791_));
AND2X2 AND2X2_1612 ( .A(_abc_40319_new_n639_), .B(_abc_40319_new_n993_), .Y(_abc_40319_new_n3792_));
AND2X2 AND2X2_1613 ( .A(_abc_40319_new_n3794_), .B(_abc_40319_new_n3581_), .Y(_abc_40319_new_n3795_));
AND2X2 AND2X2_1614 ( .A(_abc_40319_new_n3585_), .B(ADDR_REG_6_), .Y(_abc_40319_new_n3796_));
AND2X2 AND2X2_1615 ( .A(_abc_40319_new_n1029_), .B(REG2_REG_7_), .Y(_abc_40319_new_n3799_));
AND2X2 AND2X2_1616 ( .A(_abc_40319_new_n3772_), .B(_abc_40319_new_n3774_), .Y(_abc_40319_new_n3800_));
AND2X2 AND2X2_1617 ( .A(_abc_40319_new_n3801_), .B(_abc_40319_new_n3802_), .Y(_abc_40319_new_n3803_));
AND2X2 AND2X2_1618 ( .A(_abc_40319_new_n3806_), .B(_abc_40319_new_n3802_), .Y(_abc_40319_new_n3807_));
AND2X2 AND2X2_1619 ( .A(_abc_40319_new_n3808_), .B(_abc_40319_new_n3555_), .Y(_abc_40319_new_n3809_));
AND2X2 AND2X2_162 ( .A(_abc_40319_new_n856_), .B(_abc_40319_new_n863_), .Y(_abc_40319_new_n864_));
AND2X2 AND2X2_1620 ( .A(_abc_40319_new_n3805_), .B(_abc_40319_new_n3809_), .Y(_abc_40319_new_n3810_));
AND2X2 AND2X2_1621 ( .A(_abc_40319_new_n1029_), .B(REG1_REG_7_), .Y(_abc_40319_new_n3811_));
AND2X2 AND2X2_1622 ( .A(_abc_40319_new_n3784_), .B(_abc_40319_new_n3787_), .Y(_abc_40319_new_n3812_));
AND2X2 AND2X2_1623 ( .A(_abc_40319_new_n3818_), .B(_abc_40319_new_n3813_), .Y(_abc_40319_new_n3819_));
AND2X2 AND2X2_1624 ( .A(_abc_40319_new_n3820_), .B(_abc_40319_new_n629_), .Y(_abc_40319_new_n3821_));
AND2X2 AND2X2_1625 ( .A(_abc_40319_new_n3821_), .B(_abc_40319_new_n3816_), .Y(_abc_40319_new_n3822_));
AND2X2 AND2X2_1626 ( .A(_abc_40319_new_n639_), .B(_abc_40319_new_n1029_), .Y(_abc_40319_new_n3823_));
AND2X2 AND2X2_1627 ( .A(_abc_40319_new_n3825_), .B(_abc_40319_new_n3581_), .Y(_abc_40319_new_n3826_));
AND2X2 AND2X2_1628 ( .A(_abc_40319_new_n3585_), .B(ADDR_REG_7_), .Y(_abc_40319_new_n3827_));
AND2X2 AND2X2_1629 ( .A(_abc_40319_new_n639_), .B(_abc_40319_new_n1567_), .Y(_abc_40319_new_n3830_));
AND2X2 AND2X2_163 ( .A(_abc_40319_new_n705_), .B(_abc_40319_new_n865_), .Y(_abc_40319_new_n866_));
AND2X2 AND2X2_1630 ( .A(_abc_40319_new_n1567_), .B(REG2_REG_8_), .Y(_abc_40319_new_n3831_));
AND2X2 AND2X2_1631 ( .A(_abc_40319_new_n3804_), .B(_abc_40319_new_n3806_), .Y(_abc_40319_new_n3832_));
AND2X2 AND2X2_1632 ( .A(_abc_40319_new_n3833_), .B(_abc_40319_new_n3834_), .Y(_abc_40319_new_n3835_));
AND2X2 AND2X2_1633 ( .A(_abc_40319_new_n3838_), .B(_abc_40319_new_n3834_), .Y(_abc_40319_new_n3839_));
AND2X2 AND2X2_1634 ( .A(_abc_40319_new_n3840_), .B(_abc_40319_new_n3555_), .Y(_abc_40319_new_n3841_));
AND2X2 AND2X2_1635 ( .A(_abc_40319_new_n3837_), .B(_abc_40319_new_n3841_), .Y(_abc_40319_new_n3842_));
AND2X2 AND2X2_1636 ( .A(_abc_40319_new_n3815_), .B(_abc_40319_new_n3818_), .Y(_abc_40319_new_n3844_));
AND2X2 AND2X2_1637 ( .A(_abc_40319_new_n3844_), .B(_abc_40319_new_n3843_), .Y(_abc_40319_new_n3845_));
AND2X2 AND2X2_1638 ( .A(_abc_40319_new_n3848_), .B(_abc_40319_new_n1567_), .Y(_abc_40319_new_n3849_));
AND2X2 AND2X2_1639 ( .A(_abc_40319_new_n3846_), .B(_abc_40319_new_n1568_), .Y(_abc_40319_new_n3851_));
AND2X2 AND2X2_164 ( .A(_abc_40319_new_n848_), .B(_abc_40319_new_n763_), .Y(_abc_40319_new_n868_));
AND2X2 AND2X2_1640 ( .A(_abc_40319_new_n3851_), .B(_abc_40319_new_n3850_), .Y(_abc_40319_new_n3852_));
AND2X2 AND2X2_1641 ( .A(_abc_40319_new_n3853_), .B(_abc_40319_new_n629_), .Y(_abc_40319_new_n3854_));
AND2X2 AND2X2_1642 ( .A(_abc_40319_new_n3856_), .B(_abc_40319_new_n3580_), .Y(_abc_40319_new_n3857_));
AND2X2 AND2X2_1643 ( .A(_abc_40319_new_n3855_), .B(_abc_40319_new_n3579_), .Y(_abc_40319_new_n3858_));
AND2X2 AND2X2_1644 ( .A(_abc_40319_new_n3585_), .B(ADDR_REG_8_), .Y(_abc_40319_new_n3859_));
AND2X2 AND2X2_1645 ( .A(_abc_40319_new_n3579_), .B(_abc_40319_new_n3830_), .Y(_abc_40319_new_n3860_));
AND2X2 AND2X2_1646 ( .A(_abc_40319_new_n1609_), .B(REG2_REG_9_), .Y(_abc_40319_new_n3865_));
AND2X2 AND2X2_1647 ( .A(_abc_40319_new_n3866_), .B(_abc_40319_new_n3867_), .Y(_abc_40319_new_n3868_));
AND2X2 AND2X2_1648 ( .A(_abc_40319_new_n3836_), .B(_abc_40319_new_n3838_), .Y(_abc_40319_new_n3870_));
AND2X2 AND2X2_1649 ( .A(_abc_40319_new_n3871_), .B(_abc_40319_new_n3869_), .Y(_abc_40319_new_n3872_));
AND2X2 AND2X2_165 ( .A(_abc_40319_new_n865_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n869_));
AND2X2 AND2X2_1650 ( .A(_abc_40319_new_n3870_), .B(_abc_40319_new_n3868_), .Y(_abc_40319_new_n3873_));
AND2X2 AND2X2_1651 ( .A(_abc_40319_new_n3874_), .B(_abc_40319_new_n3555_), .Y(_abc_40319_new_n3875_));
AND2X2 AND2X2_1652 ( .A(_abc_40319_new_n1609_), .B(REG1_REG_9_), .Y(_abc_40319_new_n3876_));
AND2X2 AND2X2_1653 ( .A(_abc_40319_new_n3877_), .B(_abc_40319_new_n3878_), .Y(_abc_40319_new_n3879_));
AND2X2 AND2X2_1654 ( .A(_abc_40319_new_n3880_), .B(_abc_40319_new_n3879_), .Y(_abc_40319_new_n3881_));
AND2X2 AND2X2_1655 ( .A(_abc_40319_new_n3883_), .B(_abc_40319_new_n3882_), .Y(_abc_40319_new_n3884_));
AND2X2 AND2X2_1656 ( .A(_abc_40319_new_n3885_), .B(_abc_40319_new_n629_), .Y(_abc_40319_new_n3886_));
AND2X2 AND2X2_1657 ( .A(_abc_40319_new_n3887_), .B(_abc_40319_new_n3581_), .Y(_abc_40319_new_n3888_));
AND2X2 AND2X2_1658 ( .A(_abc_40319_new_n3585_), .B(ADDR_REG_9_), .Y(_abc_40319_new_n3889_));
AND2X2 AND2X2_1659 ( .A(_abc_40319_new_n639_), .B(_abc_40319_new_n1609_), .Y(_abc_40319_new_n3890_));
AND2X2 AND2X2_166 ( .A(_abc_40319_new_n872_), .B(_abc_40319_new_n873_), .Y(_abc_40319_new_n874_));
AND2X2 AND2X2_1660 ( .A(_abc_40319_new_n3579_), .B(_abc_40319_new_n3890_), .Y(_abc_40319_new_n3891_));
AND2X2 AND2X2_1661 ( .A(_abc_40319_new_n3580_), .B(_abc_40319_new_n3890_), .Y(_abc_40319_new_n3893_));
AND2X2 AND2X2_1662 ( .A(_abc_40319_new_n639_), .B(_abc_40319_new_n3897_), .Y(_abc_40319_new_n3898_));
AND2X2 AND2X2_1663 ( .A(_abc_40319_new_n3900_), .B(_abc_40319_new_n3877_), .Y(_abc_40319_new_n3901_));
AND2X2 AND2X2_1664 ( .A(_abc_40319_new_n3902_), .B(REG1_REG_10_), .Y(_abc_40319_new_n3903_));
AND2X2 AND2X2_1665 ( .A(_abc_40319_new_n3901_), .B(_abc_40319_new_n3905_), .Y(_abc_40319_new_n3906_));
AND2X2 AND2X2_1666 ( .A(_abc_40319_new_n3904_), .B(_abc_40319_new_n3907_), .Y(_abc_40319_new_n3908_));
AND2X2 AND2X2_1667 ( .A(_abc_40319_new_n3910_), .B(_abc_40319_new_n3911_), .Y(_abc_40319_new_n3912_));
AND2X2 AND2X2_1668 ( .A(_abc_40319_new_n3912_), .B(_abc_40319_new_n629_), .Y(_abc_40319_new_n3913_));
AND2X2 AND2X2_1669 ( .A(_abc_40319_new_n3914_), .B(_abc_40319_new_n3580_), .Y(_abc_40319_new_n3915_));
AND2X2 AND2X2_167 ( .A(_abc_40319_new_n875_), .B(_abc_40319_new_n871_), .Y(_abc_40319_new_n876_));
AND2X2 AND2X2_1670 ( .A(_abc_40319_new_n3579_), .B(_abc_40319_new_n629_), .Y(_abc_40319_new_n3916_));
AND2X2 AND2X2_1671 ( .A(_abc_40319_new_n3912_), .B(_abc_40319_new_n3916_), .Y(_abc_40319_new_n3917_));
AND2X2 AND2X2_1672 ( .A(_abc_40319_new_n3585_), .B(ADDR_REG_10_), .Y(_abc_40319_new_n3918_));
AND2X2 AND2X2_1673 ( .A(_abc_40319_new_n3579_), .B(_abc_40319_new_n3898_), .Y(_abc_40319_new_n3919_));
AND2X2 AND2X2_1674 ( .A(_abc_40319_new_n3897_), .B(REG2_REG_10_), .Y(_abc_40319_new_n3922_));
AND2X2 AND2X2_1675 ( .A(_abc_40319_new_n3923_), .B(_abc_40319_new_n3924_), .Y(_abc_40319_new_n3925_));
AND2X2 AND2X2_1676 ( .A(_abc_40319_new_n3871_), .B(_abc_40319_new_n3867_), .Y(_abc_40319_new_n3926_));
AND2X2 AND2X2_1677 ( .A(_abc_40319_new_n3579_), .B(_abc_40319_new_n3555_), .Y(_abc_40319_new_n3932_));
AND2X2 AND2X2_1678 ( .A(_abc_40319_new_n3580_), .B(_abc_40319_new_n3555_), .Y(_abc_40319_new_n3933_));
AND2X2 AND2X2_1679 ( .A(_abc_40319_new_n3931_), .B(_abc_40319_new_n3934_), .Y(_abc_40319_new_n3935_));
AND2X2 AND2X2_168 ( .A(_abc_40319_new_n876_), .B(_abc_40319_new_n867_), .Y(_abc_40319_new_n877_));
AND2X2 AND2X2_1680 ( .A(_abc_40319_new_n3935_), .B(_abc_40319_new_n3928_), .Y(_abc_40319_new_n3936_));
AND2X2 AND2X2_1681 ( .A(_abc_40319_new_n3940_), .B(REG1_REG_11_), .Y(_abc_40319_new_n3941_));
AND2X2 AND2X2_1682 ( .A(_abc_40319_new_n3942_), .B(_abc_40319_new_n3943_), .Y(_abc_40319_new_n3944_));
AND2X2 AND2X2_1683 ( .A(_abc_40319_new_n3904_), .B(_abc_40319_new_n3946_), .Y(_abc_40319_new_n3947_));
AND2X2 AND2X2_1684 ( .A(_abc_40319_new_n3948_), .B(_abc_40319_new_n3945_), .Y(_abc_40319_new_n3949_));
AND2X2 AND2X2_1685 ( .A(_abc_40319_new_n3947_), .B(_abc_40319_new_n3944_), .Y(_abc_40319_new_n3950_));
AND2X2 AND2X2_1686 ( .A(_abc_40319_new_n3580_), .B(_abc_40319_new_n629_), .Y(_abc_40319_new_n3952_));
AND2X2 AND2X2_1687 ( .A(_abc_40319_new_n3951_), .B(_abc_40319_new_n3953_), .Y(_abc_40319_new_n3954_));
AND2X2 AND2X2_1688 ( .A(_abc_40319_new_n3940_), .B(REG2_REG_11_), .Y(_abc_40319_new_n3955_));
AND2X2 AND2X2_1689 ( .A(_abc_40319_new_n3956_), .B(_abc_40319_new_n3957_), .Y(_abc_40319_new_n3958_));
AND2X2 AND2X2_169 ( .A(_abc_40319_new_n878_), .B(_abc_40319_new_n835_), .Y(_abc_40319_new_n879_));
AND2X2 AND2X2_1690 ( .A(_abc_40319_new_n3927_), .B(_abc_40319_new_n3924_), .Y(_abc_40319_new_n3960_));
AND2X2 AND2X2_1691 ( .A(_abc_40319_new_n3961_), .B(_abc_40319_new_n3959_), .Y(_abc_40319_new_n3962_));
AND2X2 AND2X2_1692 ( .A(_abc_40319_new_n3963_), .B(_abc_40319_new_n3958_), .Y(_abc_40319_new_n3964_));
AND2X2 AND2X2_1693 ( .A(_abc_40319_new_n3965_), .B(_abc_40319_new_n3934_), .Y(_abc_40319_new_n3966_));
AND2X2 AND2X2_1694 ( .A(_abc_40319_new_n3585_), .B(ADDR_REG_11_), .Y(_abc_40319_new_n3967_));
AND2X2 AND2X2_1695 ( .A(_abc_40319_new_n639_), .B(_abc_40319_new_n3940_), .Y(_abc_40319_new_n3969_));
AND2X2 AND2X2_1696 ( .A(_abc_40319_new_n3579_), .B(_abc_40319_new_n3969_), .Y(_abc_40319_new_n3970_));
AND2X2 AND2X2_1697 ( .A(_abc_40319_new_n3580_), .B(_abc_40319_new_n3969_), .Y(_abc_40319_new_n3971_));
AND2X2 AND2X2_1698 ( .A(_abc_40319_new_n3976_), .B(REG1_REG_12_), .Y(_abc_40319_new_n3977_));
AND2X2 AND2X2_1699 ( .A(_abc_40319_new_n3978_), .B(_abc_40319_new_n3979_), .Y(_abc_40319_new_n3980_));
AND2X2 AND2X2_17 ( .A(_abc_40319_new_n563_), .B(_abc_40319_new_n564_), .Y(_abc_40319_new_n565_));
AND2X2 AND2X2_170 ( .A(_abc_40319_new_n877_), .B(_abc_40319_new_n838_), .Y(_abc_40319_new_n880_));
AND2X2 AND2X2_1700 ( .A(_abc_40319_new_n3983_), .B(_abc_40319_new_n3942_), .Y(_abc_40319_new_n3984_));
AND2X2 AND2X2_1701 ( .A(_abc_40319_new_n3985_), .B(_abc_40319_new_n3981_), .Y(_abc_40319_new_n3986_));
AND2X2 AND2X2_1702 ( .A(_abc_40319_new_n3984_), .B(_abc_40319_new_n3980_), .Y(_abc_40319_new_n3987_));
AND2X2 AND2X2_1703 ( .A(_abc_40319_new_n3988_), .B(_abc_40319_new_n3953_), .Y(_abc_40319_new_n3989_));
AND2X2 AND2X2_1704 ( .A(_abc_40319_new_n3976_), .B(REG2_REG_12_), .Y(_abc_40319_new_n3990_));
AND2X2 AND2X2_1705 ( .A(_abc_40319_new_n3991_), .B(_abc_40319_new_n3992_), .Y(_abc_40319_new_n3993_));
AND2X2 AND2X2_1706 ( .A(_abc_40319_new_n3961_), .B(_abc_40319_new_n3957_), .Y(_abc_40319_new_n3995_));
AND2X2 AND2X2_1707 ( .A(_abc_40319_new_n3996_), .B(_abc_40319_new_n3994_), .Y(_abc_40319_new_n3997_));
AND2X2 AND2X2_1708 ( .A(_abc_40319_new_n3998_), .B(_abc_40319_new_n3993_), .Y(_abc_40319_new_n3999_));
AND2X2 AND2X2_1709 ( .A(_abc_40319_new_n4000_), .B(_abc_40319_new_n3934_), .Y(_abc_40319_new_n4001_));
AND2X2 AND2X2_171 ( .A(IR_REG_0_), .B(IR_REG_1_), .Y(_abc_40319_new_n882_));
AND2X2 AND2X2_1710 ( .A(_abc_40319_new_n3585_), .B(ADDR_REG_12_), .Y(_abc_40319_new_n4002_));
AND2X2 AND2X2_1711 ( .A(_abc_40319_new_n639_), .B(_abc_40319_new_n3976_), .Y(_abc_40319_new_n4004_));
AND2X2 AND2X2_1712 ( .A(_abc_40319_new_n3579_), .B(_abc_40319_new_n4004_), .Y(_abc_40319_new_n4005_));
AND2X2 AND2X2_1713 ( .A(_abc_40319_new_n3580_), .B(_abc_40319_new_n4004_), .Y(_abc_40319_new_n4006_));
AND2X2 AND2X2_1714 ( .A(_abc_40319_new_n4014_), .B(_abc_40319_new_n3978_), .Y(_abc_40319_new_n4015_));
AND2X2 AND2X2_1715 ( .A(_abc_40319_new_n4015_), .B(_abc_40319_new_n4012_), .Y(_abc_40319_new_n4016_));
AND2X2 AND2X2_1716 ( .A(_abc_40319_new_n4018_), .B(REG1_REG_13_), .Y(_abc_40319_new_n4019_));
AND2X2 AND2X2_1717 ( .A(_abc_40319_new_n4020_), .B(_abc_40319_new_n4017_), .Y(_abc_40319_new_n4021_));
AND2X2 AND2X2_1718 ( .A(_abc_40319_new_n4022_), .B(_abc_40319_new_n4011_), .Y(_abc_40319_new_n4023_));
AND2X2 AND2X2_1719 ( .A(_abc_40319_new_n4021_), .B(_abc_40319_new_n1651_), .Y(_abc_40319_new_n4024_));
AND2X2 AND2X2_172 ( .A(_abc_40319_new_n839_), .B(_abc_40319_new_n883_), .Y(_abc_40319_new_n884_));
AND2X2 AND2X2_1720 ( .A(_abc_40319_new_n4025_), .B(_abc_40319_new_n3953_), .Y(_abc_40319_new_n4026_));
AND2X2 AND2X2_1721 ( .A(_abc_40319_new_n4011_), .B(REG2_REG_13_), .Y(_abc_40319_new_n4027_));
AND2X2 AND2X2_1722 ( .A(_abc_40319_new_n4028_), .B(_abc_40319_new_n4029_), .Y(_abc_40319_new_n4030_));
AND2X2 AND2X2_1723 ( .A(_abc_40319_new_n3996_), .B(_abc_40319_new_n3992_), .Y(_abc_40319_new_n4031_));
AND2X2 AND2X2_1724 ( .A(_abc_40319_new_n4036_), .B(_abc_40319_new_n3934_), .Y(_abc_40319_new_n4037_));
AND2X2 AND2X2_1725 ( .A(_abc_40319_new_n4037_), .B(_abc_40319_new_n4033_), .Y(_abc_40319_new_n4038_));
AND2X2 AND2X2_1726 ( .A(_abc_40319_new_n3585_), .B(ADDR_REG_13_), .Y(_abc_40319_new_n4039_));
AND2X2 AND2X2_1727 ( .A(_abc_40319_new_n639_), .B(_abc_40319_new_n4011_), .Y(_abc_40319_new_n4040_));
AND2X2 AND2X2_1728 ( .A(_abc_40319_new_n3579_), .B(_abc_40319_new_n4040_), .Y(_abc_40319_new_n4041_));
AND2X2 AND2X2_1729 ( .A(_abc_40319_new_n3580_), .B(_abc_40319_new_n4040_), .Y(_abc_40319_new_n4043_));
AND2X2 AND2X2_173 ( .A(_abc_40319_new_n524_), .B(IR_REG_1_), .Y(_abc_40319_new_n885_));
AND2X2 AND2X2_1730 ( .A(_abc_40319_new_n4020_), .B(_abc_40319_new_n4049_), .Y(_abc_40319_new_n4050_));
AND2X2 AND2X2_1731 ( .A(_abc_40319_new_n4050_), .B(_abc_40319_new_n4048_), .Y(_abc_40319_new_n4051_));
AND2X2 AND2X2_1732 ( .A(_abc_40319_new_n4054_), .B(_abc_40319_new_n1501_), .Y(_abc_40319_new_n4055_));
AND2X2 AND2X2_1733 ( .A(_abc_40319_new_n4052_), .B(_abc_40319_new_n1502_), .Y(_abc_40319_new_n4057_));
AND2X2 AND2X2_1734 ( .A(_abc_40319_new_n4057_), .B(_abc_40319_new_n4056_), .Y(_abc_40319_new_n4058_));
AND2X2 AND2X2_1735 ( .A(_abc_40319_new_n4059_), .B(_abc_40319_new_n3953_), .Y(_abc_40319_new_n4060_));
AND2X2 AND2X2_1736 ( .A(_abc_40319_new_n1501_), .B(REG2_REG_14_), .Y(_abc_40319_new_n4061_));
AND2X2 AND2X2_1737 ( .A(_abc_40319_new_n4062_), .B(_abc_40319_new_n4063_), .Y(_abc_40319_new_n4064_));
AND2X2 AND2X2_1738 ( .A(_abc_40319_new_n4032_), .B(_abc_40319_new_n4029_), .Y(_abc_40319_new_n4066_));
AND2X2 AND2X2_1739 ( .A(_abc_40319_new_n4069_), .B(_abc_40319_new_n4070_), .Y(_abc_40319_new_n4071_));
AND2X2 AND2X2_174 ( .A(_abc_40319_new_n817_), .B(_abc_40319_new_n888_), .Y(_abc_40319_new_n889_));
AND2X2 AND2X2_1740 ( .A(_abc_40319_new_n4071_), .B(_abc_40319_new_n3932_), .Y(_abc_40319_new_n4072_));
AND2X2 AND2X2_1741 ( .A(_abc_40319_new_n3585_), .B(ADDR_REG_14_), .Y(_abc_40319_new_n4073_));
AND2X2 AND2X2_1742 ( .A(_abc_40319_new_n639_), .B(_abc_40319_new_n1501_), .Y(_abc_40319_new_n4074_));
AND2X2 AND2X2_1743 ( .A(_abc_40319_new_n3579_), .B(_abc_40319_new_n4074_), .Y(_abc_40319_new_n4075_));
AND2X2 AND2X2_1744 ( .A(_abc_40319_new_n4071_), .B(_abc_40319_new_n3555_), .Y(_abc_40319_new_n4079_));
AND2X2 AND2X2_1745 ( .A(_abc_40319_new_n4080_), .B(_abc_40319_new_n3580_), .Y(_abc_40319_new_n4081_));
AND2X2 AND2X2_1746 ( .A(_abc_40319_new_n4085_), .B(_abc_40319_new_n4084_), .Y(_abc_40319_new_n4086_));
AND2X2 AND2X2_1747 ( .A(_abc_40319_new_n4088_), .B(REG1_REG_15_), .Y(_abc_40319_new_n4089_));
AND2X2 AND2X2_1748 ( .A(_abc_40319_new_n4090_), .B(_abc_40319_new_n4087_), .Y(_abc_40319_new_n4091_));
AND2X2 AND2X2_1749 ( .A(_abc_40319_new_n4094_), .B(_abc_40319_new_n4092_), .Y(_abc_40319_new_n4095_));
AND2X2 AND2X2_175 ( .A(_abc_40319_new_n890_), .B(_abc_40319_new_n887_), .Y(_abc_40319_new_n891_));
AND2X2 AND2X2_1750 ( .A(_abc_40319_new_n4095_), .B(_abc_40319_new_n3953_), .Y(_abc_40319_new_n4096_));
AND2X2 AND2X2_1751 ( .A(_abc_40319_new_n639_), .B(_abc_40319_new_n1466_), .Y(_abc_40319_new_n4097_));
AND2X2 AND2X2_1752 ( .A(_abc_40319_new_n1466_), .B(REG2_REG_15_), .Y(_abc_40319_new_n4098_));
AND2X2 AND2X2_1753 ( .A(_abc_40319_new_n4099_), .B(_abc_40319_new_n4100_), .Y(_abc_40319_new_n4101_));
AND2X2 AND2X2_1754 ( .A(_abc_40319_new_n4067_), .B(_abc_40319_new_n4063_), .Y(_abc_40319_new_n4103_));
AND2X2 AND2X2_1755 ( .A(_abc_40319_new_n4106_), .B(_abc_40319_new_n4107_), .Y(_abc_40319_new_n4108_));
AND2X2 AND2X2_1756 ( .A(_abc_40319_new_n4108_), .B(_abc_40319_new_n3555_), .Y(_abc_40319_new_n4109_));
AND2X2 AND2X2_1757 ( .A(_abc_40319_new_n4110_), .B(_abc_40319_new_n3580_), .Y(_abc_40319_new_n4111_));
AND2X2 AND2X2_1758 ( .A(_abc_40319_new_n4108_), .B(_abc_40319_new_n3932_), .Y(_abc_40319_new_n4112_));
AND2X2 AND2X2_1759 ( .A(_abc_40319_new_n3585_), .B(ADDR_REG_15_), .Y(_abc_40319_new_n4113_));
AND2X2 AND2X2_176 ( .A(_abc_40319_new_n891_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n892_));
AND2X2 AND2X2_1760 ( .A(_abc_40319_new_n3579_), .B(_abc_40319_new_n4097_), .Y(_abc_40319_new_n4114_));
AND2X2 AND2X2_1761 ( .A(_abc_40319_new_n4120_), .B(REG1_REG_16_), .Y(_abc_40319_new_n4121_));
AND2X2 AND2X2_1762 ( .A(_abc_40319_new_n4122_), .B(_abc_40319_new_n4123_), .Y(_abc_40319_new_n4124_));
AND2X2 AND2X2_1763 ( .A(_abc_40319_new_n4090_), .B(_abc_40319_new_n4126_), .Y(_abc_40319_new_n4127_));
AND2X2 AND2X2_1764 ( .A(_abc_40319_new_n4128_), .B(_abc_40319_new_n4125_), .Y(_abc_40319_new_n4129_));
AND2X2 AND2X2_1765 ( .A(_abc_40319_new_n4127_), .B(_abc_40319_new_n4124_), .Y(_abc_40319_new_n4130_));
AND2X2 AND2X2_1766 ( .A(_abc_40319_new_n4131_), .B(_abc_40319_new_n3953_), .Y(_abc_40319_new_n4132_));
AND2X2 AND2X2_1767 ( .A(_abc_40319_new_n4120_), .B(REG2_REG_16_), .Y(_abc_40319_new_n4133_));
AND2X2 AND2X2_1768 ( .A(_abc_40319_new_n4134_), .B(_abc_40319_new_n4135_), .Y(_abc_40319_new_n4136_));
AND2X2 AND2X2_1769 ( .A(_abc_40319_new_n4104_), .B(_abc_40319_new_n4100_), .Y(_abc_40319_new_n4138_));
AND2X2 AND2X2_177 ( .A(_abc_40319_new_n736_), .B(REG0_REG_1_), .Y(_abc_40319_new_n893_));
AND2X2 AND2X2_1770 ( .A(_abc_40319_new_n4141_), .B(_abc_40319_new_n4142_), .Y(_abc_40319_new_n4143_));
AND2X2 AND2X2_1771 ( .A(_abc_40319_new_n4143_), .B(_abc_40319_new_n3932_), .Y(_abc_40319_new_n4144_));
AND2X2 AND2X2_1772 ( .A(_abc_40319_new_n639_), .B(_abc_40319_new_n4120_), .Y(_abc_40319_new_n4145_));
AND2X2 AND2X2_1773 ( .A(_abc_40319_new_n3579_), .B(_abc_40319_new_n4145_), .Y(_abc_40319_new_n4146_));
AND2X2 AND2X2_1774 ( .A(_abc_40319_new_n3585_), .B(ADDR_REG_16_), .Y(_abc_40319_new_n4147_));
AND2X2 AND2X2_1775 ( .A(_abc_40319_new_n4143_), .B(_abc_40319_new_n3555_), .Y(_abc_40319_new_n4151_));
AND2X2 AND2X2_1776 ( .A(_abc_40319_new_n4152_), .B(_abc_40319_new_n3580_), .Y(_abc_40319_new_n4153_));
AND2X2 AND2X2_1777 ( .A(_abc_40319_new_n1428_), .B(REG1_REG_17_), .Y(_abc_40319_new_n4156_));
AND2X2 AND2X2_1778 ( .A(_abc_40319_new_n4157_), .B(_abc_40319_new_n4158_), .Y(_abc_40319_new_n4159_));
AND2X2 AND2X2_1779 ( .A(_abc_40319_new_n4128_), .B(_abc_40319_new_n4123_), .Y(_abc_40319_new_n4161_));
AND2X2 AND2X2_178 ( .A(_abc_40319_new_n733_), .B(REG2_REG_1_), .Y(_abc_40319_new_n895_));
AND2X2 AND2X2_1780 ( .A(_abc_40319_new_n4162_), .B(_abc_40319_new_n4160_), .Y(_abc_40319_new_n4163_));
AND2X2 AND2X2_1781 ( .A(_abc_40319_new_n4164_), .B(_abc_40319_new_n4159_), .Y(_abc_40319_new_n4165_));
AND2X2 AND2X2_1782 ( .A(_abc_40319_new_n4166_), .B(_abc_40319_new_n3953_), .Y(_abc_40319_new_n4167_));
AND2X2 AND2X2_1783 ( .A(_abc_40319_new_n639_), .B(_abc_40319_new_n1428_), .Y(_abc_40319_new_n4168_));
AND2X2 AND2X2_1784 ( .A(_abc_40319_new_n1428_), .B(REG2_REG_17_), .Y(_abc_40319_new_n4169_));
AND2X2 AND2X2_1785 ( .A(_abc_40319_new_n4170_), .B(_abc_40319_new_n4171_), .Y(_abc_40319_new_n4172_));
AND2X2 AND2X2_1786 ( .A(_abc_40319_new_n4139_), .B(_abc_40319_new_n4135_), .Y(_abc_40319_new_n4174_));
AND2X2 AND2X2_1787 ( .A(_abc_40319_new_n4177_), .B(_abc_40319_new_n4178_), .Y(_abc_40319_new_n4179_));
AND2X2 AND2X2_1788 ( .A(_abc_40319_new_n4179_), .B(_abc_40319_new_n3555_), .Y(_abc_40319_new_n4180_));
AND2X2 AND2X2_1789 ( .A(_abc_40319_new_n4181_), .B(_abc_40319_new_n3580_), .Y(_abc_40319_new_n4182_));
AND2X2 AND2X2_179 ( .A(_abc_40319_new_n894_), .B(_abc_40319_new_n896_), .Y(_abc_40319_new_n897_));
AND2X2 AND2X2_1790 ( .A(_abc_40319_new_n4179_), .B(_abc_40319_new_n3932_), .Y(_abc_40319_new_n4183_));
AND2X2 AND2X2_1791 ( .A(_abc_40319_new_n3585_), .B(ADDR_REG_17_), .Y(_abc_40319_new_n4184_));
AND2X2 AND2X2_1792 ( .A(_abc_40319_new_n3579_), .B(_abc_40319_new_n4168_), .Y(_abc_40319_new_n4185_));
AND2X2 AND2X2_1793 ( .A(_abc_40319_new_n1359_), .B(_abc_40319_new_n4191_), .Y(_abc_40319_new_n4192_));
AND2X2 AND2X2_1794 ( .A(_abc_40319_new_n1358_), .B(REG1_REG_18_), .Y(_abc_40319_new_n4194_));
AND2X2 AND2X2_1795 ( .A(_abc_40319_new_n4193_), .B(_abc_40319_new_n4195_), .Y(_abc_40319_new_n4196_));
AND2X2 AND2X2_1796 ( .A(_abc_40319_new_n4162_), .B(_abc_40319_new_n4158_), .Y(_abc_40319_new_n4198_));
AND2X2 AND2X2_1797 ( .A(_abc_40319_new_n4199_), .B(_abc_40319_new_n4197_), .Y(_abc_40319_new_n4200_));
AND2X2 AND2X2_1798 ( .A(_abc_40319_new_n4201_), .B(_abc_40319_new_n4196_), .Y(_abc_40319_new_n4202_));
AND2X2 AND2X2_1799 ( .A(_abc_40319_new_n4203_), .B(_abc_40319_new_n629_), .Y(_abc_40319_new_n4204_));
AND2X2 AND2X2_18 ( .A(_abc_40319_new_n565_), .B(_abc_40319_new_n562_), .Y(_abc_40319_new_n566_));
AND2X2 AND2X2_180 ( .A(_abc_40319_new_n738_), .B(REG3_REG_1_), .Y(_abc_40319_new_n898_));
AND2X2 AND2X2_1800 ( .A(_abc_40319_new_n1359_), .B(_abc_40319_new_n4205_), .Y(_abc_40319_new_n4206_));
AND2X2 AND2X2_1801 ( .A(_abc_40319_new_n1358_), .B(REG2_REG_18_), .Y(_abc_40319_new_n4208_));
AND2X2 AND2X2_1802 ( .A(_abc_40319_new_n4207_), .B(_abc_40319_new_n4209_), .Y(_abc_40319_new_n4210_));
AND2X2 AND2X2_1803 ( .A(_abc_40319_new_n4175_), .B(_abc_40319_new_n4171_), .Y(_abc_40319_new_n4211_));
AND2X2 AND2X2_1804 ( .A(_abc_40319_new_n4216_), .B(_abc_40319_new_n4213_), .Y(_abc_40319_new_n4217_));
AND2X2 AND2X2_1805 ( .A(_abc_40319_new_n4217_), .B(_abc_40319_new_n3555_), .Y(_abc_40319_new_n4218_));
AND2X2 AND2X2_1806 ( .A(_abc_40319_new_n4219_), .B(_abc_40319_new_n3581_), .Y(_abc_40319_new_n4220_));
AND2X2 AND2X2_1807 ( .A(_abc_40319_new_n639_), .B(_abc_40319_new_n1358_), .Y(_abc_40319_new_n4221_));
AND2X2 AND2X2_1808 ( .A(_abc_40319_new_n3579_), .B(_abc_40319_new_n4221_), .Y(_abc_40319_new_n4222_));
AND2X2 AND2X2_1809 ( .A(_abc_40319_new_n3585_), .B(ADDR_REG_18_), .Y(_abc_40319_new_n4224_));
AND2X2 AND2X2_181 ( .A(_abc_40319_new_n722_), .B(REG1_REG_1_), .Y(_abc_40319_new_n900_));
AND2X2 AND2X2_1810 ( .A(_abc_40319_new_n3580_), .B(_abc_40319_new_n4221_), .Y(_abc_40319_new_n4225_));
AND2X2 AND2X2_1811 ( .A(_abc_40319_new_n639_), .B(_abc_40319_new_n697_), .Y(_abc_40319_new_n4229_));
AND2X2 AND2X2_1812 ( .A(_abc_40319_new_n4212_), .B(_abc_40319_new_n4207_), .Y(_abc_40319_new_n4230_));
AND2X2 AND2X2_1813 ( .A(_abc_40319_new_n698_), .B(REG2_REG_19_), .Y(_abc_40319_new_n4233_));
AND2X2 AND2X2_1814 ( .A(_abc_40319_new_n4239_), .B(_abc_40319_new_n3555_), .Y(_abc_40319_new_n4240_));
AND2X2 AND2X2_1815 ( .A(_abc_40319_new_n4240_), .B(_abc_40319_new_n4238_), .Y(_abc_40319_new_n4241_));
AND2X2 AND2X2_1816 ( .A(_abc_40319_new_n698_), .B(REG1_REG_19_), .Y(_abc_40319_new_n4242_));
AND2X2 AND2X2_1817 ( .A(_abc_40319_new_n4199_), .B(_abc_40319_new_n4193_), .Y(_abc_40319_new_n4247_));
AND2X2 AND2X2_1818 ( .A(_abc_40319_new_n4248_), .B(_abc_40319_new_n4246_), .Y(_abc_40319_new_n4249_));
AND2X2 AND2X2_1819 ( .A(_abc_40319_new_n4250_), .B(_abc_40319_new_n4245_), .Y(_abc_40319_new_n4251_));
AND2X2 AND2X2_182 ( .A(_abc_40319_new_n901_), .B(_abc_40319_new_n899_), .Y(_abc_40319_new_n902_));
AND2X2 AND2X2_1820 ( .A(_abc_40319_new_n4252_), .B(_abc_40319_new_n629_), .Y(_abc_40319_new_n4253_));
AND2X2 AND2X2_1821 ( .A(_abc_40319_new_n4255_), .B(_abc_40319_new_n3580_), .Y(_abc_40319_new_n4256_));
AND2X2 AND2X2_1822 ( .A(_abc_40319_new_n4254_), .B(_abc_40319_new_n3579_), .Y(_abc_40319_new_n4257_));
AND2X2 AND2X2_1823 ( .A(_abc_40319_new_n3585_), .B(ADDR_REG_19_), .Y(_abc_40319_new_n4258_));
AND2X2 AND2X2_1824 ( .A(_abc_40319_new_n3579_), .B(_abc_40319_new_n4229_), .Y(_abc_40319_new_n4259_));
AND2X2 AND2X2_1825 ( .A(_abc_40319_new_n752_), .B(_abc_40319_new_n1116_), .Y(_abc_40319_new_n4264_));
AND2X2 AND2X2_1826 ( .A(_abc_40319_new_n4265_), .B(_abc_40319_new_n1076_), .Y(_abc_40319_new_n4266_));
AND2X2 AND2X2_1827 ( .A(_abc_40319_new_n1108_), .B(_abc_40319_new_n4267_), .Y(_abc_40319_new_n4268_));
AND2X2 AND2X2_1828 ( .A(_abc_40319_new_n4268_), .B(_abc_40319_new_n1120_), .Y(_abc_40319_new_n4269_));
AND2X2 AND2X2_1829 ( .A(_abc_40319_new_n4269_), .B(_abc_40319_new_n4266_), .Y(_abc_40319_new_n4270_));
AND2X2 AND2X2_183 ( .A(_abc_40319_new_n897_), .B(_abc_40319_new_n902_), .Y(_abc_40319_new_n903_));
AND2X2 AND2X2_1830 ( .A(_abc_40319_new_n4271_), .B(_abc_40319_new_n4264_), .Y(_abc_40319_new_n4272_));
AND2X2 AND2X2_1831 ( .A(_abc_40319_new_n4273_), .B(_abc_40319_new_n942_), .Y(_abc_40319_new_n4274_));
AND2X2 AND2X2_1832 ( .A(_abc_40319_new_n4274_), .B(_abc_40319_new_n847_), .Y(_abc_40319_new_n4275_));
AND2X2 AND2X2_1833 ( .A(_abc_40319_new_n4275_), .B(_abc_40319_new_n819_), .Y(_abc_40319_new_n4276_));
AND2X2 AND2X2_1834 ( .A(_abc_40319_new_n4276_), .B(_abc_40319_new_n3218_), .Y(_abc_40319_new_n4277_));
AND2X2 AND2X2_1835 ( .A(_abc_40319_new_n4277_), .B(_abc_40319_new_n2605_), .Y(_abc_40319_new_n4278_));
AND2X2 AND2X2_1836 ( .A(_abc_40319_new_n4278_), .B(_abc_40319_new_n2585_), .Y(_abc_40319_new_n4279_));
AND2X2 AND2X2_1837 ( .A(_abc_40319_new_n4279_), .B(_abc_40319_new_n2578_), .Y(_abc_40319_new_n4280_));
AND2X2 AND2X2_1838 ( .A(_abc_40319_new_n4280_), .B(_abc_40319_new_n2730_), .Y(_abc_40319_new_n4281_));
AND2X2 AND2X2_1839 ( .A(_abc_40319_new_n4281_), .B(_abc_40319_new_n2714_), .Y(_abc_40319_new_n4282_));
AND2X2 AND2X2_184 ( .A(_abc_40319_new_n904_), .B(_abc_40319_new_n705_), .Y(_abc_40319_new_n905_));
AND2X2 AND2X2_1840 ( .A(_abc_40319_new_n4282_), .B(_abc_40319_new_n2703_), .Y(_abc_40319_new_n4283_));
AND2X2 AND2X2_1841 ( .A(_abc_40319_new_n4283_), .B(_abc_40319_new_n2784_), .Y(_abc_40319_new_n4284_));
AND2X2 AND2X2_1842 ( .A(_abc_40319_new_n4284_), .B(_abc_40319_new_n2762_), .Y(_abc_40319_new_n4285_));
AND2X2 AND2X2_1843 ( .A(_abc_40319_new_n4285_), .B(_abc_40319_new_n2755_), .Y(_abc_40319_new_n4286_));
AND2X2 AND2X2_1844 ( .A(_abc_40319_new_n4286_), .B(_abc_40319_new_n2809_), .Y(_abc_40319_new_n4287_));
AND2X2 AND2X2_1845 ( .A(_abc_40319_new_n4287_), .B(_abc_40319_new_n2827_), .Y(_abc_40319_new_n4288_));
AND2X2 AND2X2_1846 ( .A(_abc_40319_new_n4288_), .B(_abc_40319_new_n2844_), .Y(_abc_40319_new_n4289_));
AND2X2 AND2X2_1847 ( .A(_abc_40319_new_n4289_), .B(_abc_40319_new_n2860_), .Y(_abc_40319_new_n4290_));
AND2X2 AND2X2_1848 ( .A(_abc_40319_new_n4290_), .B(_abc_40319_new_n2877_), .Y(_abc_40319_new_n4291_));
AND2X2 AND2X2_1849 ( .A(_abc_40319_new_n4291_), .B(_abc_40319_new_n2893_), .Y(_abc_40319_new_n4292_));
AND2X2 AND2X2_185 ( .A(_abc_40319_new_n763_), .B(_abc_40319_new_n891_), .Y(_abc_40319_new_n907_));
AND2X2 AND2X2_1850 ( .A(_abc_40319_new_n4292_), .B(_abc_40319_new_n2910_), .Y(_abc_40319_new_n4293_));
AND2X2 AND2X2_1851 ( .A(_abc_40319_new_n4293_), .B(_abc_40319_new_n2926_), .Y(_abc_40319_new_n4294_));
AND2X2 AND2X2_1852 ( .A(_abc_40319_new_n4294_), .B(_abc_40319_new_n2943_), .Y(_abc_40319_new_n4295_));
AND2X2 AND2X2_1853 ( .A(_abc_40319_new_n4295_), .B(_abc_40319_new_n2959_), .Y(_abc_40319_new_n4296_));
AND2X2 AND2X2_1854 ( .A(_abc_40319_new_n4296_), .B(_abc_40319_new_n2976_), .Y(_abc_40319_new_n4297_));
AND2X2 AND2X2_1855 ( .A(_abc_40319_new_n4297_), .B(_abc_40319_new_n2992_), .Y(_abc_40319_new_n4298_));
AND2X2 AND2X2_1856 ( .A(_abc_40319_new_n4298_), .B(_abc_40319_new_n3009_), .Y(_abc_40319_new_n4299_));
AND2X2 AND2X2_1857 ( .A(_abc_40319_new_n4299_), .B(_abc_40319_new_n3025_), .Y(_abc_40319_new_n4300_));
AND2X2 AND2X2_1858 ( .A(_abc_40319_new_n4300_), .B(_abc_40319_new_n3042_), .Y(_abc_40319_new_n4301_));
AND2X2 AND2X2_1859 ( .A(_abc_40319_new_n4301_), .B(_abc_40319_new_n3059_), .Y(_abc_40319_new_n4302_));
AND2X2 AND2X2_186 ( .A(_abc_40319_new_n908_), .B(_abc_40319_new_n910_), .Y(_abc_40319_new_n911_));
AND2X2 AND2X2_1860 ( .A(_abc_40319_new_n4302_), .B(_abc_40319_new_n3169_), .Y(_abc_40319_new_n4303_));
AND2X2 AND2X2_1861 ( .A(_abc_40319_new_n4304_), .B(_abc_40319_new_n3162_), .Y(_abc_40319_new_n4305_));
AND2X2 AND2X2_1862 ( .A(_abc_40319_new_n4303_), .B(_abc_40319_new_n2553_), .Y(_abc_40319_new_n4306_));
AND2X2 AND2X2_1863 ( .A(_abc_40319_new_n4307_), .B(_abc_40319_new_n4272_), .Y(_abc_40319_new_n4308_));
AND2X2 AND2X2_1864 ( .A(_abc_40319_new_n656_), .B(_abc_40319_new_n639_), .Y(_abc_40319_new_n4310_));
AND2X2 AND2X2_1865 ( .A(_abc_40319_new_n4311_), .B(_abc_40319_new_n4310_), .Y(_abc_40319_new_n4312_));
AND2X2 AND2X2_1866 ( .A(_abc_40319_new_n2560_), .B(_abc_40319_new_n4312_), .Y(_abc_40319_new_n4313_));
AND2X2 AND2X2_1867 ( .A(_abc_40319_new_n4314_), .B(_abc_40319_new_n4315_), .Y(_abc_40319_new_n4316_));
AND2X2 AND2X2_1868 ( .A(_abc_40319_new_n4271_), .B(_abc_40319_new_n1152_), .Y(_abc_40319_new_n4317_));
AND2X2 AND2X2_1869 ( .A(_abc_40319_new_n4317_), .B(_abc_40319_new_n2553_), .Y(_abc_40319_new_n4318_));
AND2X2 AND2X2_187 ( .A(_abc_40319_new_n913_), .B(_abc_40319_new_n914_), .Y(_abc_40319_new_n915_));
AND2X2 AND2X2_1870 ( .A(_abc_40319_new_n4304_), .B(_abc_40319_new_n4322_), .Y(_abc_40319_new_n4323_));
AND2X2 AND2X2_1871 ( .A(_abc_40319_new_n4323_), .B(_abc_40319_new_n4272_), .Y(_abc_40319_new_n4324_));
AND2X2 AND2X2_1872 ( .A(_abc_40319_new_n4314_), .B(_abc_40319_new_n4325_), .Y(_abc_40319_new_n4326_));
AND2X2 AND2X2_1873 ( .A(_abc_40319_new_n4317_), .B(_abc_40319_new_n3069_), .Y(_abc_40319_new_n4327_));
AND2X2 AND2X2_1874 ( .A(_abc_40319_new_n3023_), .B(_abc_40319_new_n3025_), .Y(_abc_40319_new_n4331_));
AND2X2 AND2X2_1875 ( .A(_abc_40319_new_n2974_), .B(_abc_40319_new_n2976_), .Y(_abc_40319_new_n4333_));
AND2X2 AND2X2_1876 ( .A(_abc_40319_new_n3007_), .B(_abc_40319_new_n3009_), .Y(_abc_40319_new_n4335_));
AND2X2 AND2X2_1877 ( .A(_abc_40319_new_n2990_), .B(_abc_40319_new_n2992_), .Y(_abc_40319_new_n4337_));
AND2X2 AND2X2_1878 ( .A(_abc_40319_new_n4336_), .B(_abc_40319_new_n4338_), .Y(_abc_40319_new_n4339_));
AND2X2 AND2X2_1879 ( .A(_abc_40319_new_n4339_), .B(_abc_40319_new_n4334_), .Y(_abc_40319_new_n4340_));
AND2X2 AND2X2_188 ( .A(_abc_40319_new_n915_), .B(_abc_40319_new_n906_), .Y(_abc_40319_new_n917_));
AND2X2 AND2X2_1880 ( .A(_abc_40319_new_n4340_), .B(_abc_40319_new_n4332_), .Y(_abc_40319_new_n4341_));
AND2X2 AND2X2_1881 ( .A(_abc_40319_new_n2957_), .B(_abc_40319_new_n2959_), .Y(_abc_40319_new_n4343_));
AND2X2 AND2X2_1882 ( .A(_abc_40319_new_n1317_), .B(_abc_40319_new_n1306_), .Y(_abc_40319_new_n4344_));
AND2X2 AND2X2_1883 ( .A(_abc_40319_new_n2941_), .B(_abc_40319_new_n2943_), .Y(_abc_40319_new_n4346_));
AND2X2 AND2X2_1884 ( .A(_abc_40319_new_n1340_), .B(_abc_40319_new_n1329_), .Y(_abc_40319_new_n4347_));
AND2X2 AND2X2_1885 ( .A(_abc_40319_new_n2924_), .B(_abc_40319_new_n2926_), .Y(_abc_40319_new_n4349_));
AND2X2 AND2X2_1886 ( .A(_abc_40319_new_n1374_), .B(_abc_40319_new_n1363_), .Y(_abc_40319_new_n4351_));
AND2X2 AND2X2_1887 ( .A(_abc_40319_new_n2891_), .B(_abc_40319_new_n2893_), .Y(_abc_40319_new_n4352_));
AND2X2 AND2X2_1888 ( .A(_abc_40319_new_n4354_), .B(_abc_40319_new_n4353_), .Y(_abc_40319_new_n4355_));
AND2X2 AND2X2_1889 ( .A(_abc_40319_new_n4355_), .B(_abc_40319_new_n4350_), .Y(_abc_40319_new_n4356_));
AND2X2 AND2X2_189 ( .A(_abc_40319_new_n733_), .B(REG2_REG_0_), .Y(_abc_40319_new_n918_));
AND2X2 AND2X2_1890 ( .A(_abc_40319_new_n4356_), .B(_abc_40319_new_n4351_), .Y(_abc_40319_new_n4357_));
AND2X2 AND2X2_1891 ( .A(_abc_40319_new_n1876_), .B(_abc_40319_new_n1865_), .Y(_abc_40319_new_n4358_));
AND2X2 AND2X2_1892 ( .A(_abc_40319_new_n1828_), .B(_abc_40319_new_n1817_), .Y(_abc_40319_new_n4359_));
AND2X2 AND2X2_1893 ( .A(_abc_40319_new_n4360_), .B(_abc_40319_new_n4354_), .Y(_abc_40319_new_n4361_));
AND2X2 AND2X2_1894 ( .A(_abc_40319_new_n4363_), .B(_abc_40319_new_n4350_), .Y(_abc_40319_new_n4364_));
AND2X2 AND2X2_1895 ( .A(_abc_40319_new_n2875_), .B(_abc_40319_new_n2877_), .Y(_abc_40319_new_n4365_));
AND2X2 AND2X2_1896 ( .A(_abc_40319_new_n4356_), .B(_abc_40319_new_n4366_), .Y(_abc_40319_new_n4367_));
AND2X2 AND2X2_1897 ( .A(_abc_40319_new_n1398_), .B(_abc_40319_new_n1410_), .Y(_abc_40319_new_n4368_));
AND2X2 AND2X2_1898 ( .A(_abc_40319_new_n4369_), .B(_abc_40319_new_n2860_), .Y(_abc_40319_new_n4370_));
AND2X2 AND2X2_1899 ( .A(_abc_40319_new_n4368_), .B(_abc_40319_new_n1433_), .Y(_abc_40319_new_n4372_));
AND2X2 AND2X2_19 ( .A(_abc_40319_new_n566_), .B(_abc_40319_new_n568_), .Y(_abc_40319_new_n569_));
AND2X2 AND2X2_190 ( .A(_abc_40319_new_n736_), .B(REG0_REG_0_), .Y(_abc_40319_new_n919_));
AND2X2 AND2X2_1900 ( .A(_abc_40319_new_n4371_), .B(_abc_40319_new_n4373_), .Y(_abc_40319_new_n4374_));
AND2X2 AND2X2_1901 ( .A(_abc_40319_new_n4367_), .B(_abc_40319_new_n4375_), .Y(_abc_40319_new_n4376_));
AND2X2 AND2X2_1902 ( .A(_abc_40319_new_n1471_), .B(_abc_40319_new_n1483_), .Y(_abc_40319_new_n4379_));
AND2X2 AND2X2_1903 ( .A(_abc_40319_new_n2827_), .B(_abc_40319_new_n2825_), .Y(_abc_40319_new_n4381_));
AND2X2 AND2X2_1904 ( .A(_abc_40319_new_n1506_), .B(_abc_40319_new_n1517_), .Y(_abc_40319_new_n4382_));
AND2X2 AND2X2_1905 ( .A(_abc_40319_new_n2809_), .B(_abc_40319_new_n2807_), .Y(_abc_40319_new_n4384_));
AND2X2 AND2X2_1906 ( .A(_abc_40319_new_n2755_), .B(_abc_40319_new_n2753_), .Y(_abc_40319_new_n4385_));
AND2X2 AND2X2_1907 ( .A(_abc_40319_new_n1724_), .B(_abc_40319_new_n1735_), .Y(_abc_40319_new_n4387_));
AND2X2 AND2X2_1908 ( .A(_abc_40319_new_n2762_), .B(_abc_40319_new_n2760_), .Y(_abc_40319_new_n4388_));
AND2X2 AND2X2_1909 ( .A(_abc_40319_new_n4389_), .B(_abc_40319_new_n4386_), .Y(_abc_40319_new_n4390_));
AND2X2 AND2X2_191 ( .A(_abc_40319_new_n738_), .B(REG3_REG_0_), .Y(_abc_40319_new_n921_));
AND2X2 AND2X2_1910 ( .A(_abc_40319_new_n4390_), .B(_abc_40319_new_n4387_), .Y(_abc_40319_new_n4391_));
AND2X2 AND2X2_1911 ( .A(_abc_40319_new_n1690_), .B(_abc_40319_new_n1701_), .Y(_abc_40319_new_n4392_));
AND2X2 AND2X2_1912 ( .A(_abc_40319_new_n1655_), .B(_abc_40319_new_n1667_), .Y(_abc_40319_new_n4393_));
AND2X2 AND2X2_1913 ( .A(_abc_40319_new_n4395_), .B(_abc_40319_new_n4386_), .Y(_abc_40319_new_n4396_));
AND2X2 AND2X2_1914 ( .A(_abc_40319_new_n2784_), .B(_abc_40319_new_n2782_), .Y(_abc_40319_new_n4397_));
AND2X2 AND2X2_1915 ( .A(_abc_40319_new_n2703_), .B(_abc_40319_new_n2701_), .Y(_abc_40319_new_n4399_));
AND2X2 AND2X2_1916 ( .A(_abc_40319_new_n2714_), .B(_abc_40319_new_n2712_), .Y(_abc_40319_new_n4401_));
AND2X2 AND2X2_1917 ( .A(_abc_40319_new_n1572_), .B(_abc_40319_new_n1146_), .Y(_abc_40319_new_n4403_));
AND2X2 AND2X2_1918 ( .A(_abc_40319_new_n4400_), .B(_abc_40319_new_n4403_), .Y(_abc_40319_new_n4404_));
AND2X2 AND2X2_1919 ( .A(_abc_40319_new_n4404_), .B(_abc_40319_new_n4402_), .Y(_abc_40319_new_n4405_));
AND2X2 AND2X2_192 ( .A(_abc_40319_new_n722_), .B(REG1_REG_0_), .Y(_abc_40319_new_n922_));
AND2X2 AND2X2_1920 ( .A(_abc_40319_new_n1614_), .B(_abc_40319_new_n1625_), .Y(_abc_40319_new_n4406_));
AND2X2 AND2X2_1921 ( .A(_abc_40319_new_n1758_), .B(_abc_40319_new_n1769_), .Y(_abc_40319_new_n4407_));
AND2X2 AND2X2_1922 ( .A(_abc_40319_new_n2730_), .B(_abc_40319_new_n2728_), .Y(_abc_40319_new_n4410_));
AND2X2 AND2X2_1923 ( .A(_abc_40319_new_n2578_), .B(_abc_40319_new_n2575_), .Y(_abc_40319_new_n4412_));
AND2X2 AND2X2_1924 ( .A(_abc_40319_new_n1034_), .B(_abc_40319_new_n1046_), .Y(_abc_40319_new_n4414_));
AND2X2 AND2X2_1925 ( .A(_abc_40319_new_n998_), .B(_abc_40319_new_n1010_), .Y(_abc_40319_new_n4415_));
AND2X2 AND2X2_1926 ( .A(_abc_40319_new_n2585_), .B(_abc_40319_new_n2583_), .Y(_abc_40319_new_n4416_));
AND2X2 AND2X2_1927 ( .A(_abc_40319_new_n904_), .B(_abc_40319_new_n891_), .Y(_abc_40319_new_n4418_));
AND2X2 AND2X2_1928 ( .A(_abc_40319_new_n4273_), .B(_abc_40319_new_n903_), .Y(_abc_40319_new_n4420_));
AND2X2 AND2X2_1929 ( .A(_abc_40319_new_n924_), .B(_abc_40319_new_n930_), .Y(_abc_40319_new_n4421_));
AND2X2 AND2X2_193 ( .A(_abc_40319_new_n705_), .B(_abc_40319_new_n924_), .Y(_abc_40319_new_n925_));
AND2X2 AND2X2_1930 ( .A(_abc_40319_new_n4423_), .B(_abc_40319_new_n4419_), .Y(_abc_40319_new_n4424_));
AND2X2 AND2X2_1931 ( .A(_abc_40319_new_n3218_), .B(_abc_40319_new_n3220_), .Y(_abc_40319_new_n4426_));
AND2X2 AND2X2_1932 ( .A(_abc_40319_new_n2605_), .B(_abc_40319_new_n2603_), .Y(_abc_40319_new_n4428_));
AND2X2 AND2X2_1933 ( .A(_abc_40319_new_n4427_), .B(_abc_40319_new_n4429_), .Y(_abc_40319_new_n4430_));
AND2X2 AND2X2_1934 ( .A(_abc_40319_new_n2650_), .B(_abc_40319_new_n819_), .Y(_abc_40319_new_n4431_));
AND2X2 AND2X2_1935 ( .A(_abc_40319_new_n847_), .B(_abc_40319_new_n864_), .Y(_abc_40319_new_n4433_));
AND2X2 AND2X2_1936 ( .A(_abc_40319_new_n4432_), .B(_abc_40319_new_n4434_), .Y(_abc_40319_new_n4435_));
AND2X2 AND2X2_1937 ( .A(_abc_40319_new_n4430_), .B(_abc_40319_new_n4435_), .Y(_abc_40319_new_n4436_));
AND2X2 AND2X2_1938 ( .A(_abc_40319_new_n4436_), .B(_abc_40319_new_n4425_), .Y(_abc_40319_new_n4437_));
AND2X2 AND2X2_1939 ( .A(_abc_40319_new_n820_), .B(_abc_40319_new_n829_), .Y(_abc_40319_new_n4438_));
AND2X2 AND2X2_194 ( .A(_abc_40319_new_n817_), .B(_abc_40319_new_n927_), .Y(_abc_40319_new_n928_));
AND2X2 AND2X2_1940 ( .A(_abc_40319_new_n848_), .B(_abc_40319_new_n865_), .Y(_abc_40319_new_n4439_));
AND2X2 AND2X2_1941 ( .A(_abc_40319_new_n4432_), .B(_abc_40319_new_n4439_), .Y(_abc_40319_new_n4440_));
AND2X2 AND2X2_1942 ( .A(_abc_40319_new_n4441_), .B(_abc_40319_new_n4430_), .Y(_abc_40319_new_n4442_));
AND2X2 AND2X2_1943 ( .A(_abc_40319_new_n689_), .B(_abc_40319_new_n746_), .Y(_abc_40319_new_n4443_));
AND2X2 AND2X2_1944 ( .A(_abc_40319_new_n784_), .B(_abc_40319_new_n795_), .Y(_abc_40319_new_n4444_));
AND2X2 AND2X2_1945 ( .A(_abc_40319_new_n4429_), .B(_abc_40319_new_n4444_), .Y(_abc_40319_new_n4445_));
AND2X2 AND2X2_1946 ( .A(_abc_40319_new_n4448_), .B(_abc_40319_new_n4417_), .Y(_abc_40319_new_n4449_));
AND2X2 AND2X2_1947 ( .A(_abc_40319_new_n4451_), .B(_abc_40319_new_n4413_), .Y(_abc_40319_new_n4452_));
AND2X2 AND2X2_1948 ( .A(_abc_40319_new_n4452_), .B(_abc_40319_new_n4411_), .Y(_abc_40319_new_n4453_));
AND2X2 AND2X2_1949 ( .A(_abc_40319_new_n4453_), .B(_abc_40319_new_n4402_), .Y(_abc_40319_new_n4454_));
AND2X2 AND2X2_195 ( .A(_abc_40319_new_n929_), .B(_abc_40319_new_n926_), .Y(_abc_40319_new_n930_));
AND2X2 AND2X2_1950 ( .A(_abc_40319_new_n4455_), .B(_abc_40319_new_n4400_), .Y(_abc_40319_new_n4456_));
AND2X2 AND2X2_1951 ( .A(_abc_40319_new_n4456_), .B(_abc_40319_new_n4398_), .Y(_abc_40319_new_n4457_));
AND2X2 AND2X2_1952 ( .A(_abc_40319_new_n4457_), .B(_abc_40319_new_n4390_), .Y(_abc_40319_new_n4458_));
AND2X2 AND2X2_1953 ( .A(_abc_40319_new_n4461_), .B(_abc_40319_new_n4383_), .Y(_abc_40319_new_n4462_));
AND2X2 AND2X2_1954 ( .A(_abc_40319_new_n4463_), .B(_abc_40319_new_n4380_), .Y(_abc_40319_new_n4464_));
AND2X2 AND2X2_1955 ( .A(_abc_40319_new_n2860_), .B(_abc_40319_new_n2858_), .Y(_abc_40319_new_n4465_));
AND2X2 AND2X2_1956 ( .A(_abc_40319_new_n2844_), .B(_abc_40319_new_n2842_), .Y(_abc_40319_new_n4466_));
AND2X2 AND2X2_1957 ( .A(_abc_40319_new_n4367_), .B(_abc_40319_new_n4468_), .Y(_abc_40319_new_n4469_));
AND2X2 AND2X2_1958 ( .A(_abc_40319_new_n4471_), .B(_abc_40319_new_n4378_), .Y(_abc_40319_new_n4472_));
AND2X2 AND2X2_1959 ( .A(_abc_40319_new_n4472_), .B(_abc_40319_new_n4348_), .Y(_abc_40319_new_n4473_));
AND2X2 AND2X2_196 ( .A(_abc_40319_new_n930_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n931_));
AND2X2 AND2X2_1960 ( .A(_abc_40319_new_n4474_), .B(_abc_40319_new_n4345_), .Y(_abc_40319_new_n4475_));
AND2X2 AND2X2_1961 ( .A(_abc_40319_new_n1210_), .B(_abc_40319_new_n1180_), .Y(_abc_40319_new_n4478_));
AND2X2 AND2X2_1962 ( .A(_abc_40319_new_n1235_), .B(_abc_40319_new_n1224_), .Y(_abc_40319_new_n4479_));
AND2X2 AND2X2_1963 ( .A(_abc_40319_new_n1260_), .B(_abc_40319_new_n1249_), .Y(_abc_40319_new_n4480_));
AND2X2 AND2X2_1964 ( .A(_abc_40319_new_n4336_), .B(_abc_40319_new_n4481_), .Y(_abc_40319_new_n4482_));
AND2X2 AND2X2_1965 ( .A(_abc_40319_new_n1285_), .B(_abc_40319_new_n1274_), .Y(_abc_40319_new_n4483_));
AND2X2 AND2X2_1966 ( .A(_abc_40319_new_n4339_), .B(_abc_40319_new_n4483_), .Y(_abc_40319_new_n4484_));
AND2X2 AND2X2_1967 ( .A(_abc_40319_new_n4485_), .B(_abc_40319_new_n4332_), .Y(_abc_40319_new_n4486_));
AND2X2 AND2X2_1968 ( .A(_abc_40319_new_n4477_), .B(_abc_40319_new_n4488_), .Y(_abc_40319_new_n4489_));
AND2X2 AND2X2_1969 ( .A(_abc_40319_new_n4490_), .B(_abc_40319_new_n3250_), .Y(_abc_40319_new_n4491_));
AND2X2 AND2X2_197 ( .A(_abc_40319_new_n598_), .B(IR_REG_0_), .Y(_abc_40319_new_n932_));
AND2X2 AND2X2_1970 ( .A(_abc_40319_new_n4489_), .B(_abc_40319_new_n3249_), .Y(_abc_40319_new_n4492_));
AND2X2 AND2X2_1971 ( .A(_abc_40319_new_n4495_), .B(_abc_40319_new_n698_), .Y(_abc_40319_new_n4496_));
AND2X2 AND2X2_1972 ( .A(_abc_40319_new_n4496_), .B(_abc_40319_new_n4494_), .Y(_abc_40319_new_n4497_));
AND2X2 AND2X2_1973 ( .A(_abc_40319_new_n4493_), .B(_abc_40319_new_n4497_), .Y(_abc_40319_new_n4498_));
AND2X2 AND2X2_1974 ( .A(_abc_40319_new_n656_), .B(_abc_40319_new_n638_), .Y(_abc_40319_new_n4499_));
AND2X2 AND2X2_1975 ( .A(_abc_40319_new_n1210_), .B(_abc_40319_new_n4499_), .Y(_abc_40319_new_n4500_));
AND2X2 AND2X2_1976 ( .A(_abc_40319_new_n4503_), .B(_abc_40319_new_n3249_), .Y(_abc_40319_new_n4504_));
AND2X2 AND2X2_1977 ( .A(_abc_40319_new_n4502_), .B(_abc_40319_new_n3250_), .Y(_abc_40319_new_n4505_));
AND2X2 AND2X2_1978 ( .A(_abc_40319_new_n4506_), .B(_abc_40319_new_n4507_), .Y(_abc_40319_new_n4508_));
AND2X2 AND2X2_1979 ( .A(_abc_40319_new_n4510_), .B(_abc_40319_new_n4271_), .Y(_abc_40319_new_n4511_));
AND2X2 AND2X2_198 ( .A(_abc_40319_new_n934_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n936_));
AND2X2 AND2X2_1980 ( .A(_abc_40319_new_n4271_), .B(_abc_40319_new_n3451_), .Y(_abc_40319_new_n4512_));
AND2X2 AND2X2_1981 ( .A(_abc_40319_new_n4493_), .B(_abc_40319_new_n4512_), .Y(_abc_40319_new_n4513_));
AND2X2 AND2X2_1982 ( .A(_abc_40319_new_n4514_), .B(_abc_40319_new_n4515_), .Y(_abc_40319_new_n4516_));
AND2X2 AND2X2_1983 ( .A(_abc_40319_new_n4516_), .B(_abc_40319_new_n4272_), .Y(_abc_40319_new_n4517_));
AND2X2 AND2X2_1984 ( .A(_abc_40319_new_n4271_), .B(_abc_40319_new_n4310_), .Y(_abc_40319_new_n4518_));
AND2X2 AND2X2_1985 ( .A(_abc_40319_new_n2123_), .B(_abc_40319_new_n4518_), .Y(_abc_40319_new_n4519_));
AND2X2 AND2X2_1986 ( .A(_abc_40319_new_n1973_), .B(_abc_40319_new_n1169_), .Y(_abc_40319_new_n4520_));
AND2X2 AND2X2_1987 ( .A(_abc_40319_new_n2089_), .B(_abc_40319_new_n1152_), .Y(_abc_40319_new_n4522_));
AND2X2 AND2X2_1988 ( .A(_abc_40319_new_n4523_), .B(_abc_40319_new_n4521_), .Y(_abc_40319_new_n4524_));
AND2X2 AND2X2_1989 ( .A(_abc_40319_new_n4531_), .B(_abc_40319_new_n4340_), .Y(_abc_40319_new_n4532_));
AND2X2 AND2X2_199 ( .A(_abc_40319_new_n937_), .B(_abc_40319_new_n938_), .Y(_abc_40319_new_n939_));
AND2X2 AND2X2_1990 ( .A(_abc_40319_new_n4536_), .B(_abc_40319_new_n4534_), .Y(_abc_40319_new_n4537_));
AND2X2 AND2X2_1991 ( .A(_abc_40319_new_n4537_), .B(_abc_40319_new_n4497_), .Y(_abc_40319_new_n4538_));
AND2X2 AND2X2_1992 ( .A(_abc_40319_new_n1235_), .B(_abc_40319_new_n4499_), .Y(_abc_40319_new_n4539_));
AND2X2 AND2X2_1993 ( .A(_abc_40319_new_n4540_), .B(_abc_40319_new_n3466_), .Y(_abc_40319_new_n4541_));
AND2X2 AND2X2_1994 ( .A(_abc_40319_new_n4544_), .B(_abc_40319_new_n4507_), .Y(_abc_40319_new_n4545_));
AND2X2 AND2X2_1995 ( .A(_abc_40319_new_n4545_), .B(_abc_40319_new_n4543_), .Y(_abc_40319_new_n4546_));
AND2X2 AND2X2_1996 ( .A(_abc_40319_new_n4548_), .B(_abc_40319_new_n4271_), .Y(_abc_40319_new_n4549_));
AND2X2 AND2X2_1997 ( .A(_abc_40319_new_n4537_), .B(_abc_40319_new_n4512_), .Y(_abc_40319_new_n4550_));
AND2X2 AND2X2_1998 ( .A(_abc_40319_new_n4551_), .B(_abc_40319_new_n4552_), .Y(_abc_40319_new_n4553_));
AND2X2 AND2X2_1999 ( .A(_abc_40319_new_n4553_), .B(_abc_40319_new_n4272_), .Y(_abc_40319_new_n4554_));
AND2X2 AND2X2_2 ( .A(_abc_40319_new_n530_), .B(_abc_40319_new_n528_), .Y(_abc_40319_new_n531_));
AND2X2 AND2X2_20 ( .A(_abc_40319_new_n561_), .B(_abc_40319_new_n569_), .Y(_abc_40319_new_n570_));
AND2X2 AND2X2_200 ( .A(_abc_40319_new_n640_), .B(_abc_40319_new_n940_), .Y(_abc_40319_new_n941_));
AND2X2 AND2X2_2000 ( .A(_abc_40319_new_n1980_), .B(_abc_40319_new_n4518_), .Y(_abc_40319_new_n4555_));
AND2X2 AND2X2_2001 ( .A(_abc_40319_new_n1203_), .B(_abc_40319_new_n1169_), .Y(_abc_40319_new_n4556_));
AND2X2 AND2X2_2002 ( .A(_abc_40319_new_n1180_), .B(_abc_40319_new_n1152_), .Y(_abc_40319_new_n4558_));
AND2X2 AND2X2_2003 ( .A(_abc_40319_new_n4559_), .B(_abc_40319_new_n4557_), .Y(_abc_40319_new_n4560_));
AND2X2 AND2X2_2004 ( .A(_abc_40319_new_n4531_), .B(_abc_40319_new_n4334_), .Y(_abc_40319_new_n4567_));
AND2X2 AND2X2_2005 ( .A(_abc_40319_new_n4568_), .B(_abc_40319_new_n4338_), .Y(_abc_40319_new_n4569_));
AND2X2 AND2X2_2006 ( .A(_abc_40319_new_n4573_), .B(_abc_40319_new_n4572_), .Y(_abc_40319_new_n4574_));
AND2X2 AND2X2_2007 ( .A(_abc_40319_new_n4571_), .B(_abc_40319_new_n4577_), .Y(_abc_40319_new_n4578_));
AND2X2 AND2X2_2008 ( .A(_abc_40319_new_n4578_), .B(_abc_40319_new_n4497_), .Y(_abc_40319_new_n4579_));
AND2X2 AND2X2_2009 ( .A(_abc_40319_new_n1260_), .B(_abc_40319_new_n4499_), .Y(_abc_40319_new_n4580_));
AND2X2 AND2X2_201 ( .A(_abc_40319_new_n945_), .B(_abc_40319_new_n947_), .Y(_abc_40319_new_n948_));
AND2X2 AND2X2_2010 ( .A(_abc_40319_new_n3535_), .B(_abc_40319_new_n3379_), .Y(_abc_40319_new_n4582_));
AND2X2 AND2X2_2011 ( .A(_abc_40319_new_n4583_), .B(_abc_40319_new_n4507_), .Y(_abc_40319_new_n4584_));
AND2X2 AND2X2_2012 ( .A(_abc_40319_new_n4581_), .B(_abc_40319_new_n4584_), .Y(_abc_40319_new_n4585_));
AND2X2 AND2X2_2013 ( .A(_abc_40319_new_n4587_), .B(_abc_40319_new_n4271_), .Y(_abc_40319_new_n4588_));
AND2X2 AND2X2_2014 ( .A(_abc_40319_new_n4578_), .B(_abc_40319_new_n4512_), .Y(_abc_40319_new_n4589_));
AND2X2 AND2X2_2015 ( .A(_abc_40319_new_n4590_), .B(_abc_40319_new_n4591_), .Y(_abc_40319_new_n4592_));
AND2X2 AND2X2_2016 ( .A(_abc_40319_new_n4592_), .B(_abc_40319_new_n4272_), .Y(_abc_40319_new_n4593_));
AND2X2 AND2X2_2017 ( .A(_abc_40319_new_n1210_), .B(_abc_40319_new_n4518_), .Y(_abc_40319_new_n4594_));
AND2X2 AND2X2_2018 ( .A(_abc_40319_new_n1228_), .B(_abc_40319_new_n1169_), .Y(_abc_40319_new_n4595_));
AND2X2 AND2X2_2019 ( .A(_abc_40319_new_n1224_), .B(_abc_40319_new_n1152_), .Y(_abc_40319_new_n4597_));
AND2X2 AND2X2_202 ( .A(_abc_40319_new_n950_), .B(_abc_40319_new_n952_), .Y(_abc_40319_new_n953_));
AND2X2 AND2X2_2020 ( .A(_abc_40319_new_n4598_), .B(_abc_40319_new_n4596_), .Y(_abc_40319_new_n4599_));
AND2X2 AND2X2_2021 ( .A(_abc_40319_new_n4568_), .B(_abc_40319_new_n3258_), .Y(_abc_40319_new_n4606_));
AND2X2 AND2X2_2022 ( .A(_abc_40319_new_n4573_), .B(_abc_40319_new_n3257_), .Y(_abc_40319_new_n4607_));
AND2X2 AND2X2_2023 ( .A(_abc_40319_new_n4608_), .B(_abc_40319_new_n4497_), .Y(_abc_40319_new_n4609_));
AND2X2 AND2X2_2024 ( .A(_abc_40319_new_n1285_), .B(_abc_40319_new_n4499_), .Y(_abc_40319_new_n4610_));
AND2X2 AND2X2_2025 ( .A(_abc_40319_new_n4614_), .B(_abc_40319_new_n4507_), .Y(_abc_40319_new_n4615_));
AND2X2 AND2X2_2026 ( .A(_abc_40319_new_n4615_), .B(_abc_40319_new_n4612_), .Y(_abc_40319_new_n4616_));
AND2X2 AND2X2_2027 ( .A(_abc_40319_new_n4618_), .B(_abc_40319_new_n4271_), .Y(_abc_40319_new_n4619_));
AND2X2 AND2X2_2028 ( .A(_abc_40319_new_n4608_), .B(_abc_40319_new_n4512_), .Y(_abc_40319_new_n4620_));
AND2X2 AND2X2_2029 ( .A(_abc_40319_new_n4621_), .B(_abc_40319_new_n4622_), .Y(_abc_40319_new_n4623_));
AND2X2 AND2X2_203 ( .A(_abc_40319_new_n948_), .B(_abc_40319_new_n953_), .Y(_abc_40319_new_n954_));
AND2X2 AND2X2_2030 ( .A(_abc_40319_new_n4623_), .B(_abc_40319_new_n4272_), .Y(_abc_40319_new_n4624_));
AND2X2 AND2X2_2031 ( .A(_abc_40319_new_n1235_), .B(_abc_40319_new_n4518_), .Y(_abc_40319_new_n4625_));
AND2X2 AND2X2_2032 ( .A(_abc_40319_new_n1253_), .B(_abc_40319_new_n1169_), .Y(_abc_40319_new_n4626_));
AND2X2 AND2X2_2033 ( .A(_abc_40319_new_n1249_), .B(_abc_40319_new_n1152_), .Y(_abc_40319_new_n4628_));
AND2X2 AND2X2_2034 ( .A(_abc_40319_new_n4629_), .B(_abc_40319_new_n4627_), .Y(_abc_40319_new_n4630_));
AND2X2 AND2X2_2035 ( .A(_abc_40319_new_n4531_), .B(_abc_40319_new_n3196_), .Y(_abc_40319_new_n4637_));
AND2X2 AND2X2_2036 ( .A(_abc_40319_new_n4476_), .B(_abc_40319_new_n3195_), .Y(_abc_40319_new_n4638_));
AND2X2 AND2X2_2037 ( .A(_abc_40319_new_n4639_), .B(_abc_40319_new_n4497_), .Y(_abc_40319_new_n4640_));
AND2X2 AND2X2_2038 ( .A(_abc_40319_new_n1317_), .B(_abc_40319_new_n4499_), .Y(_abc_40319_new_n4641_));
AND2X2 AND2X2_2039 ( .A(_abc_40319_new_n3519_), .B(_abc_40319_new_n3527_), .Y(_abc_40319_new_n4642_));
AND2X2 AND2X2_204 ( .A(_abc_40319_new_n943_), .B(_abc_40319_new_n955_), .Y(_abc_40319_new_n956_));
AND2X2 AND2X2_2040 ( .A(_abc_40319_new_n4643_), .B(_abc_40319_new_n3403_), .Y(_abc_40319_new_n4644_));
AND2X2 AND2X2_2041 ( .A(_abc_40319_new_n3400_), .B(_abc_40319_new_n3474_), .Y(_abc_40319_new_n4646_));
AND2X2 AND2X2_2042 ( .A(_abc_40319_new_n4646_), .B(_abc_40319_new_n3276_), .Y(_abc_40319_new_n4647_));
AND2X2 AND2X2_2043 ( .A(_abc_40319_new_n4645_), .B(_abc_40319_new_n4647_), .Y(_abc_40319_new_n4648_));
AND2X2 AND2X2_2044 ( .A(_abc_40319_new_n3292_), .B(_abc_40319_new_n3288_), .Y(_abc_40319_new_n4649_));
AND2X2 AND2X2_2045 ( .A(_abc_40319_new_n4651_), .B(_abc_40319_new_n3400_), .Y(_abc_40319_new_n4652_));
AND2X2 AND2X2_2046 ( .A(_abc_40319_new_n3399_), .B(_abc_40319_new_n3201_), .Y(_abc_40319_new_n4653_));
AND2X2 AND2X2_2047 ( .A(_abc_40319_new_n4655_), .B(_abc_40319_new_n3276_), .Y(_abc_40319_new_n4656_));
AND2X2 AND2X2_2048 ( .A(_abc_40319_new_n4660_), .B(_abc_40319_new_n4507_), .Y(_abc_40319_new_n4661_));
AND2X2 AND2X2_2049 ( .A(_abc_40319_new_n4661_), .B(_abc_40319_new_n4659_), .Y(_abc_40319_new_n4662_));
AND2X2 AND2X2_205 ( .A(_abc_40319_new_n763_), .B(_abc_40319_new_n930_), .Y(_abc_40319_new_n958_));
AND2X2 AND2X2_2050 ( .A(_abc_40319_new_n4664_), .B(_abc_40319_new_n4271_), .Y(_abc_40319_new_n4665_));
AND2X2 AND2X2_2051 ( .A(_abc_40319_new_n4639_), .B(_abc_40319_new_n4512_), .Y(_abc_40319_new_n4666_));
AND2X2 AND2X2_2052 ( .A(_abc_40319_new_n4667_), .B(_abc_40319_new_n4668_), .Y(_abc_40319_new_n4669_));
AND2X2 AND2X2_2053 ( .A(_abc_40319_new_n4669_), .B(_abc_40319_new_n4272_), .Y(_abc_40319_new_n4670_));
AND2X2 AND2X2_2054 ( .A(_abc_40319_new_n1260_), .B(_abc_40319_new_n4518_), .Y(_abc_40319_new_n4671_));
AND2X2 AND2X2_2055 ( .A(_abc_40319_new_n1278_), .B(_abc_40319_new_n1169_), .Y(_abc_40319_new_n4672_));
AND2X2 AND2X2_2056 ( .A(_abc_40319_new_n1274_), .B(_abc_40319_new_n1152_), .Y(_abc_40319_new_n4674_));
AND2X2 AND2X2_2057 ( .A(_abc_40319_new_n4675_), .B(_abc_40319_new_n4673_), .Y(_abc_40319_new_n4676_));
AND2X2 AND2X2_2058 ( .A(_abc_40319_new_n4645_), .B(_abc_40319_new_n3474_), .Y(_abc_40319_new_n4683_));
AND2X2 AND2X2_2059 ( .A(_abc_40319_new_n4685_), .B(_abc_40319_new_n3286_), .Y(_abc_40319_new_n4686_));
AND2X2 AND2X2_206 ( .A(_abc_40319_new_n924_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n959_));
AND2X2 AND2X2_2060 ( .A(_abc_40319_new_n3262_), .B(_abc_40319_new_n3349_), .Y(_abc_40319_new_n4688_));
AND2X2 AND2X2_2061 ( .A(_abc_40319_new_n4687_), .B(_abc_40319_new_n4688_), .Y(_abc_40319_new_n4689_));
AND2X2 AND2X2_2062 ( .A(_abc_40319_new_n3261_), .B(_abc_40319_new_n3400_), .Y(_abc_40319_new_n4690_));
AND2X2 AND2X2_2063 ( .A(_abc_40319_new_n4684_), .B(_abc_40319_new_n4690_), .Y(_abc_40319_new_n4691_));
AND2X2 AND2X2_2064 ( .A(_abc_40319_new_n4692_), .B(_abc_40319_new_n3261_), .Y(_abc_40319_new_n4693_));
AND2X2 AND2X2_2065 ( .A(_abc_40319_new_n3262_), .B(_abc_40319_new_n3198_), .Y(_abc_40319_new_n4694_));
AND2X2 AND2X2_2066 ( .A(_abc_40319_new_n4697_), .B(_abc_40319_new_n4507_), .Y(_abc_40319_new_n4698_));
AND2X2 AND2X2_2067 ( .A(_abc_40319_new_n1340_), .B(_abc_40319_new_n4499_), .Y(_abc_40319_new_n4699_));
AND2X2 AND2X2_2068 ( .A(_abc_40319_new_n4700_), .B(_abc_40319_new_n3262_), .Y(_abc_40319_new_n4701_));
AND2X2 AND2X2_2069 ( .A(_abc_40319_new_n4474_), .B(_abc_40319_new_n3261_), .Y(_abc_40319_new_n4702_));
AND2X2 AND2X2_207 ( .A(_abc_40319_new_n598_), .B(REG1_REG_0_), .Y(_abc_40319_new_n961_));
AND2X2 AND2X2_2070 ( .A(_abc_40319_new_n4703_), .B(_abc_40319_new_n4497_), .Y(_abc_40319_new_n4704_));
AND2X2 AND2X2_2071 ( .A(_abc_40319_new_n4706_), .B(_abc_40319_new_n4271_), .Y(_abc_40319_new_n4707_));
AND2X2 AND2X2_2072 ( .A(_abc_40319_new_n4703_), .B(_abc_40319_new_n4512_), .Y(_abc_40319_new_n4708_));
AND2X2 AND2X2_2073 ( .A(_abc_40319_new_n4709_), .B(_abc_40319_new_n4710_), .Y(_abc_40319_new_n4711_));
AND2X2 AND2X2_2074 ( .A(_abc_40319_new_n4711_), .B(_abc_40319_new_n4272_), .Y(_abc_40319_new_n4712_));
AND2X2 AND2X2_2075 ( .A(_abc_40319_new_n4518_), .B(_abc_40319_new_n1285_), .Y(_abc_40319_new_n4713_));
AND2X2 AND2X2_2076 ( .A(_abc_40319_new_n1310_), .B(_abc_40319_new_n1169_), .Y(_abc_40319_new_n4714_));
AND2X2 AND2X2_2077 ( .A(_abc_40319_new_n1306_), .B(_abc_40319_new_n1152_), .Y(_abc_40319_new_n4716_));
AND2X2 AND2X2_2078 ( .A(_abc_40319_new_n4717_), .B(_abc_40319_new_n4715_), .Y(_abc_40319_new_n4718_));
AND2X2 AND2X2_2079 ( .A(_abc_40319_new_n4687_), .B(_abc_40319_new_n3200_), .Y(_abc_40319_new_n4725_));
AND2X2 AND2X2_208 ( .A(_abc_40319_new_n963_), .B(_abc_40319_new_n957_), .Y(_abc_40319_new_n964_));
AND2X2 AND2X2_2080 ( .A(_abc_40319_new_n4726_), .B(_abc_40319_new_n3199_), .Y(_abc_40319_new_n4727_));
AND2X2 AND2X2_2081 ( .A(_abc_40319_new_n4728_), .B(_abc_40319_new_n4507_), .Y(_abc_40319_new_n4729_));
AND2X2 AND2X2_2082 ( .A(_abc_40319_new_n1876_), .B(_abc_40319_new_n4499_), .Y(_abc_40319_new_n4730_));
AND2X2 AND2X2_2083 ( .A(_abc_40319_new_n4731_), .B(_abc_40319_new_n3200_), .Y(_abc_40319_new_n4732_));
AND2X2 AND2X2_2084 ( .A(_abc_40319_new_n4472_), .B(_abc_40319_new_n3199_), .Y(_abc_40319_new_n4733_));
AND2X2 AND2X2_2085 ( .A(_abc_40319_new_n4734_), .B(_abc_40319_new_n4497_), .Y(_abc_40319_new_n4735_));
AND2X2 AND2X2_2086 ( .A(_abc_40319_new_n4737_), .B(_abc_40319_new_n4271_), .Y(_abc_40319_new_n4738_));
AND2X2 AND2X2_2087 ( .A(_abc_40319_new_n4734_), .B(_abc_40319_new_n4512_), .Y(_abc_40319_new_n4739_));
AND2X2 AND2X2_2088 ( .A(_abc_40319_new_n4740_), .B(_abc_40319_new_n4741_), .Y(_abc_40319_new_n4742_));
AND2X2 AND2X2_2089 ( .A(_abc_40319_new_n4742_), .B(_abc_40319_new_n4272_), .Y(_abc_40319_new_n4743_));
AND2X2 AND2X2_209 ( .A(_abc_40319_new_n965_), .B(_abc_40319_new_n935_), .Y(_abc_40319_new_n966_));
AND2X2 AND2X2_2090 ( .A(_abc_40319_new_n4518_), .B(_abc_40319_new_n1317_), .Y(_abc_40319_new_n4744_));
AND2X2 AND2X2_2091 ( .A(_abc_40319_new_n1329_), .B(_abc_40319_new_n1152_), .Y(_abc_40319_new_n4746_));
AND2X2 AND2X2_2092 ( .A(_abc_40319_new_n4747_), .B(_abc_40319_new_n4745_), .Y(_abc_40319_new_n4748_));
AND2X2 AND2X2_2093 ( .A(_abc_40319_new_n1333_), .B(_abc_40319_new_n1169_), .Y(_abc_40319_new_n4749_));
AND2X2 AND2X2_2094 ( .A(_abc_40319_new_n4756_), .B(_abc_40319_new_n4468_), .Y(_abc_40319_new_n4757_));
AND2X2 AND2X2_2095 ( .A(_abc_40319_new_n4758_), .B(_abc_40319_new_n4366_), .Y(_abc_40319_new_n4759_));
AND2X2 AND2X2_2096 ( .A(_abc_40319_new_n4760_), .B(_abc_40319_new_n4355_), .Y(_abc_40319_new_n4761_));
AND2X2 AND2X2_2097 ( .A(_abc_40319_new_n4765_), .B(_abc_40319_new_n4763_), .Y(_abc_40319_new_n4766_));
AND2X2 AND2X2_2098 ( .A(_abc_40319_new_n4766_), .B(_abc_40319_new_n4497_), .Y(_abc_40319_new_n4767_));
AND2X2 AND2X2_2099 ( .A(_abc_40319_new_n1852_), .B(_abc_40319_new_n4499_), .Y(_abc_40319_new_n4768_));
AND2X2 AND2X2_21 ( .A(_abc_40319_new_n570_), .B(_abc_40319_new_n554_), .Y(_abc_40319_new_n571_));
AND2X2 AND2X2_210 ( .A(_abc_40319_new_n967_), .B(_abc_40319_new_n916_), .Y(_abc_40319_new_n968_));
AND2X2 AND2X2_2100 ( .A(_abc_40319_new_n4770_), .B(_abc_40319_new_n4507_), .Y(_abc_40319_new_n4771_));
AND2X2 AND2X2_2101 ( .A(_abc_40319_new_n4771_), .B(_abc_40319_new_n4769_), .Y(_abc_40319_new_n4772_));
AND2X2 AND2X2_2102 ( .A(_abc_40319_new_n4774_), .B(_abc_40319_new_n4271_), .Y(_abc_40319_new_n4775_));
AND2X2 AND2X2_2103 ( .A(_abc_40319_new_n4766_), .B(_abc_40319_new_n4512_), .Y(_abc_40319_new_n4776_));
AND2X2 AND2X2_2104 ( .A(_abc_40319_new_n4777_), .B(_abc_40319_new_n4778_), .Y(_abc_40319_new_n4779_));
AND2X2 AND2X2_2105 ( .A(_abc_40319_new_n4779_), .B(_abc_40319_new_n4272_), .Y(_abc_40319_new_n4780_));
AND2X2 AND2X2_2106 ( .A(_abc_40319_new_n4518_), .B(_abc_40319_new_n1340_), .Y(_abc_40319_new_n4781_));
AND2X2 AND2X2_2107 ( .A(_abc_40319_new_n1169_), .B(_abc_40319_new_n1869_), .Y(_abc_40319_new_n4782_));
AND2X2 AND2X2_2108 ( .A(_abc_40319_new_n4309_), .B(REG2_REG_21_), .Y(_abc_40319_new_n4784_));
AND2X2 AND2X2_2109 ( .A(_abc_40319_new_n1865_), .B(_abc_40319_new_n1152_), .Y(_abc_40319_new_n4785_));
AND2X2 AND2X2_211 ( .A(_abc_40319_new_n969_), .B(_abc_40319_new_n970_), .Y(_abc_40319_new_n971_));
AND2X2 AND2X2_2110 ( .A(_abc_40319_new_n4271_), .B(_abc_40319_new_n4785_), .Y(_abc_40319_new_n4786_));
AND2X2 AND2X2_2111 ( .A(_abc_40319_new_n4760_), .B(_abc_40319_new_n4353_), .Y(_abc_40319_new_n4793_));
AND2X2 AND2X2_2112 ( .A(_abc_40319_new_n4796_), .B(_abc_40319_new_n4798_), .Y(_abc_40319_new_n4799_));
AND2X2 AND2X2_2113 ( .A(_abc_40319_new_n4799_), .B(_abc_40319_new_n4497_), .Y(_abc_40319_new_n4800_));
AND2X2 AND2X2_2114 ( .A(_abc_40319_new_n1828_), .B(_abc_40319_new_n4499_), .Y(_abc_40319_new_n4801_));
AND2X2 AND2X2_2115 ( .A(_abc_40319_new_n4645_), .B(_abc_40319_new_n3472_), .Y(_abc_40319_new_n4802_));
AND2X2 AND2X2_2116 ( .A(_abc_40319_new_n4806_), .B(_abc_40319_new_n4507_), .Y(_abc_40319_new_n4807_));
AND2X2 AND2X2_2117 ( .A(_abc_40319_new_n4807_), .B(_abc_40319_new_n4804_), .Y(_abc_40319_new_n4808_));
AND2X2 AND2X2_2118 ( .A(_abc_40319_new_n4810_), .B(_abc_40319_new_n4271_), .Y(_abc_40319_new_n4811_));
AND2X2 AND2X2_2119 ( .A(_abc_40319_new_n4799_), .B(_abc_40319_new_n4512_), .Y(_abc_40319_new_n4812_));
AND2X2 AND2X2_212 ( .A(_abc_40319_new_n974_), .B(_abc_40319_new_n973_), .Y(_abc_40319_new_n975_));
AND2X2 AND2X2_2120 ( .A(_abc_40319_new_n4813_), .B(_abc_40319_new_n4814_), .Y(_abc_40319_new_n4815_));
AND2X2 AND2X2_2121 ( .A(_abc_40319_new_n4815_), .B(_abc_40319_new_n4272_), .Y(_abc_40319_new_n4816_));
AND2X2 AND2X2_2122 ( .A(_abc_40319_new_n4518_), .B(_abc_40319_new_n1876_), .Y(_abc_40319_new_n4817_));
AND2X2 AND2X2_2123 ( .A(_abc_40319_new_n1841_), .B(_abc_40319_new_n1152_), .Y(_abc_40319_new_n4818_));
AND2X2 AND2X2_2124 ( .A(_abc_40319_new_n4271_), .B(_abc_40319_new_n4818_), .Y(_abc_40319_new_n4819_));
AND2X2 AND2X2_2125 ( .A(_abc_40319_new_n4309_), .B(REG2_REG_20_), .Y(_abc_40319_new_n4820_));
AND2X2 AND2X2_2126 ( .A(_abc_40319_new_n1169_), .B(_abc_40319_new_n1846_), .Y(_abc_40319_new_n4821_));
AND2X2 AND2X2_2127 ( .A(_abc_40319_new_n4760_), .B(_abc_40319_new_n3190_), .Y(_abc_40319_new_n4829_));
AND2X2 AND2X2_2128 ( .A(_abc_40319_new_n4830_), .B(_abc_40319_new_n3189_), .Y(_abc_40319_new_n4831_));
AND2X2 AND2X2_2129 ( .A(_abc_40319_new_n4832_), .B(_abc_40319_new_n4497_), .Y(_abc_40319_new_n4833_));
AND2X2 AND2X2_213 ( .A(_abc_40319_new_n975_), .B(_abc_40319_new_n972_), .Y(_abc_40319_new_n976_));
AND2X2 AND2X2_2130 ( .A(_abc_40319_new_n1374_), .B(_abc_40319_new_n4499_), .Y(_abc_40319_new_n4834_));
AND2X2 AND2X2_2131 ( .A(_abc_40319_new_n4837_), .B(_abc_40319_new_n4507_), .Y(_abc_40319_new_n4838_));
AND2X2 AND2X2_2132 ( .A(_abc_40319_new_n4838_), .B(_abc_40319_new_n4836_), .Y(_abc_40319_new_n4839_));
AND2X2 AND2X2_2133 ( .A(_abc_40319_new_n4841_), .B(_abc_40319_new_n4271_), .Y(_abc_40319_new_n4842_));
AND2X2 AND2X2_2134 ( .A(_abc_40319_new_n4832_), .B(_abc_40319_new_n4512_), .Y(_abc_40319_new_n4843_));
AND2X2 AND2X2_2135 ( .A(_abc_40319_new_n4844_), .B(_abc_40319_new_n4845_), .Y(_abc_40319_new_n4846_));
AND2X2 AND2X2_2136 ( .A(_abc_40319_new_n4846_), .B(_abc_40319_new_n4272_), .Y(_abc_40319_new_n4847_));
AND2X2 AND2X2_2137 ( .A(_abc_40319_new_n4518_), .B(_abc_40319_new_n1852_), .Y(_abc_40319_new_n4848_));
AND2X2 AND2X2_2138 ( .A(_abc_40319_new_n4309_), .B(REG2_REG_19_), .Y(_abc_40319_new_n4849_));
AND2X2 AND2X2_2139 ( .A(_abc_40319_new_n1817_), .B(_abc_40319_new_n1152_), .Y(_abc_40319_new_n4850_));
AND2X2 AND2X2_214 ( .A(_abc_40319_new_n978_), .B(_abc_40319_new_n968_), .Y(_abc_40319_new_n979_));
AND2X2 AND2X2_2140 ( .A(_abc_40319_new_n4271_), .B(_abc_40319_new_n4850_), .Y(_abc_40319_new_n4851_));
AND2X2 AND2X2_2141 ( .A(_abc_40319_new_n1169_), .B(_abc_40319_new_n1822_), .Y(_abc_40319_new_n4852_));
AND2X2 AND2X2_2142 ( .A(_abc_40319_new_n4860_), .B(_abc_40319_new_n3153_), .Y(_abc_40319_new_n4861_));
AND2X2 AND2X2_2143 ( .A(_abc_40319_new_n4758_), .B(_abc_40319_new_n3154_), .Y(_abc_40319_new_n4862_));
AND2X2 AND2X2_2144 ( .A(_abc_40319_new_n4863_), .B(_abc_40319_new_n4497_), .Y(_abc_40319_new_n4864_));
AND2X2 AND2X2_2145 ( .A(_abc_40319_new_n1444_), .B(_abc_40319_new_n4499_), .Y(_abc_40319_new_n4865_));
AND2X2 AND2X2_2146 ( .A(_abc_40319_new_n4643_), .B(_abc_40319_new_n3402_), .Y(_abc_40319_new_n4866_));
AND2X2 AND2X2_2147 ( .A(_abc_40319_new_n4869_), .B(_abc_40319_new_n4507_), .Y(_abc_40319_new_n4870_));
AND2X2 AND2X2_2148 ( .A(_abc_40319_new_n4870_), .B(_abc_40319_new_n4868_), .Y(_abc_40319_new_n4871_));
AND2X2 AND2X2_2149 ( .A(_abc_40319_new_n4873_), .B(_abc_40319_new_n4271_), .Y(_abc_40319_new_n4874_));
AND2X2 AND2X2_215 ( .A(_abc_40319_new_n980_), .B(_abc_40319_new_n807_), .Y(_abc_40319_new_n981_));
AND2X2 AND2X2_2150 ( .A(_abc_40319_new_n4863_), .B(_abc_40319_new_n4512_), .Y(_abc_40319_new_n4875_));
AND2X2 AND2X2_2151 ( .A(_abc_40319_new_n4876_), .B(_abc_40319_new_n4877_), .Y(_abc_40319_new_n4878_));
AND2X2 AND2X2_2152 ( .A(_abc_40319_new_n4878_), .B(_abc_40319_new_n4272_), .Y(_abc_40319_new_n4879_));
AND2X2 AND2X2_2153 ( .A(_abc_40319_new_n4518_), .B(_abc_40319_new_n1828_), .Y(_abc_40319_new_n4880_));
AND2X2 AND2X2_2154 ( .A(_abc_40319_new_n4309_), .B(REG2_REG_18_), .Y(_abc_40319_new_n4881_));
AND2X2 AND2X2_2155 ( .A(_abc_40319_new_n1363_), .B(_abc_40319_new_n1152_), .Y(_abc_40319_new_n4882_));
AND2X2 AND2X2_2156 ( .A(_abc_40319_new_n4271_), .B(_abc_40319_new_n4882_), .Y(_abc_40319_new_n4883_));
AND2X2 AND2X2_2157 ( .A(_abc_40319_new_n1169_), .B(_abc_40319_new_n1368_), .Y(_abc_40319_new_n4884_));
AND2X2 AND2X2_2158 ( .A(_abc_40319_new_n4756_), .B(_abc_40319_new_n4892_), .Y(_abc_40319_new_n4893_));
AND2X2 AND2X2_2159 ( .A(_abc_40319_new_n4897_), .B(_abc_40319_new_n4895_), .Y(_abc_40319_new_n4898_));
AND2X2 AND2X2_216 ( .A(_abc_40319_new_n982_), .B(_abc_40319_new_n773_), .Y(_abc_40319_new_n983_));
AND2X2 AND2X2_2160 ( .A(_abc_40319_new_n4898_), .B(_abc_40319_new_n4497_), .Y(_abc_40319_new_n4899_));
AND2X2 AND2X2_2161 ( .A(_abc_40319_new_n1410_), .B(_abc_40319_new_n4499_), .Y(_abc_40319_new_n4900_));
AND2X2 AND2X2_2162 ( .A(_abc_40319_new_n3519_), .B(_abc_40319_new_n3524_), .Y(_abc_40319_new_n4901_));
AND2X2 AND2X2_2163 ( .A(_abc_40319_new_n4904_), .B(_abc_40319_new_n4507_), .Y(_abc_40319_new_n4905_));
AND2X2 AND2X2_2164 ( .A(_abc_40319_new_n4905_), .B(_abc_40319_new_n4903_), .Y(_abc_40319_new_n4906_));
AND2X2 AND2X2_2165 ( .A(_abc_40319_new_n4908_), .B(_abc_40319_new_n4271_), .Y(_abc_40319_new_n4909_));
AND2X2 AND2X2_2166 ( .A(_abc_40319_new_n4898_), .B(_abc_40319_new_n4512_), .Y(_abc_40319_new_n4910_));
AND2X2 AND2X2_2167 ( .A(_abc_40319_new_n4911_), .B(_abc_40319_new_n4912_), .Y(_abc_40319_new_n4913_));
AND2X2 AND2X2_2168 ( .A(_abc_40319_new_n4913_), .B(_abc_40319_new_n4272_), .Y(_abc_40319_new_n4914_));
AND2X2 AND2X2_2169 ( .A(_abc_40319_new_n1374_), .B(_abc_40319_new_n4310_), .Y(_abc_40319_new_n4915_));
AND2X2 AND2X2_217 ( .A(_abc_40319_new_n537_), .B(_abc_40319_new_n549_), .Y(_abc_40319_new_n986_));
AND2X2 AND2X2_2170 ( .A(_abc_40319_new_n4271_), .B(_abc_40319_new_n4915_), .Y(_abc_40319_new_n4916_));
AND2X2 AND2X2_2171 ( .A(_abc_40319_new_n1433_), .B(_abc_40319_new_n1152_), .Y(_abc_40319_new_n4917_));
AND2X2 AND2X2_2172 ( .A(_abc_40319_new_n4271_), .B(_abc_40319_new_n4917_), .Y(_abc_40319_new_n4918_));
AND2X2 AND2X2_2173 ( .A(_abc_40319_new_n4309_), .B(REG2_REG_17_), .Y(_abc_40319_new_n4919_));
AND2X2 AND2X2_2174 ( .A(_abc_40319_new_n1169_), .B(_abc_40319_new_n1440_), .Y(_abc_40319_new_n4920_));
AND2X2 AND2X2_2175 ( .A(_abc_40319_new_n4928_), .B(_abc_40319_new_n3476_), .Y(_abc_40319_new_n4929_));
AND2X2 AND2X2_2176 ( .A(_abc_40319_new_n4930_), .B(_abc_40319_new_n3478_), .Y(_abc_40319_new_n4931_));
AND2X2 AND2X2_2177 ( .A(_abc_40319_new_n4932_), .B(_abc_40319_new_n3231_), .Y(_abc_40319_new_n4933_));
AND2X2 AND2X2_2178 ( .A(_abc_40319_new_n4934_), .B(_abc_40319_new_n3232_), .Y(_abc_40319_new_n4935_));
AND2X2 AND2X2_2179 ( .A(_abc_40319_new_n4936_), .B(_abc_40319_new_n4507_), .Y(_abc_40319_new_n4937_));
AND2X2 AND2X2_218 ( .A(_abc_40319_new_n987_), .B(IR_REG_6_), .Y(_abc_40319_new_n988_));
AND2X2 AND2X2_2180 ( .A(_abc_40319_new_n1483_), .B(_abc_40319_new_n4499_), .Y(_abc_40319_new_n4938_));
AND2X2 AND2X2_2181 ( .A(_abc_40319_new_n4756_), .B(_abc_40319_new_n3232_), .Y(_abc_40319_new_n4939_));
AND2X2 AND2X2_2182 ( .A(_abc_40319_new_n4464_), .B(_abc_40319_new_n3231_), .Y(_abc_40319_new_n4940_));
AND2X2 AND2X2_2183 ( .A(_abc_40319_new_n4941_), .B(_abc_40319_new_n4497_), .Y(_abc_40319_new_n4942_));
AND2X2 AND2X2_2184 ( .A(_abc_40319_new_n4944_), .B(_abc_40319_new_n4271_), .Y(_abc_40319_new_n4945_));
AND2X2 AND2X2_2185 ( .A(_abc_40319_new_n4941_), .B(_abc_40319_new_n4512_), .Y(_abc_40319_new_n4946_));
AND2X2 AND2X2_2186 ( .A(_abc_40319_new_n4947_), .B(_abc_40319_new_n4948_), .Y(_abc_40319_new_n4949_));
AND2X2 AND2X2_2187 ( .A(_abc_40319_new_n4949_), .B(_abc_40319_new_n4272_), .Y(_abc_40319_new_n4950_));
AND2X2 AND2X2_2188 ( .A(_abc_40319_new_n1444_), .B(_abc_40319_new_n4310_), .Y(_abc_40319_new_n4951_));
AND2X2 AND2X2_2189 ( .A(_abc_40319_new_n4271_), .B(_abc_40319_new_n4951_), .Y(_abc_40319_new_n4952_));
AND2X2 AND2X2_219 ( .A(_abc_40319_new_n990_), .B(IR_REG_31_), .Y(_abc_40319_new_n991_));
AND2X2 AND2X2_2190 ( .A(_abc_40319_new_n1169_), .B(_abc_40319_new_n1406_), .Y(_abc_40319_new_n4953_));
AND2X2 AND2X2_2191 ( .A(_abc_40319_new_n1398_), .B(_abc_40319_new_n1152_), .Y(_abc_40319_new_n4956_));
AND2X2 AND2X2_2192 ( .A(_abc_40319_new_n4271_), .B(_abc_40319_new_n4956_), .Y(_abc_40319_new_n4957_));
AND2X2 AND2X2_2193 ( .A(_abc_40319_new_n4309_), .B(REG2_REG_16_), .Y(_abc_40319_new_n4958_));
AND2X2 AND2X2_2194 ( .A(_abc_40319_new_n4930_), .B(_abc_40319_new_n3113_), .Y(_abc_40319_new_n4964_));
AND2X2 AND2X2_2195 ( .A(_abc_40319_new_n4965_), .B(_abc_40319_new_n3114_), .Y(_abc_40319_new_n4966_));
AND2X2 AND2X2_2196 ( .A(_abc_40319_new_n4967_), .B(_abc_40319_new_n4507_), .Y(_abc_40319_new_n4968_));
AND2X2 AND2X2_2197 ( .A(_abc_40319_new_n1517_), .B(_abc_40319_new_n4499_), .Y(_abc_40319_new_n4969_));
AND2X2 AND2X2_2198 ( .A(_abc_40319_new_n4970_), .B(_abc_40319_new_n3114_), .Y(_abc_40319_new_n4971_));
AND2X2 AND2X2_2199 ( .A(_abc_40319_new_n4462_), .B(_abc_40319_new_n3113_), .Y(_abc_40319_new_n4972_));
AND2X2 AND2X2_22 ( .A(_abc_40319_new_n571_), .B(_abc_40319_new_n553_), .Y(_abc_40319_new_n572_));
AND2X2 AND2X2_220 ( .A(_abc_40319_new_n524_), .B(IR_REG_6_), .Y(_abc_40319_new_n992_));
AND2X2 AND2X2_2200 ( .A(_abc_40319_new_n4973_), .B(_abc_40319_new_n4497_), .Y(_abc_40319_new_n4974_));
AND2X2 AND2X2_2201 ( .A(_abc_40319_new_n4976_), .B(_abc_40319_new_n4271_), .Y(_abc_40319_new_n4977_));
AND2X2 AND2X2_2202 ( .A(_abc_40319_new_n4973_), .B(_abc_40319_new_n4512_), .Y(_abc_40319_new_n4978_));
AND2X2 AND2X2_2203 ( .A(_abc_40319_new_n4979_), .B(_abc_40319_new_n4980_), .Y(_abc_40319_new_n4981_));
AND2X2 AND2X2_2204 ( .A(_abc_40319_new_n4981_), .B(_abc_40319_new_n4272_), .Y(_abc_40319_new_n4982_));
AND2X2 AND2X2_2205 ( .A(_abc_40319_new_n1410_), .B(_abc_40319_new_n4310_), .Y(_abc_40319_new_n4984_));
AND2X2 AND2X2_2206 ( .A(_abc_40319_new_n1471_), .B(_abc_40319_new_n1152_), .Y(_abc_40319_new_n4985_));
AND2X2 AND2X2_2207 ( .A(_abc_40319_new_n4987_), .B(_abc_40319_new_n4983_), .Y(_abc_40319_new_n4988_));
AND2X2 AND2X2_2208 ( .A(_abc_40319_new_n1169_), .B(_abc_40319_new_n1480_), .Y(_abc_40319_new_n4989_));
AND2X2 AND2X2_2209 ( .A(_abc_40319_new_n4995_), .B(_abc_40319_new_n4996_), .Y(_abc_40319_new_n4997_));
AND2X2 AND2X2_221 ( .A(_abc_40319_new_n640_), .B(_abc_40319_new_n994_), .Y(_abc_40319_new_n995_));
AND2X2 AND2X2_2210 ( .A(_abc_40319_new_n4997_), .B(_abc_40319_new_n4507_), .Y(_abc_40319_new_n4998_));
AND2X2 AND2X2_2211 ( .A(_abc_40319_new_n1667_), .B(_abc_40319_new_n4499_), .Y(_abc_40319_new_n4999_));
AND2X2 AND2X2_2212 ( .A(_abc_40319_new_n4459_), .B(_abc_40319_new_n3147_), .Y(_abc_40319_new_n5000_));
AND2X2 AND2X2_2213 ( .A(_abc_40319_new_n4460_), .B(_abc_40319_new_n3146_), .Y(_abc_40319_new_n5001_));
AND2X2 AND2X2_2214 ( .A(_abc_40319_new_n5002_), .B(_abc_40319_new_n4497_), .Y(_abc_40319_new_n5003_));
AND2X2 AND2X2_2215 ( .A(_abc_40319_new_n5005_), .B(_abc_40319_new_n4271_), .Y(_abc_40319_new_n5006_));
AND2X2 AND2X2_2216 ( .A(_abc_40319_new_n5002_), .B(_abc_40319_new_n4512_), .Y(_abc_40319_new_n5007_));
AND2X2 AND2X2_2217 ( .A(_abc_40319_new_n5008_), .B(_abc_40319_new_n5009_), .Y(_abc_40319_new_n5010_));
AND2X2 AND2X2_2218 ( .A(_abc_40319_new_n5010_), .B(_abc_40319_new_n4272_), .Y(_abc_40319_new_n5011_));
AND2X2 AND2X2_2219 ( .A(_abc_40319_new_n1506_), .B(_abc_40319_new_n1152_), .Y(_abc_40319_new_n5012_));
AND2X2 AND2X2_222 ( .A(_abc_40319_new_n996_), .B(_abc_40319_new_n997_), .Y(_abc_40319_new_n998_));
AND2X2 AND2X2_2220 ( .A(_abc_40319_new_n1483_), .B(_abc_40319_new_n4310_), .Y(_abc_40319_new_n5013_));
AND2X2 AND2X2_2221 ( .A(_abc_40319_new_n4271_), .B(_abc_40319_new_n5014_), .Y(_abc_40319_new_n5015_));
AND2X2 AND2X2_2222 ( .A(_abc_40319_new_n4309_), .B(REG2_REG_14_), .Y(_abc_40319_new_n5016_));
AND2X2 AND2X2_2223 ( .A(_abc_40319_new_n1169_), .B(_abc_40319_new_n1513_), .Y(_abc_40319_new_n5017_));
AND2X2 AND2X2_2224 ( .A(_abc_40319_new_n5024_), .B(_abc_40319_new_n3142_), .Y(_abc_40319_new_n5025_));
AND2X2 AND2X2_2225 ( .A(_abc_40319_new_n3516_), .B(_abc_40319_new_n3143_), .Y(_abc_40319_new_n5026_));
AND2X2 AND2X2_2226 ( .A(_abc_40319_new_n5027_), .B(_abc_40319_new_n4507_), .Y(_abc_40319_new_n5028_));
AND2X2 AND2X2_2227 ( .A(_abc_40319_new_n1701_), .B(_abc_40319_new_n4499_), .Y(_abc_40319_new_n5029_));
AND2X2 AND2X2_2228 ( .A(_abc_40319_new_n5030_), .B(_abc_40319_new_n4389_), .Y(_abc_40319_new_n5031_));
AND2X2 AND2X2_2229 ( .A(_abc_40319_new_n5035_), .B(_abc_40319_new_n5033_), .Y(_abc_40319_new_n5036_));
AND2X2 AND2X2_223 ( .A(_abc_40319_new_n998_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n999_));
AND2X2 AND2X2_2230 ( .A(_abc_40319_new_n5036_), .B(_abc_40319_new_n4497_), .Y(_abc_40319_new_n5037_));
AND2X2 AND2X2_2231 ( .A(_abc_40319_new_n5039_), .B(_abc_40319_new_n4271_), .Y(_abc_40319_new_n5040_));
AND2X2 AND2X2_2232 ( .A(_abc_40319_new_n5036_), .B(_abc_40319_new_n4512_), .Y(_abc_40319_new_n5041_));
AND2X2 AND2X2_2233 ( .A(_abc_40319_new_n5042_), .B(_abc_40319_new_n5043_), .Y(_abc_40319_new_n5044_));
AND2X2 AND2X2_2234 ( .A(_abc_40319_new_n5044_), .B(_abc_40319_new_n4272_), .Y(_abc_40319_new_n5045_));
AND2X2 AND2X2_2235 ( .A(_abc_40319_new_n1517_), .B(_abc_40319_new_n4310_), .Y(_abc_40319_new_n5047_));
AND2X2 AND2X2_2236 ( .A(_abc_40319_new_n1655_), .B(_abc_40319_new_n1152_), .Y(_abc_40319_new_n5048_));
AND2X2 AND2X2_2237 ( .A(_abc_40319_new_n5050_), .B(_abc_40319_new_n5046_), .Y(_abc_40319_new_n5051_));
AND2X2 AND2X2_2238 ( .A(_abc_40319_new_n1169_), .B(_abc_40319_new_n1660_), .Y(_abc_40319_new_n5052_));
AND2X2 AND2X2_2239 ( .A(_abc_40319_new_n5058_), .B(_abc_40319_new_n3235_), .Y(_abc_40319_new_n5059_));
AND2X2 AND2X2_224 ( .A(_abc_40319_new_n740_), .B(REG3_REG_6_), .Y(_abc_40319_new_n1000_));
AND2X2 AND2X2_2240 ( .A(_abc_40319_new_n3514_), .B(_abc_40319_new_n3236_), .Y(_abc_40319_new_n5060_));
AND2X2 AND2X2_2241 ( .A(_abc_40319_new_n5061_), .B(_abc_40319_new_n4507_), .Y(_abc_40319_new_n5062_));
AND2X2 AND2X2_2242 ( .A(_abc_40319_new_n1735_), .B(_abc_40319_new_n4499_), .Y(_abc_40319_new_n5063_));
AND2X2 AND2X2_2243 ( .A(_abc_40319_new_n5030_), .B(_abc_40319_new_n3236_), .Y(_abc_40319_new_n5064_));
AND2X2 AND2X2_2244 ( .A(_abc_40319_new_n5065_), .B(_abc_40319_new_n3235_), .Y(_abc_40319_new_n5066_));
AND2X2 AND2X2_2245 ( .A(_abc_40319_new_n5067_), .B(_abc_40319_new_n4497_), .Y(_abc_40319_new_n5068_));
AND2X2 AND2X2_2246 ( .A(_abc_40319_new_n5070_), .B(_abc_40319_new_n4271_), .Y(_abc_40319_new_n5071_));
AND2X2 AND2X2_2247 ( .A(_abc_40319_new_n5067_), .B(_abc_40319_new_n4512_), .Y(_abc_40319_new_n5072_));
AND2X2 AND2X2_2248 ( .A(_abc_40319_new_n5073_), .B(_abc_40319_new_n5074_), .Y(_abc_40319_new_n5075_));
AND2X2 AND2X2_2249 ( .A(_abc_40319_new_n5075_), .B(_abc_40319_new_n4272_), .Y(_abc_40319_new_n5076_));
AND2X2 AND2X2_225 ( .A(_abc_40319_new_n1001_), .B(_abc_40319_new_n1002_), .Y(_abc_40319_new_n1003_));
AND2X2 AND2X2_2250 ( .A(_abc_40319_new_n1667_), .B(_abc_40319_new_n4310_), .Y(_abc_40319_new_n5078_));
AND2X2 AND2X2_2251 ( .A(_abc_40319_new_n1690_), .B(_abc_40319_new_n1152_), .Y(_abc_40319_new_n5079_));
AND2X2 AND2X2_2252 ( .A(_abc_40319_new_n5081_), .B(_abc_40319_new_n5077_), .Y(_abc_40319_new_n5082_));
AND2X2 AND2X2_2253 ( .A(_abc_40319_new_n1169_), .B(_abc_40319_new_n1698_), .Y(_abc_40319_new_n5083_));
AND2X2 AND2X2_2254 ( .A(_abc_40319_new_n5089_), .B(_abc_40319_new_n3510_), .Y(_abc_40319_new_n5090_));
AND2X2 AND2X2_2255 ( .A(_abc_40319_new_n5091_), .B(_abc_40319_new_n3484_), .Y(_abc_40319_new_n5092_));
AND2X2 AND2X2_2256 ( .A(_abc_40319_new_n5093_), .B(_abc_40319_new_n3226_), .Y(_abc_40319_new_n5094_));
AND2X2 AND2X2_2257 ( .A(_abc_40319_new_n5095_), .B(_abc_40319_new_n3227_), .Y(_abc_40319_new_n5096_));
AND2X2 AND2X2_2258 ( .A(_abc_40319_new_n5097_), .B(_abc_40319_new_n4507_), .Y(_abc_40319_new_n5098_));
AND2X2 AND2X2_2259 ( .A(_abc_40319_new_n1769_), .B(_abc_40319_new_n4499_), .Y(_abc_40319_new_n5099_));
AND2X2 AND2X2_226 ( .A(_abc_40319_new_n738_), .B(_abc_40319_new_n1003_), .Y(_abc_40319_new_n1004_));
AND2X2 AND2X2_2260 ( .A(_abc_40319_new_n5102_), .B(_abc_40319_new_n5100_), .Y(_abc_40319_new_n5103_));
AND2X2 AND2X2_2261 ( .A(_abc_40319_new_n5103_), .B(_abc_40319_new_n4497_), .Y(_abc_40319_new_n5104_));
AND2X2 AND2X2_2262 ( .A(_abc_40319_new_n5106_), .B(_abc_40319_new_n4271_), .Y(_abc_40319_new_n5107_));
AND2X2 AND2X2_2263 ( .A(_abc_40319_new_n5103_), .B(_abc_40319_new_n4512_), .Y(_abc_40319_new_n5108_));
AND2X2 AND2X2_2264 ( .A(_abc_40319_new_n5109_), .B(_abc_40319_new_n5110_), .Y(_abc_40319_new_n5111_));
AND2X2 AND2X2_2265 ( .A(_abc_40319_new_n5111_), .B(_abc_40319_new_n4272_), .Y(_abc_40319_new_n5112_));
AND2X2 AND2X2_2266 ( .A(_abc_40319_new_n1724_), .B(_abc_40319_new_n1152_), .Y(_abc_40319_new_n5113_));
AND2X2 AND2X2_2267 ( .A(_abc_40319_new_n1701_), .B(_abc_40319_new_n4310_), .Y(_abc_40319_new_n5114_));
AND2X2 AND2X2_2268 ( .A(_abc_40319_new_n4271_), .B(_abc_40319_new_n5115_), .Y(_abc_40319_new_n5116_));
AND2X2 AND2X2_2269 ( .A(_abc_40319_new_n4309_), .B(REG2_REG_11_), .Y(_abc_40319_new_n5117_));
AND2X2 AND2X2_227 ( .A(_abc_40319_new_n722_), .B(REG1_REG_6_), .Y(_abc_40319_new_n1005_));
AND2X2 AND2X2_2270 ( .A(_abc_40319_new_n1169_), .B(_abc_40319_new_n1732_), .Y(_abc_40319_new_n5118_));
AND2X2 AND2X2_2271 ( .A(_abc_40319_new_n5091_), .B(_abc_40319_new_n3207_), .Y(_abc_40319_new_n5125_));
AND2X2 AND2X2_2272 ( .A(_abc_40319_new_n5126_), .B(_abc_40319_new_n3208_), .Y(_abc_40319_new_n5127_));
AND2X2 AND2X2_2273 ( .A(_abc_40319_new_n5128_), .B(_abc_40319_new_n4507_), .Y(_abc_40319_new_n5129_));
AND2X2 AND2X2_2274 ( .A(_abc_40319_new_n1625_), .B(_abc_40319_new_n4499_), .Y(_abc_40319_new_n5130_));
AND2X2 AND2X2_2275 ( .A(_abc_40319_new_n5132_), .B(_abc_40319_new_n4402_), .Y(_abc_40319_new_n5133_));
AND2X2 AND2X2_2276 ( .A(_abc_40319_new_n5136_), .B(_abc_40319_new_n5134_), .Y(_abc_40319_new_n5137_));
AND2X2 AND2X2_2277 ( .A(_abc_40319_new_n5137_), .B(_abc_40319_new_n4497_), .Y(_abc_40319_new_n5138_));
AND2X2 AND2X2_2278 ( .A(_abc_40319_new_n5140_), .B(_abc_40319_new_n4271_), .Y(_abc_40319_new_n5141_));
AND2X2 AND2X2_2279 ( .A(_abc_40319_new_n5137_), .B(_abc_40319_new_n4512_), .Y(_abc_40319_new_n5142_));
AND2X2 AND2X2_228 ( .A(_abc_40319_new_n736_), .B(REG0_REG_6_), .Y(_abc_40319_new_n1007_));
AND2X2 AND2X2_2280 ( .A(_abc_40319_new_n5143_), .B(_abc_40319_new_n5144_), .Y(_abc_40319_new_n5145_));
AND2X2 AND2X2_2281 ( .A(_abc_40319_new_n5145_), .B(_abc_40319_new_n4272_), .Y(_abc_40319_new_n5146_));
AND2X2 AND2X2_2282 ( .A(_abc_40319_new_n4309_), .B(REG2_REG_10_), .Y(_abc_40319_new_n5147_));
AND2X2 AND2X2_2283 ( .A(_abc_40319_new_n1169_), .B(_abc_40319_new_n1766_), .Y(_abc_40319_new_n5148_));
AND2X2 AND2X2_2284 ( .A(_abc_40319_new_n1758_), .B(_abc_40319_new_n1152_), .Y(_abc_40319_new_n5151_));
AND2X2 AND2X2_2285 ( .A(_abc_40319_new_n4271_), .B(_abc_40319_new_n5151_), .Y(_abc_40319_new_n5152_));
AND2X2 AND2X2_2286 ( .A(_abc_40319_new_n1735_), .B(_abc_40319_new_n4310_), .Y(_abc_40319_new_n5153_));
AND2X2 AND2X2_2287 ( .A(_abc_40319_new_n4271_), .B(_abc_40319_new_n5153_), .Y(_abc_40319_new_n5154_));
AND2X2 AND2X2_2288 ( .A(_abc_40319_new_n5161_), .B(_abc_40319_new_n5160_), .Y(_abc_40319_new_n5162_));
AND2X2 AND2X2_2289 ( .A(_abc_40319_new_n5162_), .B(_abc_40319_new_n4507_), .Y(_abc_40319_new_n5163_));
AND2X2 AND2X2_229 ( .A(_abc_40319_new_n733_), .B(REG2_REG_6_), .Y(_abc_40319_new_n1008_));
AND2X2 AND2X2_2290 ( .A(_abc_40319_new_n1146_), .B(_abc_40319_new_n4499_), .Y(_abc_40319_new_n5164_));
AND2X2 AND2X2_2291 ( .A(_abc_40319_new_n5131_), .B(_abc_40319_new_n3158_), .Y(_abc_40319_new_n5165_));
AND2X2 AND2X2_2292 ( .A(_abc_40319_new_n5166_), .B(_abc_40319_new_n3157_), .Y(_abc_40319_new_n5167_));
AND2X2 AND2X2_2293 ( .A(_abc_40319_new_n5168_), .B(_abc_40319_new_n4497_), .Y(_abc_40319_new_n5169_));
AND2X2 AND2X2_2294 ( .A(_abc_40319_new_n5171_), .B(_abc_40319_new_n4271_), .Y(_abc_40319_new_n5172_));
AND2X2 AND2X2_2295 ( .A(_abc_40319_new_n5168_), .B(_abc_40319_new_n4512_), .Y(_abc_40319_new_n5173_));
AND2X2 AND2X2_2296 ( .A(_abc_40319_new_n5174_), .B(_abc_40319_new_n5175_), .Y(_abc_40319_new_n5176_));
AND2X2 AND2X2_2297 ( .A(_abc_40319_new_n5176_), .B(_abc_40319_new_n4272_), .Y(_abc_40319_new_n5177_));
AND2X2 AND2X2_2298 ( .A(_abc_40319_new_n1614_), .B(_abc_40319_new_n1152_), .Y(_abc_40319_new_n5178_));
AND2X2 AND2X2_2299 ( .A(_abc_40319_new_n1769_), .B(_abc_40319_new_n4310_), .Y(_abc_40319_new_n5179_));
AND2X2 AND2X2_23 ( .A(_abc_40319_new_n573_), .B(_abc_40319_new_n574_), .Y(_abc_40319_new_n575_));
AND2X2 AND2X2_230 ( .A(_abc_40319_new_n705_), .B(_abc_40319_new_n1010_), .Y(_abc_40319_new_n1011_));
AND2X2 AND2X2_2300 ( .A(_abc_40319_new_n4271_), .B(_abc_40319_new_n5180_), .Y(_abc_40319_new_n5181_));
AND2X2 AND2X2_2301 ( .A(_abc_40319_new_n4309_), .B(REG2_REG_9_), .Y(_abc_40319_new_n5182_));
AND2X2 AND2X2_2302 ( .A(_abc_40319_new_n1169_), .B(_abc_40319_new_n1618_), .Y(_abc_40319_new_n5183_));
AND2X2 AND2X2_2303 ( .A(_abc_40319_new_n3506_), .B(_abc_40319_new_n3316_), .Y(_abc_40319_new_n5190_));
AND2X2 AND2X2_2304 ( .A(_abc_40319_new_n5191_), .B(_abc_40319_new_n3176_), .Y(_abc_40319_new_n5192_));
AND2X2 AND2X2_2305 ( .A(_abc_40319_new_n5190_), .B(_abc_40319_new_n3177_), .Y(_abc_40319_new_n5193_));
AND2X2 AND2X2_2306 ( .A(_abc_40319_new_n5194_), .B(_abc_40319_new_n4507_), .Y(_abc_40319_new_n5195_));
AND2X2 AND2X2_2307 ( .A(_abc_40319_new_n1046_), .B(_abc_40319_new_n4499_), .Y(_abc_40319_new_n5196_));
AND2X2 AND2X2_2308 ( .A(_abc_40319_new_n5199_), .B(_abc_40319_new_n5197_), .Y(_abc_40319_new_n5200_));
AND2X2 AND2X2_2309 ( .A(_abc_40319_new_n5200_), .B(_abc_40319_new_n4497_), .Y(_abc_40319_new_n5201_));
AND2X2 AND2X2_231 ( .A(_abc_40319_new_n998_), .B(_abc_40319_new_n763_), .Y(_abc_40319_new_n1014_));
AND2X2 AND2X2_2310 ( .A(_abc_40319_new_n5203_), .B(_abc_40319_new_n4271_), .Y(_abc_40319_new_n5204_));
AND2X2 AND2X2_2311 ( .A(_abc_40319_new_n5200_), .B(_abc_40319_new_n4512_), .Y(_abc_40319_new_n5205_));
AND2X2 AND2X2_2312 ( .A(_abc_40319_new_n5206_), .B(_abc_40319_new_n5207_), .Y(_abc_40319_new_n5208_));
AND2X2 AND2X2_2313 ( .A(_abc_40319_new_n5208_), .B(_abc_40319_new_n4272_), .Y(_abc_40319_new_n5209_));
AND2X2 AND2X2_2314 ( .A(_abc_40319_new_n1572_), .B(_abc_40319_new_n1152_), .Y(_abc_40319_new_n5210_));
AND2X2 AND2X2_2315 ( .A(_abc_40319_new_n1625_), .B(_abc_40319_new_n4310_), .Y(_abc_40319_new_n5211_));
AND2X2 AND2X2_2316 ( .A(_abc_40319_new_n4271_), .B(_abc_40319_new_n5212_), .Y(_abc_40319_new_n5213_));
AND2X2 AND2X2_2317 ( .A(_abc_40319_new_n4309_), .B(REG2_REG_8_), .Y(_abc_40319_new_n5214_));
AND2X2 AND2X2_2318 ( .A(_abc_40319_new_n1169_), .B(_abc_40319_new_n1139_), .Y(_abc_40319_new_n5215_));
AND2X2 AND2X2_2319 ( .A(_abc_40319_new_n5222_), .B(_abc_40319_new_n3211_), .Y(_abc_40319_new_n5223_));
AND2X2 AND2X2_232 ( .A(_abc_40319_new_n1010_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1015_));
AND2X2 AND2X2_2320 ( .A(_abc_40319_new_n3505_), .B(_abc_40319_new_n3212_), .Y(_abc_40319_new_n5224_));
AND2X2 AND2X2_2321 ( .A(_abc_40319_new_n5225_), .B(_abc_40319_new_n4507_), .Y(_abc_40319_new_n5226_));
AND2X2 AND2X2_2322 ( .A(_abc_40319_new_n1010_), .B(_abc_40319_new_n4499_), .Y(_abc_40319_new_n5227_));
AND2X2 AND2X2_2323 ( .A(_abc_40319_new_n4450_), .B(_abc_40319_new_n3212_), .Y(_abc_40319_new_n5228_));
AND2X2 AND2X2_2324 ( .A(_abc_40319_new_n5229_), .B(_abc_40319_new_n3211_), .Y(_abc_40319_new_n5230_));
AND2X2 AND2X2_2325 ( .A(_abc_40319_new_n5231_), .B(_abc_40319_new_n4497_), .Y(_abc_40319_new_n5232_));
AND2X2 AND2X2_2326 ( .A(_abc_40319_new_n5234_), .B(_abc_40319_new_n4271_), .Y(_abc_40319_new_n5235_));
AND2X2 AND2X2_2327 ( .A(_abc_40319_new_n5231_), .B(_abc_40319_new_n4512_), .Y(_abc_40319_new_n5236_));
AND2X2 AND2X2_2328 ( .A(_abc_40319_new_n5237_), .B(_abc_40319_new_n5238_), .Y(_abc_40319_new_n5239_));
AND2X2 AND2X2_2329 ( .A(_abc_40319_new_n5239_), .B(_abc_40319_new_n4272_), .Y(_abc_40319_new_n5240_));
AND2X2 AND2X2_233 ( .A(_abc_40319_new_n1019_), .B(_abc_40319_new_n1017_), .Y(_abc_40319_new_n1020_));
AND2X2 AND2X2_2330 ( .A(_abc_40319_new_n1034_), .B(_abc_40319_new_n1152_), .Y(_abc_40319_new_n5242_));
AND2X2 AND2X2_2331 ( .A(_abc_40319_new_n1146_), .B(_abc_40319_new_n4310_), .Y(_abc_40319_new_n5243_));
AND2X2 AND2X2_2332 ( .A(_abc_40319_new_n5245_), .B(_abc_40319_new_n5241_), .Y(_abc_40319_new_n5246_));
AND2X2 AND2X2_2333 ( .A(_abc_40319_new_n1169_), .B(_abc_40319_new_n1042_), .Y(_abc_40319_new_n5247_));
AND2X2 AND2X2_2334 ( .A(_abc_40319_new_n5253_), .B(_abc_40319_new_n3496_), .Y(_abc_40319_new_n5254_));
AND2X2 AND2X2_2335 ( .A(_abc_40319_new_n5256_), .B(_abc_40319_new_n3332_), .Y(_abc_40319_new_n5257_));
AND2X2 AND2X2_2336 ( .A(_abc_40319_new_n5259_), .B(_abc_40319_new_n3215_), .Y(_abc_40319_new_n5260_));
AND2X2 AND2X2_2337 ( .A(_abc_40319_new_n5258_), .B(_abc_40319_new_n3216_), .Y(_abc_40319_new_n5261_));
AND2X2 AND2X2_2338 ( .A(_abc_40319_new_n5262_), .B(_abc_40319_new_n4507_), .Y(_abc_40319_new_n5263_));
AND2X2 AND2X2_2339 ( .A(_abc_40319_new_n746_), .B(_abc_40319_new_n4499_), .Y(_abc_40319_new_n5264_));
AND2X2 AND2X2_234 ( .A(_abc_40319_new_n985_), .B(_abc_40319_new_n1021_), .Y(_abc_40319_new_n1022_));
AND2X2 AND2X2_2340 ( .A(_abc_40319_new_n4448_), .B(_abc_40319_new_n3216_), .Y(_abc_40319_new_n5265_));
AND2X2 AND2X2_2341 ( .A(_abc_40319_new_n5266_), .B(_abc_40319_new_n3215_), .Y(_abc_40319_new_n5267_));
AND2X2 AND2X2_2342 ( .A(_abc_40319_new_n5268_), .B(_abc_40319_new_n4497_), .Y(_abc_40319_new_n5269_));
AND2X2 AND2X2_2343 ( .A(_abc_40319_new_n5271_), .B(_abc_40319_new_n4271_), .Y(_abc_40319_new_n5272_));
AND2X2 AND2X2_2344 ( .A(_abc_40319_new_n5268_), .B(_abc_40319_new_n4512_), .Y(_abc_40319_new_n5273_));
AND2X2 AND2X2_2345 ( .A(_abc_40319_new_n5274_), .B(_abc_40319_new_n5275_), .Y(_abc_40319_new_n5276_));
AND2X2 AND2X2_2346 ( .A(_abc_40319_new_n5276_), .B(_abc_40319_new_n4272_), .Y(_abc_40319_new_n5277_));
AND2X2 AND2X2_2347 ( .A(_abc_40319_new_n1046_), .B(_abc_40319_new_n4310_), .Y(_abc_40319_new_n5279_));
AND2X2 AND2X2_2348 ( .A(_abc_40319_new_n998_), .B(_abc_40319_new_n1152_), .Y(_abc_40319_new_n5280_));
AND2X2 AND2X2_2349 ( .A(_abc_40319_new_n5282_), .B(_abc_40319_new_n5278_), .Y(_abc_40319_new_n5283_));
AND2X2 AND2X2_235 ( .A(_abc_40319_new_n537_), .B(_abc_40319_new_n550_), .Y(_abc_40319_new_n1023_));
AND2X2 AND2X2_2350 ( .A(_abc_40319_new_n1169_), .B(_abc_40319_new_n1003_), .Y(_abc_40319_new_n5284_));
AND2X2 AND2X2_2351 ( .A(_abc_40319_new_n5253_), .B(_abc_40319_new_n3222_), .Y(_abc_40319_new_n5290_));
AND2X2 AND2X2_2352 ( .A(_abc_40319_new_n3495_), .B(_abc_40319_new_n3223_), .Y(_abc_40319_new_n5291_));
AND2X2 AND2X2_2353 ( .A(_abc_40319_new_n5292_), .B(_abc_40319_new_n4507_), .Y(_abc_40319_new_n5293_));
AND2X2 AND2X2_2354 ( .A(_abc_40319_new_n829_), .B(_abc_40319_new_n4499_), .Y(_abc_40319_new_n5294_));
AND2X2 AND2X2_2355 ( .A(_abc_40319_new_n4424_), .B(_abc_40319_new_n5295_), .Y(_abc_40319_new_n5296_));
AND2X2 AND2X2_2356 ( .A(_abc_40319_new_n5297_), .B(_abc_40319_new_n4435_), .Y(_abc_40319_new_n5298_));
AND2X2 AND2X2_2357 ( .A(_abc_40319_new_n5301_), .B(_abc_40319_new_n5302_), .Y(_abc_40319_new_n5303_));
AND2X2 AND2X2_2358 ( .A(_abc_40319_new_n5303_), .B(_abc_40319_new_n4497_), .Y(_abc_40319_new_n5304_));
AND2X2 AND2X2_2359 ( .A(_abc_40319_new_n5306_), .B(_abc_40319_new_n4271_), .Y(_abc_40319_new_n5307_));
AND2X2 AND2X2_236 ( .A(_abc_40319_new_n1025_), .B(_abc_40319_new_n1024_), .Y(_abc_40319_new_n1026_));
AND2X2 AND2X2_2360 ( .A(_abc_40319_new_n5303_), .B(_abc_40319_new_n4512_), .Y(_abc_40319_new_n5308_));
AND2X2 AND2X2_2361 ( .A(_abc_40319_new_n784_), .B(_abc_40319_new_n1152_), .Y(_abc_40319_new_n5310_));
AND2X2 AND2X2_2362 ( .A(_abc_40319_new_n746_), .B(_abc_40319_new_n4310_), .Y(_abc_40319_new_n5311_));
AND2X2 AND2X2_2363 ( .A(_abc_40319_new_n5313_), .B(_abc_40319_new_n5309_), .Y(_abc_40319_new_n5314_));
AND2X2 AND2X2_2364 ( .A(_abc_40319_new_n5315_), .B(_abc_40319_new_n5316_), .Y(_abc_40319_new_n5317_));
AND2X2 AND2X2_2365 ( .A(_abc_40319_new_n5317_), .B(_abc_40319_new_n4272_), .Y(_abc_40319_new_n5318_));
AND2X2 AND2X2_2366 ( .A(_abc_40319_new_n1169_), .B(_abc_40319_new_n792_), .Y(_abc_40319_new_n5319_));
AND2X2 AND2X2_2367 ( .A(_abc_40319_new_n5326_), .B(_abc_40319_new_n4507_), .Y(_abc_40319_new_n5327_));
AND2X2 AND2X2_2368 ( .A(_abc_40319_new_n5327_), .B(_abc_40319_new_n5325_), .Y(_abc_40319_new_n5328_));
AND2X2 AND2X2_2369 ( .A(_abc_40319_new_n795_), .B(_abc_40319_new_n4499_), .Y(_abc_40319_new_n5329_));
AND2X2 AND2X2_237 ( .A(_abc_40319_new_n1026_), .B(IR_REG_31_), .Y(_abc_40319_new_n1027_));
AND2X2 AND2X2_2370 ( .A(_abc_40319_new_n5299_), .B(_abc_40319_new_n4427_), .Y(_abc_40319_new_n5330_));
AND2X2 AND2X2_2371 ( .A(_abc_40319_new_n5332_), .B(_abc_40319_new_n3123_), .Y(_abc_40319_new_n5333_));
AND2X2 AND2X2_2372 ( .A(_abc_40319_new_n5331_), .B(_abc_40319_new_n3124_), .Y(_abc_40319_new_n5334_));
AND2X2 AND2X2_2373 ( .A(_abc_40319_new_n5335_), .B(_abc_40319_new_n4497_), .Y(_abc_40319_new_n5336_));
AND2X2 AND2X2_2374 ( .A(_abc_40319_new_n689_), .B(_abc_40319_new_n1152_), .Y(_abc_40319_new_n5339_));
AND2X2 AND2X2_2375 ( .A(_abc_40319_new_n1010_), .B(_abc_40319_new_n4310_), .Y(_abc_40319_new_n5340_));
AND2X2 AND2X2_2376 ( .A(_abc_40319_new_n5342_), .B(_abc_40319_new_n4271_), .Y(_abc_40319_new_n5343_));
AND2X2 AND2X2_2377 ( .A(_abc_40319_new_n5335_), .B(_abc_40319_new_n4512_), .Y(_abc_40319_new_n5344_));
AND2X2 AND2X2_2378 ( .A(_abc_40319_new_n5345_), .B(_abc_40319_new_n5346_), .Y(_abc_40319_new_n5347_));
AND2X2 AND2X2_2379 ( .A(_abc_40319_new_n5347_), .B(_abc_40319_new_n4272_), .Y(_abc_40319_new_n5348_));
AND2X2 AND2X2_238 ( .A(_abc_40319_new_n524_), .B(IR_REG_7_), .Y(_abc_40319_new_n1028_));
AND2X2 AND2X2_2380 ( .A(_abc_40319_new_n4309_), .B(REG2_REG_5_), .Y(_abc_40319_new_n5349_));
AND2X2 AND2X2_2381 ( .A(_abc_40319_new_n1169_), .B(_abc_40319_new_n743_), .Y(_abc_40319_new_n5350_));
AND2X2 AND2X2_2382 ( .A(_abc_40319_new_n5358_), .B(_abc_40319_new_n4507_), .Y(_abc_40319_new_n5359_));
AND2X2 AND2X2_2383 ( .A(_abc_40319_new_n5359_), .B(_abc_40319_new_n5356_), .Y(_abc_40319_new_n5360_));
AND2X2 AND2X2_2384 ( .A(_abc_40319_new_n865_), .B(_abc_40319_new_n4499_), .Y(_abc_40319_new_n5361_));
AND2X2 AND2X2_2385 ( .A(_abc_40319_new_n5297_), .B(_abc_40319_new_n4434_), .Y(_abc_40319_new_n5362_));
AND2X2 AND2X2_2386 ( .A(_abc_40319_new_n5364_), .B(_abc_40319_new_n5365_), .Y(_abc_40319_new_n5366_));
AND2X2 AND2X2_2387 ( .A(_abc_40319_new_n5366_), .B(_abc_40319_new_n4497_), .Y(_abc_40319_new_n5367_));
AND2X2 AND2X2_2388 ( .A(_abc_40319_new_n820_), .B(_abc_40319_new_n1152_), .Y(_abc_40319_new_n5370_));
AND2X2 AND2X2_2389 ( .A(_abc_40319_new_n795_), .B(_abc_40319_new_n4310_), .Y(_abc_40319_new_n5371_));
AND2X2 AND2X2_239 ( .A(_abc_40319_new_n640_), .B(_abc_40319_new_n1030_), .Y(_abc_40319_new_n1031_));
AND2X2 AND2X2_2390 ( .A(_abc_40319_new_n5373_), .B(_abc_40319_new_n4271_), .Y(_abc_40319_new_n5374_));
AND2X2 AND2X2_2391 ( .A(_abc_40319_new_n5366_), .B(_abc_40319_new_n4512_), .Y(_abc_40319_new_n5375_));
AND2X2 AND2X2_2392 ( .A(_abc_40319_new_n5376_), .B(_abc_40319_new_n5377_), .Y(_abc_40319_new_n5378_));
AND2X2 AND2X2_2393 ( .A(_abc_40319_new_n5378_), .B(_abc_40319_new_n4272_), .Y(_abc_40319_new_n5379_));
AND2X2 AND2X2_2394 ( .A(_abc_40319_new_n4309_), .B(REG2_REG_3_), .Y(_abc_40319_new_n5380_));
AND2X2 AND2X2_2395 ( .A(_abc_40319_new_n1169_), .B(_abc_40319_new_n826_), .Y(_abc_40319_new_n5381_));
AND2X2 AND2X2_2396 ( .A(_abc_40319_new_n4425_), .B(_abc_40319_new_n3128_), .Y(_abc_40319_new_n5388_));
AND2X2 AND2X2_2397 ( .A(_abc_40319_new_n4424_), .B(_abc_40319_new_n3127_), .Y(_abc_40319_new_n5389_));
AND2X2 AND2X2_2398 ( .A(_abc_40319_new_n5390_), .B(_abc_40319_new_n4497_), .Y(_abc_40319_new_n5391_));
AND2X2 AND2X2_2399 ( .A(_abc_40319_new_n5393_), .B(_abc_40319_new_n5394_), .Y(_abc_40319_new_n5395_));
AND2X2 AND2X2_24 ( .A(_abc_40319_new_n572_), .B(_abc_40319_new_n575_), .Y(_abc_40319_new_n576_));
AND2X2 AND2X2_240 ( .A(_abc_40319_new_n1032_), .B(_abc_40319_new_n1033_), .Y(_abc_40319_new_n1034_));
AND2X2 AND2X2_2400 ( .A(_abc_40319_new_n5395_), .B(_abc_40319_new_n4507_), .Y(_abc_40319_new_n5396_));
AND2X2 AND2X2_2401 ( .A(_abc_40319_new_n829_), .B(_abc_40319_new_n4310_), .Y(_abc_40319_new_n5397_));
AND2X2 AND2X2_2402 ( .A(_abc_40319_new_n904_), .B(_abc_40319_new_n4499_), .Y(_abc_40319_new_n5398_));
AND2X2 AND2X2_2403 ( .A(_abc_40319_new_n848_), .B(_abc_40319_new_n1152_), .Y(_abc_40319_new_n5399_));
AND2X2 AND2X2_2404 ( .A(_abc_40319_new_n752_), .B(_abc_40319_new_n671_), .Y(_abc_40319_new_n5405_));
AND2X2 AND2X2_2405 ( .A(_abc_40319_new_n5406_), .B(_abc_40319_new_n5405_), .Y(_abc_40319_new_n5407_));
AND2X2 AND2X2_2406 ( .A(_abc_40319_new_n5407_), .B(_abc_40319_new_n5404_), .Y(_abc_40319_new_n5408_));
AND2X2 AND2X2_2407 ( .A(_abc_40319_new_n5408_), .B(_abc_40319_new_n698_), .Y(_abc_40319_new_n5409_));
AND2X2 AND2X2_2408 ( .A(_abc_40319_new_n5411_), .B(_abc_40319_new_n5387_), .Y(_abc_40319_new_n5412_));
AND2X2 AND2X2_2409 ( .A(_abc_40319_new_n5390_), .B(_abc_40319_new_n4512_), .Y(_abc_40319_new_n5413_));
AND2X2 AND2X2_241 ( .A(_abc_40319_new_n1034_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1035_));
AND2X2 AND2X2_2410 ( .A(_abc_40319_new_n1169_), .B(REG3_REG_2_), .Y(_abc_40319_new_n5414_));
AND2X2 AND2X2_2411 ( .A(_abc_40319_new_n5420_), .B(_abc_40319_new_n4507_), .Y(_abc_40319_new_n5421_));
AND2X2 AND2X2_2412 ( .A(_abc_40319_new_n5419_), .B(_abc_40319_new_n5421_), .Y(_abc_40319_new_n5422_));
AND2X2 AND2X2_2413 ( .A(_abc_40319_new_n924_), .B(_abc_40319_new_n4499_), .Y(_abc_40319_new_n5423_));
AND2X2 AND2X2_2414 ( .A(_abc_40319_new_n3118_), .B(_abc_40319_new_n4422_), .Y(_abc_40319_new_n5424_));
AND2X2 AND2X2_2415 ( .A(_abc_40319_new_n3119_), .B(_abc_40319_new_n4421_), .Y(_abc_40319_new_n5425_));
AND2X2 AND2X2_2416 ( .A(_abc_40319_new_n5426_), .B(_abc_40319_new_n4497_), .Y(_abc_40319_new_n5427_));
AND2X2 AND2X2_2417 ( .A(_abc_40319_new_n5431_), .B(_abc_40319_new_n5405_), .Y(_abc_40319_new_n5432_));
AND2X2 AND2X2_2418 ( .A(_abc_40319_new_n5432_), .B(_abc_40319_new_n5430_), .Y(_abc_40319_new_n5433_));
AND2X2 AND2X2_2419 ( .A(_abc_40319_new_n5433_), .B(_abc_40319_new_n698_), .Y(_abc_40319_new_n5434_));
AND2X2 AND2X2_242 ( .A(_abc_40319_new_n736_), .B(REG0_REG_7_), .Y(_abc_40319_new_n1036_));
AND2X2 AND2X2_2420 ( .A(_abc_40319_new_n865_), .B(_abc_40319_new_n4310_), .Y(_abc_40319_new_n5435_));
AND2X2 AND2X2_2421 ( .A(_abc_40319_new_n891_), .B(_abc_40319_new_n1152_), .Y(_abc_40319_new_n5436_));
AND2X2 AND2X2_2422 ( .A(_abc_40319_new_n5439_), .B(_abc_40319_new_n4271_), .Y(_abc_40319_new_n5440_));
AND2X2 AND2X2_2423 ( .A(_abc_40319_new_n5426_), .B(_abc_40319_new_n4512_), .Y(_abc_40319_new_n5441_));
AND2X2 AND2X2_2424 ( .A(_abc_40319_new_n4309_), .B(REG2_REG_1_), .Y(_abc_40319_new_n5442_));
AND2X2 AND2X2_2425 ( .A(_abc_40319_new_n1169_), .B(REG3_REG_1_), .Y(_abc_40319_new_n5443_));
AND2X2 AND2X2_2426 ( .A(_abc_40319_new_n3137_), .B(_abc_40319_new_n5448_), .Y(_abc_40319_new_n5449_));
AND2X2 AND2X2_2427 ( .A(_abc_40319_new_n904_), .B(_abc_40319_new_n4310_), .Y(_abc_40319_new_n5450_));
AND2X2 AND2X2_2428 ( .A(_abc_40319_new_n930_), .B(_abc_40319_new_n5452_), .Y(_abc_40319_new_n5453_));
AND2X2 AND2X2_2429 ( .A(_abc_40319_new_n5455_), .B(_abc_40319_new_n5456_), .Y(_abc_40319_new_n5457_));
AND2X2 AND2X2_243 ( .A(_abc_40319_new_n733_), .B(REG2_REG_7_), .Y(_abc_40319_new_n1037_));
AND2X2 AND2X2_2430 ( .A(_abc_40319_new_n4512_), .B(_abc_40319_new_n3137_), .Y(_abc_40319_new_n5458_));
AND2X2 AND2X2_2431 ( .A(_abc_40319_new_n1169_), .B(REG3_REG_0_), .Y(_abc_40319_new_n5459_));
AND2X2 AND2X2_2432 ( .A(IR_REG_31_), .B(STATE_REG), .Y(_abc_40319_new_n5463_));
AND2X2 AND2X2_2433 ( .A(_abc_40319_new_n711_), .B(_abc_40319_new_n5463_), .Y(_abc_40319_new_n5464_));
AND2X2 AND2X2_2434 ( .A(n1336), .B(DATAI_31_), .Y(_abc_40319_new_n5465_));
AND2X2 AND2X2_2435 ( .A(_abc_40319_new_n1120_), .B(_abc_40319_new_n1072_), .Y(_abc_40319_new_n5468_));
AND2X2 AND2X2_2436 ( .A(_abc_40319_new_n5469_), .B(nRESET_G), .Y(_abc_40319_new_n5470_));
AND2X2 AND2X2_2437 ( .A(_abc_40319_new_n5470_), .B(D_REG_31_), .Y(n493));
AND2X2 AND2X2_2438 ( .A(_abc_40319_new_n5470_), .B(D_REG_30_), .Y(n488));
AND2X2 AND2X2_2439 ( .A(_abc_40319_new_n5470_), .B(D_REG_29_), .Y(n483));
AND2X2 AND2X2_244 ( .A(_abc_40319_new_n1000_), .B(REG3_REG_7_), .Y(_abc_40319_new_n1039_));
AND2X2 AND2X2_2440 ( .A(_abc_40319_new_n5470_), .B(D_REG_28_), .Y(n478));
AND2X2 AND2X2_2441 ( .A(_abc_40319_new_n5470_), .B(D_REG_27_), .Y(n473));
AND2X2 AND2X2_2442 ( .A(_abc_40319_new_n5470_), .B(D_REG_26_), .Y(n468));
AND2X2 AND2X2_2443 ( .A(_abc_40319_new_n5470_), .B(D_REG_25_), .Y(n463));
AND2X2 AND2X2_2444 ( .A(_abc_40319_new_n5470_), .B(D_REG_24_), .Y(n458));
AND2X2 AND2X2_2445 ( .A(_abc_40319_new_n5470_), .B(D_REG_23_), .Y(n453));
AND2X2 AND2X2_2446 ( .A(_abc_40319_new_n5470_), .B(D_REG_22_), .Y(n448));
AND2X2 AND2X2_2447 ( .A(_abc_40319_new_n5470_), .B(D_REG_21_), .Y(n443));
AND2X2 AND2X2_2448 ( .A(_abc_40319_new_n5470_), .B(D_REG_20_), .Y(n438));
AND2X2 AND2X2_2449 ( .A(_abc_40319_new_n5470_), .B(D_REG_19_), .Y(n433));
AND2X2 AND2X2_245 ( .A(_abc_40319_new_n1040_), .B(_abc_40319_new_n1041_), .Y(_abc_40319_new_n1042_));
AND2X2 AND2X2_2450 ( .A(_abc_40319_new_n5470_), .B(D_REG_18_), .Y(n428));
AND2X2 AND2X2_2451 ( .A(_abc_40319_new_n5470_), .B(D_REG_17_), .Y(n423));
AND2X2 AND2X2_2452 ( .A(_abc_40319_new_n5470_), .B(D_REG_16_), .Y(n418));
AND2X2 AND2X2_2453 ( .A(_abc_40319_new_n5470_), .B(D_REG_15_), .Y(n413));
AND2X2 AND2X2_2454 ( .A(_abc_40319_new_n5470_), .B(D_REG_14_), .Y(n408));
AND2X2 AND2X2_2455 ( .A(_abc_40319_new_n5470_), .B(D_REG_13_), .Y(n403));
AND2X2 AND2X2_2456 ( .A(_abc_40319_new_n5470_), .B(D_REG_12_), .Y(n398));
AND2X2 AND2X2_2457 ( .A(_abc_40319_new_n5470_), .B(D_REG_11_), .Y(n393));
AND2X2 AND2X2_2458 ( .A(_abc_40319_new_n5470_), .B(D_REG_10_), .Y(n388));
AND2X2 AND2X2_2459 ( .A(_abc_40319_new_n5470_), .B(D_REG_9_), .Y(n383));
AND2X2 AND2X2_246 ( .A(_abc_40319_new_n738_), .B(_abc_40319_new_n1042_), .Y(_abc_40319_new_n1043_));
AND2X2 AND2X2_2460 ( .A(_abc_40319_new_n5470_), .B(D_REG_8_), .Y(n378));
AND2X2 AND2X2_2461 ( .A(_abc_40319_new_n5470_), .B(D_REG_7_), .Y(n373));
AND2X2 AND2X2_2462 ( .A(_abc_40319_new_n5470_), .B(D_REG_6_), .Y(n368));
AND2X2 AND2X2_2463 ( .A(_abc_40319_new_n5470_), .B(D_REG_5_), .Y(n363));
AND2X2 AND2X2_2464 ( .A(_abc_40319_new_n5470_), .B(D_REG_4_), .Y(n358));
AND2X2 AND2X2_2465 ( .A(_abc_40319_new_n5470_), .B(D_REG_3_), .Y(n353));
AND2X2 AND2X2_2466 ( .A(_abc_40319_new_n5470_), .B(D_REG_2_), .Y(n348));
AND2X2 AND2X2_2467 ( .A(_abc_40319_new_n727_), .B(_abc_40319_new_n5463_), .Y(_abc_40319_new_n5501_));
AND2X2 AND2X2_2468 ( .A(_abc_40319_new_n524_), .B(STATE_REG), .Y(_abc_40319_new_n5502_));
AND2X2 AND2X2_2469 ( .A(_abc_40319_new_n5502_), .B(IR_REG_30_), .Y(_abc_40319_new_n5503_));
AND2X2 AND2X2_247 ( .A(_abc_40319_new_n722_), .B(REG1_REG_7_), .Y(_abc_40319_new_n1044_));
AND2X2 AND2X2_2470 ( .A(n1336), .B(DATAI_30_), .Y(_abc_40319_new_n5504_));
AND2X2 AND2X2_2471 ( .A(_abc_40319_new_n718_), .B(_abc_40319_new_n5463_), .Y(_abc_40319_new_n5508_));
AND2X2 AND2X2_2472 ( .A(_abc_40319_new_n5502_), .B(IR_REG_29_), .Y(_abc_40319_new_n5509_));
AND2X2 AND2X2_2473 ( .A(n1336), .B(DATAI_29_), .Y(_abc_40319_new_n5510_));
AND2X2 AND2X2_2474 ( .A(_abc_40319_new_n636_), .B(_abc_40319_new_n5463_), .Y(_abc_40319_new_n5514_));
AND2X2 AND2X2_2475 ( .A(_abc_40319_new_n5502_), .B(IR_REG_28_), .Y(_abc_40319_new_n5515_));
AND2X2 AND2X2_2476 ( .A(n1336), .B(DATAI_28_), .Y(_abc_40319_new_n5516_));
AND2X2 AND2X2_2477 ( .A(_abc_40319_new_n625_), .B(_abc_40319_new_n5463_), .Y(_abc_40319_new_n5520_));
AND2X2 AND2X2_2478 ( .A(n1336), .B(DATAI_27_), .Y(_abc_40319_new_n5521_));
AND2X2 AND2X2_2479 ( .A(_abc_40319_new_n5502_), .B(IR_REG_27_), .Y(_abc_40319_new_n5522_));
AND2X2 AND2X2_248 ( .A(_abc_40319_new_n705_), .B(_abc_40319_new_n1046_), .Y(_abc_40319_new_n1047_));
AND2X2 AND2X2_2480 ( .A(_abc_40319_new_n580_), .B(_abc_40319_new_n5463_), .Y(_abc_40319_new_n5526_));
AND2X2 AND2X2_2481 ( .A(n1336), .B(DATAI_26_), .Y(_abc_40319_new_n5527_));
AND2X2 AND2X2_2482 ( .A(_abc_40319_new_n5502_), .B(IR_REG_26_), .Y(_abc_40319_new_n5528_));
AND2X2 AND2X2_2483 ( .A(_abc_40319_new_n586_), .B(_abc_40319_new_n5463_), .Y(_abc_40319_new_n5532_));
AND2X2 AND2X2_2484 ( .A(n1336), .B(DATAI_25_), .Y(_abc_40319_new_n5533_));
AND2X2 AND2X2_2485 ( .A(_abc_40319_new_n5502_), .B(IR_REG_25_), .Y(_abc_40319_new_n5534_));
AND2X2 AND2X2_2486 ( .A(_abc_40319_new_n594_), .B(_abc_40319_new_n5463_), .Y(_abc_40319_new_n5538_));
AND2X2 AND2X2_2487 ( .A(n1336), .B(DATAI_24_), .Y(_abc_40319_new_n5539_));
AND2X2 AND2X2_2488 ( .A(_abc_40319_new_n5502_), .B(IR_REG_24_), .Y(_abc_40319_new_n5540_));
AND2X2 AND2X2_2489 ( .A(n1336), .B(DATAI_23_), .Y(_abc_40319_new_n5544_));
AND2X2 AND2X2_249 ( .A(_abc_40319_new_n1034_), .B(_abc_40319_new_n763_), .Y(_abc_40319_new_n1050_));
AND2X2 AND2X2_2490 ( .A(_abc_40319_new_n5547_), .B(_abc_40319_new_n5463_), .Y(_abc_40319_new_n5548_));
AND2X2 AND2X2_2491 ( .A(n1336), .B(DATAI_22_), .Y(_abc_40319_new_n5549_));
AND2X2 AND2X2_2492 ( .A(_abc_40319_new_n5502_), .B(IR_REG_22_), .Y(_abc_40319_new_n5550_));
AND2X2 AND2X2_2493 ( .A(_abc_40319_new_n652_), .B(_abc_40319_new_n5463_), .Y(_abc_40319_new_n5554_));
AND2X2 AND2X2_2494 ( .A(n1336), .B(DATAI_21_), .Y(_abc_40319_new_n5555_));
AND2X2 AND2X2_2495 ( .A(_abc_40319_new_n5502_), .B(IR_REG_21_), .Y(_abc_40319_new_n5556_));
AND2X2 AND2X2_2496 ( .A(_abc_40319_new_n668_), .B(_abc_40319_new_n5463_), .Y(_abc_40319_new_n5560_));
AND2X2 AND2X2_2497 ( .A(n1336), .B(DATAI_20_), .Y(_abc_40319_new_n5561_));
AND2X2 AND2X2_2498 ( .A(_abc_40319_new_n5502_), .B(IR_REG_20_), .Y(_abc_40319_new_n5562_));
AND2X2 AND2X2_2499 ( .A(_abc_40319_new_n695_), .B(_abc_40319_new_n5463_), .Y(_abc_40319_new_n5566_));
AND2X2 AND2X2_25 ( .A(_abc_40319_new_n576_), .B(_abc_40319_new_n525_), .Y(_abc_40319_new_n578_));
AND2X2 AND2X2_250 ( .A(_abc_40319_new_n1046_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1051_));
AND2X2 AND2X2_2500 ( .A(n1336), .B(DATAI_19_), .Y(_abc_40319_new_n5567_));
AND2X2 AND2X2_2501 ( .A(_abc_40319_new_n5502_), .B(IR_REG_19_), .Y(_abc_40319_new_n5568_));
AND2X2 AND2X2_2502 ( .A(_abc_40319_new_n1355_), .B(_abc_40319_new_n5463_), .Y(_abc_40319_new_n5572_));
AND2X2 AND2X2_2503 ( .A(n1336), .B(DATAI_18_), .Y(_abc_40319_new_n5573_));
AND2X2 AND2X2_2504 ( .A(_abc_40319_new_n5502_), .B(IR_REG_18_), .Y(_abc_40319_new_n5574_));
AND2X2 AND2X2_2505 ( .A(_abc_40319_new_n1425_), .B(_abc_40319_new_n5463_), .Y(_abc_40319_new_n5578_));
AND2X2 AND2X2_2506 ( .A(n1336), .B(DATAI_17_), .Y(_abc_40319_new_n5579_));
AND2X2 AND2X2_2507 ( .A(_abc_40319_new_n5502_), .B(IR_REG_17_), .Y(_abc_40319_new_n5580_));
AND2X2 AND2X2_2508 ( .A(_abc_40319_new_n5584_), .B(_abc_40319_new_n5463_), .Y(_abc_40319_new_n5585_));
AND2X2 AND2X2_2509 ( .A(n1336), .B(DATAI_16_), .Y(_abc_40319_new_n5586_));
AND2X2 AND2X2_251 ( .A(_abc_40319_new_n1055_), .B(_abc_40319_new_n1053_), .Y(_abc_40319_new_n1056_));
AND2X2 AND2X2_2510 ( .A(_abc_40319_new_n5502_), .B(IR_REG_16_), .Y(_abc_40319_new_n5587_));
AND2X2 AND2X2_2511 ( .A(_abc_40319_new_n1463_), .B(_abc_40319_new_n5463_), .Y(_abc_40319_new_n5591_));
AND2X2 AND2X2_2512 ( .A(n1336), .B(DATAI_15_), .Y(_abc_40319_new_n5592_));
AND2X2 AND2X2_2513 ( .A(_abc_40319_new_n5502_), .B(IR_REG_15_), .Y(_abc_40319_new_n5593_));
AND2X2 AND2X2_2514 ( .A(_abc_40319_new_n1498_), .B(_abc_40319_new_n5463_), .Y(_abc_40319_new_n5597_));
AND2X2 AND2X2_2515 ( .A(n1336), .B(DATAI_14_), .Y(_abc_40319_new_n5598_));
AND2X2 AND2X2_2516 ( .A(_abc_40319_new_n5502_), .B(IR_REG_14_), .Y(_abc_40319_new_n5599_));
AND2X2 AND2X2_2517 ( .A(_abc_40319_new_n5603_), .B(_abc_40319_new_n5463_), .Y(_abc_40319_new_n5604_));
AND2X2 AND2X2_2518 ( .A(_abc_40319_new_n5502_), .B(IR_REG_13_), .Y(_abc_40319_new_n5605_));
AND2X2 AND2X2_2519 ( .A(n1336), .B(DATAI_13_), .Y(_abc_40319_new_n5606_));
AND2X2 AND2X2_252 ( .A(_abc_40319_new_n1020_), .B(_abc_40319_new_n1013_), .Y(_abc_40319_new_n1059_));
AND2X2 AND2X2_2520 ( .A(_abc_40319_new_n5610_), .B(_abc_40319_new_n5463_), .Y(_abc_40319_new_n5611_));
AND2X2 AND2X2_2521 ( .A(_abc_40319_new_n5502_), .B(IR_REG_12_), .Y(_abc_40319_new_n5612_));
AND2X2 AND2X2_2522 ( .A(n1336), .B(DATAI_12_), .Y(_abc_40319_new_n5613_));
AND2X2 AND2X2_2523 ( .A(_abc_40319_new_n5617_), .B(_abc_40319_new_n5463_), .Y(_abc_40319_new_n5618_));
AND2X2 AND2X2_2524 ( .A(_abc_40319_new_n5502_), .B(IR_REG_11_), .Y(_abc_40319_new_n5619_));
AND2X2 AND2X2_2525 ( .A(n1336), .B(DATAI_11_), .Y(_abc_40319_new_n5620_));
AND2X2 AND2X2_2526 ( .A(_abc_40319_new_n5624_), .B(_abc_40319_new_n5463_), .Y(_abc_40319_new_n5625_));
AND2X2 AND2X2_2527 ( .A(n1336), .B(DATAI_10_), .Y(_abc_40319_new_n5626_));
AND2X2 AND2X2_2528 ( .A(_abc_40319_new_n5502_), .B(IR_REG_10_), .Y(_abc_40319_new_n5627_));
AND2X2 AND2X2_2529 ( .A(_abc_40319_new_n1607_), .B(_abc_40319_new_n5463_), .Y(_abc_40319_new_n5631_));
AND2X2 AND2X2_253 ( .A(_abc_40319_new_n1056_), .B(_abc_40319_new_n1049_), .Y(_abc_40319_new_n1060_));
AND2X2 AND2X2_2530 ( .A(n1336), .B(DATAI_9_), .Y(_abc_40319_new_n5632_));
AND2X2 AND2X2_2531 ( .A(_abc_40319_new_n5502_), .B(IR_REG_9_), .Y(_abc_40319_new_n5633_));
AND2X2 AND2X2_2532 ( .A(_abc_40319_new_n1564_), .B(_abc_40319_new_n5463_), .Y(_abc_40319_new_n5637_));
AND2X2 AND2X2_2533 ( .A(n1336), .B(DATAI_8_), .Y(_abc_40319_new_n5638_));
AND2X2 AND2X2_2534 ( .A(_abc_40319_new_n5502_), .B(IR_REG_8_), .Y(_abc_40319_new_n5639_));
AND2X2 AND2X2_2535 ( .A(_abc_40319_new_n1026_), .B(_abc_40319_new_n5463_), .Y(_abc_40319_new_n5643_));
AND2X2 AND2X2_2536 ( .A(n1336), .B(DATAI_7_), .Y(_abc_40319_new_n5644_));
AND2X2 AND2X2_2537 ( .A(_abc_40319_new_n5502_), .B(IR_REG_7_), .Y(_abc_40319_new_n5645_));
AND2X2 AND2X2_2538 ( .A(_abc_40319_new_n990_), .B(_abc_40319_new_n5463_), .Y(_abc_40319_new_n5649_));
AND2X2 AND2X2_2539 ( .A(n1336), .B(DATAI_6_), .Y(_abc_40319_new_n5650_));
AND2X2 AND2X2_254 ( .A(_abc_40319_new_n1065_), .B(B_REG), .Y(_abc_40319_new_n1066_));
AND2X2 AND2X2_2540 ( .A(_abc_40319_new_n5502_), .B(IR_REG_6_), .Y(_abc_40319_new_n5651_));
AND2X2 AND2X2_2541 ( .A(_abc_40319_new_n681_), .B(_abc_40319_new_n5463_), .Y(_abc_40319_new_n5655_));
AND2X2 AND2X2_2542 ( .A(n1336), .B(DATAI_5_), .Y(_abc_40319_new_n5656_));
AND2X2 AND2X2_2543 ( .A(_abc_40319_new_n5502_), .B(IR_REG_5_), .Y(_abc_40319_new_n5657_));
AND2X2 AND2X2_2544 ( .A(_abc_40319_new_n776_), .B(_abc_40319_new_n5463_), .Y(_abc_40319_new_n5661_));
AND2X2 AND2X2_2545 ( .A(n1336), .B(DATAI_4_), .Y(_abc_40319_new_n5662_));
AND2X2 AND2X2_2546 ( .A(_abc_40319_new_n5502_), .B(IR_REG_4_), .Y(_abc_40319_new_n5663_));
AND2X2 AND2X2_2547 ( .A(_abc_40319_new_n810_), .B(_abc_40319_new_n5463_), .Y(_abc_40319_new_n5667_));
AND2X2 AND2X2_2548 ( .A(n1336), .B(DATAI_3_), .Y(_abc_40319_new_n5668_));
AND2X2 AND2X2_2549 ( .A(_abc_40319_new_n5502_), .B(IR_REG_3_), .Y(_abc_40319_new_n5669_));
AND2X2 AND2X2_255 ( .A(_abc_40319_new_n1066_), .B(_abc_40319_new_n1064_), .Y(_abc_40319_new_n1067_));
AND2X2 AND2X2_2550 ( .A(_abc_40319_new_n674_), .B(_abc_40319_new_n5463_), .Y(_abc_40319_new_n5674_));
AND2X2 AND2X2_2551 ( .A(_abc_40319_new_n5674_), .B(_abc_40319_new_n5673_), .Y(_abc_40319_new_n5675_));
AND2X2 AND2X2_2552 ( .A(_abc_40319_new_n5502_), .B(IR_REG_2_), .Y(_abc_40319_new_n5676_));
AND2X2 AND2X2_2553 ( .A(n1336), .B(DATAI_2_), .Y(_abc_40319_new_n5677_));
AND2X2 AND2X2_2554 ( .A(_abc_40319_new_n886_), .B(STATE_REG), .Y(_abc_40319_new_n5681_));
AND2X2 AND2X2_2555 ( .A(n1336), .B(DATAI_1_), .Y(_abc_40319_new_n5682_));
AND2X2 AND2X2_2556 ( .A(n1336), .B(DATAI_0_), .Y(_abc_40319_new_n5685_));
AND2X2 AND2X2_2557 ( .A(IR_REG_0_), .B(STATE_REG), .Y(_abc_40319_new_n5686_));
AND2X2 AND2X2_2558 ( .A(_abc_40319_new_n3452_), .B(_abc_40319_new_n670_), .Y(_abc_40319_new_n5689_));
AND2X2 AND2X2_2559 ( .A(_abc_40319_new_n5693_), .B(_abc_40319_new_n5690_), .Y(_abc_40319_new_n5694_));
AND2X2 AND2X2_256 ( .A(_abc_40319_new_n596_), .B(_abc_40319_new_n1069_), .Y(_abc_40319_new_n1070_));
AND2X2 AND2X2_2560 ( .A(_abc_40319_new_n5694_), .B(_abc_40319_new_n5689_), .Y(_abc_40319_new_n5695_));
AND2X2 AND2X2_2561 ( .A(_abc_40319_new_n3040_), .B(_abc_40319_new_n3042_), .Y(_abc_40319_new_n5696_));
AND2X2 AND2X2_2562 ( .A(_abc_40319_new_n1980_), .B(_abc_40319_new_n2089_), .Y(_abc_40319_new_n5697_));
AND2X2 AND2X2_2563 ( .A(_abc_40319_new_n4489_), .B(_abc_40319_new_n5698_), .Y(_abc_40319_new_n5699_));
AND2X2 AND2X2_2564 ( .A(_abc_40319_new_n5703_), .B(_abc_40319_new_n5701_), .Y(_abc_40319_new_n5704_));
AND2X2 AND2X2_2565 ( .A(_abc_40319_new_n5704_), .B(_abc_40319_new_n4497_), .Y(_abc_40319_new_n5705_));
AND2X2 AND2X2_2566 ( .A(_abc_40319_new_n5694_), .B(_abc_40319_new_n5706_), .Y(_abc_40319_new_n5707_));
AND2X2 AND2X2_2567 ( .A(_abc_40319_new_n3075_), .B(_abc_40319_new_n4312_), .Y(_abc_40319_new_n5708_));
AND2X2 AND2X2_2568 ( .A(_abc_40319_new_n1980_), .B(_abc_40319_new_n4499_), .Y(_abc_40319_new_n5709_));
AND2X2 AND2X2_2569 ( .A(_abc_40319_new_n5713_), .B(_abc_40319_new_n4271_), .Y(_abc_40319_new_n5714_));
AND2X2 AND2X2_257 ( .A(_abc_40319_new_n1068_), .B(_abc_40319_new_n1064_), .Y(_abc_40319_new_n1074_));
AND2X2 AND2X2_2570 ( .A(_abc_40319_new_n5704_), .B(_abc_40319_new_n4512_), .Y(_abc_40319_new_n5715_));
AND2X2 AND2X2_2571 ( .A(_abc_40319_new_n5716_), .B(_abc_40319_new_n5717_), .Y(_abc_40319_new_n5718_));
AND2X2 AND2X2_2572 ( .A(_abc_40319_new_n5718_), .B(_abc_40319_new_n4272_), .Y(_abc_40319_new_n5719_));
AND2X2 AND2X2_2573 ( .A(_abc_40319_new_n1970_), .B(_abc_40319_new_n1169_), .Y(_abc_40319_new_n5720_));
AND2X2 AND2X2_2574 ( .A(_abc_40319_new_n3051_), .B(_abc_40319_new_n1152_), .Y(_abc_40319_new_n5721_));
AND2X2 AND2X2_2575 ( .A(_abc_40319_new_n4271_), .B(_abc_40319_new_n5721_), .Y(_abc_40319_new_n5722_));
AND2X2 AND2X2_2576 ( .A(_abc_40319_new_n4309_), .B(REG2_REG_29_), .Y(_abc_40319_new_n5723_));
AND2X2 AND2X2_2577 ( .A(_abc_40319_new_n1064_), .B(_abc_40319_new_n582_), .Y(_abc_40319_new_n5730_));
AND2X2 AND2X2_2578 ( .A(_abc_40319_new_n5468_), .B(_abc_40319_new_n5731_), .Y(_abc_40319_new_n5732_));
AND2X2 AND2X2_2579 ( .A(_abc_40319_new_n5469_), .B(D_REG_0_), .Y(_abc_40319_new_n5733_));
AND2X2 AND2X2_258 ( .A(_abc_40319_new_n1073_), .B(_abc_40319_new_n1075_), .Y(_abc_40319_new_n1076_));
AND2X2 AND2X2_2580 ( .A(_abc_40319_new_n5469_), .B(D_REG_1_), .Y(_abc_40319_new_n5736_));
AND2X2 AND2X2_2581 ( .A(_abc_40319_new_n5468_), .B(_abc_40319_new_n1075_), .Y(_abc_40319_new_n5737_));
AND2X2 AND2X2_2582 ( .A(_abc_40319_new_n5740_), .B(_abc_40319_new_n5741_), .Y(_abc_40319_new_n5742_));
AND2X2 AND2X2_2583 ( .A(_abc_40319_new_n4269_), .B(_abc_40319_new_n5742_), .Y(_abc_40319_new_n5743_));
AND2X2 AND2X2_2584 ( .A(_abc_40319_new_n5743_), .B(_abc_40319_new_n4265_), .Y(_abc_40319_new_n5744_));
AND2X2 AND2X2_2585 ( .A(_abc_40319_new_n4799_), .B(_abc_40319_new_n1167_), .Y(_abc_40319_new_n5745_));
AND2X2 AND2X2_2586 ( .A(_abc_40319_new_n4815_), .B(_abc_40319_new_n5405_), .Y(_abc_40319_new_n5746_));
AND2X2 AND2X2_2587 ( .A(_abc_40319_new_n1876_), .B(_abc_40319_new_n4310_), .Y(_abc_40319_new_n5747_));
AND2X2 AND2X2_2588 ( .A(_abc_40319_new_n5751_), .B(_abc_40319_new_n5744_), .Y(_abc_40319_new_n5752_));
AND2X2 AND2X2_2589 ( .A(_abc_40319_new_n5753_), .B(REG0_REG_20_), .Y(_abc_40319_new_n5754_));
AND2X2 AND2X2_259 ( .A(_abc_40319_new_n1077_), .B(_abc_40319_new_n1106_), .Y(_abc_40319_new_n1107_));
AND2X2 AND2X2_2590 ( .A(_abc_40319_new_n3137_), .B(_abc_40319_new_n1167_), .Y(_abc_40319_new_n5757_));
AND2X2 AND2X2_2591 ( .A(_abc_40319_new_n930_), .B(_abc_40319_new_n752_), .Y(_abc_40319_new_n5758_));
AND2X2 AND2X2_2592 ( .A(_abc_40319_new_n5760_), .B(_abc_40319_new_n5744_), .Y(_abc_40319_new_n5761_));
AND2X2 AND2X2_2593 ( .A(_abc_40319_new_n5753_), .B(REG0_REG_0_), .Y(_abc_40319_new_n5762_));
AND2X2 AND2X2_2594 ( .A(_abc_40319_new_n5426_), .B(_abc_40319_new_n1167_), .Y(_abc_40319_new_n5765_));
AND2X2 AND2X2_2595 ( .A(_abc_40319_new_n5768_), .B(_abc_40319_new_n5744_), .Y(_abc_40319_new_n5769_));
AND2X2 AND2X2_2596 ( .A(_abc_40319_new_n5753_), .B(REG0_REG_1_), .Y(_abc_40319_new_n5770_));
AND2X2 AND2X2_2597 ( .A(_abc_40319_new_n5390_), .B(_abc_40319_new_n1167_), .Y(_abc_40319_new_n5773_));
AND2X2 AND2X2_2598 ( .A(_abc_40319_new_n5775_), .B(_abc_40319_new_n5744_), .Y(_abc_40319_new_n5776_));
AND2X2 AND2X2_2599 ( .A(_abc_40319_new_n5753_), .B(REG0_REG_2_), .Y(_abc_40319_new_n5777_));
AND2X2 AND2X2_26 ( .A(_abc_40319_new_n579_), .B(_abc_40319_new_n577_), .Y(_abc_40319_new_n580_));
AND2X2 AND2X2_260 ( .A(_abc_40319_new_n1068_), .B(_abc_40319_new_n1065_), .Y(_abc_40319_new_n1110_));
AND2X2 AND2X2_2600 ( .A(_abc_40319_new_n5366_), .B(_abc_40319_new_n1167_), .Y(_abc_40319_new_n5780_));
AND2X2 AND2X2_2601 ( .A(_abc_40319_new_n5378_), .B(_abc_40319_new_n5405_), .Y(_abc_40319_new_n5781_));
AND2X2 AND2X2_2602 ( .A(_abc_40319_new_n5784_), .B(_abc_40319_new_n5744_), .Y(_abc_40319_new_n5785_));
AND2X2 AND2X2_2603 ( .A(_abc_40319_new_n5753_), .B(REG0_REG_3_), .Y(_abc_40319_new_n5786_));
AND2X2 AND2X2_2604 ( .A(_abc_40319_new_n5303_), .B(_abc_40319_new_n1167_), .Y(_abc_40319_new_n5789_));
AND2X2 AND2X2_2605 ( .A(_abc_40319_new_n5317_), .B(_abc_40319_new_n5405_), .Y(_abc_40319_new_n5790_));
AND2X2 AND2X2_2606 ( .A(_abc_40319_new_n5793_), .B(_abc_40319_new_n5744_), .Y(_abc_40319_new_n5794_));
AND2X2 AND2X2_2607 ( .A(_abc_40319_new_n5753_), .B(REG0_REG_4_), .Y(_abc_40319_new_n5795_));
AND2X2 AND2X2_2608 ( .A(_abc_40319_new_n5335_), .B(_abc_40319_new_n1167_), .Y(_abc_40319_new_n5798_));
AND2X2 AND2X2_2609 ( .A(_abc_40319_new_n5347_), .B(_abc_40319_new_n5405_), .Y(_abc_40319_new_n5799_));
AND2X2 AND2X2_261 ( .A(_abc_40319_new_n1109_), .B(_abc_40319_new_n1111_), .Y(_abc_40319_new_n1112_));
AND2X2 AND2X2_2610 ( .A(_abc_40319_new_n5802_), .B(_abc_40319_new_n5744_), .Y(_abc_40319_new_n5803_));
AND2X2 AND2X2_2611 ( .A(_abc_40319_new_n5753_), .B(REG0_REG_5_), .Y(_abc_40319_new_n5804_));
AND2X2 AND2X2_2612 ( .A(_abc_40319_new_n5276_), .B(_abc_40319_new_n5405_), .Y(_abc_40319_new_n5807_));
AND2X2 AND2X2_2613 ( .A(_abc_40319_new_n5268_), .B(_abc_40319_new_n1167_), .Y(_abc_40319_new_n5809_));
AND2X2 AND2X2_2614 ( .A(_abc_40319_new_n5811_), .B(_abc_40319_new_n5744_), .Y(_abc_40319_new_n5812_));
AND2X2 AND2X2_2615 ( .A(_abc_40319_new_n5753_), .B(REG0_REG_6_), .Y(_abc_40319_new_n5813_));
AND2X2 AND2X2_2616 ( .A(_abc_40319_new_n5231_), .B(_abc_40319_new_n1167_), .Y(_abc_40319_new_n5816_));
AND2X2 AND2X2_2617 ( .A(_abc_40319_new_n5239_), .B(_abc_40319_new_n5405_), .Y(_abc_40319_new_n5817_));
AND2X2 AND2X2_2618 ( .A(_abc_40319_new_n5820_), .B(_abc_40319_new_n5744_), .Y(_abc_40319_new_n5821_));
AND2X2 AND2X2_2619 ( .A(_abc_40319_new_n5753_), .B(REG0_REG_7_), .Y(_abc_40319_new_n5822_));
AND2X2 AND2X2_262 ( .A(_abc_40319_new_n1108_), .B(_abc_40319_new_n1112_), .Y(_abc_40319_new_n1113_));
AND2X2 AND2X2_2620 ( .A(_abc_40319_new_n5200_), .B(_abc_40319_new_n1167_), .Y(_abc_40319_new_n5825_));
AND2X2 AND2X2_2621 ( .A(_abc_40319_new_n5208_), .B(_abc_40319_new_n5405_), .Y(_abc_40319_new_n5826_));
AND2X2 AND2X2_2622 ( .A(_abc_40319_new_n5829_), .B(_abc_40319_new_n5744_), .Y(_abc_40319_new_n5830_));
AND2X2 AND2X2_2623 ( .A(_abc_40319_new_n5753_), .B(REG0_REG_8_), .Y(_abc_40319_new_n5831_));
AND2X2 AND2X2_2624 ( .A(_abc_40319_new_n5168_), .B(_abc_40319_new_n1167_), .Y(_abc_40319_new_n5834_));
AND2X2 AND2X2_2625 ( .A(_abc_40319_new_n5176_), .B(_abc_40319_new_n5405_), .Y(_abc_40319_new_n5835_));
AND2X2 AND2X2_2626 ( .A(_abc_40319_new_n5838_), .B(_abc_40319_new_n5744_), .Y(_abc_40319_new_n5839_));
AND2X2 AND2X2_2627 ( .A(_abc_40319_new_n5753_), .B(REG0_REG_9_), .Y(_abc_40319_new_n5840_));
AND2X2 AND2X2_2628 ( .A(_abc_40319_new_n5137_), .B(_abc_40319_new_n1167_), .Y(_abc_40319_new_n5843_));
AND2X2 AND2X2_2629 ( .A(_abc_40319_new_n5145_), .B(_abc_40319_new_n5405_), .Y(_abc_40319_new_n5844_));
AND2X2 AND2X2_263 ( .A(_abc_40319_new_n1113_), .B(_abc_40319_new_n1076_), .Y(_abc_40319_new_n1114_));
AND2X2 AND2X2_2630 ( .A(_abc_40319_new_n5848_), .B(_abc_40319_new_n5744_), .Y(_abc_40319_new_n5849_));
AND2X2 AND2X2_2631 ( .A(_abc_40319_new_n5753_), .B(REG0_REG_10_), .Y(_abc_40319_new_n5850_));
AND2X2 AND2X2_2632 ( .A(_abc_40319_new_n5103_), .B(_abc_40319_new_n1167_), .Y(_abc_40319_new_n5853_));
AND2X2 AND2X2_2633 ( .A(_abc_40319_new_n5111_), .B(_abc_40319_new_n5405_), .Y(_abc_40319_new_n5854_));
AND2X2 AND2X2_2634 ( .A(_abc_40319_new_n5857_), .B(_abc_40319_new_n5744_), .Y(_abc_40319_new_n5858_));
AND2X2 AND2X2_2635 ( .A(_abc_40319_new_n5753_), .B(REG0_REG_11_), .Y(_abc_40319_new_n5859_));
AND2X2 AND2X2_2636 ( .A(_abc_40319_new_n5067_), .B(_abc_40319_new_n1167_), .Y(_abc_40319_new_n5862_));
AND2X2 AND2X2_2637 ( .A(_abc_40319_new_n5075_), .B(_abc_40319_new_n5405_), .Y(_abc_40319_new_n5863_));
AND2X2 AND2X2_2638 ( .A(_abc_40319_new_n5867_), .B(_abc_40319_new_n5744_), .Y(_abc_40319_new_n5868_));
AND2X2 AND2X2_2639 ( .A(_abc_40319_new_n5753_), .B(REG0_REG_12_), .Y(_abc_40319_new_n5869_));
AND2X2 AND2X2_264 ( .A(_abc_40319_new_n671_), .B(_abc_40319_new_n698_), .Y(_abc_40319_new_n1116_));
AND2X2 AND2X2_2640 ( .A(_abc_40319_new_n5036_), .B(_abc_40319_new_n1167_), .Y(_abc_40319_new_n5872_));
AND2X2 AND2X2_2641 ( .A(_abc_40319_new_n5044_), .B(_abc_40319_new_n5405_), .Y(_abc_40319_new_n5873_));
AND2X2 AND2X2_2642 ( .A(_abc_40319_new_n5877_), .B(_abc_40319_new_n5744_), .Y(_abc_40319_new_n5878_));
AND2X2 AND2X2_2643 ( .A(_abc_40319_new_n5753_), .B(REG0_REG_13_), .Y(_abc_40319_new_n5879_));
AND2X2 AND2X2_2644 ( .A(_abc_40319_new_n5010_), .B(_abc_40319_new_n5405_), .Y(_abc_40319_new_n5882_));
AND2X2 AND2X2_2645 ( .A(_abc_40319_new_n5002_), .B(_abc_40319_new_n1167_), .Y(_abc_40319_new_n5884_));
AND2X2 AND2X2_2646 ( .A(_abc_40319_new_n5886_), .B(_abc_40319_new_n5744_), .Y(_abc_40319_new_n5887_));
AND2X2 AND2X2_2647 ( .A(_abc_40319_new_n5753_), .B(REG0_REG_14_), .Y(_abc_40319_new_n5888_));
AND2X2 AND2X2_2648 ( .A(_abc_40319_new_n4973_), .B(_abc_40319_new_n1167_), .Y(_abc_40319_new_n5891_));
AND2X2 AND2X2_2649 ( .A(_abc_40319_new_n4981_), .B(_abc_40319_new_n5405_), .Y(_abc_40319_new_n5892_));
AND2X2 AND2X2_265 ( .A(_abc_40319_new_n1117_), .B(_abc_40319_new_n1115_), .Y(_abc_40319_new_n1118_));
AND2X2 AND2X2_2650 ( .A(_abc_40319_new_n5896_), .B(_abc_40319_new_n5744_), .Y(_abc_40319_new_n5897_));
AND2X2 AND2X2_2651 ( .A(_abc_40319_new_n5753_), .B(REG0_REG_15_), .Y(_abc_40319_new_n5898_));
AND2X2 AND2X2_2652 ( .A(_abc_40319_new_n4941_), .B(_abc_40319_new_n1167_), .Y(_abc_40319_new_n5901_));
AND2X2 AND2X2_2653 ( .A(_abc_40319_new_n4949_), .B(_abc_40319_new_n5405_), .Y(_abc_40319_new_n5902_));
AND2X2 AND2X2_2654 ( .A(_abc_40319_new_n5906_), .B(_abc_40319_new_n5744_), .Y(_abc_40319_new_n5907_));
AND2X2 AND2X2_2655 ( .A(_abc_40319_new_n5753_), .B(REG0_REG_16_), .Y(_abc_40319_new_n5908_));
AND2X2 AND2X2_2656 ( .A(_abc_40319_new_n4913_), .B(_abc_40319_new_n5405_), .Y(_abc_40319_new_n5911_));
AND2X2 AND2X2_2657 ( .A(_abc_40319_new_n4898_), .B(_abc_40319_new_n1167_), .Y(_abc_40319_new_n5914_));
AND2X2 AND2X2_2658 ( .A(_abc_40319_new_n5916_), .B(_abc_40319_new_n5744_), .Y(_abc_40319_new_n5917_));
AND2X2 AND2X2_2659 ( .A(_abc_40319_new_n5753_), .B(REG0_REG_17_), .Y(_abc_40319_new_n5918_));
AND2X2 AND2X2_266 ( .A(_abc_40319_new_n663_), .B(_abc_40319_new_n613_), .Y(_abc_40319_new_n1119_));
AND2X2 AND2X2_2660 ( .A(_abc_40319_new_n4863_), .B(_abc_40319_new_n1167_), .Y(_abc_40319_new_n5921_));
AND2X2 AND2X2_2661 ( .A(_abc_40319_new_n4878_), .B(_abc_40319_new_n5405_), .Y(_abc_40319_new_n5922_));
AND2X2 AND2X2_2662 ( .A(_abc_40319_new_n1828_), .B(_abc_40319_new_n4310_), .Y(_abc_40319_new_n5923_));
AND2X2 AND2X2_2663 ( .A(_abc_40319_new_n5927_), .B(_abc_40319_new_n5744_), .Y(_abc_40319_new_n5928_));
AND2X2 AND2X2_2664 ( .A(_abc_40319_new_n5753_), .B(REG0_REG_18_), .Y(_abc_40319_new_n5929_));
AND2X2 AND2X2_2665 ( .A(_abc_40319_new_n4832_), .B(_abc_40319_new_n1167_), .Y(_abc_40319_new_n5932_));
AND2X2 AND2X2_2666 ( .A(_abc_40319_new_n4846_), .B(_abc_40319_new_n5405_), .Y(_abc_40319_new_n5933_));
AND2X2 AND2X2_2667 ( .A(_abc_40319_new_n1852_), .B(_abc_40319_new_n4310_), .Y(_abc_40319_new_n5934_));
AND2X2 AND2X2_2668 ( .A(_abc_40319_new_n5938_), .B(_abc_40319_new_n5744_), .Y(_abc_40319_new_n5939_));
AND2X2 AND2X2_2669 ( .A(_abc_40319_new_n5753_), .B(REG0_REG_19_), .Y(_abc_40319_new_n5940_));
AND2X2 AND2X2_267 ( .A(_abc_40319_new_n1119_), .B(STATE_REG), .Y(_abc_40319_new_n1120_));
AND2X2 AND2X2_2670 ( .A(_abc_40319_new_n4779_), .B(_abc_40319_new_n5405_), .Y(_abc_40319_new_n5943_));
AND2X2 AND2X2_2671 ( .A(_abc_40319_new_n1340_), .B(_abc_40319_new_n4310_), .Y(_abc_40319_new_n5944_));
AND2X2 AND2X2_2672 ( .A(_abc_40319_new_n4766_), .B(_abc_40319_new_n1167_), .Y(_abc_40319_new_n5947_));
AND2X2 AND2X2_2673 ( .A(_abc_40319_new_n5949_), .B(_abc_40319_new_n5744_), .Y(_abc_40319_new_n5950_));
AND2X2 AND2X2_2674 ( .A(_abc_40319_new_n5753_), .B(REG0_REG_21_), .Y(_abc_40319_new_n5951_));
AND2X2 AND2X2_2675 ( .A(_abc_40319_new_n4734_), .B(_abc_40319_new_n1167_), .Y(_abc_40319_new_n5954_));
AND2X2 AND2X2_2676 ( .A(_abc_40319_new_n4742_), .B(_abc_40319_new_n5405_), .Y(_abc_40319_new_n5955_));
AND2X2 AND2X2_2677 ( .A(_abc_40319_new_n1317_), .B(_abc_40319_new_n4310_), .Y(_abc_40319_new_n5956_));
AND2X2 AND2X2_2678 ( .A(_abc_40319_new_n5960_), .B(_abc_40319_new_n5744_), .Y(_abc_40319_new_n5961_));
AND2X2 AND2X2_2679 ( .A(_abc_40319_new_n5753_), .B(REG0_REG_22_), .Y(_abc_40319_new_n5962_));
AND2X2 AND2X2_268 ( .A(_abc_40319_new_n1120_), .B(_abc_40319_new_n1118_), .Y(_abc_40319_new_n1121_));
AND2X2 AND2X2_2680 ( .A(_abc_40319_new_n4703_), .B(_abc_40319_new_n1167_), .Y(_abc_40319_new_n5965_));
AND2X2 AND2X2_2681 ( .A(_abc_40319_new_n4711_), .B(_abc_40319_new_n5405_), .Y(_abc_40319_new_n5966_));
AND2X2 AND2X2_2682 ( .A(_abc_40319_new_n1285_), .B(_abc_40319_new_n4310_), .Y(_abc_40319_new_n5967_));
AND2X2 AND2X2_2683 ( .A(_abc_40319_new_n5971_), .B(_abc_40319_new_n5744_), .Y(_abc_40319_new_n5972_));
AND2X2 AND2X2_2684 ( .A(_abc_40319_new_n5753_), .B(REG0_REG_23_), .Y(_abc_40319_new_n5973_));
AND2X2 AND2X2_2685 ( .A(_abc_40319_new_n4639_), .B(_abc_40319_new_n1167_), .Y(_abc_40319_new_n5976_));
AND2X2 AND2X2_2686 ( .A(_abc_40319_new_n4669_), .B(_abc_40319_new_n5405_), .Y(_abc_40319_new_n5977_));
AND2X2 AND2X2_2687 ( .A(_abc_40319_new_n1260_), .B(_abc_40319_new_n4310_), .Y(_abc_40319_new_n5978_));
AND2X2 AND2X2_2688 ( .A(_abc_40319_new_n5982_), .B(_abc_40319_new_n5744_), .Y(_abc_40319_new_n5983_));
AND2X2 AND2X2_2689 ( .A(_abc_40319_new_n5753_), .B(REG0_REG_24_), .Y(_abc_40319_new_n5984_));
AND2X2 AND2X2_269 ( .A(_abc_40319_new_n1114_), .B(_abc_40319_new_n1121_), .Y(_abc_40319_new_n1122_));
AND2X2 AND2X2_2690 ( .A(_abc_40319_new_n4608_), .B(_abc_40319_new_n1167_), .Y(_abc_40319_new_n5987_));
AND2X2 AND2X2_2691 ( .A(_abc_40319_new_n4623_), .B(_abc_40319_new_n5405_), .Y(_abc_40319_new_n5988_));
AND2X2 AND2X2_2692 ( .A(_abc_40319_new_n1235_), .B(_abc_40319_new_n4310_), .Y(_abc_40319_new_n5989_));
AND2X2 AND2X2_2693 ( .A(_abc_40319_new_n5993_), .B(_abc_40319_new_n5744_), .Y(_abc_40319_new_n5994_));
AND2X2 AND2X2_2694 ( .A(_abc_40319_new_n5753_), .B(REG0_REG_25_), .Y(_abc_40319_new_n5995_));
AND2X2 AND2X2_2695 ( .A(_abc_40319_new_n4578_), .B(_abc_40319_new_n1167_), .Y(_abc_40319_new_n5998_));
AND2X2 AND2X2_2696 ( .A(_abc_40319_new_n4592_), .B(_abc_40319_new_n5405_), .Y(_abc_40319_new_n5999_));
AND2X2 AND2X2_2697 ( .A(_abc_40319_new_n1210_), .B(_abc_40319_new_n4310_), .Y(_abc_40319_new_n6000_));
AND2X2 AND2X2_2698 ( .A(_abc_40319_new_n6004_), .B(_abc_40319_new_n5744_), .Y(_abc_40319_new_n6005_));
AND2X2 AND2X2_2699 ( .A(_abc_40319_new_n5753_), .B(REG0_REG_26_), .Y(_abc_40319_new_n6006_));
AND2X2 AND2X2_27 ( .A(_abc_40319_new_n581_), .B(_abc_40319_new_n527_), .Y(_abc_40319_new_n582_));
AND2X2 AND2X2_270 ( .A(_abc_40319_new_n984_), .B(_abc_40319_new_n1123_), .Y(_abc_40319_new_n1124_));
AND2X2 AND2X2_2700 ( .A(_abc_40319_new_n4537_), .B(_abc_40319_new_n1167_), .Y(_abc_40319_new_n6009_));
AND2X2 AND2X2_2701 ( .A(_abc_40319_new_n4553_), .B(_abc_40319_new_n5405_), .Y(_abc_40319_new_n6010_));
AND2X2 AND2X2_2702 ( .A(_abc_40319_new_n1980_), .B(_abc_40319_new_n4310_), .Y(_abc_40319_new_n6011_));
AND2X2 AND2X2_2703 ( .A(_abc_40319_new_n6015_), .B(_abc_40319_new_n5744_), .Y(_abc_40319_new_n6016_));
AND2X2 AND2X2_2704 ( .A(_abc_40319_new_n5753_), .B(REG0_REG_27_), .Y(_abc_40319_new_n6017_));
AND2X2 AND2X2_2705 ( .A(_abc_40319_new_n4493_), .B(_abc_40319_new_n1167_), .Y(_abc_40319_new_n6020_));
AND2X2 AND2X2_2706 ( .A(_abc_40319_new_n4516_), .B(_abc_40319_new_n5405_), .Y(_abc_40319_new_n6021_));
AND2X2 AND2X2_2707 ( .A(_abc_40319_new_n2123_), .B(_abc_40319_new_n4310_), .Y(_abc_40319_new_n6022_));
AND2X2 AND2X2_2708 ( .A(_abc_40319_new_n6026_), .B(_abc_40319_new_n5744_), .Y(_abc_40319_new_n6027_));
AND2X2 AND2X2_2709 ( .A(_abc_40319_new_n5753_), .B(REG0_REG_28_), .Y(_abc_40319_new_n6028_));
AND2X2 AND2X2_271 ( .A(_abc_40319_new_n1126_), .B(_abc_40319_new_n1057_), .Y(_abc_40319_new_n1127_));
AND2X2 AND2X2_2710 ( .A(_abc_40319_new_n5704_), .B(_abc_40319_new_n1167_), .Y(_abc_40319_new_n6031_));
AND2X2 AND2X2_2711 ( .A(_abc_40319_new_n5718_), .B(_abc_40319_new_n5405_), .Y(_abc_40319_new_n6032_));
AND2X2 AND2X2_2712 ( .A(_abc_40319_new_n6036_), .B(_abc_40319_new_n5744_), .Y(_abc_40319_new_n6037_));
AND2X2 AND2X2_2713 ( .A(_abc_40319_new_n5753_), .B(REG0_REG_29_), .Y(_abc_40319_new_n6038_));
AND2X2 AND2X2_2714 ( .A(_abc_40319_new_n4323_), .B(_abc_40319_new_n5405_), .Y(_abc_40319_new_n6041_));
AND2X2 AND2X2_2715 ( .A(_abc_40319_new_n3069_), .B(_abc_40319_new_n1152_), .Y(_abc_40319_new_n6042_));
AND2X2 AND2X2_2716 ( .A(_abc_40319_new_n6044_), .B(_abc_40319_new_n5744_), .Y(_abc_40319_new_n6045_));
AND2X2 AND2X2_2717 ( .A(_abc_40319_new_n5753_), .B(REG0_REG_30_), .Y(_abc_40319_new_n6046_));
AND2X2 AND2X2_2718 ( .A(_abc_40319_new_n4307_), .B(_abc_40319_new_n5405_), .Y(_abc_40319_new_n6049_));
AND2X2 AND2X2_2719 ( .A(_abc_40319_new_n2553_), .B(_abc_40319_new_n1152_), .Y(_abc_40319_new_n6050_));
AND2X2 AND2X2_272 ( .A(_abc_40319_new_n1129_), .B(_abc_40319_new_n1122_), .Y(_abc_40319_new_n1130_));
AND2X2 AND2X2_2720 ( .A(_abc_40319_new_n6052_), .B(_abc_40319_new_n5744_), .Y(_abc_40319_new_n6053_));
AND2X2 AND2X2_2721 ( .A(_abc_40319_new_n5753_), .B(REG0_REG_31_), .Y(_abc_40319_new_n6054_));
AND2X2 AND2X2_2722 ( .A(_abc_40319_new_n5743_), .B(_abc_40319_new_n1112_), .Y(_abc_40319_new_n6057_));
AND2X2 AND2X2_2723 ( .A(_abc_40319_new_n5760_), .B(_abc_40319_new_n6057_), .Y(_abc_40319_new_n6058_));
AND2X2 AND2X2_2724 ( .A(_abc_40319_new_n6059_), .B(REG1_REG_0_), .Y(_abc_40319_new_n6060_));
AND2X2 AND2X2_2725 ( .A(_abc_40319_new_n5768_), .B(_abc_40319_new_n6057_), .Y(_abc_40319_new_n6063_));
AND2X2 AND2X2_2726 ( .A(_abc_40319_new_n6059_), .B(REG1_REG_1_), .Y(_abc_40319_new_n6064_));
AND2X2 AND2X2_2727 ( .A(_abc_40319_new_n5775_), .B(_abc_40319_new_n6057_), .Y(_abc_40319_new_n6067_));
AND2X2 AND2X2_2728 ( .A(_abc_40319_new_n6059_), .B(REG1_REG_2_), .Y(_abc_40319_new_n6068_));
AND2X2 AND2X2_2729 ( .A(_abc_40319_new_n5784_), .B(_abc_40319_new_n6057_), .Y(_abc_40319_new_n6071_));
AND2X2 AND2X2_273 ( .A(_abc_40319_new_n1130_), .B(_abc_40319_new_n1063_), .Y(_abc_40319_new_n1131_));
AND2X2 AND2X2_2730 ( .A(_abc_40319_new_n6059_), .B(REG1_REG_3_), .Y(_abc_40319_new_n6072_));
AND2X2 AND2X2_2731 ( .A(_abc_40319_new_n5793_), .B(_abc_40319_new_n6057_), .Y(_abc_40319_new_n6075_));
AND2X2 AND2X2_2732 ( .A(_abc_40319_new_n6059_), .B(REG1_REG_4_), .Y(_abc_40319_new_n6076_));
AND2X2 AND2X2_2733 ( .A(_abc_40319_new_n5802_), .B(_abc_40319_new_n6057_), .Y(_abc_40319_new_n6079_));
AND2X2 AND2X2_2734 ( .A(_abc_40319_new_n6059_), .B(REG1_REG_5_), .Y(_abc_40319_new_n6080_));
AND2X2 AND2X2_2735 ( .A(_abc_40319_new_n5811_), .B(_abc_40319_new_n6057_), .Y(_abc_40319_new_n6083_));
AND2X2 AND2X2_2736 ( .A(_abc_40319_new_n6059_), .B(REG1_REG_6_), .Y(_abc_40319_new_n6084_));
AND2X2 AND2X2_2737 ( .A(_abc_40319_new_n5820_), .B(_abc_40319_new_n6057_), .Y(_abc_40319_new_n6087_));
AND2X2 AND2X2_2738 ( .A(_abc_40319_new_n6059_), .B(REG1_REG_7_), .Y(_abc_40319_new_n6088_));
AND2X2 AND2X2_2739 ( .A(_abc_40319_new_n5829_), .B(_abc_40319_new_n6057_), .Y(_abc_40319_new_n6091_));
AND2X2 AND2X2_274 ( .A(_abc_40319_new_n672_), .B(_abc_40319_new_n699_), .Y(_abc_40319_new_n1132_));
AND2X2 AND2X2_2740 ( .A(_abc_40319_new_n6059_), .B(REG1_REG_8_), .Y(_abc_40319_new_n6092_));
AND2X2 AND2X2_2741 ( .A(_abc_40319_new_n5838_), .B(_abc_40319_new_n6057_), .Y(_abc_40319_new_n6095_));
AND2X2 AND2X2_2742 ( .A(_abc_40319_new_n6059_), .B(REG1_REG_9_), .Y(_abc_40319_new_n6096_));
AND2X2 AND2X2_2743 ( .A(_abc_40319_new_n5848_), .B(_abc_40319_new_n6057_), .Y(_abc_40319_new_n6099_));
AND2X2 AND2X2_2744 ( .A(_abc_40319_new_n6059_), .B(REG1_REG_10_), .Y(_abc_40319_new_n6100_));
AND2X2 AND2X2_2745 ( .A(_abc_40319_new_n5857_), .B(_abc_40319_new_n6057_), .Y(_abc_40319_new_n6103_));
AND2X2 AND2X2_2746 ( .A(_abc_40319_new_n6059_), .B(REG1_REG_11_), .Y(_abc_40319_new_n6104_));
AND2X2 AND2X2_2747 ( .A(_abc_40319_new_n5867_), .B(_abc_40319_new_n6057_), .Y(_abc_40319_new_n6107_));
AND2X2 AND2X2_2748 ( .A(_abc_40319_new_n6059_), .B(REG1_REG_12_), .Y(_abc_40319_new_n6108_));
AND2X2 AND2X2_2749 ( .A(_abc_40319_new_n5877_), .B(_abc_40319_new_n6057_), .Y(_abc_40319_new_n6111_));
AND2X2 AND2X2_275 ( .A(_abc_40319_new_n1120_), .B(_abc_40319_new_n1132_), .Y(_abc_40319_new_n1133_));
AND2X2 AND2X2_2750 ( .A(_abc_40319_new_n6059_), .B(REG1_REG_13_), .Y(_abc_40319_new_n6112_));
AND2X2 AND2X2_2751 ( .A(_abc_40319_new_n5886_), .B(_abc_40319_new_n6057_), .Y(_abc_40319_new_n6115_));
AND2X2 AND2X2_2752 ( .A(_abc_40319_new_n6059_), .B(REG1_REG_14_), .Y(_abc_40319_new_n6116_));
AND2X2 AND2X2_2753 ( .A(_abc_40319_new_n5896_), .B(_abc_40319_new_n6057_), .Y(_abc_40319_new_n6119_));
AND2X2 AND2X2_2754 ( .A(_abc_40319_new_n6059_), .B(REG1_REG_15_), .Y(_abc_40319_new_n6120_));
AND2X2 AND2X2_2755 ( .A(_abc_40319_new_n5906_), .B(_abc_40319_new_n6057_), .Y(_abc_40319_new_n6123_));
AND2X2 AND2X2_2756 ( .A(_abc_40319_new_n6059_), .B(REG1_REG_16_), .Y(_abc_40319_new_n6124_));
AND2X2 AND2X2_2757 ( .A(_abc_40319_new_n5916_), .B(_abc_40319_new_n6057_), .Y(_abc_40319_new_n6127_));
AND2X2 AND2X2_2758 ( .A(_abc_40319_new_n6059_), .B(REG1_REG_17_), .Y(_abc_40319_new_n6128_));
AND2X2 AND2X2_2759 ( .A(_abc_40319_new_n5927_), .B(_abc_40319_new_n6057_), .Y(_abc_40319_new_n6131_));
AND2X2 AND2X2_276 ( .A(_abc_40319_new_n1114_), .B(_abc_40319_new_n638_), .Y(_abc_40319_new_n1134_));
AND2X2 AND2X2_2760 ( .A(_abc_40319_new_n6059_), .B(REG1_REG_18_), .Y(_abc_40319_new_n6132_));
AND2X2 AND2X2_2761 ( .A(_abc_40319_new_n5938_), .B(_abc_40319_new_n6057_), .Y(_abc_40319_new_n6135_));
AND2X2 AND2X2_2762 ( .A(_abc_40319_new_n6059_), .B(REG1_REG_19_), .Y(_abc_40319_new_n6136_));
AND2X2 AND2X2_2763 ( .A(_abc_40319_new_n5751_), .B(_abc_40319_new_n6057_), .Y(_abc_40319_new_n6139_));
AND2X2 AND2X2_2764 ( .A(_abc_40319_new_n6059_), .B(REG1_REG_20_), .Y(_abc_40319_new_n6140_));
AND2X2 AND2X2_2765 ( .A(_abc_40319_new_n5949_), .B(_abc_40319_new_n6057_), .Y(_abc_40319_new_n6143_));
AND2X2 AND2X2_2766 ( .A(_abc_40319_new_n6059_), .B(REG1_REG_21_), .Y(_abc_40319_new_n6144_));
AND2X2 AND2X2_2767 ( .A(_abc_40319_new_n5960_), .B(_abc_40319_new_n6057_), .Y(_abc_40319_new_n6147_));
AND2X2 AND2X2_2768 ( .A(_abc_40319_new_n6059_), .B(REG1_REG_22_), .Y(_abc_40319_new_n6148_));
AND2X2 AND2X2_2769 ( .A(_abc_40319_new_n5971_), .B(_abc_40319_new_n6057_), .Y(_abc_40319_new_n6151_));
AND2X2 AND2X2_277 ( .A(_abc_40319_new_n1134_), .B(_abc_40319_new_n1010_), .Y(_abc_40319_new_n1135_));
AND2X2 AND2X2_2770 ( .A(_abc_40319_new_n6059_), .B(REG1_REG_23_), .Y(_abc_40319_new_n6152_));
AND2X2 AND2X2_2771 ( .A(_abc_40319_new_n5982_), .B(_abc_40319_new_n6057_), .Y(_abc_40319_new_n6155_));
AND2X2 AND2X2_2772 ( .A(_abc_40319_new_n6059_), .B(REG1_REG_24_), .Y(_abc_40319_new_n6156_));
AND2X2 AND2X2_2773 ( .A(_abc_40319_new_n5993_), .B(_abc_40319_new_n6057_), .Y(_abc_40319_new_n6159_));
AND2X2 AND2X2_2774 ( .A(_abc_40319_new_n6059_), .B(REG1_REG_25_), .Y(_abc_40319_new_n6160_));
AND2X2 AND2X2_2775 ( .A(_abc_40319_new_n6004_), .B(_abc_40319_new_n6057_), .Y(_abc_40319_new_n6163_));
AND2X2 AND2X2_2776 ( .A(_abc_40319_new_n6059_), .B(REG1_REG_26_), .Y(_abc_40319_new_n6164_));
AND2X2 AND2X2_2777 ( .A(_abc_40319_new_n6015_), .B(_abc_40319_new_n6057_), .Y(_abc_40319_new_n6167_));
AND2X2 AND2X2_2778 ( .A(_abc_40319_new_n6059_), .B(REG1_REG_27_), .Y(_abc_40319_new_n6168_));
AND2X2 AND2X2_2779 ( .A(_abc_40319_new_n6026_), .B(_abc_40319_new_n6057_), .Y(_abc_40319_new_n6171_));
AND2X2 AND2X2_278 ( .A(_abc_40319_new_n1039_), .B(REG3_REG_8_), .Y(_abc_40319_new_n1137_));
AND2X2 AND2X2_2780 ( .A(_abc_40319_new_n6059_), .B(REG1_REG_28_), .Y(_abc_40319_new_n6172_));
AND2X2 AND2X2_2781 ( .A(_abc_40319_new_n6036_), .B(_abc_40319_new_n6057_), .Y(_abc_40319_new_n6175_));
AND2X2 AND2X2_2782 ( .A(_abc_40319_new_n6059_), .B(REG1_REG_29_), .Y(_abc_40319_new_n6176_));
AND2X2 AND2X2_2783 ( .A(_abc_40319_new_n6044_), .B(_abc_40319_new_n6057_), .Y(_abc_40319_new_n6179_));
AND2X2 AND2X2_2784 ( .A(_abc_40319_new_n6059_), .B(REG1_REG_30_), .Y(_abc_40319_new_n6180_));
AND2X2 AND2X2_2785 ( .A(_abc_40319_new_n6052_), .B(_abc_40319_new_n6057_), .Y(_abc_40319_new_n6183_));
AND2X2 AND2X2_2786 ( .A(_abc_40319_new_n6059_), .B(REG1_REG_31_), .Y(_abc_40319_new_n6184_));
AND2X2 AND2X2_2787 ( .A(_abc_40319_new_n924_), .B(n1345), .Y(_abc_40319_new_n6187_));
AND2X2 AND2X2_2788 ( .A(_abc_40319_new_n6188_), .B(DATAO_REG_0_), .Y(_abc_40319_new_n6189_));
AND2X2 AND2X2_2789 ( .A(_abc_40319_new_n904_), .B(n1345), .Y(_abc_40319_new_n6192_));
AND2X2 AND2X2_279 ( .A(_abc_40319_new_n1138_), .B(_abc_40319_new_n1136_), .Y(_abc_40319_new_n1139_));
AND2X2 AND2X2_2790 ( .A(_abc_40319_new_n6188_), .B(DATAO_REG_1_), .Y(_abc_40319_new_n6193_));
AND2X2 AND2X2_2791 ( .A(_abc_40319_new_n865_), .B(n1345), .Y(_abc_40319_new_n6196_));
AND2X2 AND2X2_2792 ( .A(_abc_40319_new_n6188_), .B(DATAO_REG_2_), .Y(_abc_40319_new_n6197_));
AND2X2 AND2X2_2793 ( .A(_abc_40319_new_n829_), .B(n1345), .Y(_abc_40319_new_n6200_));
AND2X2 AND2X2_2794 ( .A(_abc_40319_new_n6188_), .B(DATAO_REG_3_), .Y(_abc_40319_new_n6201_));
AND2X2 AND2X2_2795 ( .A(_abc_40319_new_n795_), .B(n1345), .Y(_abc_40319_new_n6204_));
AND2X2 AND2X2_2796 ( .A(_abc_40319_new_n6188_), .B(DATAO_REG_4_), .Y(_abc_40319_new_n6205_));
AND2X2 AND2X2_2797 ( .A(_abc_40319_new_n746_), .B(n1345), .Y(_abc_40319_new_n6208_));
AND2X2 AND2X2_2798 ( .A(_abc_40319_new_n6188_), .B(DATAO_REG_5_), .Y(_abc_40319_new_n6209_));
AND2X2 AND2X2_2799 ( .A(_abc_40319_new_n1010_), .B(n1345), .Y(_abc_40319_new_n6212_));
AND2X2 AND2X2_28 ( .A(_abc_40319_new_n572_), .B(_abc_40319_new_n573_), .Y(_abc_40319_new_n584_));
AND2X2 AND2X2_280 ( .A(_abc_40319_new_n738_), .B(_abc_40319_new_n1139_), .Y(_abc_40319_new_n1140_));
AND2X2 AND2X2_2800 ( .A(_abc_40319_new_n6188_), .B(DATAO_REG_6_), .Y(_abc_40319_new_n6213_));
AND2X2 AND2X2_2801 ( .A(_abc_40319_new_n1046_), .B(n1345), .Y(_abc_40319_new_n6216_));
AND2X2 AND2X2_2802 ( .A(_abc_40319_new_n6188_), .B(DATAO_REG_7_), .Y(_abc_40319_new_n6217_));
AND2X2 AND2X2_2803 ( .A(_abc_40319_new_n1146_), .B(n1345), .Y(_abc_40319_new_n6220_));
AND2X2 AND2X2_2804 ( .A(_abc_40319_new_n6188_), .B(DATAO_REG_8_), .Y(_abc_40319_new_n6221_));
AND2X2 AND2X2_2805 ( .A(_abc_40319_new_n1625_), .B(n1345), .Y(_abc_40319_new_n6224_));
AND2X2 AND2X2_2806 ( .A(_abc_40319_new_n6188_), .B(DATAO_REG_9_), .Y(_abc_40319_new_n6225_));
AND2X2 AND2X2_2807 ( .A(_abc_40319_new_n1769_), .B(n1345), .Y(_abc_40319_new_n6228_));
AND2X2 AND2X2_2808 ( .A(_abc_40319_new_n6188_), .B(DATAO_REG_10_), .Y(_abc_40319_new_n6229_));
AND2X2 AND2X2_2809 ( .A(_abc_40319_new_n1735_), .B(n1345), .Y(_abc_40319_new_n6232_));
AND2X2 AND2X2_281 ( .A(_abc_40319_new_n722_), .B(REG1_REG_8_), .Y(_abc_40319_new_n1141_));
AND2X2 AND2X2_2810 ( .A(_abc_40319_new_n6188_), .B(DATAO_REG_11_), .Y(_abc_40319_new_n6233_));
AND2X2 AND2X2_2811 ( .A(_abc_40319_new_n1701_), .B(n1345), .Y(_abc_40319_new_n6236_));
AND2X2 AND2X2_2812 ( .A(_abc_40319_new_n6188_), .B(DATAO_REG_12_), .Y(_abc_40319_new_n6237_));
AND2X2 AND2X2_2813 ( .A(_abc_40319_new_n1667_), .B(n1345), .Y(_abc_40319_new_n6240_));
AND2X2 AND2X2_2814 ( .A(_abc_40319_new_n6188_), .B(DATAO_REG_13_), .Y(_abc_40319_new_n6241_));
AND2X2 AND2X2_2815 ( .A(_abc_40319_new_n1517_), .B(n1345), .Y(_abc_40319_new_n6244_));
AND2X2 AND2X2_2816 ( .A(_abc_40319_new_n6188_), .B(DATAO_REG_14_), .Y(_abc_40319_new_n6245_));
AND2X2 AND2X2_2817 ( .A(_abc_40319_new_n1483_), .B(n1345), .Y(_abc_40319_new_n6248_));
AND2X2 AND2X2_2818 ( .A(_abc_40319_new_n6188_), .B(DATAO_REG_15_), .Y(_abc_40319_new_n6249_));
AND2X2 AND2X2_2819 ( .A(_abc_40319_new_n1410_), .B(n1345), .Y(_abc_40319_new_n6252_));
AND2X2 AND2X2_282 ( .A(_abc_40319_new_n736_), .B(REG0_REG_8_), .Y(_abc_40319_new_n1143_));
AND2X2 AND2X2_2820 ( .A(_abc_40319_new_n6188_), .B(DATAO_REG_16_), .Y(_abc_40319_new_n6253_));
AND2X2 AND2X2_2821 ( .A(_abc_40319_new_n1444_), .B(n1345), .Y(_abc_40319_new_n6256_));
AND2X2 AND2X2_2822 ( .A(_abc_40319_new_n6188_), .B(DATAO_REG_17_), .Y(_abc_40319_new_n6257_));
AND2X2 AND2X2_2823 ( .A(_abc_40319_new_n1374_), .B(n1345), .Y(_abc_40319_new_n6260_));
AND2X2 AND2X2_2824 ( .A(_abc_40319_new_n6188_), .B(DATAO_REG_18_), .Y(_abc_40319_new_n6261_));
AND2X2 AND2X2_2825 ( .A(_abc_40319_new_n1828_), .B(n1345), .Y(_abc_40319_new_n6264_));
AND2X2 AND2X2_2826 ( .A(_abc_40319_new_n6188_), .B(DATAO_REG_19_), .Y(_abc_40319_new_n6265_));
AND2X2 AND2X2_2827 ( .A(_abc_40319_new_n1852_), .B(n1345), .Y(_abc_40319_new_n6268_));
AND2X2 AND2X2_2828 ( .A(_abc_40319_new_n6188_), .B(DATAO_REG_20_), .Y(_abc_40319_new_n6269_));
AND2X2 AND2X2_2829 ( .A(_abc_40319_new_n1876_), .B(n1345), .Y(_abc_40319_new_n6272_));
AND2X2 AND2X2_283 ( .A(_abc_40319_new_n733_), .B(REG2_REG_8_), .Y(_abc_40319_new_n1144_));
AND2X2 AND2X2_2830 ( .A(_abc_40319_new_n6188_), .B(DATAO_REG_21_), .Y(_abc_40319_new_n6273_));
AND2X2 AND2X2_2831 ( .A(_abc_40319_new_n1340_), .B(n1345), .Y(_abc_40319_new_n6276_));
AND2X2 AND2X2_2832 ( .A(_abc_40319_new_n6188_), .B(DATAO_REG_22_), .Y(_abc_40319_new_n6277_));
AND2X2 AND2X2_2833 ( .A(_abc_40319_new_n1317_), .B(n1345), .Y(_abc_40319_new_n6280_));
AND2X2 AND2X2_2834 ( .A(_abc_40319_new_n6188_), .B(DATAO_REG_23_), .Y(_abc_40319_new_n6281_));
AND2X2 AND2X2_2835 ( .A(_abc_40319_new_n1285_), .B(n1345), .Y(_abc_40319_new_n6284_));
AND2X2 AND2X2_2836 ( .A(_abc_40319_new_n6188_), .B(DATAO_REG_24_), .Y(_abc_40319_new_n6285_));
AND2X2 AND2X2_2837 ( .A(_abc_40319_new_n1260_), .B(n1345), .Y(_abc_40319_new_n6288_));
AND2X2 AND2X2_2838 ( .A(_abc_40319_new_n6188_), .B(DATAO_REG_25_), .Y(_abc_40319_new_n6289_));
AND2X2 AND2X2_2839 ( .A(_abc_40319_new_n1235_), .B(n1345), .Y(_abc_40319_new_n6292_));
AND2X2 AND2X2_284 ( .A(_abc_40319_new_n1114_), .B(_abc_40319_new_n639_), .Y(_abc_40319_new_n1147_));
AND2X2 AND2X2_2840 ( .A(_abc_40319_new_n6188_), .B(DATAO_REG_26_), .Y(_abc_40319_new_n6293_));
AND2X2 AND2X2_2841 ( .A(_abc_40319_new_n1210_), .B(n1345), .Y(_abc_40319_new_n6296_));
AND2X2 AND2X2_2842 ( .A(_abc_40319_new_n6188_), .B(DATAO_REG_27_), .Y(_abc_40319_new_n6297_));
AND2X2 AND2X2_2843 ( .A(_abc_40319_new_n1980_), .B(n1345), .Y(_abc_40319_new_n6300_));
AND2X2 AND2X2_2844 ( .A(_abc_40319_new_n6188_), .B(DATAO_REG_28_), .Y(_abc_40319_new_n6301_));
AND2X2 AND2X2_2845 ( .A(_abc_40319_new_n2123_), .B(n1345), .Y(_abc_40319_new_n6304_));
AND2X2 AND2X2_2846 ( .A(_abc_40319_new_n6188_), .B(DATAO_REG_29_), .Y(_abc_40319_new_n6305_));
AND2X2 AND2X2_2847 ( .A(_abc_40319_new_n3075_), .B(n1345), .Y(_abc_40319_new_n6308_));
AND2X2 AND2X2_2848 ( .A(_abc_40319_new_n6188_), .B(DATAO_REG_30_), .Y(_abc_40319_new_n6309_));
AND2X2 AND2X2_2849 ( .A(_abc_40319_new_n2560_), .B(n1345), .Y(_abc_40319_new_n6312_));
AND2X2 AND2X2_285 ( .A(_abc_40319_new_n1147_), .B(_abc_40319_new_n1146_), .Y(_abc_40319_new_n1148_));
AND2X2 AND2X2_2850 ( .A(_abc_40319_new_n6188_), .B(DATAO_REG_31_), .Y(_abc_40319_new_n6313_));
AND2X2 AND2X2_286 ( .A(_abc_40319_new_n1149_), .B(_abc_40319_new_n1133_), .Y(_abc_40319_new_n1150_));
AND2X2 AND2X2_287 ( .A(_abc_40319_new_n752_), .B(_abc_40319_new_n670_), .Y(_abc_40319_new_n1152_));
AND2X2 AND2X2_288 ( .A(_abc_40319_new_n1120_), .B(_abc_40319_new_n1152_), .Y(_abc_40319_new_n1153_));
AND2X2 AND2X2_289 ( .A(_abc_40319_new_n1118_), .B(STATE_REG), .Y(_abc_40319_new_n1154_));
AND2X2 AND2X2_29 ( .A(_abc_40319_new_n585_), .B(_abc_40319_new_n583_), .Y(_abc_40319_new_n586_));
AND2X2 AND2X2_290 ( .A(_abc_40319_new_n1151_), .B(_abc_40319_new_n1155_), .Y(_abc_40319_new_n1156_));
AND2X2 AND2X2_291 ( .A(_abc_40319_new_n1158_), .B(_abc_40319_new_n656_), .Y(_abc_40319_new_n1159_));
AND2X2 AND2X2_292 ( .A(_abc_40319_new_n1160_), .B(STATE_REG), .Y(_abc_40319_new_n1161_));
AND2X2 AND2X2_293 ( .A(_abc_40319_new_n1151_), .B(_abc_40319_new_n1133_), .Y(_abc_40319_new_n1163_));
AND2X2 AND2X2_294 ( .A(_abc_40319_new_n1164_), .B(_abc_40319_new_n1042_), .Y(_abc_40319_new_n1165_));
AND2X2 AND2X2_295 ( .A(_abc_40319_new_n645_), .B(_abc_40319_new_n697_), .Y(_abc_40319_new_n1166_));
AND2X2 AND2X2_296 ( .A(_abc_40319_new_n1166_), .B(_abc_40319_new_n671_), .Y(_abc_40319_new_n1167_));
AND2X2 AND2X2_297 ( .A(_abc_40319_new_n1167_), .B(_abc_40319_new_n751_), .Y(_abc_40319_new_n1168_));
AND2X2 AND2X2_298 ( .A(_abc_40319_new_n1120_), .B(_abc_40319_new_n1168_), .Y(_abc_40319_new_n1169_));
AND2X2 AND2X2_299 ( .A(_abc_40319_new_n1114_), .B(_abc_40319_new_n1153_), .Y(_abc_40319_new_n1170_));
AND2X2 AND2X2_3 ( .A(_abc_40319_new_n533_), .B(_abc_40319_new_n534_), .Y(_abc_40319_new_n535_));
AND2X2 AND2X2_30 ( .A(_abc_40319_new_n586_), .B(IR_REG_31_), .Y(_abc_40319_new_n587_));
AND2X2 AND2X2_300 ( .A(_abc_40319_new_n1171_), .B(_abc_40319_new_n1034_), .Y(_abc_40319_new_n1172_));
AND2X2 AND2X2_301 ( .A(n1336), .B(REG3_REG_7_), .Y(_abc_40319_new_n1174_));
AND2X2 AND2X2_302 ( .A(_abc_40319_new_n817_), .B(DATAI_27_), .Y(_abc_40319_new_n1180_));
AND2X2 AND2X2_303 ( .A(_abc_40319_new_n1180_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1181_));
AND2X2 AND2X2_304 ( .A(_abc_40319_new_n1137_), .B(REG3_REG_9_), .Y(_abc_40319_new_n1182_));
AND2X2 AND2X2_305 ( .A(_abc_40319_new_n1182_), .B(REG3_REG_10_), .Y(_abc_40319_new_n1183_));
AND2X2 AND2X2_306 ( .A(_abc_40319_new_n1183_), .B(REG3_REG_11_), .Y(_abc_40319_new_n1184_));
AND2X2 AND2X2_307 ( .A(REG3_REG_12_), .B(REG3_REG_13_), .Y(_abc_40319_new_n1185_));
AND2X2 AND2X2_308 ( .A(_abc_40319_new_n1184_), .B(_abc_40319_new_n1185_), .Y(_abc_40319_new_n1186_));
AND2X2 AND2X2_309 ( .A(REG3_REG_14_), .B(REG3_REG_15_), .Y(_abc_40319_new_n1187_));
AND2X2 AND2X2_31 ( .A(_abc_40319_new_n524_), .B(IR_REG_25_), .Y(_abc_40319_new_n588_));
AND2X2 AND2X2_310 ( .A(_abc_40319_new_n1186_), .B(_abc_40319_new_n1187_), .Y(_abc_40319_new_n1188_));
AND2X2 AND2X2_311 ( .A(REG3_REG_16_), .B(REG3_REG_17_), .Y(_abc_40319_new_n1189_));
AND2X2 AND2X2_312 ( .A(_abc_40319_new_n1188_), .B(_abc_40319_new_n1189_), .Y(_abc_40319_new_n1190_));
AND2X2 AND2X2_313 ( .A(_abc_40319_new_n1190_), .B(REG3_REG_18_), .Y(_abc_40319_new_n1191_));
AND2X2 AND2X2_314 ( .A(_abc_40319_new_n1191_), .B(REG3_REG_19_), .Y(_abc_40319_new_n1192_));
AND2X2 AND2X2_315 ( .A(_abc_40319_new_n1192_), .B(REG3_REG_20_), .Y(_abc_40319_new_n1193_));
AND2X2 AND2X2_316 ( .A(_abc_40319_new_n1193_), .B(REG3_REG_21_), .Y(_abc_40319_new_n1194_));
AND2X2 AND2X2_317 ( .A(_abc_40319_new_n1194_), .B(REG3_REG_22_), .Y(_abc_40319_new_n1195_));
AND2X2 AND2X2_318 ( .A(_abc_40319_new_n1195_), .B(REG3_REG_23_), .Y(_abc_40319_new_n1196_));
AND2X2 AND2X2_319 ( .A(_abc_40319_new_n1196_), .B(REG3_REG_24_), .Y(_abc_40319_new_n1197_));
AND2X2 AND2X2_32 ( .A(_abc_40319_new_n573_), .B(_abc_40319_new_n524_), .Y(_abc_40319_new_n590_));
AND2X2 AND2X2_320 ( .A(_abc_40319_new_n1197_), .B(REG3_REG_25_), .Y(_abc_40319_new_n1198_));
AND2X2 AND2X2_321 ( .A(_abc_40319_new_n1198_), .B(REG3_REG_26_), .Y(_abc_40319_new_n1199_));
AND2X2 AND2X2_322 ( .A(_abc_40319_new_n1199_), .B(REG3_REG_27_), .Y(_abc_40319_new_n1201_));
AND2X2 AND2X2_323 ( .A(_abc_40319_new_n1202_), .B(_abc_40319_new_n1200_), .Y(_abc_40319_new_n1203_));
AND2X2 AND2X2_324 ( .A(_abc_40319_new_n1203_), .B(_abc_40319_new_n738_), .Y(_abc_40319_new_n1204_));
AND2X2 AND2X2_325 ( .A(_abc_40319_new_n736_), .B(REG0_REG_27_), .Y(_abc_40319_new_n1205_));
AND2X2 AND2X2_326 ( .A(_abc_40319_new_n722_), .B(REG1_REG_27_), .Y(_abc_40319_new_n1206_));
AND2X2 AND2X2_327 ( .A(_abc_40319_new_n733_), .B(REG2_REG_27_), .Y(_abc_40319_new_n1207_));
AND2X2 AND2X2_328 ( .A(_abc_40319_new_n1210_), .B(_abc_40319_new_n705_), .Y(_abc_40319_new_n1211_));
AND2X2 AND2X2_329 ( .A(_abc_40319_new_n763_), .B(_abc_40319_new_n1180_), .Y(_abc_40319_new_n1213_));
AND2X2 AND2X2_33 ( .A(_abc_40319_new_n592_), .B(_abc_40319_new_n593_), .Y(_abc_40319_new_n594_));
AND2X2 AND2X2_330 ( .A(_abc_40319_new_n1210_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1214_));
AND2X2 AND2X2_331 ( .A(_abc_40319_new_n1216_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1217_));
AND2X2 AND2X2_332 ( .A(_abc_40319_new_n1215_), .B(_abc_40319_new_n768_), .Y(_abc_40319_new_n1218_));
AND2X2 AND2X2_333 ( .A(_abc_40319_new_n1219_), .B(_abc_40319_new_n1212_), .Y(_abc_40319_new_n1220_));
AND2X2 AND2X2_334 ( .A(_abc_40319_new_n1221_), .B(_abc_40319_new_n1222_), .Y(_abc_40319_new_n1223_));
AND2X2 AND2X2_335 ( .A(_abc_40319_new_n817_), .B(DATAI_26_), .Y(_abc_40319_new_n1224_));
AND2X2 AND2X2_336 ( .A(_abc_40319_new_n1224_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1225_));
AND2X2 AND2X2_337 ( .A(_abc_40319_new_n1226_), .B(_abc_40319_new_n1227_), .Y(_abc_40319_new_n1228_));
AND2X2 AND2X2_338 ( .A(_abc_40319_new_n1228_), .B(_abc_40319_new_n738_), .Y(_abc_40319_new_n1229_));
AND2X2 AND2X2_339 ( .A(_abc_40319_new_n733_), .B(REG2_REG_26_), .Y(_abc_40319_new_n1230_));
AND2X2 AND2X2_34 ( .A(_abc_40319_new_n595_), .B(_abc_40319_new_n591_), .Y(_abc_40319_new_n596_));
AND2X2 AND2X2_340 ( .A(_abc_40319_new_n736_), .B(REG0_REG_26_), .Y(_abc_40319_new_n1231_));
AND2X2 AND2X2_341 ( .A(_abc_40319_new_n722_), .B(REG1_REG_26_), .Y(_abc_40319_new_n1232_));
AND2X2 AND2X2_342 ( .A(_abc_40319_new_n1235_), .B(_abc_40319_new_n705_), .Y(_abc_40319_new_n1236_));
AND2X2 AND2X2_343 ( .A(_abc_40319_new_n763_), .B(_abc_40319_new_n1224_), .Y(_abc_40319_new_n1239_));
AND2X2 AND2X2_344 ( .A(_abc_40319_new_n1235_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1240_));
AND2X2 AND2X2_345 ( .A(_abc_40319_new_n1242_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1243_));
AND2X2 AND2X2_346 ( .A(_abc_40319_new_n1241_), .B(_abc_40319_new_n768_), .Y(_abc_40319_new_n1244_));
AND2X2 AND2X2_347 ( .A(_abc_40319_new_n1246_), .B(_abc_40319_new_n1238_), .Y(_abc_40319_new_n1247_));
AND2X2 AND2X2_348 ( .A(_abc_40319_new_n817_), .B(DATAI_25_), .Y(_abc_40319_new_n1249_));
AND2X2 AND2X2_349 ( .A(_abc_40319_new_n1249_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1250_));
AND2X2 AND2X2_35 ( .A(_abc_40319_new_n589_), .B(_abc_40319_new_n596_), .Y(_abc_40319_new_n597_));
AND2X2 AND2X2_350 ( .A(_abc_40319_new_n1251_), .B(_abc_40319_new_n1252_), .Y(_abc_40319_new_n1253_));
AND2X2 AND2X2_351 ( .A(_abc_40319_new_n1253_), .B(_abc_40319_new_n738_), .Y(_abc_40319_new_n1254_));
AND2X2 AND2X2_352 ( .A(_abc_40319_new_n722_), .B(REG1_REG_25_), .Y(_abc_40319_new_n1255_));
AND2X2 AND2X2_353 ( .A(_abc_40319_new_n736_), .B(REG0_REG_25_), .Y(_abc_40319_new_n1256_));
AND2X2 AND2X2_354 ( .A(_abc_40319_new_n733_), .B(REG2_REG_25_), .Y(_abc_40319_new_n1257_));
AND2X2 AND2X2_355 ( .A(_abc_40319_new_n1260_), .B(_abc_40319_new_n705_), .Y(_abc_40319_new_n1261_));
AND2X2 AND2X2_356 ( .A(_abc_40319_new_n763_), .B(_abc_40319_new_n1249_), .Y(_abc_40319_new_n1264_));
AND2X2 AND2X2_357 ( .A(_abc_40319_new_n1260_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1265_));
AND2X2 AND2X2_358 ( .A(_abc_40319_new_n1267_), .B(_abc_40319_new_n768_), .Y(_abc_40319_new_n1268_));
AND2X2 AND2X2_359 ( .A(_abc_40319_new_n1266_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1269_));
AND2X2 AND2X2_36 ( .A(_abc_40319_new_n597_), .B(_abc_40319_new_n582_), .Y(_abc_40319_new_n598_));
AND2X2 AND2X2_360 ( .A(_abc_40319_new_n1270_), .B(_abc_40319_new_n1263_), .Y(_abc_40319_new_n1271_));
AND2X2 AND2X2_361 ( .A(_abc_40319_new_n1248_), .B(_abc_40319_new_n1272_), .Y(_abc_40319_new_n1273_));
AND2X2 AND2X2_362 ( .A(_abc_40319_new_n817_), .B(DATAI_24_), .Y(_abc_40319_new_n1274_));
AND2X2 AND2X2_363 ( .A(_abc_40319_new_n1274_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1275_));
AND2X2 AND2X2_364 ( .A(_abc_40319_new_n1276_), .B(_abc_40319_new_n1277_), .Y(_abc_40319_new_n1278_));
AND2X2 AND2X2_365 ( .A(_abc_40319_new_n1278_), .B(_abc_40319_new_n738_), .Y(_abc_40319_new_n1279_));
AND2X2 AND2X2_366 ( .A(_abc_40319_new_n722_), .B(REG1_REG_24_), .Y(_abc_40319_new_n1280_));
AND2X2 AND2X2_367 ( .A(_abc_40319_new_n736_), .B(REG0_REG_24_), .Y(_abc_40319_new_n1281_));
AND2X2 AND2X2_368 ( .A(_abc_40319_new_n733_), .B(REG2_REG_24_), .Y(_abc_40319_new_n1282_));
AND2X2 AND2X2_369 ( .A(_abc_40319_new_n1285_), .B(_abc_40319_new_n705_), .Y(_abc_40319_new_n1286_));
AND2X2 AND2X2_37 ( .A(_abc_40319_new_n524_), .B(IR_REG_23_), .Y(_abc_40319_new_n599_));
AND2X2 AND2X2_370 ( .A(_abc_40319_new_n763_), .B(_abc_40319_new_n1274_), .Y(_abc_40319_new_n1288_));
AND2X2 AND2X2_371 ( .A(_abc_40319_new_n1285_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1289_));
AND2X2 AND2X2_372 ( .A(_abc_40319_new_n1291_), .B(_abc_40319_new_n768_), .Y(_abc_40319_new_n1292_));
AND2X2 AND2X2_373 ( .A(_abc_40319_new_n1290_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1293_));
AND2X2 AND2X2_374 ( .A(_abc_40319_new_n1295_), .B(_abc_40319_new_n1287_), .Y(_abc_40319_new_n1296_));
AND2X2 AND2X2_375 ( .A(_abc_40319_new_n1273_), .B(_abc_40319_new_n1296_), .Y(_abc_40319_new_n1297_));
AND2X2 AND2X2_376 ( .A(_abc_40319_new_n1245_), .B(_abc_40319_new_n1237_), .Y(_abc_40319_new_n1299_));
AND2X2 AND2X2_377 ( .A(_abc_40319_new_n1300_), .B(_abc_40319_new_n1301_), .Y(_abc_40319_new_n1302_));
AND2X2 AND2X2_378 ( .A(_abc_40319_new_n1298_), .B(_abc_40319_new_n1302_), .Y(_abc_40319_new_n1303_));
AND2X2 AND2X2_379 ( .A(_abc_40319_new_n817_), .B(DATAI_23_), .Y(_abc_40319_new_n1306_));
AND2X2 AND2X2_38 ( .A(_abc_40319_new_n553_), .B(_abc_40319_new_n561_), .Y(_abc_40319_new_n601_));
AND2X2 AND2X2_380 ( .A(_abc_40319_new_n1306_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1307_));
AND2X2 AND2X2_381 ( .A(_abc_40319_new_n1308_), .B(_abc_40319_new_n1309_), .Y(_abc_40319_new_n1310_));
AND2X2 AND2X2_382 ( .A(_abc_40319_new_n1310_), .B(_abc_40319_new_n738_), .Y(_abc_40319_new_n1311_));
AND2X2 AND2X2_383 ( .A(_abc_40319_new_n736_), .B(REG0_REG_23_), .Y(_abc_40319_new_n1312_));
AND2X2 AND2X2_384 ( .A(_abc_40319_new_n722_), .B(REG1_REG_23_), .Y(_abc_40319_new_n1313_));
AND2X2 AND2X2_385 ( .A(_abc_40319_new_n733_), .B(REG2_REG_23_), .Y(_abc_40319_new_n1314_));
AND2X2 AND2X2_386 ( .A(_abc_40319_new_n1317_), .B(_abc_40319_new_n705_), .Y(_abc_40319_new_n1318_));
AND2X2 AND2X2_387 ( .A(_abc_40319_new_n763_), .B(_abc_40319_new_n1306_), .Y(_abc_40319_new_n1320_));
AND2X2 AND2X2_388 ( .A(_abc_40319_new_n1317_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1321_));
AND2X2 AND2X2_389 ( .A(_abc_40319_new_n1325_), .B(_abc_40319_new_n1323_), .Y(_abc_40319_new_n1326_));
AND2X2 AND2X2_39 ( .A(_abc_40319_new_n607_), .B(_abc_40319_new_n554_), .Y(_abc_40319_new_n608_));
AND2X2 AND2X2_390 ( .A(_abc_40319_new_n1326_), .B(_abc_40319_new_n1319_), .Y(_abc_40319_new_n1327_));
AND2X2 AND2X2_391 ( .A(_abc_40319_new_n817_), .B(DATAI_22_), .Y(_abc_40319_new_n1329_));
AND2X2 AND2X2_392 ( .A(_abc_40319_new_n1329_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1330_));
AND2X2 AND2X2_393 ( .A(_abc_40319_new_n1331_), .B(_abc_40319_new_n1332_), .Y(_abc_40319_new_n1333_));
AND2X2 AND2X2_394 ( .A(_abc_40319_new_n1333_), .B(_abc_40319_new_n738_), .Y(_abc_40319_new_n1334_));
AND2X2 AND2X2_395 ( .A(_abc_40319_new_n736_), .B(REG0_REG_22_), .Y(_abc_40319_new_n1335_));
AND2X2 AND2X2_396 ( .A(_abc_40319_new_n722_), .B(REG1_REG_22_), .Y(_abc_40319_new_n1336_));
AND2X2 AND2X2_397 ( .A(_abc_40319_new_n733_), .B(REG2_REG_22_), .Y(_abc_40319_new_n1337_));
AND2X2 AND2X2_398 ( .A(_abc_40319_new_n1340_), .B(_abc_40319_new_n705_), .Y(_abc_40319_new_n1341_));
AND2X2 AND2X2_399 ( .A(_abc_40319_new_n763_), .B(_abc_40319_new_n1329_), .Y(_abc_40319_new_n1343_));
AND2X2 AND2X2_4 ( .A(_abc_40319_new_n535_), .B(_abc_40319_new_n532_), .Y(_abc_40319_new_n536_));
AND2X2 AND2X2_40 ( .A(_abc_40319_new_n609_), .B(IR_REG_23_), .Y(_abc_40319_new_n610_));
AND2X2 AND2X2_400 ( .A(_abc_40319_new_n1340_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1344_));
AND2X2 AND2X2_401 ( .A(_abc_40319_new_n1346_), .B(_abc_40319_new_n768_), .Y(_abc_40319_new_n1347_));
AND2X2 AND2X2_402 ( .A(_abc_40319_new_n1345_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1348_));
AND2X2 AND2X2_403 ( .A(_abc_40319_new_n1350_), .B(_abc_40319_new_n1342_), .Y(_abc_40319_new_n1351_));
AND2X2 AND2X2_404 ( .A(_abc_40319_new_n602_), .B(IR_REG_18_), .Y(_abc_40319_new_n1353_));
AND2X2 AND2X2_405 ( .A(_abc_40319_new_n1355_), .B(IR_REG_31_), .Y(_abc_40319_new_n1356_));
AND2X2 AND2X2_406 ( .A(_abc_40319_new_n524_), .B(IR_REG_18_), .Y(_abc_40319_new_n1357_));
AND2X2 AND2X2_407 ( .A(_abc_40319_new_n640_), .B(_abc_40319_new_n1359_), .Y(_abc_40319_new_n1360_));
AND2X2 AND2X2_408 ( .A(_abc_40319_new_n1361_), .B(_abc_40319_new_n1362_), .Y(_abc_40319_new_n1363_));
AND2X2 AND2X2_409 ( .A(_abc_40319_new_n1363_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1364_));
AND2X2 AND2X2_41 ( .A(_abc_40319_new_n612_), .B(_abc_40319_new_n600_), .Y(_abc_40319_new_n613_));
AND2X2 AND2X2_410 ( .A(_abc_40319_new_n722_), .B(REG1_REG_18_), .Y(_abc_40319_new_n1365_));
AND2X2 AND2X2_411 ( .A(_abc_40319_new_n1366_), .B(_abc_40319_new_n1367_), .Y(_abc_40319_new_n1368_));
AND2X2 AND2X2_412 ( .A(_abc_40319_new_n738_), .B(_abc_40319_new_n1368_), .Y(_abc_40319_new_n1369_));
AND2X2 AND2X2_413 ( .A(_abc_40319_new_n733_), .B(REG2_REG_18_), .Y(_abc_40319_new_n1370_));
AND2X2 AND2X2_414 ( .A(_abc_40319_new_n736_), .B(REG0_REG_18_), .Y(_abc_40319_new_n1371_));
AND2X2 AND2X2_415 ( .A(_abc_40319_new_n1374_), .B(_abc_40319_new_n705_), .Y(_abc_40319_new_n1375_));
AND2X2 AND2X2_416 ( .A(_abc_40319_new_n1363_), .B(_abc_40319_new_n763_), .Y(_abc_40319_new_n1377_));
AND2X2 AND2X2_417 ( .A(_abc_40319_new_n1374_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1378_));
AND2X2 AND2X2_418 ( .A(_abc_40319_new_n1380_), .B(_abc_40319_new_n768_), .Y(_abc_40319_new_n1381_));
AND2X2 AND2X2_419 ( .A(_abc_40319_new_n1379_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1382_));
AND2X2 AND2X2_42 ( .A(_abc_40319_new_n598_), .B(_abc_40319_new_n613_), .Y(_abc_40319_new_n614_));
AND2X2 AND2X2_420 ( .A(_abc_40319_new_n1384_), .B(_abc_40319_new_n1376_), .Y(_abc_40319_new_n1385_));
AND2X2 AND2X2_421 ( .A(_abc_40319_new_n524_), .B(_abc_40319_new_n556_), .Y(_abc_40319_new_n1387_));
AND2X2 AND2X2_422 ( .A(_abc_40319_new_n553_), .B(_abc_40319_new_n560_), .Y(_abc_40319_new_n1388_));
AND2X2 AND2X2_423 ( .A(_abc_40319_new_n553_), .B(_abc_40319_new_n559_), .Y(_abc_40319_new_n1389_));
AND2X2 AND2X2_424 ( .A(_abc_40319_new_n1390_), .B(IR_REG_16_), .Y(_abc_40319_new_n1391_));
AND2X2 AND2X2_425 ( .A(_abc_40319_new_n1392_), .B(IR_REG_31_), .Y(_abc_40319_new_n1393_));
AND2X2 AND2X2_426 ( .A(_abc_40319_new_n640_), .B(_abc_40319_new_n1394_), .Y(_abc_40319_new_n1395_));
AND2X2 AND2X2_427 ( .A(_abc_40319_new_n1396_), .B(_abc_40319_new_n1397_), .Y(_abc_40319_new_n1398_));
AND2X2 AND2X2_428 ( .A(_abc_40319_new_n1398_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1399_));
AND2X2 AND2X2_429 ( .A(_abc_40319_new_n736_), .B(REG0_REG_16_), .Y(_abc_40319_new_n1400_));
AND2X2 AND2X2_43 ( .A(_abc_40319_new_n614_), .B(STATE_REG), .Y(_abc_40319_new_n615_));
AND2X2 AND2X2_430 ( .A(_abc_40319_new_n733_), .B(REG2_REG_16_), .Y(_abc_40319_new_n1401_));
AND2X2 AND2X2_431 ( .A(_abc_40319_new_n1188_), .B(REG3_REG_16_), .Y(_abc_40319_new_n1404_));
AND2X2 AND2X2_432 ( .A(_abc_40319_new_n1405_), .B(_abc_40319_new_n1403_), .Y(_abc_40319_new_n1406_));
AND2X2 AND2X2_433 ( .A(_abc_40319_new_n738_), .B(_abc_40319_new_n1406_), .Y(_abc_40319_new_n1407_));
AND2X2 AND2X2_434 ( .A(_abc_40319_new_n722_), .B(REG1_REG_16_), .Y(_abc_40319_new_n1408_));
AND2X2 AND2X2_435 ( .A(_abc_40319_new_n705_), .B(_abc_40319_new_n1410_), .Y(_abc_40319_new_n1411_));
AND2X2 AND2X2_436 ( .A(_abc_40319_new_n1398_), .B(_abc_40319_new_n763_), .Y(_abc_40319_new_n1414_));
AND2X2 AND2X2_437 ( .A(_abc_40319_new_n1410_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1415_));
AND2X2 AND2X2_438 ( .A(_abc_40319_new_n1419_), .B(_abc_40319_new_n1417_), .Y(_abc_40319_new_n1420_));
AND2X2 AND2X2_439 ( .A(_abc_40319_new_n1421_), .B(_abc_40319_new_n1413_), .Y(_abc_40319_new_n1422_));
AND2X2 AND2X2_44 ( .A(_abc_40319_new_n615_), .B(_abc_40319_new_n523_), .Y(n1345));
AND2X2 AND2X2_440 ( .A(_abc_40319_new_n1424_), .B(_abc_40319_new_n602_), .Y(_abc_40319_new_n1425_));
AND2X2 AND2X2_441 ( .A(_abc_40319_new_n1425_), .B(IR_REG_31_), .Y(_abc_40319_new_n1426_));
AND2X2 AND2X2_442 ( .A(_abc_40319_new_n524_), .B(IR_REG_17_), .Y(_abc_40319_new_n1427_));
AND2X2 AND2X2_443 ( .A(_abc_40319_new_n640_), .B(_abc_40319_new_n1429_), .Y(_abc_40319_new_n1430_));
AND2X2 AND2X2_444 ( .A(_abc_40319_new_n1431_), .B(_abc_40319_new_n1432_), .Y(_abc_40319_new_n1433_));
AND2X2 AND2X2_445 ( .A(_abc_40319_new_n1433_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1434_));
AND2X2 AND2X2_446 ( .A(_abc_40319_new_n736_), .B(REG0_REG_17_), .Y(_abc_40319_new_n1435_));
AND2X2 AND2X2_447 ( .A(_abc_40319_new_n722_), .B(REG1_REG_17_), .Y(_abc_40319_new_n1436_));
AND2X2 AND2X2_448 ( .A(_abc_40319_new_n1439_), .B(_abc_40319_new_n1438_), .Y(_abc_40319_new_n1440_));
AND2X2 AND2X2_449 ( .A(_abc_40319_new_n738_), .B(_abc_40319_new_n1440_), .Y(_abc_40319_new_n1441_));
AND2X2 AND2X2_45 ( .A(_abc_40319_new_n617_), .B(_abc_40319_new_n523_), .Y(n1336));
AND2X2 AND2X2_450 ( .A(_abc_40319_new_n733_), .B(REG2_REG_17_), .Y(_abc_40319_new_n1442_));
AND2X2 AND2X2_451 ( .A(_abc_40319_new_n705_), .B(_abc_40319_new_n1444_), .Y(_abc_40319_new_n1445_));
AND2X2 AND2X2_452 ( .A(_abc_40319_new_n1433_), .B(_abc_40319_new_n763_), .Y(_abc_40319_new_n1448_));
AND2X2 AND2X2_453 ( .A(_abc_40319_new_n1444_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1449_));
AND2X2 AND2X2_454 ( .A(_abc_40319_new_n1453_), .B(_abc_40319_new_n1451_), .Y(_abc_40319_new_n1454_));
AND2X2 AND2X2_455 ( .A(_abc_40319_new_n1455_), .B(_abc_40319_new_n1447_), .Y(_abc_40319_new_n1456_));
AND2X2 AND2X2_456 ( .A(_abc_40319_new_n1423_), .B(_abc_40319_new_n1457_), .Y(_abc_40319_new_n1458_));
AND2X2 AND2X2_457 ( .A(_abc_40319_new_n553_), .B(_abc_40319_new_n558_), .Y(_abc_40319_new_n1459_));
AND2X2 AND2X2_458 ( .A(_abc_40319_new_n1460_), .B(IR_REG_15_), .Y(_abc_40319_new_n1461_));
AND2X2 AND2X2_459 ( .A(_abc_40319_new_n1463_), .B(IR_REG_31_), .Y(_abc_40319_new_n1464_));
AND2X2 AND2X2_46 ( .A(_abc_40319_new_n579_), .B(IR_REG_27_), .Y(_abc_40319_new_n619_));
AND2X2 AND2X2_460 ( .A(_abc_40319_new_n524_), .B(IR_REG_15_), .Y(_abc_40319_new_n1465_));
AND2X2 AND2X2_461 ( .A(_abc_40319_new_n640_), .B(_abc_40319_new_n1467_), .Y(_abc_40319_new_n1468_));
AND2X2 AND2X2_462 ( .A(_abc_40319_new_n1469_), .B(_abc_40319_new_n1470_), .Y(_abc_40319_new_n1471_));
AND2X2 AND2X2_463 ( .A(_abc_40319_new_n1471_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1472_));
AND2X2 AND2X2_464 ( .A(_abc_40319_new_n722_), .B(REG1_REG_15_), .Y(_abc_40319_new_n1473_));
AND2X2 AND2X2_465 ( .A(_abc_40319_new_n733_), .B(REG2_REG_15_), .Y(_abc_40319_new_n1474_));
AND2X2 AND2X2_466 ( .A(_abc_40319_new_n736_), .B(REG0_REG_15_), .Y(_abc_40319_new_n1476_));
AND2X2 AND2X2_467 ( .A(_abc_40319_new_n1186_), .B(REG3_REG_14_), .Y(_abc_40319_new_n1478_));
AND2X2 AND2X2_468 ( .A(_abc_40319_new_n1479_), .B(_abc_40319_new_n1477_), .Y(_abc_40319_new_n1480_));
AND2X2 AND2X2_469 ( .A(_abc_40319_new_n738_), .B(_abc_40319_new_n1480_), .Y(_abc_40319_new_n1481_));
AND2X2 AND2X2_47 ( .A(_abc_40319_new_n575_), .B(_abc_40319_new_n525_), .Y(_abc_40319_new_n621_));
AND2X2 AND2X2_470 ( .A(_abc_40319_new_n705_), .B(_abc_40319_new_n1483_), .Y(_abc_40319_new_n1484_));
AND2X2 AND2X2_471 ( .A(_abc_40319_new_n1471_), .B(_abc_40319_new_n763_), .Y(_abc_40319_new_n1486_));
AND2X2 AND2X2_472 ( .A(_abc_40319_new_n1483_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1487_));
AND2X2 AND2X2_473 ( .A(_abc_40319_new_n1491_), .B(_abc_40319_new_n1489_), .Y(_abc_40319_new_n1492_));
AND2X2 AND2X2_474 ( .A(_abc_40319_new_n1492_), .B(_abc_40319_new_n1485_), .Y(_abc_40319_new_n1493_));
AND2X2 AND2X2_475 ( .A(_abc_40319_new_n1495_), .B(IR_REG_14_), .Y(_abc_40319_new_n1496_));
AND2X2 AND2X2_476 ( .A(_abc_40319_new_n1498_), .B(IR_REG_31_), .Y(_abc_40319_new_n1499_));
AND2X2 AND2X2_477 ( .A(_abc_40319_new_n524_), .B(IR_REG_14_), .Y(_abc_40319_new_n1500_));
AND2X2 AND2X2_478 ( .A(_abc_40319_new_n640_), .B(_abc_40319_new_n1502_), .Y(_abc_40319_new_n1503_));
AND2X2 AND2X2_479 ( .A(_abc_40319_new_n1504_), .B(_abc_40319_new_n1505_), .Y(_abc_40319_new_n1506_));
AND2X2 AND2X2_48 ( .A(_abc_40319_new_n621_), .B(_abc_40319_new_n620_), .Y(_abc_40319_new_n622_));
AND2X2 AND2X2_480 ( .A(_abc_40319_new_n1506_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1507_));
AND2X2 AND2X2_481 ( .A(_abc_40319_new_n736_), .B(REG0_REG_14_), .Y(_abc_40319_new_n1508_));
AND2X2 AND2X2_482 ( .A(_abc_40319_new_n733_), .B(REG2_REG_14_), .Y(_abc_40319_new_n1509_));
AND2X2 AND2X2_483 ( .A(_abc_40319_new_n1511_), .B(_abc_40319_new_n1512_), .Y(_abc_40319_new_n1513_));
AND2X2 AND2X2_484 ( .A(_abc_40319_new_n738_), .B(_abc_40319_new_n1513_), .Y(_abc_40319_new_n1514_));
AND2X2 AND2X2_485 ( .A(_abc_40319_new_n722_), .B(REG1_REG_14_), .Y(_abc_40319_new_n1515_));
AND2X2 AND2X2_486 ( .A(_abc_40319_new_n705_), .B(_abc_40319_new_n1517_), .Y(_abc_40319_new_n1518_));
AND2X2 AND2X2_487 ( .A(_abc_40319_new_n1506_), .B(_abc_40319_new_n763_), .Y(_abc_40319_new_n1520_));
AND2X2 AND2X2_488 ( .A(_abc_40319_new_n1517_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1521_));
AND2X2 AND2X2_489 ( .A(_abc_40319_new_n1525_), .B(_abc_40319_new_n1523_), .Y(_abc_40319_new_n1526_));
AND2X2 AND2X2_49 ( .A(_abc_40319_new_n572_), .B(_abc_40319_new_n622_), .Y(_abc_40319_new_n623_));
AND2X2 AND2X2_490 ( .A(_abc_40319_new_n1526_), .B(_abc_40319_new_n1519_), .Y(_abc_40319_new_n1527_));
AND2X2 AND2X2_491 ( .A(_abc_40319_new_n1531_), .B(_abc_40319_new_n970_), .Y(_abc_40319_new_n1532_));
AND2X2 AND2X2_492 ( .A(_abc_40319_new_n1533_), .B(_abc_40319_new_n1534_), .Y(_abc_40319_new_n1535_));
AND2X2 AND2X2_493 ( .A(_abc_40319_new_n1538_), .B(_abc_40319_new_n1539_), .Y(_abc_40319_new_n1540_));
AND2X2 AND2X2_494 ( .A(_abc_40319_new_n1540_), .B(_abc_40319_new_n1537_), .Y(_abc_40319_new_n1541_));
AND2X2 AND2X2_495 ( .A(_abc_40319_new_n1544_), .B(_abc_40319_new_n1545_), .Y(_abc_40319_new_n1546_));
AND2X2 AND2X2_496 ( .A(_abc_40319_new_n1543_), .B(_abc_40319_new_n1546_), .Y(_abc_40319_new_n1547_));
AND2X2 AND2X2_497 ( .A(_abc_40319_new_n1547_), .B(_abc_40319_new_n768_), .Y(_abc_40319_new_n1548_));
AND2X2 AND2X2_498 ( .A(_abc_40319_new_n1551_), .B(_abc_40319_new_n1549_), .Y(_abc_40319_new_n1552_));
AND2X2 AND2X2_499 ( .A(_abc_40319_new_n1553_), .B(_abc_40319_new_n1542_), .Y(_abc_40319_new_n1554_));
AND2X2 AND2X2_5 ( .A(_abc_40319_new_n531_), .B(_abc_40319_new_n536_), .Y(_abc_40319_new_n537_));
AND2X2 AND2X2_50 ( .A(_abc_40319_new_n625_), .B(IR_REG_31_), .Y(_abc_40319_new_n626_));
AND2X2 AND2X2_500 ( .A(_abc_40319_new_n1555_), .B(_abc_40319_new_n1536_), .Y(_abc_40319_new_n1556_));
AND2X2 AND2X2_501 ( .A(_abc_40319_new_n1557_), .B(_abc_40319_new_n1535_), .Y(_abc_40319_new_n1558_));
AND2X2 AND2X2_502 ( .A(_abc_40319_new_n1559_), .B(_abc_40319_new_n1529_), .Y(_abc_40319_new_n1560_));
AND2X2 AND2X2_503 ( .A(_abc_40319_new_n1023_), .B(_abc_40319_new_n546_), .Y(_abc_40319_new_n1561_));
AND2X2 AND2X2_504 ( .A(_abc_40319_new_n1024_), .B(IR_REG_8_), .Y(_abc_40319_new_n1562_));
AND2X2 AND2X2_505 ( .A(_abc_40319_new_n1564_), .B(IR_REG_31_), .Y(_abc_40319_new_n1565_));
AND2X2 AND2X2_506 ( .A(_abc_40319_new_n524_), .B(IR_REG_8_), .Y(_abc_40319_new_n1566_));
AND2X2 AND2X2_507 ( .A(_abc_40319_new_n640_), .B(_abc_40319_new_n1568_), .Y(_abc_40319_new_n1569_));
AND2X2 AND2X2_508 ( .A(_abc_40319_new_n1570_), .B(_abc_40319_new_n1571_), .Y(_abc_40319_new_n1572_));
AND2X2 AND2X2_509 ( .A(_abc_40319_new_n1572_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1573_));
AND2X2 AND2X2_51 ( .A(_abc_40319_new_n524_), .B(IR_REG_27_), .Y(_abc_40319_new_n627_));
AND2X2 AND2X2_510 ( .A(_abc_40319_new_n705_), .B(_abc_40319_new_n1146_), .Y(_abc_40319_new_n1574_));
AND2X2 AND2X2_511 ( .A(_abc_40319_new_n1572_), .B(_abc_40319_new_n763_), .Y(_abc_40319_new_n1577_));
AND2X2 AND2X2_512 ( .A(_abc_40319_new_n1146_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1578_));
AND2X2 AND2X2_513 ( .A(_abc_40319_new_n1582_), .B(_abc_40319_new_n1580_), .Y(_abc_40319_new_n1583_));
AND2X2 AND2X2_514 ( .A(_abc_40319_new_n1584_), .B(_abc_40319_new_n1576_), .Y(_abc_40319_new_n1585_));
AND2X2 AND2X2_515 ( .A(_abc_40319_new_n1587_), .B(_abc_40319_new_n773_), .Y(_abc_40319_new_n1588_));
AND2X2 AND2X2_516 ( .A(_abc_40319_new_n1588_), .B(_abc_40319_new_n1586_), .Y(_abc_40319_new_n1589_));
AND2X2 AND2X2_517 ( .A(_abc_40319_new_n1583_), .B(_abc_40319_new_n1575_), .Y(_abc_40319_new_n1592_));
AND2X2 AND2X2_518 ( .A(_abc_40319_new_n1021_), .B(_abc_40319_new_n1057_), .Y(_abc_40319_new_n1596_));
AND2X2 AND2X2_519 ( .A(_abc_40319_new_n1595_), .B(_abc_40319_new_n1597_), .Y(_abc_40319_new_n1598_));
AND2X2 AND2X2_52 ( .A(_abc_40319_new_n524_), .B(_abc_40319_new_n630_), .Y(_abc_40319_new_n631_));
AND2X2 AND2X2_520 ( .A(_abc_40319_new_n1598_), .B(_abc_40319_new_n1593_), .Y(_abc_40319_new_n1599_));
AND2X2 AND2X2_521 ( .A(_abc_40319_new_n1591_), .B(_abc_40319_new_n1600_), .Y(_abc_40319_new_n1601_));
AND2X2 AND2X2_522 ( .A(_abc_40319_new_n524_), .B(_abc_40319_new_n545_), .Y(_abc_40319_new_n1602_));
AND2X2 AND2X2_523 ( .A(_abc_40319_new_n537_), .B(_abc_40319_new_n551_), .Y(_abc_40319_new_n1604_));
AND2X2 AND2X2_524 ( .A(_abc_40319_new_n1606_), .B(_abc_40319_new_n1605_), .Y(_abc_40319_new_n1607_));
AND2X2 AND2X2_525 ( .A(_abc_40319_new_n1608_), .B(_abc_40319_new_n1603_), .Y(_abc_40319_new_n1609_));
AND2X2 AND2X2_526 ( .A(_abc_40319_new_n640_), .B(_abc_40319_new_n1610_), .Y(_abc_40319_new_n1611_));
AND2X2 AND2X2_527 ( .A(_abc_40319_new_n1612_), .B(_abc_40319_new_n1613_), .Y(_abc_40319_new_n1614_));
AND2X2 AND2X2_528 ( .A(_abc_40319_new_n1614_), .B(_abc_40319_new_n763_), .Y(_abc_40319_new_n1615_));
AND2X2 AND2X2_529 ( .A(_abc_40319_new_n1616_), .B(_abc_40319_new_n1617_), .Y(_abc_40319_new_n1618_));
AND2X2 AND2X2_53 ( .A(_abc_40319_new_n623_), .B(_abc_40319_new_n630_), .Y(_abc_40319_new_n633_));
AND2X2 AND2X2_530 ( .A(_abc_40319_new_n738_), .B(_abc_40319_new_n1618_), .Y(_abc_40319_new_n1619_));
AND2X2 AND2X2_531 ( .A(_abc_40319_new_n722_), .B(REG1_REG_9_), .Y(_abc_40319_new_n1620_));
AND2X2 AND2X2_532 ( .A(_abc_40319_new_n736_), .B(REG0_REG_9_), .Y(_abc_40319_new_n1622_));
AND2X2 AND2X2_533 ( .A(_abc_40319_new_n733_), .B(REG2_REG_9_), .Y(_abc_40319_new_n1623_));
AND2X2 AND2X2_534 ( .A(_abc_40319_new_n1625_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1626_));
AND2X2 AND2X2_535 ( .A(_abc_40319_new_n1630_), .B(_abc_40319_new_n1628_), .Y(_abc_40319_new_n1631_));
AND2X2 AND2X2_536 ( .A(_abc_40319_new_n1601_), .B(_abc_40319_new_n1632_), .Y(_abc_40319_new_n1633_));
AND2X2 AND2X2_537 ( .A(_abc_40319_new_n982_), .B(_abc_40319_new_n1589_), .Y(_abc_40319_new_n1635_));
AND2X2 AND2X2_538 ( .A(_abc_40319_new_n1637_), .B(_abc_40319_new_n1631_), .Y(_abc_40319_new_n1638_));
AND2X2 AND2X2_539 ( .A(_abc_40319_new_n1614_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1639_));
AND2X2 AND2X2_54 ( .A(_abc_40319_new_n634_), .B(_abc_40319_new_n635_), .Y(_abc_40319_new_n636_));
AND2X2 AND2X2_540 ( .A(_abc_40319_new_n705_), .B(_abc_40319_new_n1625_), .Y(_abc_40319_new_n1640_));
AND2X2 AND2X2_541 ( .A(_abc_40319_new_n1642_), .B(_abc_40319_new_n1634_), .Y(_abc_40319_new_n1643_));
AND2X2 AND2X2_542 ( .A(_abc_40319_new_n524_), .B(_abc_40319_new_n541_), .Y(_abc_40319_new_n1644_));
AND2X2 AND2X2_543 ( .A(_abc_40319_new_n1604_), .B(_abc_40319_new_n542_), .Y(_abc_40319_new_n1645_));
AND2X2 AND2X2_544 ( .A(_abc_40319_new_n1645_), .B(_abc_40319_new_n540_), .Y(_abc_40319_new_n1646_));
AND2X2 AND2X2_545 ( .A(_abc_40319_new_n1647_), .B(IR_REG_13_), .Y(_abc_40319_new_n1648_));
AND2X2 AND2X2_546 ( .A(_abc_40319_new_n1649_), .B(IR_REG_31_), .Y(_abc_40319_new_n1650_));
AND2X2 AND2X2_547 ( .A(_abc_40319_new_n640_), .B(_abc_40319_new_n1651_), .Y(_abc_40319_new_n1652_));
AND2X2 AND2X2_548 ( .A(_abc_40319_new_n1653_), .B(_abc_40319_new_n1654_), .Y(_abc_40319_new_n1655_));
AND2X2 AND2X2_549 ( .A(_abc_40319_new_n1655_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1656_));
AND2X2 AND2X2_55 ( .A(_abc_40319_new_n637_), .B(_abc_40319_new_n632_), .Y(_abc_40319_new_n638_));
AND2X2 AND2X2_550 ( .A(_abc_40319_new_n1184_), .B(REG3_REG_12_), .Y(_abc_40319_new_n1658_));
AND2X2 AND2X2_551 ( .A(_abc_40319_new_n1659_), .B(_abc_40319_new_n1657_), .Y(_abc_40319_new_n1660_));
AND2X2 AND2X2_552 ( .A(_abc_40319_new_n738_), .B(_abc_40319_new_n1660_), .Y(_abc_40319_new_n1661_));
AND2X2 AND2X2_553 ( .A(_abc_40319_new_n722_), .B(REG1_REG_13_), .Y(_abc_40319_new_n1662_));
AND2X2 AND2X2_554 ( .A(_abc_40319_new_n736_), .B(REG0_REG_13_), .Y(_abc_40319_new_n1664_));
AND2X2 AND2X2_555 ( .A(_abc_40319_new_n733_), .B(REG2_REG_13_), .Y(_abc_40319_new_n1665_));
AND2X2 AND2X2_556 ( .A(_abc_40319_new_n705_), .B(_abc_40319_new_n1667_), .Y(_abc_40319_new_n1668_));
AND2X2 AND2X2_557 ( .A(_abc_40319_new_n1655_), .B(_abc_40319_new_n763_), .Y(_abc_40319_new_n1671_));
AND2X2 AND2X2_558 ( .A(_abc_40319_new_n1667_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1672_));
AND2X2 AND2X2_559 ( .A(_abc_40319_new_n1676_), .B(_abc_40319_new_n1674_), .Y(_abc_40319_new_n1677_));
AND2X2 AND2X2_56 ( .A(_abc_40319_new_n629_), .B(_abc_40319_new_n639_), .Y(_abc_40319_new_n640_));
AND2X2 AND2X2_560 ( .A(_abc_40319_new_n1677_), .B(_abc_40319_new_n1670_), .Y(_abc_40319_new_n1678_));
AND2X2 AND2X2_561 ( .A(_abc_40319_new_n524_), .B(_abc_40319_new_n538_), .Y(_abc_40319_new_n1680_));
AND2X2 AND2X2_562 ( .A(_abc_40319_new_n1645_), .B(_abc_40319_new_n539_), .Y(_abc_40319_new_n1681_));
AND2X2 AND2X2_563 ( .A(_abc_40319_new_n1682_), .B(IR_REG_12_), .Y(_abc_40319_new_n1683_));
AND2X2 AND2X2_564 ( .A(_abc_40319_new_n1684_), .B(IR_REG_31_), .Y(_abc_40319_new_n1685_));
AND2X2 AND2X2_565 ( .A(_abc_40319_new_n640_), .B(_abc_40319_new_n1686_), .Y(_abc_40319_new_n1687_));
AND2X2 AND2X2_566 ( .A(_abc_40319_new_n1688_), .B(_abc_40319_new_n1689_), .Y(_abc_40319_new_n1690_));
AND2X2 AND2X2_567 ( .A(_abc_40319_new_n1690_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1691_));
AND2X2 AND2X2_568 ( .A(_abc_40319_new_n722_), .B(REG1_REG_12_), .Y(_abc_40319_new_n1692_));
AND2X2 AND2X2_569 ( .A(_abc_40319_new_n733_), .B(REG2_REG_12_), .Y(_abc_40319_new_n1693_));
AND2X2 AND2X2_57 ( .A(_abc_40319_new_n524_), .B(_abc_40319_new_n554_), .Y(_abc_40319_new_n641_));
AND2X2 AND2X2_570 ( .A(_abc_40319_new_n736_), .B(REG0_REG_12_), .Y(_abc_40319_new_n1695_));
AND2X2 AND2X2_571 ( .A(_abc_40319_new_n1696_), .B(_abc_40319_new_n1697_), .Y(_abc_40319_new_n1698_));
AND2X2 AND2X2_572 ( .A(_abc_40319_new_n738_), .B(_abc_40319_new_n1698_), .Y(_abc_40319_new_n1699_));
AND2X2 AND2X2_573 ( .A(_abc_40319_new_n705_), .B(_abc_40319_new_n1701_), .Y(_abc_40319_new_n1702_));
AND2X2 AND2X2_574 ( .A(_abc_40319_new_n1690_), .B(_abc_40319_new_n763_), .Y(_abc_40319_new_n1705_));
AND2X2 AND2X2_575 ( .A(_abc_40319_new_n1701_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1706_));
AND2X2 AND2X2_576 ( .A(_abc_40319_new_n1710_), .B(_abc_40319_new_n1708_), .Y(_abc_40319_new_n1711_));
AND2X2 AND2X2_577 ( .A(_abc_40319_new_n1711_), .B(_abc_40319_new_n1704_), .Y(_abc_40319_new_n1712_));
AND2X2 AND2X2_578 ( .A(_abc_40319_new_n1679_), .B(_abc_40319_new_n1713_), .Y(_abc_40319_new_n1714_));
AND2X2 AND2X2_579 ( .A(_abc_40319_new_n524_), .B(_abc_40319_new_n539_), .Y(_abc_40319_new_n1715_));
AND2X2 AND2X2_58 ( .A(_abc_40319_new_n606_), .B(IR_REG_22_), .Y(_abc_40319_new_n642_));
AND2X2 AND2X2_580 ( .A(_abc_40319_new_n1716_), .B(IR_REG_11_), .Y(_abc_40319_new_n1717_));
AND2X2 AND2X2_581 ( .A(_abc_40319_new_n1718_), .B(IR_REG_31_), .Y(_abc_40319_new_n1719_));
AND2X2 AND2X2_582 ( .A(_abc_40319_new_n640_), .B(_abc_40319_new_n1720_), .Y(_abc_40319_new_n1721_));
AND2X2 AND2X2_583 ( .A(_abc_40319_new_n1722_), .B(_abc_40319_new_n1723_), .Y(_abc_40319_new_n1724_));
AND2X2 AND2X2_584 ( .A(_abc_40319_new_n1724_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1725_));
AND2X2 AND2X2_585 ( .A(_abc_40319_new_n722_), .B(REG1_REG_11_), .Y(_abc_40319_new_n1726_));
AND2X2 AND2X2_586 ( .A(_abc_40319_new_n733_), .B(REG2_REG_11_), .Y(_abc_40319_new_n1727_));
AND2X2 AND2X2_587 ( .A(_abc_40319_new_n736_), .B(REG0_REG_11_), .Y(_abc_40319_new_n1729_));
AND2X2 AND2X2_588 ( .A(_abc_40319_new_n1730_), .B(_abc_40319_new_n1731_), .Y(_abc_40319_new_n1732_));
AND2X2 AND2X2_589 ( .A(_abc_40319_new_n738_), .B(_abc_40319_new_n1732_), .Y(_abc_40319_new_n1733_));
AND2X2 AND2X2_59 ( .A(_abc_40319_new_n643_), .B(IR_REG_31_), .Y(_abc_40319_new_n644_));
AND2X2 AND2X2_590 ( .A(_abc_40319_new_n705_), .B(_abc_40319_new_n1735_), .Y(_abc_40319_new_n1736_));
AND2X2 AND2X2_591 ( .A(_abc_40319_new_n1724_), .B(_abc_40319_new_n763_), .Y(_abc_40319_new_n1739_));
AND2X2 AND2X2_592 ( .A(_abc_40319_new_n1735_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1740_));
AND2X2 AND2X2_593 ( .A(_abc_40319_new_n1744_), .B(_abc_40319_new_n1742_), .Y(_abc_40319_new_n1745_));
AND2X2 AND2X2_594 ( .A(_abc_40319_new_n1746_), .B(_abc_40319_new_n1738_), .Y(_abc_40319_new_n1747_));
AND2X2 AND2X2_595 ( .A(_abc_40319_new_n1714_), .B(_abc_40319_new_n1748_), .Y(_abc_40319_new_n1749_));
AND2X2 AND2X2_596 ( .A(_abc_40319_new_n524_), .B(_abc_40319_new_n542_), .Y(_abc_40319_new_n1750_));
AND2X2 AND2X2_597 ( .A(_abc_40319_new_n1605_), .B(IR_REG_10_), .Y(_abc_40319_new_n1751_));
AND2X2 AND2X2_598 ( .A(_abc_40319_new_n1752_), .B(IR_REG_31_), .Y(_abc_40319_new_n1753_));
AND2X2 AND2X2_599 ( .A(_abc_40319_new_n640_), .B(_abc_40319_new_n1754_), .Y(_abc_40319_new_n1755_));
AND2X2 AND2X2_6 ( .A(_abc_40319_new_n538_), .B(_abc_40319_new_n539_), .Y(_abc_40319_new_n540_));
AND2X2 AND2X2_60 ( .A(_abc_40319_new_n601_), .B(_abc_40319_new_n647_), .Y(_abc_40319_new_n648_));
AND2X2 AND2X2_600 ( .A(_abc_40319_new_n1756_), .B(_abc_40319_new_n1757_), .Y(_abc_40319_new_n1758_));
AND2X2 AND2X2_601 ( .A(_abc_40319_new_n1758_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1759_));
AND2X2 AND2X2_602 ( .A(_abc_40319_new_n722_), .B(REG1_REG_10_), .Y(_abc_40319_new_n1760_));
AND2X2 AND2X2_603 ( .A(_abc_40319_new_n733_), .B(REG2_REG_10_), .Y(_abc_40319_new_n1761_));
AND2X2 AND2X2_604 ( .A(_abc_40319_new_n736_), .B(REG0_REG_10_), .Y(_abc_40319_new_n1763_));
AND2X2 AND2X2_605 ( .A(_abc_40319_new_n1764_), .B(_abc_40319_new_n1765_), .Y(_abc_40319_new_n1766_));
AND2X2 AND2X2_606 ( .A(_abc_40319_new_n738_), .B(_abc_40319_new_n1766_), .Y(_abc_40319_new_n1767_));
AND2X2 AND2X2_607 ( .A(_abc_40319_new_n705_), .B(_abc_40319_new_n1769_), .Y(_abc_40319_new_n1770_));
AND2X2 AND2X2_608 ( .A(_abc_40319_new_n1758_), .B(_abc_40319_new_n763_), .Y(_abc_40319_new_n1773_));
AND2X2 AND2X2_609 ( .A(_abc_40319_new_n1769_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1774_));
AND2X2 AND2X2_61 ( .A(_abc_40319_new_n648_), .B(_abc_40319_new_n562_), .Y(_abc_40319_new_n649_));
AND2X2 AND2X2_610 ( .A(_abc_40319_new_n1778_), .B(_abc_40319_new_n1776_), .Y(_abc_40319_new_n1779_));
AND2X2 AND2X2_611 ( .A(_abc_40319_new_n1780_), .B(_abc_40319_new_n1772_), .Y(_abc_40319_new_n1781_));
AND2X2 AND2X2_612 ( .A(_abc_40319_new_n1749_), .B(_abc_40319_new_n1782_), .Y(_abc_40319_new_n1783_));
AND2X2 AND2X2_613 ( .A(_abc_40319_new_n1643_), .B(_abc_40319_new_n1783_), .Y(_abc_40319_new_n1784_));
AND2X2 AND2X2_614 ( .A(_abc_40319_new_n1779_), .B(_abc_40319_new_n1771_), .Y(_abc_40319_new_n1785_));
AND2X2 AND2X2_615 ( .A(_abc_40319_new_n1749_), .B(_abc_40319_new_n1785_), .Y(_abc_40319_new_n1786_));
AND2X2 AND2X2_616 ( .A(_abc_40319_new_n1745_), .B(_abc_40319_new_n1737_), .Y(_abc_40319_new_n1788_));
AND2X2 AND2X2_617 ( .A(_abc_40319_new_n1714_), .B(_abc_40319_new_n1788_), .Y(_abc_40319_new_n1789_));
AND2X2 AND2X2_618 ( .A(_abc_40319_new_n1791_), .B(_abc_40319_new_n1792_), .Y(_abc_40319_new_n1793_));
AND2X2 AND2X2_619 ( .A(_abc_40319_new_n1790_), .B(_abc_40319_new_n1793_), .Y(_abc_40319_new_n1794_));
AND2X2 AND2X2_62 ( .A(_abc_40319_new_n649_), .B(_abc_40319_new_n563_), .Y(_abc_40319_new_n650_));
AND2X2 AND2X2_620 ( .A(_abc_40319_new_n1795_), .B(_abc_40319_new_n1787_), .Y(_abc_40319_new_n1796_));
AND2X2 AND2X2_621 ( .A(_abc_40319_new_n1798_), .B(_abc_40319_new_n1528_), .Y(_abc_40319_new_n1799_));
AND2X2 AND2X2_622 ( .A(_abc_40319_new_n1800_), .B(_abc_40319_new_n1494_), .Y(_abc_40319_new_n1801_));
AND2X2 AND2X2_623 ( .A(_abc_40319_new_n1802_), .B(_abc_40319_new_n1458_), .Y(_abc_40319_new_n1803_));
AND2X2 AND2X2_624 ( .A(_abc_40319_new_n1420_), .B(_abc_40319_new_n1412_), .Y(_abc_40319_new_n1804_));
AND2X2 AND2X2_625 ( .A(_abc_40319_new_n1454_), .B(_abc_40319_new_n1446_), .Y(_abc_40319_new_n1806_));
AND2X2 AND2X2_626 ( .A(_abc_40319_new_n1805_), .B(_abc_40319_new_n1807_), .Y(_abc_40319_new_n1808_));
AND2X2 AND2X2_627 ( .A(_abc_40319_new_n1811_), .B(_abc_40319_new_n1386_), .Y(_abc_40319_new_n1812_));
AND2X2 AND2X2_628 ( .A(_abc_40319_new_n640_), .B(_abc_40319_new_n698_), .Y(_abc_40319_new_n1814_));
AND2X2 AND2X2_629 ( .A(_abc_40319_new_n1815_), .B(_abc_40319_new_n1816_), .Y(_abc_40319_new_n1817_));
AND2X2 AND2X2_63 ( .A(_abc_40319_new_n651_), .B(_abc_40319_new_n606_), .Y(_abc_40319_new_n652_));
AND2X2 AND2X2_630 ( .A(_abc_40319_new_n1817_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1818_));
AND2X2 AND2X2_631 ( .A(_abc_40319_new_n722_), .B(REG1_REG_19_), .Y(_abc_40319_new_n1819_));
AND2X2 AND2X2_632 ( .A(_abc_40319_new_n1820_), .B(_abc_40319_new_n1821_), .Y(_abc_40319_new_n1822_));
AND2X2 AND2X2_633 ( .A(_abc_40319_new_n1822_), .B(_abc_40319_new_n738_), .Y(_abc_40319_new_n1823_));
AND2X2 AND2X2_634 ( .A(_abc_40319_new_n733_), .B(REG2_REG_19_), .Y(_abc_40319_new_n1824_));
AND2X2 AND2X2_635 ( .A(_abc_40319_new_n736_), .B(REG0_REG_19_), .Y(_abc_40319_new_n1825_));
AND2X2 AND2X2_636 ( .A(_abc_40319_new_n1828_), .B(_abc_40319_new_n705_), .Y(_abc_40319_new_n1829_));
AND2X2 AND2X2_637 ( .A(_abc_40319_new_n1817_), .B(_abc_40319_new_n763_), .Y(_abc_40319_new_n1832_));
AND2X2 AND2X2_638 ( .A(_abc_40319_new_n1828_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1833_));
AND2X2 AND2X2_639 ( .A(_abc_40319_new_n1835_), .B(_abc_40319_new_n768_), .Y(_abc_40319_new_n1836_));
AND2X2 AND2X2_64 ( .A(_abc_40319_new_n652_), .B(IR_REG_31_), .Y(_abc_40319_new_n653_));
AND2X2 AND2X2_640 ( .A(_abc_40319_new_n1834_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1837_));
AND2X2 AND2X2_641 ( .A(_abc_40319_new_n1838_), .B(_abc_40319_new_n1831_), .Y(_abc_40319_new_n1839_));
AND2X2 AND2X2_642 ( .A(_abc_40319_new_n817_), .B(DATAI_20_), .Y(_abc_40319_new_n1841_));
AND2X2 AND2X2_643 ( .A(_abc_40319_new_n1841_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1842_));
AND2X2 AND2X2_644 ( .A(_abc_40319_new_n722_), .B(REG1_REG_20_), .Y(_abc_40319_new_n1843_));
AND2X2 AND2X2_645 ( .A(_abc_40319_new_n1844_), .B(_abc_40319_new_n1845_), .Y(_abc_40319_new_n1846_));
AND2X2 AND2X2_646 ( .A(_abc_40319_new_n1846_), .B(_abc_40319_new_n738_), .Y(_abc_40319_new_n1847_));
AND2X2 AND2X2_647 ( .A(_abc_40319_new_n733_), .B(REG2_REG_20_), .Y(_abc_40319_new_n1848_));
AND2X2 AND2X2_648 ( .A(_abc_40319_new_n736_), .B(REG0_REG_20_), .Y(_abc_40319_new_n1849_));
AND2X2 AND2X2_649 ( .A(_abc_40319_new_n1852_), .B(_abc_40319_new_n705_), .Y(_abc_40319_new_n1853_));
AND2X2 AND2X2_65 ( .A(_abc_40319_new_n524_), .B(IR_REG_21_), .Y(_abc_40319_new_n654_));
AND2X2 AND2X2_650 ( .A(_abc_40319_new_n763_), .B(_abc_40319_new_n1841_), .Y(_abc_40319_new_n1856_));
AND2X2 AND2X2_651 ( .A(_abc_40319_new_n1852_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1857_));
AND2X2 AND2X2_652 ( .A(_abc_40319_new_n1859_), .B(_abc_40319_new_n768_), .Y(_abc_40319_new_n1860_));
AND2X2 AND2X2_653 ( .A(_abc_40319_new_n1858_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1861_));
AND2X2 AND2X2_654 ( .A(_abc_40319_new_n1862_), .B(_abc_40319_new_n1855_), .Y(_abc_40319_new_n1863_));
AND2X2 AND2X2_655 ( .A(_abc_40319_new_n817_), .B(DATAI_21_), .Y(_abc_40319_new_n1865_));
AND2X2 AND2X2_656 ( .A(_abc_40319_new_n1865_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1866_));
AND2X2 AND2X2_657 ( .A(_abc_40319_new_n1867_), .B(_abc_40319_new_n1868_), .Y(_abc_40319_new_n1869_));
AND2X2 AND2X2_658 ( .A(_abc_40319_new_n1869_), .B(_abc_40319_new_n738_), .Y(_abc_40319_new_n1870_));
AND2X2 AND2X2_659 ( .A(_abc_40319_new_n736_), .B(REG0_REG_21_), .Y(_abc_40319_new_n1871_));
AND2X2 AND2X2_66 ( .A(_abc_40319_new_n655_), .B(_abc_40319_new_n646_), .Y(_abc_40319_new_n656_));
AND2X2 AND2X2_660 ( .A(_abc_40319_new_n722_), .B(REG1_REG_21_), .Y(_abc_40319_new_n1872_));
AND2X2 AND2X2_661 ( .A(_abc_40319_new_n733_), .B(REG2_REG_21_), .Y(_abc_40319_new_n1873_));
AND2X2 AND2X2_662 ( .A(_abc_40319_new_n1876_), .B(_abc_40319_new_n705_), .Y(_abc_40319_new_n1877_));
AND2X2 AND2X2_663 ( .A(_abc_40319_new_n763_), .B(_abc_40319_new_n1865_), .Y(_abc_40319_new_n1880_));
AND2X2 AND2X2_664 ( .A(_abc_40319_new_n1876_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n1881_));
AND2X2 AND2X2_665 ( .A(_abc_40319_new_n1883_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1884_));
AND2X2 AND2X2_666 ( .A(_abc_40319_new_n1882_), .B(_abc_40319_new_n768_), .Y(_abc_40319_new_n1885_));
AND2X2 AND2X2_667 ( .A(_abc_40319_new_n1887_), .B(_abc_40319_new_n1879_), .Y(_abc_40319_new_n1888_));
AND2X2 AND2X2_668 ( .A(_abc_40319_new_n1889_), .B(_abc_40319_new_n1864_), .Y(_abc_40319_new_n1890_));
AND2X2 AND2X2_669 ( .A(_abc_40319_new_n1890_), .B(_abc_40319_new_n1840_), .Y(_abc_40319_new_n1891_));
AND2X2 AND2X2_67 ( .A(_abc_40319_new_n657_), .B(_abc_40319_new_n613_), .Y(_abc_40319_new_n658_));
AND2X2 AND2X2_670 ( .A(_abc_40319_new_n1813_), .B(_abc_40319_new_n1891_), .Y(_abc_40319_new_n1892_));
AND2X2 AND2X2_671 ( .A(_abc_40319_new_n1890_), .B(_abc_40319_new_n1894_), .Y(_abc_40319_new_n1895_));
AND2X2 AND2X2_672 ( .A(_abc_40319_new_n1886_), .B(_abc_40319_new_n1878_), .Y(_abc_40319_new_n1897_));
AND2X2 AND2X2_673 ( .A(_abc_40319_new_n1898_), .B(_abc_40319_new_n1899_), .Y(_abc_40319_new_n1900_));
AND2X2 AND2X2_674 ( .A(_abc_40319_new_n1896_), .B(_abc_40319_new_n1900_), .Y(_abc_40319_new_n1901_));
AND2X2 AND2X2_675 ( .A(_abc_40319_new_n1904_), .B(_abc_40319_new_n1352_), .Y(_abc_40319_new_n1905_));
AND2X2 AND2X2_676 ( .A(_abc_40319_new_n1906_), .B(_abc_40319_new_n1328_), .Y(_abc_40319_new_n1907_));
AND2X2 AND2X2_677 ( .A(_abc_40319_new_n1273_), .B(_abc_40319_new_n1909_), .Y(_abc_40319_new_n1910_));
AND2X2 AND2X2_678 ( .A(_abc_40319_new_n1908_), .B(_abc_40319_new_n1910_), .Y(_abc_40319_new_n1911_));
AND2X2 AND2X2_679 ( .A(_abc_40319_new_n1928_), .B(_abc_40319_new_n1926_), .Y(_abc_40319_new_n1929_));
AND2X2 AND2X2_68 ( .A(STATE_REG), .B(nRESET_G), .Y(_abc_40319_new_n660_));
AND2X2 AND2X2_680 ( .A(_abc_40319_new_n1931_), .B(_abc_40319_new_n1796_), .Y(_abc_40319_new_n1932_));
AND2X2 AND2X2_681 ( .A(_abc_40319_new_n1933_), .B(_abc_40319_new_n1924_), .Y(_abc_40319_new_n1934_));
AND2X2 AND2X2_682 ( .A(_abc_40319_new_n1935_), .B(_abc_40319_new_n1922_), .Y(_abc_40319_new_n1936_));
AND2X2 AND2X2_683 ( .A(_abc_40319_new_n1937_), .B(_abc_40319_new_n1809_), .Y(_abc_40319_new_n1938_));
AND2X2 AND2X2_684 ( .A(_abc_40319_new_n1939_), .B(_abc_40319_new_n1919_), .Y(_abc_40319_new_n1940_));
AND2X2 AND2X2_685 ( .A(_abc_40319_new_n1942_), .B(_abc_40319_new_n1902_), .Y(_abc_40319_new_n1943_));
AND2X2 AND2X2_686 ( .A(_abc_40319_new_n1944_), .B(_abc_40319_new_n1917_), .Y(_abc_40319_new_n1945_));
AND2X2 AND2X2_687 ( .A(_abc_40319_new_n1946_), .B(_abc_40319_new_n1915_), .Y(_abc_40319_new_n1947_));
AND2X2 AND2X2_688 ( .A(_abc_40319_new_n1949_), .B(_abc_40319_new_n1304_), .Y(_abc_40319_new_n1950_));
AND2X2 AND2X2_689 ( .A(_abc_40319_new_n1951_), .B(_abc_40319_new_n1122_), .Y(_abc_40319_new_n1952_));
AND2X2 AND2X2_69 ( .A(_abc_40319_new_n659_), .B(_abc_40319_new_n660_), .Y(_abc_40319_new_n661_));
AND2X2 AND2X2_690 ( .A(_abc_40319_new_n1952_), .B(_abc_40319_new_n1913_), .Y(_abc_40319_new_n1953_));
AND2X2 AND2X2_691 ( .A(_abc_40319_new_n1235_), .B(_abc_40319_new_n1134_), .Y(_abc_40319_new_n1954_));
AND2X2 AND2X2_692 ( .A(_abc_40319_new_n1658_), .B(REG3_REG_13_), .Y(_abc_40319_new_n1955_));
AND2X2 AND2X2_693 ( .A(_abc_40319_new_n1955_), .B(REG3_REG_14_), .Y(_abc_40319_new_n1956_));
AND2X2 AND2X2_694 ( .A(_abc_40319_new_n1956_), .B(REG3_REG_15_), .Y(_abc_40319_new_n1957_));
AND2X2 AND2X2_695 ( .A(_abc_40319_new_n1957_), .B(REG3_REG_16_), .Y(_abc_40319_new_n1958_));
AND2X2 AND2X2_696 ( .A(_abc_40319_new_n1958_), .B(REG3_REG_17_), .Y(_abc_40319_new_n1959_));
AND2X2 AND2X2_697 ( .A(_abc_40319_new_n1959_), .B(REG3_REG_18_), .Y(_abc_40319_new_n1960_));
AND2X2 AND2X2_698 ( .A(_abc_40319_new_n1960_), .B(REG3_REG_19_), .Y(_abc_40319_new_n1961_));
AND2X2 AND2X2_699 ( .A(_abc_40319_new_n1961_), .B(REG3_REG_20_), .Y(_abc_40319_new_n1962_));
AND2X2 AND2X2_7 ( .A(_abc_40319_new_n541_), .B(_abc_40319_new_n542_), .Y(_abc_40319_new_n543_));
AND2X2 AND2X2_70 ( .A(_abc_40319_new_n524_), .B(_abc_40319_new_n563_), .Y(_abc_40319_new_n664_));
AND2X2 AND2X2_700 ( .A(_abc_40319_new_n1962_), .B(REG3_REG_21_), .Y(_abc_40319_new_n1963_));
AND2X2 AND2X2_701 ( .A(_abc_40319_new_n1963_), .B(REG3_REG_22_), .Y(_abc_40319_new_n1964_));
AND2X2 AND2X2_702 ( .A(_abc_40319_new_n1964_), .B(REG3_REG_23_), .Y(_abc_40319_new_n1965_));
AND2X2 AND2X2_703 ( .A(_abc_40319_new_n1965_), .B(REG3_REG_24_), .Y(_abc_40319_new_n1966_));
AND2X2 AND2X2_704 ( .A(_abc_40319_new_n1966_), .B(REG3_REG_25_), .Y(_abc_40319_new_n1967_));
AND2X2 AND2X2_705 ( .A(_abc_40319_new_n1967_), .B(REG3_REG_26_), .Y(_abc_40319_new_n1968_));
AND2X2 AND2X2_706 ( .A(_abc_40319_new_n1968_), .B(REG3_REG_27_), .Y(_abc_40319_new_n1969_));
AND2X2 AND2X2_707 ( .A(_abc_40319_new_n1969_), .B(REG3_REG_28_), .Y(_abc_40319_new_n1970_));
AND2X2 AND2X2_708 ( .A(_abc_40319_new_n1971_), .B(_abc_40319_new_n1972_), .Y(_abc_40319_new_n1973_));
AND2X2 AND2X2_709 ( .A(_abc_40319_new_n1973_), .B(_abc_40319_new_n738_), .Y(_abc_40319_new_n1974_));
AND2X2 AND2X2_71 ( .A(_abc_40319_new_n666_), .B(_abc_40319_new_n667_), .Y(_abc_40319_new_n668_));
AND2X2 AND2X2_710 ( .A(_abc_40319_new_n736_), .B(REG0_REG_28_), .Y(_abc_40319_new_n1975_));
AND2X2 AND2X2_711 ( .A(_abc_40319_new_n722_), .B(REG1_REG_28_), .Y(_abc_40319_new_n1976_));
AND2X2 AND2X2_712 ( .A(_abc_40319_new_n733_), .B(REG2_REG_28_), .Y(_abc_40319_new_n1977_));
AND2X2 AND2X2_713 ( .A(_abc_40319_new_n1980_), .B(_abc_40319_new_n1147_), .Y(_abc_40319_new_n1981_));
AND2X2 AND2X2_714 ( .A(_abc_40319_new_n1982_), .B(_abc_40319_new_n1133_), .Y(_abc_40319_new_n1983_));
AND2X2 AND2X2_715 ( .A(_abc_40319_new_n1164_), .B(_abc_40319_new_n1203_), .Y(_abc_40319_new_n1984_));
AND2X2 AND2X2_716 ( .A(_abc_40319_new_n1171_), .B(_abc_40319_new_n1180_), .Y(_abc_40319_new_n1985_));
AND2X2 AND2X2_717 ( .A(n1336), .B(REG3_REG_27_), .Y(_abc_40319_new_n1986_));
AND2X2 AND2X2_718 ( .A(_abc_40319_new_n1924_), .B(_abc_40319_new_n1528_), .Y(_abc_40319_new_n1992_));
AND2X2 AND2X2_719 ( .A(_abc_40319_new_n1995_), .B(_abc_40319_new_n1122_), .Y(_abc_40319_new_n1996_));
AND2X2 AND2X2_72 ( .A(_abc_40319_new_n669_), .B(_abc_40319_new_n665_), .Y(_abc_40319_new_n670_));
AND2X2 AND2X2_720 ( .A(_abc_40319_new_n1996_), .B(_abc_40319_new_n1994_), .Y(_abc_40319_new_n1997_));
AND2X2 AND2X2_721 ( .A(_abc_40319_new_n1134_), .B(_abc_40319_new_n1667_), .Y(_abc_40319_new_n1998_));
AND2X2 AND2X2_722 ( .A(_abc_40319_new_n1147_), .B(_abc_40319_new_n1483_), .Y(_abc_40319_new_n1999_));
AND2X2 AND2X2_723 ( .A(_abc_40319_new_n2000_), .B(_abc_40319_new_n1133_), .Y(_abc_40319_new_n2001_));
AND2X2 AND2X2_724 ( .A(_abc_40319_new_n1164_), .B(_abc_40319_new_n1513_), .Y(_abc_40319_new_n2002_));
AND2X2 AND2X2_725 ( .A(_abc_40319_new_n1171_), .B(_abc_40319_new_n1506_), .Y(_abc_40319_new_n2003_));
AND2X2 AND2X2_726 ( .A(n1336), .B(REG3_REG_14_), .Y(_abc_40319_new_n2004_));
AND2X2 AND2X2_727 ( .A(_abc_40319_new_n1915_), .B(_abc_40319_new_n1328_), .Y(_abc_40319_new_n2010_));
AND2X2 AND2X2_728 ( .A(_abc_40319_new_n2013_), .B(_abc_40319_new_n1122_), .Y(_abc_40319_new_n2014_));
AND2X2 AND2X2_729 ( .A(_abc_40319_new_n2014_), .B(_abc_40319_new_n2012_), .Y(_abc_40319_new_n2015_));
AND2X2 AND2X2_73 ( .A(_abc_40319_new_n671_), .B(_abc_40319_new_n655_), .Y(_abc_40319_new_n672_));
AND2X2 AND2X2_730 ( .A(_abc_40319_new_n1134_), .B(_abc_40319_new_n1340_), .Y(_abc_40319_new_n2016_));
AND2X2 AND2X2_731 ( .A(_abc_40319_new_n1285_), .B(_abc_40319_new_n1147_), .Y(_abc_40319_new_n2017_));
AND2X2 AND2X2_732 ( .A(_abc_40319_new_n2018_), .B(_abc_40319_new_n1133_), .Y(_abc_40319_new_n2019_));
AND2X2 AND2X2_733 ( .A(_abc_40319_new_n1164_), .B(_abc_40319_new_n1310_), .Y(_abc_40319_new_n2020_));
AND2X2 AND2X2_734 ( .A(_abc_40319_new_n1171_), .B(_abc_40319_new_n1306_), .Y(_abc_40319_new_n2021_));
AND2X2 AND2X2_735 ( .A(n1336), .B(REG3_REG_23_), .Y(_abc_40319_new_n2022_));
AND2X2 AND2X2_736 ( .A(_abc_40319_new_n1782_), .B(_abc_40319_new_n2028_), .Y(_abc_40319_new_n2029_));
AND2X2 AND2X2_737 ( .A(_abc_40319_new_n2032_), .B(_abc_40319_new_n1122_), .Y(_abc_40319_new_n2033_));
AND2X2 AND2X2_738 ( .A(_abc_40319_new_n2033_), .B(_abc_40319_new_n2031_), .Y(_abc_40319_new_n2034_));
AND2X2 AND2X2_739 ( .A(_abc_40319_new_n1134_), .B(_abc_40319_new_n1625_), .Y(_abc_40319_new_n2035_));
AND2X2 AND2X2_74 ( .A(_abc_40319_new_n663_), .B(_abc_40319_new_n672_), .Y(_abc_40319_new_n673_));
AND2X2 AND2X2_740 ( .A(_abc_40319_new_n1147_), .B(_abc_40319_new_n1735_), .Y(_abc_40319_new_n2036_));
AND2X2 AND2X2_741 ( .A(_abc_40319_new_n2037_), .B(_abc_40319_new_n1133_), .Y(_abc_40319_new_n2038_));
AND2X2 AND2X2_742 ( .A(_abc_40319_new_n1164_), .B(_abc_40319_new_n1766_), .Y(_abc_40319_new_n2039_));
AND2X2 AND2X2_743 ( .A(_abc_40319_new_n1171_), .B(_abc_40319_new_n1758_), .Y(_abc_40319_new_n2040_));
AND2X2 AND2X2_744 ( .A(n1336), .B(REG3_REG_10_), .Y(_abc_40319_new_n2041_));
AND2X2 AND2X2_745 ( .A(_abc_40319_new_n835_), .B(_abc_40319_new_n838_), .Y(_abc_40319_new_n2047_));
AND2X2 AND2X2_746 ( .A(_abc_40319_new_n968_), .B(_abc_40319_new_n2049_), .Y(_abc_40319_new_n2050_));
AND2X2 AND2X2_747 ( .A(_abc_40319_new_n2055_), .B(_abc_40319_new_n1122_), .Y(_abc_40319_new_n2056_));
AND2X2 AND2X2_748 ( .A(_abc_40319_new_n2056_), .B(_abc_40319_new_n2053_), .Y(_abc_40319_new_n2057_));
AND2X2 AND2X2_749 ( .A(_abc_40319_new_n1134_), .B(_abc_40319_new_n865_), .Y(_abc_40319_new_n2058_));
AND2X2 AND2X2_75 ( .A(_abc_40319_new_n676_), .B(_abc_40319_new_n534_), .Y(_abc_40319_new_n677_));
AND2X2 AND2X2_750 ( .A(_abc_40319_new_n1147_), .B(_abc_40319_new_n795_), .Y(_abc_40319_new_n2059_));
AND2X2 AND2X2_751 ( .A(_abc_40319_new_n2060_), .B(_abc_40319_new_n1133_), .Y(_abc_40319_new_n2061_));
AND2X2 AND2X2_752 ( .A(_abc_40319_new_n1171_), .B(_abc_40319_new_n820_), .Y(_abc_40319_new_n2062_));
AND2X2 AND2X2_753 ( .A(n1336), .B(REG3_REG_3_), .Y(_abc_40319_new_n2063_));
AND2X2 AND2X2_754 ( .A(_abc_40319_new_n1164_), .B(_abc_40319_new_n826_), .Y(_abc_40319_new_n2066_));
AND2X2 AND2X2_755 ( .A(_abc_40319_new_n1840_), .B(_abc_40319_new_n1893_), .Y(_abc_40319_new_n2070_));
AND2X2 AND2X2_756 ( .A(_abc_40319_new_n2073_), .B(_abc_40319_new_n1122_), .Y(_abc_40319_new_n2074_));
AND2X2 AND2X2_757 ( .A(_abc_40319_new_n2074_), .B(_abc_40319_new_n2072_), .Y(_abc_40319_new_n2075_));
AND2X2 AND2X2_758 ( .A(_abc_40319_new_n1134_), .B(_abc_40319_new_n1374_), .Y(_abc_40319_new_n2076_));
AND2X2 AND2X2_759 ( .A(_abc_40319_new_n1147_), .B(_abc_40319_new_n1852_), .Y(_abc_40319_new_n2077_));
AND2X2 AND2X2_76 ( .A(_abc_40319_new_n678_), .B(IR_REG_5_), .Y(_abc_40319_new_n679_));
AND2X2 AND2X2_760 ( .A(_abc_40319_new_n2078_), .B(_abc_40319_new_n1133_), .Y(_abc_40319_new_n2079_));
AND2X2 AND2X2_761 ( .A(_abc_40319_new_n1164_), .B(_abc_40319_new_n1822_), .Y(_abc_40319_new_n2080_));
AND2X2 AND2X2_762 ( .A(_abc_40319_new_n1171_), .B(_abc_40319_new_n1817_), .Y(_abc_40319_new_n2081_));
AND2X2 AND2X2_763 ( .A(n1336), .B(REG3_REG_19_), .Y(_abc_40319_new_n2082_));
AND2X2 AND2X2_764 ( .A(_abc_40319_new_n817_), .B(DATAI_28_), .Y(_abc_40319_new_n2089_));
AND2X2 AND2X2_765 ( .A(_abc_40319_new_n2089_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n2090_));
AND2X2 AND2X2_766 ( .A(_abc_40319_new_n1980_), .B(_abc_40319_new_n705_), .Y(_abc_40319_new_n2091_));
AND2X2 AND2X2_767 ( .A(_abc_40319_new_n763_), .B(_abc_40319_new_n2089_), .Y(_abc_40319_new_n2093_));
AND2X2 AND2X2_768 ( .A(_abc_40319_new_n1980_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n2094_));
AND2X2 AND2X2_769 ( .A(_abc_40319_new_n2096_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n2097_));
AND2X2 AND2X2_77 ( .A(_abc_40319_new_n681_), .B(IR_REG_31_), .Y(_abc_40319_new_n682_));
AND2X2 AND2X2_770 ( .A(_abc_40319_new_n2095_), .B(_abc_40319_new_n768_), .Y(_abc_40319_new_n2098_));
AND2X2 AND2X2_771 ( .A(_abc_40319_new_n2103_), .B(_abc_40319_new_n2100_), .Y(_abc_40319_new_n2104_));
AND2X2 AND2X2_772 ( .A(_abc_40319_new_n2105_), .B(_abc_40319_new_n1222_), .Y(_abc_40319_new_n2106_));
AND2X2 AND2X2_773 ( .A(_abc_40319_new_n2088_), .B(_abc_40319_new_n2106_), .Y(_abc_40319_new_n2107_));
AND2X2 AND2X2_774 ( .A(_abc_40319_new_n2104_), .B(_abc_40319_new_n1221_), .Y(_abc_40319_new_n2110_));
AND2X2 AND2X2_775 ( .A(_abc_40319_new_n2109_), .B(_abc_40319_new_n2110_), .Y(_abc_40319_new_n2111_));
AND2X2 AND2X2_776 ( .A(_abc_40319_new_n2112_), .B(_abc_40319_new_n1122_), .Y(_abc_40319_new_n2113_));
AND2X2 AND2X2_777 ( .A(_abc_40319_new_n1210_), .B(_abc_40319_new_n1134_), .Y(_abc_40319_new_n2114_));
AND2X2 AND2X2_778 ( .A(_abc_40319_new_n722_), .B(REG1_REG_29_), .Y(_abc_40319_new_n2115_));
AND2X2 AND2X2_779 ( .A(_abc_40319_new_n736_), .B(REG0_REG_29_), .Y(_abc_40319_new_n2116_));
AND2X2 AND2X2_78 ( .A(_abc_40319_new_n524_), .B(IR_REG_5_), .Y(_abc_40319_new_n683_));
AND2X2 AND2X2_780 ( .A(_abc_40319_new_n733_), .B(REG2_REG_29_), .Y(_abc_40319_new_n2117_));
AND2X2 AND2X2_781 ( .A(REG3_REG_27_), .B(REG3_REG_28_), .Y(_abc_40319_new_n2118_));
AND2X2 AND2X2_782 ( .A(_abc_40319_new_n1199_), .B(_abc_40319_new_n2118_), .Y(_abc_40319_new_n2119_));
AND2X2 AND2X2_783 ( .A(_abc_40319_new_n2119_), .B(_abc_40319_new_n738_), .Y(_abc_40319_new_n2120_));
AND2X2 AND2X2_784 ( .A(_abc_40319_new_n2123_), .B(_abc_40319_new_n1147_), .Y(_abc_40319_new_n2124_));
AND2X2 AND2X2_785 ( .A(_abc_40319_new_n2125_), .B(_abc_40319_new_n1133_), .Y(_abc_40319_new_n2126_));
AND2X2 AND2X2_786 ( .A(_abc_40319_new_n1973_), .B(_abc_40319_new_n1164_), .Y(_abc_40319_new_n2127_));
AND2X2 AND2X2_787 ( .A(_abc_40319_new_n1171_), .B(_abc_40319_new_n2089_), .Y(_abc_40319_new_n2128_));
AND2X2 AND2X2_788 ( .A(n1336), .B(REG3_REG_28_), .Y(_abc_40319_new_n2129_));
AND2X2 AND2X2_789 ( .A(_abc_40319_new_n1586_), .B(_abc_40319_new_n1593_), .Y(_abc_40319_new_n2135_));
AND2X2 AND2X2_79 ( .A(_abc_40319_new_n640_), .B(_abc_40319_new_n685_), .Y(_abc_40319_new_n686_));
AND2X2 AND2X2_790 ( .A(_abc_40319_new_n982_), .B(_abc_40319_new_n1588_), .Y(_abc_40319_new_n2136_));
AND2X2 AND2X2_791 ( .A(_abc_40319_new_n2137_), .B(_abc_40319_new_n1598_), .Y(_abc_40319_new_n2138_));
AND2X2 AND2X2_792 ( .A(_abc_40319_new_n2142_), .B(_abc_40319_new_n1122_), .Y(_abc_40319_new_n2143_));
AND2X2 AND2X2_793 ( .A(_abc_40319_new_n2143_), .B(_abc_40319_new_n2140_), .Y(_abc_40319_new_n2144_));
AND2X2 AND2X2_794 ( .A(_abc_40319_new_n1134_), .B(_abc_40319_new_n1046_), .Y(_abc_40319_new_n2145_));
AND2X2 AND2X2_795 ( .A(_abc_40319_new_n1147_), .B(_abc_40319_new_n1625_), .Y(_abc_40319_new_n2146_));
AND2X2 AND2X2_796 ( .A(_abc_40319_new_n2147_), .B(_abc_40319_new_n1133_), .Y(_abc_40319_new_n2148_));
AND2X2 AND2X2_797 ( .A(_abc_40319_new_n1164_), .B(_abc_40319_new_n1139_), .Y(_abc_40319_new_n2149_));
AND2X2 AND2X2_798 ( .A(_abc_40319_new_n1171_), .B(_abc_40319_new_n1572_), .Y(_abc_40319_new_n2150_));
AND2X2 AND2X2_799 ( .A(n1336), .B(REG3_REG_8_), .Y(_abc_40319_new_n2151_));
AND2X2 AND2X2_8 ( .A(_abc_40319_new_n540_), .B(_abc_40319_new_n543_), .Y(_abc_40319_new_n544_));
AND2X2 AND2X2_80 ( .A(_abc_40319_new_n687_), .B(_abc_40319_new_n688_), .Y(_abc_40319_new_n689_));
AND2X2 AND2X2_800 ( .A(_abc_40319_new_n1536_), .B(_abc_40319_new_n916_), .Y(_abc_40319_new_n2158_));
AND2X2 AND2X2_801 ( .A(_abc_40319_new_n2159_), .B(_abc_40319_new_n1122_), .Y(_abc_40319_new_n2160_));
AND2X2 AND2X2_802 ( .A(_abc_40319_new_n2160_), .B(_abc_40319_new_n2157_), .Y(_abc_40319_new_n2161_));
AND2X2 AND2X2_803 ( .A(_abc_40319_new_n1134_), .B(_abc_40319_new_n924_), .Y(_abc_40319_new_n2162_));
AND2X2 AND2X2_804 ( .A(_abc_40319_new_n1147_), .B(_abc_40319_new_n865_), .Y(_abc_40319_new_n2163_));
AND2X2 AND2X2_805 ( .A(_abc_40319_new_n2164_), .B(_abc_40319_new_n1133_), .Y(_abc_40319_new_n2165_));
AND2X2 AND2X2_806 ( .A(_abc_40319_new_n1171_), .B(_abc_40319_new_n891_), .Y(_abc_40319_new_n2166_));
AND2X2 AND2X2_807 ( .A(n1336), .B(REG3_REG_1_), .Y(_abc_40319_new_n2167_));
AND2X2 AND2X2_808 ( .A(_abc_40319_new_n1164_), .B(REG3_REG_1_), .Y(_abc_40319_new_n2170_));
AND2X2 AND2X2_809 ( .A(_abc_40319_new_n1813_), .B(_abc_40319_new_n1840_), .Y(_abc_40319_new_n2174_));
AND2X2 AND2X2_81 ( .A(_abc_40319_new_n689_), .B(_abc_40319_new_n673_), .Y(_abc_40319_new_n690_));
AND2X2 AND2X2_810 ( .A(_abc_40319_new_n2176_), .B(_abc_40319_new_n1899_), .Y(_abc_40319_new_n2177_));
AND2X2 AND2X2_811 ( .A(_abc_40319_new_n2175_), .B(_abc_40319_new_n1864_), .Y(_abc_40319_new_n2181_));
AND2X2 AND2X2_812 ( .A(_abc_40319_new_n1889_), .B(_abc_40319_new_n1898_), .Y(_abc_40319_new_n2183_));
AND2X2 AND2X2_813 ( .A(_abc_40319_new_n2185_), .B(_abc_40319_new_n1122_), .Y(_abc_40319_new_n2186_));
AND2X2 AND2X2_814 ( .A(_abc_40319_new_n2186_), .B(_abc_40319_new_n2180_), .Y(_abc_40319_new_n2187_));
AND2X2 AND2X2_815 ( .A(_abc_40319_new_n1147_), .B(_abc_40319_new_n1340_), .Y(_abc_40319_new_n2188_));
AND2X2 AND2X2_816 ( .A(_abc_40319_new_n1134_), .B(_abc_40319_new_n1852_), .Y(_abc_40319_new_n2189_));
AND2X2 AND2X2_817 ( .A(_abc_40319_new_n1151_), .B(_abc_40319_new_n1869_), .Y(_abc_40319_new_n2190_));
AND2X2 AND2X2_818 ( .A(_abc_40319_new_n2192_), .B(_abc_40319_new_n1133_), .Y(_abc_40319_new_n2193_));
AND2X2 AND2X2_819 ( .A(_abc_40319_new_n1162_), .B(_abc_40319_new_n1869_), .Y(_abc_40319_new_n2194_));
AND2X2 AND2X2_82 ( .A(_abc_40319_new_n524_), .B(_abc_40319_new_n562_), .Y(_abc_40319_new_n691_));
AND2X2 AND2X2_820 ( .A(_abc_40319_new_n1171_), .B(_abc_40319_new_n1865_), .Y(_abc_40319_new_n2195_));
AND2X2 AND2X2_821 ( .A(n1336), .B(REG3_REG_21_), .Y(_abc_40319_new_n2196_));
AND2X2 AND2X2_822 ( .A(_abc_40319_new_n1713_), .B(_abc_40319_new_n1791_), .Y(_abc_40319_new_n2202_));
AND2X2 AND2X2_823 ( .A(_abc_40319_new_n1643_), .B(_abc_40319_new_n1782_), .Y(_abc_40319_new_n2203_));
AND2X2 AND2X2_824 ( .A(_abc_40319_new_n2204_), .B(_abc_40319_new_n1748_), .Y(_abc_40319_new_n2205_));
AND2X2 AND2X2_825 ( .A(_abc_40319_new_n2210_), .B(_abc_40319_new_n1122_), .Y(_abc_40319_new_n2211_));
AND2X2 AND2X2_826 ( .A(_abc_40319_new_n2211_), .B(_abc_40319_new_n2207_), .Y(_abc_40319_new_n2212_));
AND2X2 AND2X2_827 ( .A(_abc_40319_new_n1134_), .B(_abc_40319_new_n1735_), .Y(_abc_40319_new_n2213_));
AND2X2 AND2X2_828 ( .A(_abc_40319_new_n1147_), .B(_abc_40319_new_n1667_), .Y(_abc_40319_new_n2214_));
AND2X2 AND2X2_829 ( .A(_abc_40319_new_n2215_), .B(_abc_40319_new_n1133_), .Y(_abc_40319_new_n2216_));
AND2X2 AND2X2_83 ( .A(_abc_40319_new_n693_), .B(_abc_40319_new_n694_), .Y(_abc_40319_new_n695_));
AND2X2 AND2X2_830 ( .A(_abc_40319_new_n1164_), .B(_abc_40319_new_n1698_), .Y(_abc_40319_new_n2217_));
AND2X2 AND2X2_831 ( .A(_abc_40319_new_n1171_), .B(_abc_40319_new_n1690_), .Y(_abc_40319_new_n2218_));
AND2X2 AND2X2_832 ( .A(n1336), .B(REG3_REG_12_), .Y(_abc_40319_new_n2219_));
AND2X2 AND2X2_833 ( .A(_abc_40319_new_n1272_), .B(_abc_40319_new_n1301_), .Y(_abc_40319_new_n2225_));
AND2X2 AND2X2_834 ( .A(_abc_40319_new_n1908_), .B(_abc_40319_new_n1909_), .Y(_abc_40319_new_n2226_));
AND2X2 AND2X2_835 ( .A(_abc_40319_new_n2231_), .B(_abc_40319_new_n1122_), .Y(_abc_40319_new_n2232_));
AND2X2 AND2X2_836 ( .A(_abc_40319_new_n2232_), .B(_abc_40319_new_n2228_), .Y(_abc_40319_new_n2233_));
AND2X2 AND2X2_837 ( .A(_abc_40319_new_n1285_), .B(_abc_40319_new_n1134_), .Y(_abc_40319_new_n2234_));
AND2X2 AND2X2_838 ( .A(_abc_40319_new_n1235_), .B(_abc_40319_new_n1147_), .Y(_abc_40319_new_n2235_));
AND2X2 AND2X2_839 ( .A(_abc_40319_new_n2236_), .B(_abc_40319_new_n1133_), .Y(_abc_40319_new_n2237_));
AND2X2 AND2X2_84 ( .A(_abc_40319_new_n696_), .B(_abc_40319_new_n692_), .Y(_abc_40319_new_n697_));
AND2X2 AND2X2_840 ( .A(_abc_40319_new_n1164_), .B(_abc_40319_new_n1253_), .Y(_abc_40319_new_n2238_));
AND2X2 AND2X2_841 ( .A(_abc_40319_new_n1171_), .B(_abc_40319_new_n1249_), .Y(_abc_40319_new_n2239_));
AND2X2 AND2X2_842 ( .A(n1336), .B(REG3_REG_25_), .Y(_abc_40319_new_n2240_));
AND2X2 AND2X2_843 ( .A(_abc_40319_new_n1423_), .B(_abc_40319_new_n1805_), .Y(_abc_40319_new_n2246_));
AND2X2 AND2X2_844 ( .A(_abc_40319_new_n2249_), .B(_abc_40319_new_n1122_), .Y(_abc_40319_new_n2250_));
AND2X2 AND2X2_845 ( .A(_abc_40319_new_n2250_), .B(_abc_40319_new_n2248_), .Y(_abc_40319_new_n2251_));
AND2X2 AND2X2_846 ( .A(_abc_40319_new_n1134_), .B(_abc_40319_new_n1483_), .Y(_abc_40319_new_n2252_));
AND2X2 AND2X2_847 ( .A(_abc_40319_new_n1147_), .B(_abc_40319_new_n1444_), .Y(_abc_40319_new_n2253_));
AND2X2 AND2X2_848 ( .A(_abc_40319_new_n2254_), .B(_abc_40319_new_n1133_), .Y(_abc_40319_new_n2255_));
AND2X2 AND2X2_849 ( .A(_abc_40319_new_n1171_), .B(_abc_40319_new_n1398_), .Y(_abc_40319_new_n2256_));
AND2X2 AND2X2_85 ( .A(_abc_40319_new_n646_), .B(_abc_40319_new_n698_), .Y(_abc_40319_new_n699_));
AND2X2 AND2X2_850 ( .A(n1336), .B(REG3_REG_16_), .Y(_abc_40319_new_n2257_));
AND2X2 AND2X2_851 ( .A(_abc_40319_new_n1164_), .B(_abc_40319_new_n1406_), .Y(_abc_40319_new_n2260_));
AND2X2 AND2X2_852 ( .A(_abc_40319_new_n1594_), .B(_abc_40319_new_n773_), .Y(_abc_40319_new_n2264_));
AND2X2 AND2X2_853 ( .A(_abc_40319_new_n2267_), .B(_abc_40319_new_n1122_), .Y(_abc_40319_new_n2268_));
AND2X2 AND2X2_854 ( .A(_abc_40319_new_n2268_), .B(_abc_40319_new_n2266_), .Y(_abc_40319_new_n2269_));
AND2X2 AND2X2_855 ( .A(_abc_40319_new_n1134_), .B(_abc_40319_new_n795_), .Y(_abc_40319_new_n2270_));
AND2X2 AND2X2_856 ( .A(_abc_40319_new_n1147_), .B(_abc_40319_new_n1010_), .Y(_abc_40319_new_n2271_));
AND2X2 AND2X2_857 ( .A(_abc_40319_new_n2272_), .B(_abc_40319_new_n1133_), .Y(_abc_40319_new_n2273_));
AND2X2 AND2X2_858 ( .A(_abc_40319_new_n1171_), .B(_abc_40319_new_n689_), .Y(_abc_40319_new_n2274_));
AND2X2 AND2X2_859 ( .A(n1336), .B(REG3_REG_5_), .Y(_abc_40319_new_n2275_));
AND2X2 AND2X2_86 ( .A(_abc_40319_new_n701_), .B(_abc_40319_new_n702_), .Y(_abc_40319_new_n703_));
AND2X2 AND2X2_860 ( .A(_abc_40319_new_n1164_), .B(_abc_40319_new_n743_), .Y(_abc_40319_new_n2278_));
AND2X2 AND2X2_861 ( .A(_abc_40319_new_n1802_), .B(_abc_40319_new_n1423_), .Y(_abc_40319_new_n2282_));
AND2X2 AND2X2_862 ( .A(_abc_40319_new_n1457_), .B(_abc_40319_new_n1807_), .Y(_abc_40319_new_n2283_));
AND2X2 AND2X2_863 ( .A(_abc_40319_new_n1936_), .B(_abc_40319_new_n1805_), .Y(_abc_40319_new_n2286_));
AND2X2 AND2X2_864 ( .A(_abc_40319_new_n2288_), .B(_abc_40319_new_n1122_), .Y(_abc_40319_new_n2289_));
AND2X2 AND2X2_865 ( .A(_abc_40319_new_n2289_), .B(_abc_40319_new_n2285_), .Y(_abc_40319_new_n2290_));
AND2X2 AND2X2_866 ( .A(_abc_40319_new_n1134_), .B(_abc_40319_new_n1410_), .Y(_abc_40319_new_n2291_));
AND2X2 AND2X2_867 ( .A(_abc_40319_new_n1147_), .B(_abc_40319_new_n1374_), .Y(_abc_40319_new_n2292_));
AND2X2 AND2X2_868 ( .A(_abc_40319_new_n2293_), .B(_abc_40319_new_n1133_), .Y(_abc_40319_new_n2294_));
AND2X2 AND2X2_869 ( .A(_abc_40319_new_n1171_), .B(_abc_40319_new_n1433_), .Y(_abc_40319_new_n2295_));
AND2X2 AND2X2_87 ( .A(_abc_40319_new_n524_), .B(_abc_40319_new_n706_), .Y(_abc_40319_new_n707_));
AND2X2 AND2X2_870 ( .A(n1336), .B(REG3_REG_17_), .Y(_abc_40319_new_n2296_));
AND2X2 AND2X2_871 ( .A(_abc_40319_new_n1164_), .B(_abc_40319_new_n1440_), .Y(_abc_40319_new_n2299_));
AND2X2 AND2X2_872 ( .A(_abc_40319_new_n2303_), .B(_abc_40319_new_n1909_), .Y(_abc_40319_new_n2304_));
AND2X2 AND2X2_873 ( .A(_abc_40319_new_n2307_), .B(_abc_40319_new_n1122_), .Y(_abc_40319_new_n2308_));
AND2X2 AND2X2_874 ( .A(_abc_40319_new_n2308_), .B(_abc_40319_new_n2306_), .Y(_abc_40319_new_n2309_));
AND2X2 AND2X2_875 ( .A(_abc_40319_new_n1317_), .B(_abc_40319_new_n1134_), .Y(_abc_40319_new_n2310_));
AND2X2 AND2X2_876 ( .A(_abc_40319_new_n1260_), .B(_abc_40319_new_n1147_), .Y(_abc_40319_new_n2311_));
AND2X2 AND2X2_877 ( .A(_abc_40319_new_n2312_), .B(_abc_40319_new_n1133_), .Y(_abc_40319_new_n2313_));
AND2X2 AND2X2_878 ( .A(_abc_40319_new_n1164_), .B(_abc_40319_new_n1278_), .Y(_abc_40319_new_n2314_));
AND2X2 AND2X2_879 ( .A(_abc_40319_new_n1171_), .B(_abc_40319_new_n1274_), .Y(_abc_40319_new_n2315_));
AND2X2 AND2X2_88 ( .A(_abc_40319_new_n630_), .B(_abc_40319_new_n708_), .Y(_abc_40319_new_n709_));
AND2X2 AND2X2_880 ( .A(n1336), .B(REG3_REG_24_), .Y(_abc_40319_new_n2316_));
AND2X2 AND2X2_881 ( .A(_abc_40319_new_n1529_), .B(_abc_40319_new_n807_), .Y(_abc_40319_new_n2322_));
AND2X2 AND2X2_882 ( .A(_abc_40319_new_n2325_), .B(_abc_40319_new_n1122_), .Y(_abc_40319_new_n2326_));
AND2X2 AND2X2_883 ( .A(_abc_40319_new_n2326_), .B(_abc_40319_new_n2324_), .Y(_abc_40319_new_n2327_));
AND2X2 AND2X2_884 ( .A(_abc_40319_new_n1134_), .B(_abc_40319_new_n829_), .Y(_abc_40319_new_n2328_));
AND2X2 AND2X2_885 ( .A(_abc_40319_new_n1147_), .B(_abc_40319_new_n746_), .Y(_abc_40319_new_n2329_));
AND2X2 AND2X2_886 ( .A(_abc_40319_new_n2330_), .B(_abc_40319_new_n1133_), .Y(_abc_40319_new_n2331_));
AND2X2 AND2X2_887 ( .A(_abc_40319_new_n1171_), .B(_abc_40319_new_n784_), .Y(_abc_40319_new_n2332_));
AND2X2 AND2X2_888 ( .A(n1336), .B(REG3_REG_4_), .Y(_abc_40319_new_n2333_));
AND2X2 AND2X2_889 ( .A(_abc_40319_new_n1164_), .B(_abc_40319_new_n792_), .Y(_abc_40319_new_n2336_));
AND2X2 AND2X2_89 ( .A(_abc_40319_new_n623_), .B(_abc_40319_new_n709_), .Y(_abc_40319_new_n710_));
AND2X2 AND2X2_890 ( .A(_abc_40319_new_n1926_), .B(_abc_40319_new_n1634_), .Y(_abc_40319_new_n2341_));
AND2X2 AND2X2_891 ( .A(_abc_40319_new_n2342_), .B(_abc_40319_new_n2340_), .Y(_abc_40319_new_n2343_));
AND2X2 AND2X2_892 ( .A(_abc_40319_new_n2343_), .B(_abc_40319_new_n1122_), .Y(_abc_40319_new_n2344_));
AND2X2 AND2X2_893 ( .A(_abc_40319_new_n1134_), .B(_abc_40319_new_n1146_), .Y(_abc_40319_new_n2345_));
AND2X2 AND2X2_894 ( .A(_abc_40319_new_n1147_), .B(_abc_40319_new_n1769_), .Y(_abc_40319_new_n2346_));
AND2X2 AND2X2_895 ( .A(_abc_40319_new_n2347_), .B(_abc_40319_new_n1133_), .Y(_abc_40319_new_n2348_));
AND2X2 AND2X2_896 ( .A(_abc_40319_new_n1164_), .B(_abc_40319_new_n1618_), .Y(_abc_40319_new_n2349_));
AND2X2 AND2X2_897 ( .A(_abc_40319_new_n1171_), .B(_abc_40319_new_n1614_), .Y(_abc_40319_new_n2350_));
AND2X2 AND2X2_898 ( .A(n1336), .B(REG3_REG_9_), .Y(_abc_40319_new_n2351_));
AND2X2 AND2X2_899 ( .A(_abc_40319_new_n1542_), .B(_abc_40319_new_n935_), .Y(_abc_40319_new_n2357_));
AND2X2 AND2X2_9 ( .A(_abc_40319_new_n545_), .B(_abc_40319_new_n546_), .Y(_abc_40319_new_n547_));
AND2X2 AND2X2_90 ( .A(_abc_40319_new_n710_), .B(_abc_40319_new_n706_), .Y(_abc_40319_new_n711_));
AND2X2 AND2X2_900 ( .A(_abc_40319_new_n2359_), .B(_abc_40319_new_n2360_), .Y(_abc_40319_new_n2361_));
AND2X2 AND2X2_901 ( .A(_abc_40319_new_n2361_), .B(_abc_40319_new_n1122_), .Y(_abc_40319_new_n2362_));
AND2X2 AND2X2_902 ( .A(n1336), .B(REG3_REG_0_), .Y(_abc_40319_new_n2363_));
AND2X2 AND2X2_903 ( .A(_abc_40319_new_n1171_), .B(_abc_40319_new_n930_), .Y(_abc_40319_new_n2365_));
AND2X2 AND2X2_904 ( .A(_abc_40319_new_n904_), .B(_abc_40319_new_n1133_), .Y(_abc_40319_new_n2366_));
AND2X2 AND2X2_905 ( .A(_abc_40319_new_n1147_), .B(_abc_40319_new_n2366_), .Y(_abc_40319_new_n2367_));
AND2X2 AND2X2_906 ( .A(_abc_40319_new_n1164_), .B(REG3_REG_0_), .Y(_abc_40319_new_n2369_));
AND2X2 AND2X2_907 ( .A(_abc_40319_new_n1864_), .B(_abc_40319_new_n1899_), .Y(_abc_40319_new_n2373_));
AND2X2 AND2X2_908 ( .A(_abc_40319_new_n2376_), .B(_abc_40319_new_n1122_), .Y(_abc_40319_new_n2377_));
AND2X2 AND2X2_909 ( .A(_abc_40319_new_n2377_), .B(_abc_40319_new_n2375_), .Y(_abc_40319_new_n2378_));
AND2X2 AND2X2_91 ( .A(_abc_40319_new_n712_), .B(IR_REG_30_), .Y(_abc_40319_new_n713_));
AND2X2 AND2X2_910 ( .A(_abc_40319_new_n1134_), .B(_abc_40319_new_n1828_), .Y(_abc_40319_new_n2379_));
AND2X2 AND2X2_911 ( .A(_abc_40319_new_n1147_), .B(_abc_40319_new_n1876_), .Y(_abc_40319_new_n2380_));
AND2X2 AND2X2_912 ( .A(_abc_40319_new_n2381_), .B(_abc_40319_new_n1133_), .Y(_abc_40319_new_n2382_));
AND2X2 AND2X2_913 ( .A(_abc_40319_new_n1171_), .B(_abc_40319_new_n1841_), .Y(_abc_40319_new_n2383_));
AND2X2 AND2X2_914 ( .A(n1336), .B(REG3_REG_20_), .Y(_abc_40319_new_n2384_));
AND2X2 AND2X2_915 ( .A(_abc_40319_new_n1164_), .B(_abc_40319_new_n1846_), .Y(_abc_40319_new_n2387_));
AND2X2 AND2X2_916 ( .A(_abc_40319_new_n2209_), .B(_abc_40319_new_n1791_), .Y(_abc_40319_new_n2391_));
AND2X2 AND2X2_917 ( .A(_abc_40319_new_n2206_), .B(_abc_40319_new_n1713_), .Y(_abc_40319_new_n2396_));
AND2X2 AND2X2_918 ( .A(_abc_40319_new_n1679_), .B(_abc_40319_new_n1792_), .Y(_abc_40319_new_n2398_));
AND2X2 AND2X2_919 ( .A(_abc_40319_new_n2400_), .B(_abc_40319_new_n1122_), .Y(_abc_40319_new_n2401_));
AND2X2 AND2X2_92 ( .A(_abc_40319_new_n714_), .B(IR_REG_31_), .Y(_abc_40319_new_n715_));
AND2X2 AND2X2_920 ( .A(_abc_40319_new_n2401_), .B(_abc_40319_new_n2395_), .Y(_abc_40319_new_n2402_));
AND2X2 AND2X2_921 ( .A(_abc_40319_new_n1147_), .B(_abc_40319_new_n1517_), .Y(_abc_40319_new_n2403_));
AND2X2 AND2X2_922 ( .A(_abc_40319_new_n1134_), .B(_abc_40319_new_n1701_), .Y(_abc_40319_new_n2404_));
AND2X2 AND2X2_923 ( .A(_abc_40319_new_n1151_), .B(_abc_40319_new_n1660_), .Y(_abc_40319_new_n2405_));
AND2X2 AND2X2_924 ( .A(_abc_40319_new_n2407_), .B(_abc_40319_new_n1133_), .Y(_abc_40319_new_n2408_));
AND2X2 AND2X2_925 ( .A(_abc_40319_new_n1162_), .B(_abc_40319_new_n1660_), .Y(_abc_40319_new_n2409_));
AND2X2 AND2X2_926 ( .A(_abc_40319_new_n1171_), .B(_abc_40319_new_n1655_), .Y(_abc_40319_new_n2410_));
AND2X2 AND2X2_927 ( .A(n1336), .B(REG3_REG_13_), .Y(_abc_40319_new_n2411_));
AND2X2 AND2X2_928 ( .A(_abc_40319_new_n1917_), .B(_abc_40319_new_n1352_), .Y(_abc_40319_new_n2417_));
AND2X2 AND2X2_929 ( .A(_abc_40319_new_n2420_), .B(_abc_40319_new_n1122_), .Y(_abc_40319_new_n2421_));
AND2X2 AND2X2_93 ( .A(_abc_40319_new_n717_), .B(_abc_40319_new_n712_), .Y(_abc_40319_new_n718_));
AND2X2 AND2X2_930 ( .A(_abc_40319_new_n2421_), .B(_abc_40319_new_n2418_), .Y(_abc_40319_new_n2422_));
AND2X2 AND2X2_931 ( .A(_abc_40319_new_n1134_), .B(_abc_40319_new_n1876_), .Y(_abc_40319_new_n2423_));
AND2X2 AND2X2_932 ( .A(_abc_40319_new_n1317_), .B(_abc_40319_new_n1147_), .Y(_abc_40319_new_n2424_));
AND2X2 AND2X2_933 ( .A(_abc_40319_new_n2425_), .B(_abc_40319_new_n1133_), .Y(_abc_40319_new_n2426_));
AND2X2 AND2X2_934 ( .A(_abc_40319_new_n1164_), .B(_abc_40319_new_n1333_), .Y(_abc_40319_new_n2427_));
AND2X2 AND2X2_935 ( .A(_abc_40319_new_n1171_), .B(_abc_40319_new_n1329_), .Y(_abc_40319_new_n2428_));
AND2X2 AND2X2_936 ( .A(n1336), .B(REG3_REG_22_), .Y(_abc_40319_new_n2429_));
AND2X2 AND2X2_937 ( .A(_abc_40319_new_n2439_), .B(_abc_40319_new_n1122_), .Y(_abc_40319_new_n2440_));
AND2X2 AND2X2_938 ( .A(_abc_40319_new_n2440_), .B(_abc_40319_new_n2437_), .Y(_abc_40319_new_n2441_));
AND2X2 AND2X2_939 ( .A(_abc_40319_new_n1134_), .B(_abc_40319_new_n1769_), .Y(_abc_40319_new_n2442_));
AND2X2 AND2X2_94 ( .A(_abc_40319_new_n718_), .B(IR_REG_31_), .Y(_abc_40319_new_n719_));
AND2X2 AND2X2_940 ( .A(_abc_40319_new_n1147_), .B(_abc_40319_new_n1701_), .Y(_abc_40319_new_n2443_));
AND2X2 AND2X2_941 ( .A(_abc_40319_new_n2444_), .B(_abc_40319_new_n1133_), .Y(_abc_40319_new_n2445_));
AND2X2 AND2X2_942 ( .A(_abc_40319_new_n1171_), .B(_abc_40319_new_n1724_), .Y(_abc_40319_new_n2446_));
AND2X2 AND2X2_943 ( .A(n1336), .B(REG3_REG_11_), .Y(_abc_40319_new_n2447_));
AND2X2 AND2X2_944 ( .A(_abc_40319_new_n1164_), .B(_abc_40319_new_n1732_), .Y(_abc_40319_new_n2450_));
AND2X2 AND2X2_945 ( .A(_abc_40319_new_n2049_), .B(_abc_40319_new_n1531_), .Y(_abc_40319_new_n2454_));
AND2X2 AND2X2_946 ( .A(_abc_40319_new_n2457_), .B(_abc_40319_new_n1122_), .Y(_abc_40319_new_n2458_));
AND2X2 AND2X2_947 ( .A(_abc_40319_new_n2458_), .B(_abc_40319_new_n2456_), .Y(_abc_40319_new_n2459_));
AND2X2 AND2X2_948 ( .A(_abc_40319_new_n1134_), .B(_abc_40319_new_n904_), .Y(_abc_40319_new_n2460_));
AND2X2 AND2X2_949 ( .A(_abc_40319_new_n1147_), .B(_abc_40319_new_n829_), .Y(_abc_40319_new_n2461_));
AND2X2 AND2X2_95 ( .A(_abc_40319_new_n524_), .B(IR_REG_29_), .Y(_abc_40319_new_n720_));
AND2X2 AND2X2_950 ( .A(_abc_40319_new_n2462_), .B(_abc_40319_new_n1133_), .Y(_abc_40319_new_n2463_));
AND2X2 AND2X2_951 ( .A(_abc_40319_new_n1164_), .B(REG3_REG_2_), .Y(_abc_40319_new_n2464_));
AND2X2 AND2X2_952 ( .A(_abc_40319_new_n1171_), .B(_abc_40319_new_n848_), .Y(_abc_40319_new_n2465_));
AND2X2 AND2X2_953 ( .A(n1336), .B(REG3_REG_2_), .Y(_abc_40319_new_n2466_));
AND2X2 AND2X2_954 ( .A(_abc_40319_new_n1919_), .B(_abc_40319_new_n1386_), .Y(_abc_40319_new_n2472_));
AND2X2 AND2X2_955 ( .A(_abc_40319_new_n2475_), .B(_abc_40319_new_n1122_), .Y(_abc_40319_new_n2476_));
AND2X2 AND2X2_956 ( .A(_abc_40319_new_n2476_), .B(_abc_40319_new_n2473_), .Y(_abc_40319_new_n2477_));
AND2X2 AND2X2_957 ( .A(_abc_40319_new_n1134_), .B(_abc_40319_new_n1444_), .Y(_abc_40319_new_n2478_));
AND2X2 AND2X2_958 ( .A(_abc_40319_new_n1147_), .B(_abc_40319_new_n1828_), .Y(_abc_40319_new_n2479_));
AND2X2 AND2X2_959 ( .A(_abc_40319_new_n2480_), .B(_abc_40319_new_n1133_), .Y(_abc_40319_new_n2481_));
AND2X2 AND2X2_96 ( .A(_abc_40319_new_n716_), .B(_abc_40319_new_n721_), .Y(_abc_40319_new_n722_));
AND2X2 AND2X2_960 ( .A(_abc_40319_new_n1164_), .B(_abc_40319_new_n1368_), .Y(_abc_40319_new_n2482_));
AND2X2 AND2X2_961 ( .A(_abc_40319_new_n1171_), .B(_abc_40319_new_n1363_), .Y(_abc_40319_new_n2483_));
AND2X2 AND2X2_962 ( .A(n1336), .B(REG3_REG_18_), .Y(_abc_40319_new_n2484_));
AND2X2 AND2X2_963 ( .A(_abc_40319_new_n1123_), .B(_abc_40319_new_n1021_), .Y(_abc_40319_new_n2490_));
AND2X2 AND2X2_964 ( .A(_abc_40319_new_n2493_), .B(_abc_40319_new_n1122_), .Y(_abc_40319_new_n2494_));
AND2X2 AND2X2_965 ( .A(_abc_40319_new_n2494_), .B(_abc_40319_new_n2492_), .Y(_abc_40319_new_n2495_));
AND2X2 AND2X2_966 ( .A(_abc_40319_new_n1134_), .B(_abc_40319_new_n746_), .Y(_abc_40319_new_n2496_));
AND2X2 AND2X2_967 ( .A(_abc_40319_new_n1147_), .B(_abc_40319_new_n1046_), .Y(_abc_40319_new_n2497_));
AND2X2 AND2X2_968 ( .A(_abc_40319_new_n2498_), .B(_abc_40319_new_n1133_), .Y(_abc_40319_new_n2499_));
AND2X2 AND2X2_969 ( .A(_abc_40319_new_n1164_), .B(_abc_40319_new_n1003_), .Y(_abc_40319_new_n2500_));
AND2X2 AND2X2_97 ( .A(_abc_40319_new_n722_), .B(REG1_REG_5_), .Y(_abc_40319_new_n723_));
AND2X2 AND2X2_970 ( .A(_abc_40319_new_n1171_), .B(_abc_40319_new_n998_), .Y(_abc_40319_new_n2501_));
AND2X2 AND2X2_971 ( .A(n1336), .B(REG3_REG_6_), .Y(_abc_40319_new_n2502_));
AND2X2 AND2X2_972 ( .A(_abc_40319_new_n2230_), .B(_abc_40319_new_n1301_), .Y(_abc_40319_new_n2508_));
AND2X2 AND2X2_973 ( .A(_abc_40319_new_n2227_), .B(_abc_40319_new_n1272_), .Y(_abc_40319_new_n2512_));
AND2X2 AND2X2_974 ( .A(_abc_40319_new_n1248_), .B(_abc_40319_new_n1300_), .Y(_abc_40319_new_n2514_));
AND2X2 AND2X2_975 ( .A(_abc_40319_new_n2516_), .B(_abc_40319_new_n1122_), .Y(_abc_40319_new_n2517_));
AND2X2 AND2X2_976 ( .A(_abc_40319_new_n2517_), .B(_abc_40319_new_n2511_), .Y(_abc_40319_new_n2518_));
AND2X2 AND2X2_977 ( .A(_abc_40319_new_n1260_), .B(_abc_40319_new_n1134_), .Y(_abc_40319_new_n2519_));
AND2X2 AND2X2_978 ( .A(_abc_40319_new_n1210_), .B(_abc_40319_new_n1147_), .Y(_abc_40319_new_n2520_));
AND2X2 AND2X2_979 ( .A(_abc_40319_new_n2521_), .B(_abc_40319_new_n1133_), .Y(_abc_40319_new_n2522_));
AND2X2 AND2X2_98 ( .A(_abc_40319_new_n725_), .B(_abc_40319_new_n726_), .Y(_abc_40319_new_n727_));
AND2X2 AND2X2_980 ( .A(_abc_40319_new_n1164_), .B(_abc_40319_new_n1228_), .Y(_abc_40319_new_n2523_));
AND2X2 AND2X2_981 ( .A(_abc_40319_new_n1171_), .B(_abc_40319_new_n1224_), .Y(_abc_40319_new_n2524_));
AND2X2 AND2X2_982 ( .A(n1336), .B(REG3_REG_26_), .Y(_abc_40319_new_n2525_));
AND2X2 AND2X2_983 ( .A(_abc_40319_new_n1922_), .B(_abc_40319_new_n1494_), .Y(_abc_40319_new_n2531_));
AND2X2 AND2X2_984 ( .A(_abc_40319_new_n2534_), .B(_abc_40319_new_n1122_), .Y(_abc_40319_new_n2535_));
AND2X2 AND2X2_985 ( .A(_abc_40319_new_n2535_), .B(_abc_40319_new_n2533_), .Y(_abc_40319_new_n2536_));
AND2X2 AND2X2_986 ( .A(_abc_40319_new_n1134_), .B(_abc_40319_new_n1517_), .Y(_abc_40319_new_n2537_));
AND2X2 AND2X2_987 ( .A(_abc_40319_new_n1147_), .B(_abc_40319_new_n1410_), .Y(_abc_40319_new_n2538_));
AND2X2 AND2X2_988 ( .A(_abc_40319_new_n2539_), .B(_abc_40319_new_n1133_), .Y(_abc_40319_new_n2540_));
AND2X2 AND2X2_989 ( .A(_abc_40319_new_n1171_), .B(_abc_40319_new_n1471_), .Y(_abc_40319_new_n2541_));
AND2X2 AND2X2_99 ( .A(_abc_40319_new_n728_), .B(_abc_40319_new_n724_), .Y(_abc_40319_new_n729_));
AND2X2 AND2X2_990 ( .A(n1336), .B(REG3_REG_15_), .Y(_abc_40319_new_n2542_));
AND2X2 AND2X2_991 ( .A(_abc_40319_new_n1164_), .B(_abc_40319_new_n1480_), .Y(_abc_40319_new_n2545_));
AND2X2 AND2X2_992 ( .A(_abc_40319_new_n2549_), .B(STATE_REG), .Y(_abc_40319_new_n2550_));
AND2X2 AND2X2_993 ( .A(_abc_40319_new_n671_), .B(_abc_40319_new_n646_), .Y(_abc_40319_new_n2551_));
AND2X2 AND2X2_994 ( .A(_abc_40319_new_n2551_), .B(_abc_40319_new_n2549_), .Y(_abc_40319_new_n2552_));
AND2X2 AND2X2_995 ( .A(_abc_40319_new_n817_), .B(DATAI_31_), .Y(_abc_40319_new_n2553_));
AND2X2 AND2X2_996 ( .A(_abc_40319_new_n2553_), .B(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2554_));
AND2X2 AND2X2_997 ( .A(_abc_40319_new_n736_), .B(REG0_REG_31_), .Y(_abc_40319_new_n2556_));
AND2X2 AND2X2_998 ( .A(_abc_40319_new_n733_), .B(REG2_REG_31_), .Y(_abc_40319_new_n2557_));
AND2X2 AND2X2_999 ( .A(_abc_40319_new_n722_), .B(REG1_REG_31_), .Y(_abc_40319_new_n2558_));
DFFPOSX1 DFFPOSX1_1 ( .CLK(clock), .D(n978), .Q(ADDR_REG_19_));
DFFPOSX1 DFFPOSX1_10 ( .CLK(clock), .D(n1014), .Q(ADDR_REG_10_));
DFFPOSX1 DFFPOSX1_100 ( .CLK(clock), .D(n403), .Q(D_REG_13_));
DFFPOSX1 DFFPOSX1_101 ( .CLK(clock), .D(n408), .Q(D_REG_14_));
DFFPOSX1 DFFPOSX1_102 ( .CLK(clock), .D(n413), .Q(D_REG_15_));
DFFPOSX1 DFFPOSX1_103 ( .CLK(clock), .D(n418), .Q(D_REG_16_));
DFFPOSX1 DFFPOSX1_104 ( .CLK(clock), .D(n423), .Q(D_REG_17_));
DFFPOSX1 DFFPOSX1_105 ( .CLK(clock), .D(n428), .Q(D_REG_18_));
DFFPOSX1 DFFPOSX1_106 ( .CLK(clock), .D(n433), .Q(D_REG_19_));
DFFPOSX1 DFFPOSX1_107 ( .CLK(clock), .D(n438), .Q(D_REG_20_));
DFFPOSX1 DFFPOSX1_108 ( .CLK(clock), .D(n443), .Q(D_REG_21_));
DFFPOSX1 DFFPOSX1_109 ( .CLK(clock), .D(n448), .Q(D_REG_22_));
DFFPOSX1 DFFPOSX1_11 ( .CLK(clock), .D(n1018), .Q(ADDR_REG_9_));
DFFPOSX1 DFFPOSX1_110 ( .CLK(clock), .D(n453), .Q(D_REG_23_));
DFFPOSX1 DFFPOSX1_111 ( .CLK(clock), .D(n458), .Q(D_REG_24_));
DFFPOSX1 DFFPOSX1_112 ( .CLK(clock), .D(n463), .Q(D_REG_25_));
DFFPOSX1 DFFPOSX1_113 ( .CLK(clock), .D(n468), .Q(D_REG_26_));
DFFPOSX1 DFFPOSX1_114 ( .CLK(clock), .D(n473), .Q(D_REG_27_));
DFFPOSX1 DFFPOSX1_115 ( .CLK(clock), .D(n478), .Q(D_REG_28_));
DFFPOSX1 DFFPOSX1_116 ( .CLK(clock), .D(n483), .Q(D_REG_29_));
DFFPOSX1 DFFPOSX1_117 ( .CLK(clock), .D(n488), .Q(D_REG_30_));
DFFPOSX1 DFFPOSX1_118 ( .CLK(clock), .D(n493), .Q(D_REG_31_));
DFFPOSX1 DFFPOSX1_119 ( .CLK(clock), .D(n498), .Q(REG0_REG_0_));
DFFPOSX1 DFFPOSX1_12 ( .CLK(clock), .D(n1022), .Q(ADDR_REG_8_));
DFFPOSX1 DFFPOSX1_120 ( .CLK(clock), .D(n503), .Q(REG0_REG_1_));
DFFPOSX1 DFFPOSX1_121 ( .CLK(clock), .D(n508), .Q(REG0_REG_2_));
DFFPOSX1 DFFPOSX1_122 ( .CLK(clock), .D(n513), .Q(REG0_REG_3_));
DFFPOSX1 DFFPOSX1_123 ( .CLK(clock), .D(n518), .Q(REG0_REG_4_));
DFFPOSX1 DFFPOSX1_124 ( .CLK(clock), .D(n523), .Q(REG0_REG_5_));
DFFPOSX1 DFFPOSX1_125 ( .CLK(clock), .D(n528), .Q(REG0_REG_6_));
DFFPOSX1 DFFPOSX1_126 ( .CLK(clock), .D(n533), .Q(REG0_REG_7_));
DFFPOSX1 DFFPOSX1_127 ( .CLK(clock), .D(n538), .Q(REG0_REG_8_));
DFFPOSX1 DFFPOSX1_128 ( .CLK(clock), .D(n543), .Q(REG0_REG_9_));
DFFPOSX1 DFFPOSX1_129 ( .CLK(clock), .D(n548), .Q(REG0_REG_10_));
DFFPOSX1 DFFPOSX1_13 ( .CLK(clock), .D(n1026), .Q(ADDR_REG_7_));
DFFPOSX1 DFFPOSX1_130 ( .CLK(clock), .D(n553), .Q(REG0_REG_11_));
DFFPOSX1 DFFPOSX1_131 ( .CLK(clock), .D(n558), .Q(REG0_REG_12_));
DFFPOSX1 DFFPOSX1_132 ( .CLK(clock), .D(n563), .Q(REG0_REG_13_));
DFFPOSX1 DFFPOSX1_133 ( .CLK(clock), .D(n568), .Q(REG0_REG_14_));
DFFPOSX1 DFFPOSX1_134 ( .CLK(clock), .D(n573), .Q(REG0_REG_15_));
DFFPOSX1 DFFPOSX1_135 ( .CLK(clock), .D(n578), .Q(REG0_REG_16_));
DFFPOSX1 DFFPOSX1_136 ( .CLK(clock), .D(n583), .Q(REG0_REG_17_));
DFFPOSX1 DFFPOSX1_137 ( .CLK(clock), .D(n588), .Q(REG0_REG_18_));
DFFPOSX1 DFFPOSX1_138 ( .CLK(clock), .D(n593), .Q(REG0_REG_19_));
DFFPOSX1 DFFPOSX1_139 ( .CLK(clock), .D(n598), .Q(REG0_REG_20_));
DFFPOSX1 DFFPOSX1_14 ( .CLK(clock), .D(n1030), .Q(ADDR_REG_6_));
DFFPOSX1 DFFPOSX1_140 ( .CLK(clock), .D(n603), .Q(REG0_REG_21_));
DFFPOSX1 DFFPOSX1_141 ( .CLK(clock), .D(n608), .Q(REG0_REG_22_));
DFFPOSX1 DFFPOSX1_142 ( .CLK(clock), .D(n613), .Q(REG0_REG_23_));
DFFPOSX1 DFFPOSX1_143 ( .CLK(clock), .D(n618), .Q(REG0_REG_24_));
DFFPOSX1 DFFPOSX1_144 ( .CLK(clock), .D(n623), .Q(REG0_REG_25_));
DFFPOSX1 DFFPOSX1_145 ( .CLK(clock), .D(n628), .Q(REG0_REG_26_));
DFFPOSX1 DFFPOSX1_146 ( .CLK(clock), .D(n633), .Q(REG0_REG_27_));
DFFPOSX1 DFFPOSX1_147 ( .CLK(clock), .D(n638), .Q(REG0_REG_28_));
DFFPOSX1 DFFPOSX1_148 ( .CLK(clock), .D(n643), .Q(REG0_REG_29_));
DFFPOSX1 DFFPOSX1_149 ( .CLK(clock), .D(n648), .Q(REG0_REG_30_));
DFFPOSX1 DFFPOSX1_15 ( .CLK(clock), .D(n1034), .Q(ADDR_REG_5_));
DFFPOSX1 DFFPOSX1_150 ( .CLK(clock), .D(n653), .Q(REG0_REG_31_));
DFFPOSX1 DFFPOSX1_151 ( .CLK(clock), .D(n658), .Q(REG1_REG_0_));
DFFPOSX1 DFFPOSX1_152 ( .CLK(clock), .D(n663), .Q(REG1_REG_1_));
DFFPOSX1 DFFPOSX1_153 ( .CLK(clock), .D(n668), .Q(REG1_REG_2_));
DFFPOSX1 DFFPOSX1_154 ( .CLK(clock), .D(n673), .Q(REG1_REG_3_));
DFFPOSX1 DFFPOSX1_155 ( .CLK(clock), .D(n678), .Q(REG1_REG_4_));
DFFPOSX1 DFFPOSX1_156 ( .CLK(clock), .D(n683), .Q(REG1_REG_5_));
DFFPOSX1 DFFPOSX1_157 ( .CLK(clock), .D(n688), .Q(REG1_REG_6_));
DFFPOSX1 DFFPOSX1_158 ( .CLK(clock), .D(n693), .Q(REG1_REG_7_));
DFFPOSX1 DFFPOSX1_159 ( .CLK(clock), .D(n698), .Q(REG1_REG_8_));
DFFPOSX1 DFFPOSX1_16 ( .CLK(clock), .D(n1038), .Q(ADDR_REG_4_));
DFFPOSX1 DFFPOSX1_160 ( .CLK(clock), .D(n703), .Q(REG1_REG_9_));
DFFPOSX1 DFFPOSX1_161 ( .CLK(clock), .D(n708), .Q(REG1_REG_10_));
DFFPOSX1 DFFPOSX1_162 ( .CLK(clock), .D(n713), .Q(REG1_REG_11_));
DFFPOSX1 DFFPOSX1_163 ( .CLK(clock), .D(n718), .Q(REG1_REG_12_));
DFFPOSX1 DFFPOSX1_164 ( .CLK(clock), .D(n723), .Q(REG1_REG_13_));
DFFPOSX1 DFFPOSX1_165 ( .CLK(clock), .D(n728), .Q(REG1_REG_14_));
DFFPOSX1 DFFPOSX1_166 ( .CLK(clock), .D(n733), .Q(REG1_REG_15_));
DFFPOSX1 DFFPOSX1_167 ( .CLK(clock), .D(n738), .Q(REG1_REG_16_));
DFFPOSX1 DFFPOSX1_168 ( .CLK(clock), .D(n743), .Q(REG1_REG_17_));
DFFPOSX1 DFFPOSX1_169 ( .CLK(clock), .D(n748), .Q(REG1_REG_18_));
DFFPOSX1 DFFPOSX1_17 ( .CLK(clock), .D(n1042), .Q(ADDR_REG_3_));
DFFPOSX1 DFFPOSX1_170 ( .CLK(clock), .D(n753), .Q(REG1_REG_19_));
DFFPOSX1 DFFPOSX1_171 ( .CLK(clock), .D(n758), .Q(REG1_REG_20_));
DFFPOSX1 DFFPOSX1_172 ( .CLK(clock), .D(n763), .Q(REG1_REG_21_));
DFFPOSX1 DFFPOSX1_173 ( .CLK(clock), .D(n768), .Q(REG1_REG_22_));
DFFPOSX1 DFFPOSX1_174 ( .CLK(clock), .D(n773), .Q(REG1_REG_23_));
DFFPOSX1 DFFPOSX1_175 ( .CLK(clock), .D(n778), .Q(REG1_REG_24_));
DFFPOSX1 DFFPOSX1_176 ( .CLK(clock), .D(n783), .Q(REG1_REG_25_));
DFFPOSX1 DFFPOSX1_177 ( .CLK(clock), .D(n788), .Q(REG1_REG_26_));
DFFPOSX1 DFFPOSX1_178 ( .CLK(clock), .D(n793), .Q(REG1_REG_27_));
DFFPOSX1 DFFPOSX1_179 ( .CLK(clock), .D(n798), .Q(REG1_REG_28_));
DFFPOSX1 DFFPOSX1_18 ( .CLK(clock), .D(n1046), .Q(ADDR_REG_2_));
DFFPOSX1 DFFPOSX1_180 ( .CLK(clock), .D(n803), .Q(REG1_REG_29_));
DFFPOSX1 DFFPOSX1_181 ( .CLK(clock), .D(n808), .Q(REG1_REG_30_));
DFFPOSX1 DFFPOSX1_182 ( .CLK(clock), .D(n813), .Q(REG1_REG_31_));
DFFPOSX1 DFFPOSX1_183 ( .CLK(clock), .D(n818), .Q(REG2_REG_0_));
DFFPOSX1 DFFPOSX1_184 ( .CLK(clock), .D(n823), .Q(REG2_REG_1_));
DFFPOSX1 DFFPOSX1_185 ( .CLK(clock), .D(n828), .Q(REG2_REG_2_));
DFFPOSX1 DFFPOSX1_186 ( .CLK(clock), .D(n833), .Q(REG2_REG_3_));
DFFPOSX1 DFFPOSX1_187 ( .CLK(clock), .D(n838), .Q(REG2_REG_4_));
DFFPOSX1 DFFPOSX1_188 ( .CLK(clock), .D(n843), .Q(REG2_REG_5_));
DFFPOSX1 DFFPOSX1_189 ( .CLK(clock), .D(n848), .Q(REG2_REG_6_));
DFFPOSX1 DFFPOSX1_19 ( .CLK(clock), .D(n1050), .Q(ADDR_REG_1_));
DFFPOSX1 DFFPOSX1_190 ( .CLK(clock), .D(n853), .Q(REG2_REG_7_));
DFFPOSX1 DFFPOSX1_191 ( .CLK(clock), .D(n858), .Q(REG2_REG_8_));
DFFPOSX1 DFFPOSX1_192 ( .CLK(clock), .D(n863), .Q(REG2_REG_9_));
DFFPOSX1 DFFPOSX1_193 ( .CLK(clock), .D(n868), .Q(REG2_REG_10_));
DFFPOSX1 DFFPOSX1_194 ( .CLK(clock), .D(n873), .Q(REG2_REG_11_));
DFFPOSX1 DFFPOSX1_195 ( .CLK(clock), .D(n878), .Q(REG2_REG_12_));
DFFPOSX1 DFFPOSX1_196 ( .CLK(clock), .D(n883), .Q(REG2_REG_13_));
DFFPOSX1 DFFPOSX1_197 ( .CLK(clock), .D(n888), .Q(REG2_REG_14_));
DFFPOSX1 DFFPOSX1_198 ( .CLK(clock), .D(n893), .Q(REG2_REG_15_));
DFFPOSX1 DFFPOSX1_199 ( .CLK(clock), .D(n898), .Q(REG2_REG_16_));
DFFPOSX1 DFFPOSX1_2 ( .CLK(clock), .D(n986), .Q(ADDR_REG_17_));
DFFPOSX1 DFFPOSX1_20 ( .CLK(clock), .D(n1054), .Q(ADDR_REG_0_));
DFFPOSX1 DFFPOSX1_200 ( .CLK(clock), .D(n903), .Q(REG2_REG_17_));
DFFPOSX1 DFFPOSX1_201 ( .CLK(clock), .D(n908), .Q(REG2_REG_18_));
DFFPOSX1 DFFPOSX1_202 ( .CLK(clock), .D(n913), .Q(REG2_REG_19_));
DFFPOSX1 DFFPOSX1_203 ( .CLK(clock), .D(n918), .Q(REG2_REG_20_));
DFFPOSX1 DFFPOSX1_204 ( .CLK(clock), .D(n923), .Q(REG2_REG_21_));
DFFPOSX1 DFFPOSX1_205 ( .CLK(clock), .D(n928), .Q(REG2_REG_22_));
DFFPOSX1 DFFPOSX1_206 ( .CLK(clock), .D(n933), .Q(REG2_REG_23_));
DFFPOSX1 DFFPOSX1_207 ( .CLK(clock), .D(n938), .Q(REG2_REG_24_));
DFFPOSX1 DFFPOSX1_208 ( .CLK(clock), .D(n943), .Q(REG2_REG_25_));
DFFPOSX1 DFFPOSX1_209 ( .CLK(clock), .D(n948), .Q(REG2_REG_26_));
DFFPOSX1 DFFPOSX1_21 ( .CLK(clock), .D(n1182), .Q(DATAO_REG_31_));
DFFPOSX1 DFFPOSX1_210 ( .CLK(clock), .D(n953), .Q(REG2_REG_27_));
DFFPOSX1 DFFPOSX1_211 ( .CLK(clock), .D(n958), .Q(REG2_REG_28_));
DFFPOSX1 DFFPOSX1_212 ( .CLK(clock), .D(n963), .Q(REG2_REG_29_));
DFFPOSX1 DFFPOSX1_213 ( .CLK(clock), .D(n968), .Q(REG2_REG_30_));
DFFPOSX1 DFFPOSX1_214 ( .CLK(clock), .D(n973), .Q(REG2_REG_31_));
DFFPOSX1 DFFPOSX1_215 ( .CLK(clock), .D(n1186), .Q(B_REG));
DFFPOSX1 DFFPOSX1_216 ( .CLK(clock), .D(n1191), .Q(REG3_REG_15_));
DFFPOSX1 DFFPOSX1_217 ( .CLK(clock), .D(n1196), .Q(REG3_REG_26_));
DFFPOSX1 DFFPOSX1_218 ( .CLK(clock), .D(n1201), .Q(REG3_REG_6_));
DFFPOSX1 DFFPOSX1_219 ( .CLK(clock), .D(n1206), .Q(REG3_REG_18_));
DFFPOSX1 DFFPOSX1_22 ( .CLK(clock), .D(n1178), .Q(DATAO_REG_30_));
DFFPOSX1 DFFPOSX1_220 ( .CLK(clock), .D(n1211), .Q(REG3_REG_2_));
DFFPOSX1 DFFPOSX1_221 ( .CLK(clock), .D(n1216), .Q(REG3_REG_11_));
DFFPOSX1 DFFPOSX1_222 ( .CLK(clock), .D(n1221), .Q(REG3_REG_22_));
DFFPOSX1 DFFPOSX1_223 ( .CLK(clock), .D(n1226), .Q(REG3_REG_13_));
DFFPOSX1 DFFPOSX1_224 ( .CLK(clock), .D(n1231), .Q(REG3_REG_20_));
DFFPOSX1 DFFPOSX1_225 ( .CLK(clock), .D(n1236), .Q(REG3_REG_0_));
DFFPOSX1 DFFPOSX1_226 ( .CLK(clock), .D(n1241), .Q(REG3_REG_9_));
DFFPOSX1 DFFPOSX1_227 ( .CLK(clock), .D(n1246), .Q(REG3_REG_4_));
DFFPOSX1 DFFPOSX1_228 ( .CLK(clock), .D(n1251), .Q(REG3_REG_24_));
DFFPOSX1 DFFPOSX1_229 ( .CLK(clock), .D(n1256), .Q(REG3_REG_17_));
DFFPOSX1 DFFPOSX1_23 ( .CLK(clock), .D(n1174), .Q(DATAO_REG_29_));
DFFPOSX1 DFFPOSX1_230 ( .CLK(clock), .D(n1261), .Q(REG3_REG_5_));
DFFPOSX1 DFFPOSX1_231 ( .CLK(clock), .D(n1266), .Q(REG3_REG_16_));
DFFPOSX1 DFFPOSX1_232 ( .CLK(clock), .D(n1271), .Q(REG3_REG_25_));
DFFPOSX1 DFFPOSX1_233 ( .CLK(clock), .D(n1276), .Q(REG3_REG_12_));
DFFPOSX1 DFFPOSX1_234 ( .CLK(clock), .D(n1281), .Q(REG3_REG_21_));
DFFPOSX1 DFFPOSX1_235 ( .CLK(clock), .D(n1286), .Q(REG3_REG_1_));
DFFPOSX1 DFFPOSX1_236 ( .CLK(clock), .D(n1291), .Q(REG3_REG_8_));
DFFPOSX1 DFFPOSX1_237 ( .CLK(clock), .D(n1296), .Q(REG3_REG_28_));
DFFPOSX1 DFFPOSX1_238 ( .CLK(clock), .D(n1301), .Q(REG3_REG_19_));
DFFPOSX1 DFFPOSX1_239 ( .CLK(clock), .D(n1306), .Q(REG3_REG_3_));
DFFPOSX1 DFFPOSX1_24 ( .CLK(clock), .D(n1170), .Q(DATAO_REG_28_));
DFFPOSX1 DFFPOSX1_240 ( .CLK(clock), .D(n1311), .Q(REG3_REG_10_));
DFFPOSX1 DFFPOSX1_241 ( .CLK(clock), .D(n1316), .Q(REG3_REG_23_));
DFFPOSX1 DFFPOSX1_242 ( .CLK(clock), .D(n1321), .Q(REG3_REG_14_));
DFFPOSX1 DFFPOSX1_243 ( .CLK(clock), .D(n1326), .Q(REG3_REG_27_));
DFFPOSX1 DFFPOSX1_244 ( .CLK(clock), .D(n1331), .Q(REG3_REG_7_));
DFFPOSX1 DFFPOSX1_245 ( .CLK(clock), .D(n1336), .Q(STATE_REG));
DFFPOSX1 DFFPOSX1_25 ( .CLK(clock), .D(n1166), .Q(DATAO_REG_27_));
DFFPOSX1 DFFPOSX1_26 ( .CLK(clock), .D(n1162), .Q(DATAO_REG_26_));
DFFPOSX1 DFFPOSX1_27 ( .CLK(clock), .D(n1158), .Q(DATAO_REG_25_));
DFFPOSX1 DFFPOSX1_28 ( .CLK(clock), .D(n1154), .Q(DATAO_REG_24_));
DFFPOSX1 DFFPOSX1_29 ( .CLK(clock), .D(n1150), .Q(DATAO_REG_23_));
DFFPOSX1 DFFPOSX1_3 ( .CLK(clock), .D(n998), .Q(ADDR_REG_14_));
DFFPOSX1 DFFPOSX1_30 ( .CLK(clock), .D(n1146), .Q(DATAO_REG_22_));
DFFPOSX1 DFFPOSX1_31 ( .CLK(clock), .D(n1142), .Q(DATAO_REG_21_));
DFFPOSX1 DFFPOSX1_32 ( .CLK(clock), .D(n1138), .Q(DATAO_REG_20_));
DFFPOSX1 DFFPOSX1_33 ( .CLK(clock), .D(n1134), .Q(DATAO_REG_19_));
DFFPOSX1 DFFPOSX1_34 ( .CLK(clock), .D(n1130), .Q(DATAO_REG_18_));
DFFPOSX1 DFFPOSX1_35 ( .CLK(clock), .D(n1126), .Q(DATAO_REG_17_));
DFFPOSX1 DFFPOSX1_36 ( .CLK(clock), .D(n1122), .Q(DATAO_REG_16_));
DFFPOSX1 DFFPOSX1_37 ( .CLK(clock), .D(n1118), .Q(DATAO_REG_15_));
DFFPOSX1 DFFPOSX1_38 ( .CLK(clock), .D(n1114), .Q(DATAO_REG_14_));
DFFPOSX1 DFFPOSX1_39 ( .CLK(clock), .D(n1110), .Q(DATAO_REG_13_));
DFFPOSX1 DFFPOSX1_4 ( .CLK(clock), .D(n990), .Q(ADDR_REG_16_));
DFFPOSX1 DFFPOSX1_40 ( .CLK(clock), .D(n1106), .Q(DATAO_REG_12_));
DFFPOSX1 DFFPOSX1_41 ( .CLK(clock), .D(n1102), .Q(DATAO_REG_11_));
DFFPOSX1 DFFPOSX1_42 ( .CLK(clock), .D(n1098), .Q(DATAO_REG_10_));
DFFPOSX1 DFFPOSX1_43 ( .CLK(clock), .D(n1094), .Q(DATAO_REG_9_));
DFFPOSX1 DFFPOSX1_44 ( .CLK(clock), .D(n1090), .Q(DATAO_REG_8_));
DFFPOSX1 DFFPOSX1_45 ( .CLK(clock), .D(n1086), .Q(DATAO_REG_7_));
DFFPOSX1 DFFPOSX1_46 ( .CLK(clock), .D(n1082), .Q(DATAO_REG_6_));
DFFPOSX1 DFFPOSX1_47 ( .CLK(clock), .D(n1078), .Q(DATAO_REG_5_));
DFFPOSX1 DFFPOSX1_48 ( .CLK(clock), .D(n1074), .Q(DATAO_REG_4_));
DFFPOSX1 DFFPOSX1_49 ( .CLK(clock), .D(n1070), .Q(DATAO_REG_3_));
DFFPOSX1 DFFPOSX1_5 ( .CLK(clock), .D(n994), .Q(ADDR_REG_15_));
DFFPOSX1 DFFPOSX1_50 ( .CLK(clock), .D(n1066), .Q(DATAO_REG_2_));
DFFPOSX1 DFFPOSX1_51 ( .CLK(clock), .D(n1062), .Q(DATAO_REG_1_));
DFFPOSX1 DFFPOSX1_52 ( .CLK(clock), .D(n1058), .Q(DATAO_REG_0_));
DFFPOSX1 DFFPOSX1_53 ( .CLK(clock), .D(n1341), .Q(RD_REG));
DFFPOSX1 DFFPOSX1_54 ( .CLK(clock), .D(n1345), .Q(WR_REG));
DFFPOSX1 DFFPOSX1_55 ( .CLK(clock), .D(n178), .Q(IR_REG_0_));
DFFPOSX1 DFFPOSX1_56 ( .CLK(clock), .D(n183), .Q(IR_REG_1_));
DFFPOSX1 DFFPOSX1_57 ( .CLK(clock), .D(n188), .Q(IR_REG_2_));
DFFPOSX1 DFFPOSX1_58 ( .CLK(clock), .D(n193), .Q(IR_REG_3_));
DFFPOSX1 DFFPOSX1_59 ( .CLK(clock), .D(n198), .Q(IR_REG_4_));
DFFPOSX1 DFFPOSX1_6 ( .CLK(clock), .D(n982), .Q(ADDR_REG_18_));
DFFPOSX1 DFFPOSX1_60 ( .CLK(clock), .D(n203), .Q(IR_REG_5_));
DFFPOSX1 DFFPOSX1_61 ( .CLK(clock), .D(n208), .Q(IR_REG_6_));
DFFPOSX1 DFFPOSX1_62 ( .CLK(clock), .D(n213), .Q(IR_REG_7_));
DFFPOSX1 DFFPOSX1_63 ( .CLK(clock), .D(n218), .Q(IR_REG_8_));
DFFPOSX1 DFFPOSX1_64 ( .CLK(clock), .D(n223), .Q(IR_REG_9_));
DFFPOSX1 DFFPOSX1_65 ( .CLK(clock), .D(n228), .Q(IR_REG_10_));
DFFPOSX1 DFFPOSX1_66 ( .CLK(clock), .D(n233), .Q(IR_REG_11_));
DFFPOSX1 DFFPOSX1_67 ( .CLK(clock), .D(n238), .Q(IR_REG_12_));
DFFPOSX1 DFFPOSX1_68 ( .CLK(clock), .D(n243), .Q(IR_REG_13_));
DFFPOSX1 DFFPOSX1_69 ( .CLK(clock), .D(n248), .Q(IR_REG_14_));
DFFPOSX1 DFFPOSX1_7 ( .CLK(clock), .D(n1002), .Q(ADDR_REG_13_));
DFFPOSX1 DFFPOSX1_70 ( .CLK(clock), .D(n253), .Q(IR_REG_15_));
DFFPOSX1 DFFPOSX1_71 ( .CLK(clock), .D(n258), .Q(IR_REG_16_));
DFFPOSX1 DFFPOSX1_72 ( .CLK(clock), .D(n263), .Q(IR_REG_17_));
DFFPOSX1 DFFPOSX1_73 ( .CLK(clock), .D(n268), .Q(IR_REG_18_));
DFFPOSX1 DFFPOSX1_74 ( .CLK(clock), .D(n273), .Q(IR_REG_19_));
DFFPOSX1 DFFPOSX1_75 ( .CLK(clock), .D(n278), .Q(IR_REG_20_));
DFFPOSX1 DFFPOSX1_76 ( .CLK(clock), .D(n283), .Q(IR_REG_21_));
DFFPOSX1 DFFPOSX1_77 ( .CLK(clock), .D(n288), .Q(IR_REG_22_));
DFFPOSX1 DFFPOSX1_78 ( .CLK(clock), .D(n293), .Q(IR_REG_23_));
DFFPOSX1 DFFPOSX1_79 ( .CLK(clock), .D(n298), .Q(IR_REG_24_));
DFFPOSX1 DFFPOSX1_8 ( .CLK(clock), .D(n1006), .Q(ADDR_REG_12_));
DFFPOSX1 DFFPOSX1_80 ( .CLK(clock), .D(n303), .Q(IR_REG_25_));
DFFPOSX1 DFFPOSX1_81 ( .CLK(clock), .D(n308), .Q(IR_REG_26_));
DFFPOSX1 DFFPOSX1_82 ( .CLK(clock), .D(n313), .Q(IR_REG_27_));
DFFPOSX1 DFFPOSX1_83 ( .CLK(clock), .D(n318), .Q(IR_REG_28_));
DFFPOSX1 DFFPOSX1_84 ( .CLK(clock), .D(n323), .Q(IR_REG_29_));
DFFPOSX1 DFFPOSX1_85 ( .CLK(clock), .D(n328), .Q(IR_REG_30_));
DFFPOSX1 DFFPOSX1_86 ( .CLK(clock), .D(n333), .Q(IR_REG_31_));
DFFPOSX1 DFFPOSX1_87 ( .CLK(clock), .D(n338), .Q(D_REG_0_));
DFFPOSX1 DFFPOSX1_88 ( .CLK(clock), .D(n343), .Q(D_REG_1_));
DFFPOSX1 DFFPOSX1_89 ( .CLK(clock), .D(n348), .Q(D_REG_2_));
DFFPOSX1 DFFPOSX1_9 ( .CLK(clock), .D(n1010), .Q(ADDR_REG_11_));
DFFPOSX1 DFFPOSX1_90 ( .CLK(clock), .D(n353), .Q(D_REG_3_));
DFFPOSX1 DFFPOSX1_91 ( .CLK(clock), .D(n358), .Q(D_REG_4_));
DFFPOSX1 DFFPOSX1_92 ( .CLK(clock), .D(n363), .Q(D_REG_5_));
DFFPOSX1 DFFPOSX1_93 ( .CLK(clock), .D(n368), .Q(D_REG_6_));
DFFPOSX1 DFFPOSX1_94 ( .CLK(clock), .D(n373), .Q(D_REG_7_));
DFFPOSX1 DFFPOSX1_95 ( .CLK(clock), .D(n378), .Q(D_REG_8_));
DFFPOSX1 DFFPOSX1_96 ( .CLK(clock), .D(n383), .Q(D_REG_9_));
DFFPOSX1 DFFPOSX1_97 ( .CLK(clock), .D(n388), .Q(D_REG_10_));
DFFPOSX1 DFFPOSX1_98 ( .CLK(clock), .D(n393), .Q(D_REG_11_));
DFFPOSX1 DFFPOSX1_99 ( .CLK(clock), .D(n398), .Q(D_REG_12_));
INVX1 INVX1_1 ( .A(RESET_G), .Y(_abc_40319_new_n523_));
INVX1 INVX1_10 ( .A(IR_REG_12_), .Y(_abc_40319_new_n538_));
INVX1 INVX1_100 ( .A(DATAI_1_), .Y(_abc_40319_new_n888_));
INVX1 INVX1_101 ( .A(_abc_40319_new_n889_), .Y(_abc_40319_new_n890_));
INVX1 INVX1_102 ( .A(_abc_40319_new_n893_), .Y(_abc_40319_new_n894_));
INVX1 INVX1_103 ( .A(_abc_40319_new_n895_), .Y(_abc_40319_new_n896_));
INVX1 INVX1_104 ( .A(_abc_40319_new_n898_), .Y(_abc_40319_new_n899_));
INVX1 INVX1_105 ( .A(_abc_40319_new_n900_), .Y(_abc_40319_new_n901_));
INVX1 INVX1_106 ( .A(_abc_40319_new_n903_), .Y(_abc_40319_new_n904_));
INVX1 INVX1_107 ( .A(_abc_40319_new_n907_), .Y(_abc_40319_new_n908_));
INVX1 INVX1_108 ( .A(_abc_40319_new_n673_), .Y(_abc_40319_new_n909_));
INVX1 INVX1_109 ( .A(_abc_40319_new_n911_), .Y(_abc_40319_new_n912_));
INVX1 INVX1_11 ( .A(IR_REG_11_), .Y(_abc_40319_new_n539_));
INVX1 INVX1_110 ( .A(DATAI_0_), .Y(_abc_40319_new_n927_));
INVX1 INVX1_111 ( .A(_abc_40319_new_n928_), .Y(_abc_40319_new_n929_));
INVX1 INVX1_112 ( .A(_abc_40319_new_n758_), .Y(_abc_40319_new_n937_));
INVX1 INVX1_113 ( .A(IR_REG_0_), .Y(_abc_40319_new_n940_));
INVX1 INVX1_114 ( .A(REG2_REG_0_), .Y(_abc_40319_new_n944_));
INVX1 INVX1_115 ( .A(REG0_REG_0_), .Y(_abc_40319_new_n946_));
INVX1 INVX1_116 ( .A(REG3_REG_0_), .Y(_abc_40319_new_n949_));
INVX1 INVX1_117 ( .A(REG1_REG_0_), .Y(_abc_40319_new_n951_));
INVX1 INVX1_118 ( .A(_abc_40319_new_n835_), .Y(_abc_40319_new_n969_));
INVX1 INVX1_119 ( .A(_abc_40319_new_n838_), .Y(_abc_40319_new_n970_));
INVX1 INVX1_12 ( .A(IR_REG_13_), .Y(_abc_40319_new_n541_));
INVX1 INVX1_120 ( .A(_abc_40319_new_n867_), .Y(_abc_40319_new_n972_));
INVX1 INVX1_121 ( .A(_abc_40319_new_n977_), .Y(_abc_40319_new_n978_));
INVX1 INVX1_122 ( .A(_abc_40319_new_n984_), .Y(_abc_40319_new_n985_));
INVX1 INVX1_123 ( .A(_abc_40319_new_n537_), .Y(_abc_40319_new_n987_));
INVX1 INVX1_124 ( .A(_abc_40319_new_n989_), .Y(_abc_40319_new_n990_));
INVX1 INVX1_125 ( .A(_abc_40319_new_n993_), .Y(_abc_40319_new_n994_));
INVX1 INVX1_126 ( .A(_abc_40319_new_n995_), .Y(_abc_40319_new_n996_));
INVX1 INVX1_127 ( .A(_abc_40319_new_n1000_), .Y(_abc_40319_new_n1001_));
INVX1 INVX1_128 ( .A(_abc_40319_new_n1012_), .Y(_abc_40319_new_n1013_));
INVX1 INVX1_129 ( .A(_abc_40319_new_n1016_), .Y(_abc_40319_new_n1018_));
INVX1 INVX1_13 ( .A(IR_REG_10_), .Y(_abc_40319_new_n542_));
INVX1 INVX1_130 ( .A(_abc_40319_new_n1023_), .Y(_abc_40319_new_n1024_));
INVX1 INVX1_131 ( .A(_abc_40319_new_n1029_), .Y(_abc_40319_new_n1030_));
INVX1 INVX1_132 ( .A(_abc_40319_new_n1031_), .Y(_abc_40319_new_n1032_));
INVX1 INVX1_133 ( .A(_abc_40319_new_n1039_), .Y(_abc_40319_new_n1040_));
INVX1 INVX1_134 ( .A(_abc_40319_new_n1048_), .Y(_abc_40319_new_n1049_));
INVX1 INVX1_135 ( .A(_abc_40319_new_n1052_), .Y(_abc_40319_new_n1054_));
INVX1 INVX1_136 ( .A(_abc_40319_new_n1057_), .Y(_abc_40319_new_n1058_));
INVX1 INVX1_137 ( .A(_abc_40319_new_n589_), .Y(_abc_40319_new_n1064_));
INVX1 INVX1_138 ( .A(_abc_40319_new_n596_), .Y(_abc_40319_new_n1065_));
INVX1 INVX1_139 ( .A(_abc_40319_new_n582_), .Y(_abc_40319_new_n1068_));
INVX1 INVX1_14 ( .A(IR_REG_9_), .Y(_abc_40319_new_n545_));
INVX1 INVX1_140 ( .A(B_REG), .Y(_abc_40319_new_n1069_));
INVX1 INVX1_141 ( .A(_abc_40319_new_n1074_), .Y(_abc_40319_new_n1075_));
INVX1 INVX1_142 ( .A(_abc_40319_new_n1072_), .Y(_abc_40319_new_n1077_));
INVX1 INVX1_143 ( .A(_abc_40319_new_n1107_), .Y(_abc_40319_new_n1108_));
INVX1 INVX1_144 ( .A(_abc_40319_new_n1110_), .Y(_abc_40319_new_n1111_));
INVX1 INVX1_145 ( .A(_abc_40319_new_n656_), .Y(_abc_40319_new_n1115_));
INVX1 INVX1_146 ( .A(_abc_40319_new_n1059_), .Y(_abc_40319_new_n1123_));
INVX1 INVX1_147 ( .A(_abc_40319_new_n1021_), .Y(_abc_40319_new_n1125_));
INVX1 INVX1_148 ( .A(_abc_40319_new_n1060_), .Y(_abc_40319_new_n1126_));
INVX1 INVX1_149 ( .A(_abc_40319_new_n1137_), .Y(_abc_40319_new_n1138_));
INVX1 INVX1_15 ( .A(IR_REG_8_), .Y(_abc_40319_new_n546_));
INVX1 INVX1_150 ( .A(_abc_40319_new_n1114_), .Y(_abc_40319_new_n1151_));
INVX1 INVX1_151 ( .A(_abc_40319_new_n1119_), .Y(_abc_40319_new_n1157_));
INVX1 INVX1_152 ( .A(_abc_40319_new_n1116_), .Y(_abc_40319_new_n1158_));
INVX1 INVX1_153 ( .A(nRESET_G), .Y(_abc_40319_new_n1173_));
INVX1 INVX1_154 ( .A(_abc_40319_new_n1201_), .Y(_abc_40319_new_n1202_));
INVX1 INVX1_155 ( .A(_abc_40319_new_n1215_), .Y(_abc_40319_new_n1216_));
INVX1 INVX1_156 ( .A(_abc_40319_new_n1220_), .Y(_abc_40319_new_n1221_));
INVX1 INVX1_157 ( .A(_abc_40319_new_n1199_), .Y(_abc_40319_new_n1226_));
INVX1 INVX1_158 ( .A(_abc_40319_new_n1237_), .Y(_abc_40319_new_n1238_));
INVX1 INVX1_159 ( .A(_abc_40319_new_n1241_), .Y(_abc_40319_new_n1242_));
INVX1 INVX1_16 ( .A(IR_REG_7_), .Y(_abc_40319_new_n548_));
INVX1 INVX1_160 ( .A(_abc_40319_new_n1245_), .Y(_abc_40319_new_n1246_));
INVX1 INVX1_161 ( .A(_abc_40319_new_n1247_), .Y(_abc_40319_new_n1248_));
INVX1 INVX1_162 ( .A(_abc_40319_new_n1198_), .Y(_abc_40319_new_n1251_));
INVX1 INVX1_163 ( .A(_abc_40319_new_n1262_), .Y(_abc_40319_new_n1263_));
INVX1 INVX1_164 ( .A(_abc_40319_new_n1266_), .Y(_abc_40319_new_n1267_));
INVX1 INVX1_165 ( .A(_abc_40319_new_n1271_), .Y(_abc_40319_new_n1272_));
INVX1 INVX1_166 ( .A(_abc_40319_new_n1197_), .Y(_abc_40319_new_n1276_));
INVX1 INVX1_167 ( .A(_abc_40319_new_n1290_), .Y(_abc_40319_new_n1291_));
INVX1 INVX1_168 ( .A(_abc_40319_new_n1294_), .Y(_abc_40319_new_n1295_));
INVX1 INVX1_169 ( .A(_abc_40319_new_n1297_), .Y(_abc_40319_new_n1298_));
INVX1 INVX1_17 ( .A(IR_REG_6_), .Y(_abc_40319_new_n549_));
INVX1 INVX1_170 ( .A(_abc_40319_new_n1299_), .Y(_abc_40319_new_n1300_));
INVX1 INVX1_171 ( .A(_abc_40319_new_n1304_), .Y(_abc_40319_new_n1305_));
INVX1 INVX1_172 ( .A(_abc_40319_new_n1196_), .Y(_abc_40319_new_n1308_));
INVX1 INVX1_173 ( .A(_abc_40319_new_n1322_), .Y(_abc_40319_new_n1324_));
INVX1 INVX1_174 ( .A(_abc_40319_new_n1195_), .Y(_abc_40319_new_n1331_));
INVX1 INVX1_175 ( .A(_abc_40319_new_n1345_), .Y(_abc_40319_new_n1346_));
INVX1 INVX1_176 ( .A(_abc_40319_new_n1349_), .Y(_abc_40319_new_n1350_));
INVX1 INVX1_177 ( .A(_abc_40319_new_n1354_), .Y(_abc_40319_new_n1355_));
INVX1 INVX1_178 ( .A(_abc_40319_new_n1358_), .Y(_abc_40319_new_n1359_));
INVX1 INVX1_179 ( .A(_abc_40319_new_n1360_), .Y(_abc_40319_new_n1361_));
INVX1 INVX1_18 ( .A(IR_REG_22_), .Y(_abc_40319_new_n554_));
INVX1 INVX1_180 ( .A(_abc_40319_new_n1191_), .Y(_abc_40319_new_n1366_));
INVX1 INVX1_181 ( .A(_abc_40319_new_n1379_), .Y(_abc_40319_new_n1380_));
INVX1 INVX1_182 ( .A(_abc_40319_new_n1383_), .Y(_abc_40319_new_n1384_));
INVX1 INVX1_183 ( .A(_abc_40319_new_n1389_), .Y(_abc_40319_new_n1390_));
INVX1 INVX1_184 ( .A(_abc_40319_new_n1395_), .Y(_abc_40319_new_n1396_));
INVX1 INVX1_185 ( .A(_abc_40319_new_n1404_), .Y(_abc_40319_new_n1405_));
INVX1 INVX1_186 ( .A(_abc_40319_new_n1412_), .Y(_abc_40319_new_n1413_));
INVX1 INVX1_187 ( .A(_abc_40319_new_n1416_), .Y(_abc_40319_new_n1418_));
INVX1 INVX1_188 ( .A(_abc_40319_new_n1420_), .Y(_abc_40319_new_n1421_));
INVX1 INVX1_189 ( .A(_abc_40319_new_n1422_), .Y(_abc_40319_new_n1423_));
INVX1 INVX1_19 ( .A(IR_REG_17_), .Y(_abc_40319_new_n555_));
INVX1 INVX1_190 ( .A(_abc_40319_new_n1428_), .Y(_abc_40319_new_n1429_));
INVX1 INVX1_191 ( .A(_abc_40319_new_n1430_), .Y(_abc_40319_new_n1431_));
INVX1 INVX1_192 ( .A(_abc_40319_new_n1190_), .Y(_abc_40319_new_n1438_));
INVX1 INVX1_193 ( .A(_abc_40319_new_n1446_), .Y(_abc_40319_new_n1447_));
INVX1 INVX1_194 ( .A(_abc_40319_new_n1450_), .Y(_abc_40319_new_n1452_));
INVX1 INVX1_195 ( .A(_abc_40319_new_n1454_), .Y(_abc_40319_new_n1455_));
INVX1 INVX1_196 ( .A(_abc_40319_new_n1456_), .Y(_abc_40319_new_n1457_));
INVX1 INVX1_197 ( .A(_abc_40319_new_n1459_), .Y(_abc_40319_new_n1460_));
INVX1 INVX1_198 ( .A(_abc_40319_new_n1462_), .Y(_abc_40319_new_n1463_));
INVX1 INVX1_199 ( .A(_abc_40319_new_n1466_), .Y(_abc_40319_new_n1467_));
INVX1 INVX1_2 ( .A(IR_REG_31_), .Y(_abc_40319_new_n524_));
INVX1 INVX1_20 ( .A(IR_REG_16_), .Y(_abc_40319_new_n556_));
INVX1 INVX1_200 ( .A(_abc_40319_new_n1468_), .Y(_abc_40319_new_n1469_));
INVX1 INVX1_201 ( .A(_abc_40319_new_n1188_), .Y(_abc_40319_new_n1477_));
INVX1 INVX1_202 ( .A(_abc_40319_new_n1488_), .Y(_abc_40319_new_n1490_));
INVX1 INVX1_203 ( .A(_abc_40319_new_n553_), .Y(_abc_40319_new_n1495_));
INVX1 INVX1_204 ( .A(_abc_40319_new_n1497_), .Y(_abc_40319_new_n1498_));
INVX1 INVX1_205 ( .A(_abc_40319_new_n1501_), .Y(_abc_40319_new_n1502_));
INVX1 INVX1_206 ( .A(_abc_40319_new_n1503_), .Y(_abc_40319_new_n1504_));
INVX1 INVX1_207 ( .A(_abc_40319_new_n1478_), .Y(_abc_40319_new_n1511_));
INVX1 INVX1_208 ( .A(_abc_40319_new_n1522_), .Y(_abc_40319_new_n1524_));
INVX1 INVX1_209 ( .A(_abc_40319_new_n806_), .Y(_abc_40319_new_n1529_));
INVX1 INVX1_21 ( .A(IR_REG_15_), .Y(_abc_40319_new_n557_));
INVX1 INVX1_210 ( .A(_abc_40319_new_n807_), .Y(_abc_40319_new_n1530_));
INVX1 INVX1_211 ( .A(_abc_40319_new_n880_), .Y(_abc_40319_new_n1534_));
INVX1 INVX1_212 ( .A(_abc_40319_new_n917_), .Y(_abc_40319_new_n1536_));
INVX1 INVX1_213 ( .A(_abc_40319_new_n906_), .Y(_abc_40319_new_n1537_));
INVX1 INVX1_214 ( .A(_abc_40319_new_n936_), .Y(_abc_40319_new_n1542_));
INVX1 INVX1_215 ( .A(_abc_40319_new_n925_), .Y(_abc_40319_new_n1543_));
INVX1 INVX1_216 ( .A(_abc_40319_new_n932_), .Y(_abc_40319_new_n1545_));
INVX1 INVX1_217 ( .A(_abc_40319_new_n962_), .Y(_abc_40319_new_n1550_));
INVX1 INVX1_218 ( .A(_abc_40319_new_n1563_), .Y(_abc_40319_new_n1564_));
INVX1 INVX1_219 ( .A(_abc_40319_new_n1567_), .Y(_abc_40319_new_n1568_));
INVX1 INVX1_22 ( .A(IR_REG_14_), .Y(_abc_40319_new_n558_));
INVX1 INVX1_220 ( .A(_abc_40319_new_n1569_), .Y(_abc_40319_new_n1570_));
INVX1 INVX1_221 ( .A(_abc_40319_new_n1575_), .Y(_abc_40319_new_n1576_));
INVX1 INVX1_222 ( .A(_abc_40319_new_n1579_), .Y(_abc_40319_new_n1581_));
INVX1 INVX1_223 ( .A(_abc_40319_new_n1583_), .Y(_abc_40319_new_n1584_));
INVX1 INVX1_224 ( .A(_abc_40319_new_n1585_), .Y(_abc_40319_new_n1586_));
INVX1 INVX1_225 ( .A(_abc_40319_new_n1061_), .Y(_abc_40319_new_n1587_));
INVX1 INVX1_226 ( .A(_abc_40319_new_n1589_), .Y(_abc_40319_new_n1590_));
INVX1 INVX1_227 ( .A(_abc_40319_new_n1592_), .Y(_abc_40319_new_n1593_));
INVX1 INVX1_228 ( .A(_abc_40319_new_n772_), .Y(_abc_40319_new_n1594_));
INVX1 INVX1_229 ( .A(_abc_40319_new_n1602_), .Y(_abc_40319_new_n1603_));
INVX1 INVX1_23 ( .A(IR_REG_19_), .Y(_abc_40319_new_n562_));
INVX1 INVX1_230 ( .A(_abc_40319_new_n1604_), .Y(_abc_40319_new_n1605_));
INVX1 INVX1_231 ( .A(_abc_40319_new_n1609_), .Y(_abc_40319_new_n1610_));
INVX1 INVX1_232 ( .A(_abc_40319_new_n1611_), .Y(_abc_40319_new_n1612_));
INVX1 INVX1_233 ( .A(_abc_40319_new_n1182_), .Y(_abc_40319_new_n1616_));
INVX1 INVX1_234 ( .A(_abc_40319_new_n1627_), .Y(_abc_40319_new_n1629_));
INVX1 INVX1_235 ( .A(_abc_40319_new_n1631_), .Y(_abc_40319_new_n1632_));
INVX1 INVX1_236 ( .A(_abc_40319_new_n1633_), .Y(_abc_40319_new_n1634_));
INVX1 INVX1_237 ( .A(_abc_40319_new_n1600_), .Y(_abc_40319_new_n1636_));
INVX1 INVX1_238 ( .A(_abc_40319_new_n1646_), .Y(_abc_40319_new_n1647_));
INVX1 INVX1_239 ( .A(_abc_40319_new_n1652_), .Y(_abc_40319_new_n1653_));
INVX1 INVX1_24 ( .A(IR_REG_20_), .Y(_abc_40319_new_n563_));
INVX1 INVX1_240 ( .A(_abc_40319_new_n1186_), .Y(_abc_40319_new_n1657_));
INVX1 INVX1_241 ( .A(_abc_40319_new_n1669_), .Y(_abc_40319_new_n1670_));
INVX1 INVX1_242 ( .A(_abc_40319_new_n1673_), .Y(_abc_40319_new_n1675_));
INVX1 INVX1_243 ( .A(_abc_40319_new_n1678_), .Y(_abc_40319_new_n1679_));
INVX1 INVX1_244 ( .A(_abc_40319_new_n1681_), .Y(_abc_40319_new_n1682_));
INVX1 INVX1_245 ( .A(_abc_40319_new_n1687_), .Y(_abc_40319_new_n1688_));
INVX1 INVX1_246 ( .A(_abc_40319_new_n1658_), .Y(_abc_40319_new_n1696_));
INVX1 INVX1_247 ( .A(_abc_40319_new_n1703_), .Y(_abc_40319_new_n1704_));
INVX1 INVX1_248 ( .A(_abc_40319_new_n1707_), .Y(_abc_40319_new_n1709_));
INVX1 INVX1_249 ( .A(_abc_40319_new_n1712_), .Y(_abc_40319_new_n1713_));
INVX1 INVX1_25 ( .A(IR_REG_21_), .Y(_abc_40319_new_n564_));
INVX1 INVX1_250 ( .A(_abc_40319_new_n1645_), .Y(_abc_40319_new_n1716_));
INVX1 INVX1_251 ( .A(_abc_40319_new_n1721_), .Y(_abc_40319_new_n1722_));
INVX1 INVX1_252 ( .A(_abc_40319_new_n1184_), .Y(_abc_40319_new_n1730_));
INVX1 INVX1_253 ( .A(_abc_40319_new_n1737_), .Y(_abc_40319_new_n1738_));
INVX1 INVX1_254 ( .A(_abc_40319_new_n1741_), .Y(_abc_40319_new_n1743_));
INVX1 INVX1_255 ( .A(_abc_40319_new_n1745_), .Y(_abc_40319_new_n1746_));
INVX1 INVX1_256 ( .A(_abc_40319_new_n1747_), .Y(_abc_40319_new_n1748_));
INVX1 INVX1_257 ( .A(_abc_40319_new_n1755_), .Y(_abc_40319_new_n1756_));
INVX1 INVX1_258 ( .A(_abc_40319_new_n1183_), .Y(_abc_40319_new_n1764_));
INVX1 INVX1_259 ( .A(_abc_40319_new_n1771_), .Y(_abc_40319_new_n1772_));
INVX1 INVX1_26 ( .A(_abc_40319_new_n567_), .Y(_abc_40319_new_n568_));
INVX1 INVX1_260 ( .A(_abc_40319_new_n1775_), .Y(_abc_40319_new_n1777_));
INVX1 INVX1_261 ( .A(_abc_40319_new_n1779_), .Y(_abc_40319_new_n1780_));
INVX1 INVX1_262 ( .A(_abc_40319_new_n1781_), .Y(_abc_40319_new_n1782_));
INVX1 INVX1_263 ( .A(_abc_40319_new_n1786_), .Y(_abc_40319_new_n1787_));
INVX1 INVX1_264 ( .A(_abc_40319_new_n1789_), .Y(_abc_40319_new_n1790_));
INVX1 INVX1_265 ( .A(_abc_40319_new_n1796_), .Y(_abc_40319_new_n1797_));
INVX1 INVX1_266 ( .A(_abc_40319_new_n1804_), .Y(_abc_40319_new_n1805_));
INVX1 INVX1_267 ( .A(_abc_40319_new_n1806_), .Y(_abc_40319_new_n1807_));
INVX1 INVX1_268 ( .A(_abc_40319_new_n1809_), .Y(_abc_40319_new_n1810_));
INVX1 INVX1_269 ( .A(_abc_40319_new_n1814_), .Y(_abc_40319_new_n1815_));
INVX1 INVX1_27 ( .A(IR_REG_24_), .Y(_abc_40319_new_n573_));
INVX1 INVX1_270 ( .A(_abc_40319_new_n1192_), .Y(_abc_40319_new_n1820_));
INVX1 INVX1_271 ( .A(_abc_40319_new_n1830_), .Y(_abc_40319_new_n1831_));
INVX1 INVX1_272 ( .A(_abc_40319_new_n1834_), .Y(_abc_40319_new_n1835_));
INVX1 INVX1_273 ( .A(_abc_40319_new_n1839_), .Y(_abc_40319_new_n1840_));
INVX1 INVX1_274 ( .A(_abc_40319_new_n1193_), .Y(_abc_40319_new_n1844_));
INVX1 INVX1_275 ( .A(_abc_40319_new_n1854_), .Y(_abc_40319_new_n1855_));
INVX1 INVX1_276 ( .A(_abc_40319_new_n1858_), .Y(_abc_40319_new_n1859_));
INVX1 INVX1_277 ( .A(_abc_40319_new_n1863_), .Y(_abc_40319_new_n1864_));
INVX1 INVX1_278 ( .A(_abc_40319_new_n1194_), .Y(_abc_40319_new_n1867_));
INVX1 INVX1_279 ( .A(_abc_40319_new_n1878_), .Y(_abc_40319_new_n1879_));
INVX1 INVX1_28 ( .A(IR_REG_25_), .Y(_abc_40319_new_n574_));
INVX1 INVX1_280 ( .A(_abc_40319_new_n1882_), .Y(_abc_40319_new_n1883_));
INVX1 INVX1_281 ( .A(_abc_40319_new_n1886_), .Y(_abc_40319_new_n1887_));
INVX1 INVX1_282 ( .A(_abc_40319_new_n1888_), .Y(_abc_40319_new_n1889_));
INVX1 INVX1_283 ( .A(_abc_40319_new_n1893_), .Y(_abc_40319_new_n1894_));
INVX1 INVX1_284 ( .A(_abc_40319_new_n1895_), .Y(_abc_40319_new_n1896_));
INVX1 INVX1_285 ( .A(_abc_40319_new_n1897_), .Y(_abc_40319_new_n1898_));
INVX1 INVX1_286 ( .A(_abc_40319_new_n1902_), .Y(_abc_40319_new_n1903_));
INVX1 INVX1_287 ( .A(_abc_40319_new_n1223_), .Y(_abc_40319_new_n1914_));
INVX1 INVX1_288 ( .A(_abc_40319_new_n1327_), .Y(_abc_40319_new_n1915_));
INVX1 INVX1_289 ( .A(_abc_40319_new_n1328_), .Y(_abc_40319_new_n1916_));
INVX1 INVX1_29 ( .A(_abc_40319_new_n578_), .Y(_abc_40319_new_n579_));
INVX1 INVX1_290 ( .A(_abc_40319_new_n1351_), .Y(_abc_40319_new_n1917_));
INVX1 INVX1_291 ( .A(_abc_40319_new_n1352_), .Y(_abc_40319_new_n1918_));
INVX1 INVX1_292 ( .A(_abc_40319_new_n1385_), .Y(_abc_40319_new_n1919_));
INVX1 INVX1_293 ( .A(_abc_40319_new_n1386_), .Y(_abc_40319_new_n1920_));
INVX1 INVX1_294 ( .A(_abc_40319_new_n1458_), .Y(_abc_40319_new_n1921_));
INVX1 INVX1_295 ( .A(_abc_40319_new_n1493_), .Y(_abc_40319_new_n1922_));
INVX1 INVX1_296 ( .A(_abc_40319_new_n1494_), .Y(_abc_40319_new_n1923_));
INVX1 INVX1_297 ( .A(_abc_40319_new_n1527_), .Y(_abc_40319_new_n1924_));
INVX1 INVX1_298 ( .A(_abc_40319_new_n1528_), .Y(_abc_40319_new_n1925_));
INVX1 INVX1_299 ( .A(_abc_40319_new_n1638_), .Y(_abc_40319_new_n1926_));
INVX1 INVX1_3 ( .A(IR_REG_26_), .Y(_abc_40319_new_n525_));
INVX1 INVX1_30 ( .A(_abc_40319_new_n576_), .Y(_abc_40319_new_n583_));
INVX1 INVX1_300 ( .A(_abc_40319_new_n1641_), .Y(_abc_40319_new_n1927_));
INVX1 INVX1_301 ( .A(_abc_40319_new_n1783_), .Y(_abc_40319_new_n1930_));
INVX1 INVX1_302 ( .A(_abc_40319_new_n1891_), .Y(_abc_40319_new_n1941_));
INVX1 INVX1_303 ( .A(_abc_40319_new_n1910_), .Y(_abc_40319_new_n1948_));
INVX1 INVX1_304 ( .A(_abc_40319_new_n1970_), .Y(_abc_40319_new_n1971_));
INVX1 INVX1_305 ( .A(_abc_40319_new_n1992_), .Y(_abc_40319_new_n1993_));
INVX1 INVX1_306 ( .A(_abc_40319_new_n2010_), .Y(_abc_40319_new_n2011_));
INVX1 INVX1_307 ( .A(_abc_40319_new_n1785_), .Y(_abc_40319_new_n2028_));
INVX1 INVX1_308 ( .A(_abc_40319_new_n2029_), .Y(_abc_40319_new_n2030_));
INVX1 INVX1_309 ( .A(_abc_40319_new_n976_), .Y(_abc_40319_new_n2049_));
INVX1 INVX1_31 ( .A(_abc_40319_new_n590_), .Y(_abc_40319_new_n591_));
INVX1 INVX1_310 ( .A(_abc_40319_new_n2051_), .Y(_abc_40319_new_n2052_));
INVX1 INVX1_311 ( .A(_abc_40319_new_n2048_), .Y(_abc_40319_new_n2054_));
INVX1 INVX1_312 ( .A(_abc_40319_new_n2070_), .Y(_abc_40319_new_n2071_));
INVX1 INVX1_313 ( .A(_abc_40319_new_n2095_), .Y(_abc_40319_new_n2096_));
INVX1 INVX1_314 ( .A(_abc_40319_new_n2092_), .Y(_abc_40319_new_n2101_));
INVX1 INVX1_315 ( .A(_abc_40319_new_n2099_), .Y(_abc_40319_new_n2102_));
INVX1 INVX1_316 ( .A(_abc_40319_new_n2104_), .Y(_abc_40319_new_n2105_));
INVX1 INVX1_317 ( .A(_abc_40319_new_n1222_), .Y(_abc_40319_new_n2108_));
INVX1 INVX1_318 ( .A(_abc_40319_new_n2136_), .Y(_abc_40319_new_n2137_));
INVX1 INVX1_319 ( .A(_abc_40319_new_n2138_), .Y(_abc_40319_new_n2139_));
INVX1 INVX1_32 ( .A(_abc_40319_new_n584_), .Y(_abc_40319_new_n592_));
INVX1 INVX1_320 ( .A(_abc_40319_new_n2135_), .Y(_abc_40319_new_n2141_));
INVX1 INVX1_321 ( .A(_abc_40319_new_n2175_), .Y(_abc_40319_new_n2176_));
INVX1 INVX1_322 ( .A(_abc_40319_new_n1890_), .Y(_abc_40319_new_n2178_));
INVX1 INVX1_323 ( .A(_abc_40319_new_n1899_), .Y(_abc_40319_new_n2182_));
INVX1 INVX1_324 ( .A(_abc_40319_new_n2202_), .Y(_abc_40319_new_n2208_));
INVX1 INVX1_325 ( .A(_abc_40319_new_n2206_), .Y(_abc_40319_new_n2209_));
INVX1 INVX1_326 ( .A(_abc_40319_new_n2225_), .Y(_abc_40319_new_n2229_));
INVX1 INVX1_327 ( .A(_abc_40319_new_n2227_), .Y(_abc_40319_new_n2230_));
INVX1 INVX1_328 ( .A(_abc_40319_new_n2246_), .Y(_abc_40319_new_n2247_));
INVX1 INVX1_329 ( .A(_abc_40319_new_n2264_), .Y(_abc_40319_new_n2265_));
INVX1 INVX1_33 ( .A(_abc_40319_new_n599_), .Y(_abc_40319_new_n600_));
INVX1 INVX1_330 ( .A(_abc_40319_new_n1296_), .Y(_abc_40319_new_n2303_));
INVX1 INVX1_331 ( .A(_abc_40319_new_n2304_), .Y(_abc_40319_new_n2305_));
INVX1 INVX1_332 ( .A(_abc_40319_new_n2322_), .Y(_abc_40319_new_n2323_));
INVX1 INVX1_333 ( .A(_abc_40319_new_n2357_), .Y(_abc_40319_new_n2358_));
INVX1 INVX1_334 ( .A(_abc_40319_new_n2373_), .Y(_abc_40319_new_n2374_));
INVX1 INVX1_335 ( .A(_abc_40319_new_n1714_), .Y(_abc_40319_new_n2392_));
INVX1 INVX1_336 ( .A(_abc_40319_new_n1792_), .Y(_abc_40319_new_n2393_));
INVX1 INVX1_337 ( .A(_abc_40319_new_n1791_), .Y(_abc_40319_new_n2397_));
INVX1 INVX1_338 ( .A(_abc_40319_new_n2417_), .Y(_abc_40319_new_n2419_));
INVX1 INVX1_339 ( .A(_abc_40319_new_n2204_), .Y(_abc_40319_new_n2435_));
INVX1 INVX1_34 ( .A(_abc_40319_new_n601_), .Y(_abc_40319_new_n602_));
INVX1 INVX1_340 ( .A(_abc_40319_new_n2436_), .Y(_abc_40319_new_n2438_));
INVX1 INVX1_341 ( .A(_abc_40319_new_n2454_), .Y(_abc_40319_new_n2455_));
INVX1 INVX1_342 ( .A(_abc_40319_new_n2472_), .Y(_abc_40319_new_n2474_));
INVX1 INVX1_343 ( .A(_abc_40319_new_n2490_), .Y(_abc_40319_new_n2491_));
INVX1 INVX1_344 ( .A(_abc_40319_new_n1273_), .Y(_abc_40319_new_n2509_));
INVX1 INVX1_345 ( .A(_abc_40319_new_n1301_), .Y(_abc_40319_new_n2513_));
INVX1 INVX1_346 ( .A(_abc_40319_new_n2531_), .Y(_abc_40319_new_n2532_));
INVX1 INVX1_347 ( .A(_abc_40319_new_n613_), .Y(_abc_40319_new_n2549_));
INVX1 INVX1_348 ( .A(_abc_40319_new_n2551_), .Y(_abc_40319_new_n2555_));
INVX1 INVX1_349 ( .A(_abc_40319_new_n2565_), .Y(_abc_40319_new_n2566_));
INVX1 INVX1_35 ( .A(_abc_40319_new_n565_), .Y(_abc_40319_new_n603_));
INVX1 INVX1_350 ( .A(_abc_40319_new_n2567_), .Y(_abc_40319_new_n2568_));
INVX1 INVX1_351 ( .A(_abc_40319_new_n2573_), .Y(_abc_40319_new_n2574_));
INVX1 INVX1_352 ( .A(_abc_40319_new_n1046_), .Y(_abc_40319_new_n2575_));
INVX1 INVX1_353 ( .A(_abc_40319_new_n1034_), .Y(_abc_40319_new_n2578_));
INVX1 INVX1_354 ( .A(_abc_40319_new_n2580_), .Y(_abc_40319_new_n2581_));
INVX1 INVX1_355 ( .A(_abc_40319_new_n1010_), .Y(_abc_40319_new_n2583_));
INVX1 INVX1_356 ( .A(_abc_40319_new_n998_), .Y(_abc_40319_new_n2585_));
INVX1 INVX1_357 ( .A(_abc_40319_new_n2587_), .Y(_abc_40319_new_n2588_));
INVX1 INVX1_358 ( .A(_abc_40319_new_n2593_), .Y(_abc_40319_new_n2594_));
INVX1 INVX1_359 ( .A(_abc_40319_new_n2596_), .Y(_abc_40319_new_n2597_));
INVX1 INVX1_36 ( .A(_abc_40319_new_n606_), .Y(_abc_40319_new_n607_));
INVX1 INVX1_360 ( .A(_abc_40319_new_n746_), .Y(_abc_40319_new_n2603_));
INVX1 INVX1_361 ( .A(_abc_40319_new_n689_), .Y(_abc_40319_new_n2605_));
INVX1 INVX1_362 ( .A(_abc_40319_new_n2609_), .Y(_abc_40319_new_n2610_));
INVX1 INVX1_363 ( .A(_abc_40319_new_n2552_), .Y(_abc_40319_new_n2611_));
INVX1 INVX1_364 ( .A(_abc_40319_new_n2613_), .Y(_abc_40319_new_n2614_));
INVX1 INVX1_365 ( .A(_abc_40319_new_n2617_), .Y(_abc_40319_new_n2618_));
INVX1 INVX1_366 ( .A(_abc_40319_new_n2622_), .Y(_abc_40319_new_n2623_));
INVX1 INVX1_367 ( .A(_abc_40319_new_n2634_), .Y(_abc_40319_new_n2635_));
INVX1 INVX1_368 ( .A(_abc_40319_new_n2638_), .Y(_abc_40319_new_n2639_));
INVX1 INVX1_369 ( .A(_abc_40319_new_n829_), .Y(_abc_40319_new_n2650_));
INVX1 INVX1_37 ( .A(_abc_40319_new_n608_), .Y(_abc_40319_new_n609_));
INVX1 INVX1_370 ( .A(_abc_40319_new_n2576_), .Y(_abc_40319_new_n2656_));
INVX1 INVX1_371 ( .A(_abc_40319_new_n2665_), .Y(_abc_40319_new_n2666_));
INVX1 INVX1_372 ( .A(_abc_40319_new_n2667_), .Y(_abc_40319_new_n2668_));
INVX1 INVX1_373 ( .A(_abc_40319_new_n2642_), .Y(_abc_40319_new_n2675_));
INVX1 INVX1_374 ( .A(_abc_40319_new_n2644_), .Y(_abc_40319_new_n2677_));
INVX1 INVX1_375 ( .A(_abc_40319_new_n2680_), .Y(_abc_40319_new_n2681_));
INVX1 INVX1_376 ( .A(_abc_40319_new_n2621_), .Y(_abc_40319_new_n2688_));
INVX1 INVX1_377 ( .A(_abc_40319_new_n1769_), .Y(_abc_40319_new_n2701_));
INVX1 INVX1_378 ( .A(_abc_40319_new_n1758_), .Y(_abc_40319_new_n2703_));
INVX1 INVX1_379 ( .A(_abc_40319_new_n1625_), .Y(_abc_40319_new_n2712_));
INVX1 INVX1_38 ( .A(STATE_REG), .Y(_abc_40319_new_n617_));
INVX1 INVX1_380 ( .A(_abc_40319_new_n1614_), .Y(_abc_40319_new_n2714_));
INVX1 INVX1_381 ( .A(_abc_40319_new_n2718_), .Y(_abc_40319_new_n2719_));
INVX1 INVX1_382 ( .A(_abc_40319_new_n1146_), .Y(_abc_40319_new_n2728_));
INVX1 INVX1_383 ( .A(_abc_40319_new_n1572_), .Y(_abc_40319_new_n2730_));
INVX1 INVX1_384 ( .A(_abc_40319_new_n2734_), .Y(_abc_40319_new_n2735_));
INVX1 INVX1_385 ( .A(_abc_40319_new_n2739_), .Y(_abc_40319_new_n2740_));
INVX1 INVX1_386 ( .A(_abc_40319_new_n2751_), .Y(_abc_40319_new_n2752_));
INVX1 INVX1_387 ( .A(_abc_40319_new_n1667_), .Y(_abc_40319_new_n2753_));
INVX1 INVX1_388 ( .A(_abc_40319_new_n1655_), .Y(_abc_40319_new_n2755_));
INVX1 INVX1_389 ( .A(_abc_40319_new_n2757_), .Y(_abc_40319_new_n2758_));
INVX1 INVX1_39 ( .A(IR_REG_27_), .Y(_abc_40319_new_n620_));
INVX1 INVX1_390 ( .A(_abc_40319_new_n1701_), .Y(_abc_40319_new_n2760_));
INVX1 INVX1_391 ( .A(_abc_40319_new_n1690_), .Y(_abc_40319_new_n2762_));
INVX1 INVX1_392 ( .A(_abc_40319_new_n2764_), .Y(_abc_40319_new_n2765_));
INVX1 INVX1_393 ( .A(_abc_40319_new_n2770_), .Y(_abc_40319_new_n2771_));
INVX1 INVX1_394 ( .A(_abc_40319_new_n2773_), .Y(_abc_40319_new_n2774_));
INVX1 INVX1_395 ( .A(_abc_40319_new_n2780_), .Y(_abc_40319_new_n2781_));
INVX1 INVX1_396 ( .A(_abc_40319_new_n1735_), .Y(_abc_40319_new_n2782_));
INVX1 INVX1_397 ( .A(_abc_40319_new_n1724_), .Y(_abc_40319_new_n2784_));
INVX1 INVX1_398 ( .A(_abc_40319_new_n2786_), .Y(_abc_40319_new_n2787_));
INVX1 INVX1_399 ( .A(_abc_40319_new_n2788_), .Y(_abc_40319_new_n2789_));
INVX1 INVX1_4 ( .A(_abc_40319_new_n526_), .Y(_abc_40319_new_n527_));
INVX1 INVX1_40 ( .A(_abc_40319_new_n624_), .Y(_abc_40319_new_n625_));
INVX1 INVX1_400 ( .A(_abc_40319_new_n2793_), .Y(_abc_40319_new_n2794_));
INVX1 INVX1_401 ( .A(_abc_40319_new_n2759_), .Y(_abc_40319_new_n2798_));
INVX1 INVX1_402 ( .A(_abc_40319_new_n1517_), .Y(_abc_40319_new_n2807_));
INVX1 INVX1_403 ( .A(_abc_40319_new_n1506_), .Y(_abc_40319_new_n2809_));
INVX1 INVX1_404 ( .A(_abc_40319_new_n2815_), .Y(_abc_40319_new_n2816_));
INVX1 INVX1_405 ( .A(_abc_40319_new_n2823_), .Y(_abc_40319_new_n2824_));
INVX1 INVX1_406 ( .A(_abc_40319_new_n1483_), .Y(_abc_40319_new_n2825_));
INVX1 INVX1_407 ( .A(_abc_40319_new_n1471_), .Y(_abc_40319_new_n2827_));
INVX1 INVX1_408 ( .A(_abc_40319_new_n2829_), .Y(_abc_40319_new_n2830_));
INVX1 INVX1_409 ( .A(_abc_40319_new_n2831_), .Y(_abc_40319_new_n2832_));
INVX1 INVX1_41 ( .A(_abc_40319_new_n628_), .Y(_abc_40319_new_n629_));
INVX1 INVX1_410 ( .A(_abc_40319_new_n2833_), .Y(_abc_40319_new_n2834_));
INVX1 INVX1_411 ( .A(_abc_40319_new_n1410_), .Y(_abc_40319_new_n2842_));
INVX1 INVX1_412 ( .A(_abc_40319_new_n1398_), .Y(_abc_40319_new_n2844_));
INVX1 INVX1_413 ( .A(_abc_40319_new_n2848_), .Y(_abc_40319_new_n2849_));
INVX1 INVX1_414 ( .A(_abc_40319_new_n2856_), .Y(_abc_40319_new_n2857_));
INVX1 INVX1_415 ( .A(_abc_40319_new_n1444_), .Y(_abc_40319_new_n2858_));
INVX1 INVX1_416 ( .A(_abc_40319_new_n1433_), .Y(_abc_40319_new_n2860_));
INVX1 INVX1_417 ( .A(_abc_40319_new_n2862_), .Y(_abc_40319_new_n2863_));
INVX1 INVX1_418 ( .A(_abc_40319_new_n2864_), .Y(_abc_40319_new_n2865_));
INVX1 INVX1_419 ( .A(_abc_40319_new_n2866_), .Y(_abc_40319_new_n2867_));
INVX1 INVX1_42 ( .A(IR_REG_28_), .Y(_abc_40319_new_n630_));
INVX1 INVX1_420 ( .A(_abc_40319_new_n1374_), .Y(_abc_40319_new_n2875_));
INVX1 INVX1_421 ( .A(_abc_40319_new_n1363_), .Y(_abc_40319_new_n2877_));
INVX1 INVX1_422 ( .A(_abc_40319_new_n2881_), .Y(_abc_40319_new_n2882_));
INVX1 INVX1_423 ( .A(_abc_40319_new_n2889_), .Y(_abc_40319_new_n2890_));
INVX1 INVX1_424 ( .A(_abc_40319_new_n1828_), .Y(_abc_40319_new_n2891_));
INVX1 INVX1_425 ( .A(_abc_40319_new_n1817_), .Y(_abc_40319_new_n2893_));
INVX1 INVX1_426 ( .A(_abc_40319_new_n2895_), .Y(_abc_40319_new_n2896_));
INVX1 INVX1_427 ( .A(_abc_40319_new_n2897_), .Y(_abc_40319_new_n2898_));
INVX1 INVX1_428 ( .A(_abc_40319_new_n2899_), .Y(_abc_40319_new_n2900_));
INVX1 INVX1_429 ( .A(_abc_40319_new_n1852_), .Y(_abc_40319_new_n2908_));
INVX1 INVX1_43 ( .A(_abc_40319_new_n631_), .Y(_abc_40319_new_n632_));
INVX1 INVX1_430 ( .A(_abc_40319_new_n1841_), .Y(_abc_40319_new_n2910_));
INVX1 INVX1_431 ( .A(_abc_40319_new_n2914_), .Y(_abc_40319_new_n2915_));
INVX1 INVX1_432 ( .A(_abc_40319_new_n2922_), .Y(_abc_40319_new_n2923_));
INVX1 INVX1_433 ( .A(_abc_40319_new_n1876_), .Y(_abc_40319_new_n2924_));
INVX1 INVX1_434 ( .A(_abc_40319_new_n1865_), .Y(_abc_40319_new_n2926_));
INVX1 INVX1_435 ( .A(_abc_40319_new_n2928_), .Y(_abc_40319_new_n2929_));
INVX1 INVX1_436 ( .A(_abc_40319_new_n2930_), .Y(_abc_40319_new_n2931_));
INVX1 INVX1_437 ( .A(_abc_40319_new_n2932_), .Y(_abc_40319_new_n2933_));
INVX1 INVX1_438 ( .A(_abc_40319_new_n1340_), .Y(_abc_40319_new_n2941_));
INVX1 INVX1_439 ( .A(_abc_40319_new_n1329_), .Y(_abc_40319_new_n2943_));
INVX1 INVX1_44 ( .A(_abc_40319_new_n633_), .Y(_abc_40319_new_n634_));
INVX1 INVX1_440 ( .A(_abc_40319_new_n2947_), .Y(_abc_40319_new_n2948_));
INVX1 INVX1_441 ( .A(_abc_40319_new_n2955_), .Y(_abc_40319_new_n2956_));
INVX1 INVX1_442 ( .A(_abc_40319_new_n1317_), .Y(_abc_40319_new_n2957_));
INVX1 INVX1_443 ( .A(_abc_40319_new_n1306_), .Y(_abc_40319_new_n2959_));
INVX1 INVX1_444 ( .A(_abc_40319_new_n2961_), .Y(_abc_40319_new_n2962_));
INVX1 INVX1_445 ( .A(_abc_40319_new_n2963_), .Y(_abc_40319_new_n2964_));
INVX1 INVX1_446 ( .A(_abc_40319_new_n2965_), .Y(_abc_40319_new_n2966_));
INVX1 INVX1_447 ( .A(_abc_40319_new_n1285_), .Y(_abc_40319_new_n2974_));
INVX1 INVX1_448 ( .A(_abc_40319_new_n1274_), .Y(_abc_40319_new_n2976_));
INVX1 INVX1_449 ( .A(_abc_40319_new_n2980_), .Y(_abc_40319_new_n2981_));
INVX1 INVX1_45 ( .A(_abc_40319_new_n638_), .Y(_abc_40319_new_n639_));
INVX1 INVX1_450 ( .A(_abc_40319_new_n2988_), .Y(_abc_40319_new_n2989_));
INVX1 INVX1_451 ( .A(_abc_40319_new_n1260_), .Y(_abc_40319_new_n2990_));
INVX1 INVX1_452 ( .A(_abc_40319_new_n1249_), .Y(_abc_40319_new_n2992_));
INVX1 INVX1_453 ( .A(_abc_40319_new_n2994_), .Y(_abc_40319_new_n2995_));
INVX1 INVX1_454 ( .A(_abc_40319_new_n2996_), .Y(_abc_40319_new_n2997_));
INVX1 INVX1_455 ( .A(_abc_40319_new_n2998_), .Y(_abc_40319_new_n2999_));
INVX1 INVX1_456 ( .A(_abc_40319_new_n1235_), .Y(_abc_40319_new_n3007_));
INVX1 INVX1_457 ( .A(_abc_40319_new_n1224_), .Y(_abc_40319_new_n3009_));
INVX1 INVX1_458 ( .A(_abc_40319_new_n3013_), .Y(_abc_40319_new_n3014_));
INVX1 INVX1_459 ( .A(_abc_40319_new_n3021_), .Y(_abc_40319_new_n3022_));
INVX1 INVX1_46 ( .A(_abc_40319_new_n645_), .Y(_abc_40319_new_n646_));
INVX1 INVX1_460 ( .A(_abc_40319_new_n1210_), .Y(_abc_40319_new_n3023_));
INVX1 INVX1_461 ( .A(_abc_40319_new_n1180_), .Y(_abc_40319_new_n3025_));
INVX1 INVX1_462 ( .A(_abc_40319_new_n3027_), .Y(_abc_40319_new_n3028_));
INVX1 INVX1_463 ( .A(_abc_40319_new_n3029_), .Y(_abc_40319_new_n3030_));
INVX1 INVX1_464 ( .A(_abc_40319_new_n3031_), .Y(_abc_40319_new_n3032_));
INVX1 INVX1_465 ( .A(_abc_40319_new_n1980_), .Y(_abc_40319_new_n3040_));
INVX1 INVX1_466 ( .A(_abc_40319_new_n2089_), .Y(_abc_40319_new_n3042_));
INVX1 INVX1_467 ( .A(_abc_40319_new_n3046_), .Y(_abc_40319_new_n3047_));
INVX1 INVX1_468 ( .A(_abc_40319_new_n3055_), .Y(_abc_40319_new_n3056_));
INVX1 INVX1_469 ( .A(_abc_40319_new_n2123_), .Y(_abc_40319_new_n3057_));
INVX1 INVX1_47 ( .A(IR_REG_18_), .Y(_abc_40319_new_n647_));
INVX1 INVX1_470 ( .A(_abc_40319_new_n3051_), .Y(_abc_40319_new_n3059_));
INVX1 INVX1_471 ( .A(_abc_40319_new_n3061_), .Y(_abc_40319_new_n3062_));
INVX1 INVX1_472 ( .A(_abc_40319_new_n3063_), .Y(_abc_40319_new_n3064_));
INVX1 INVX1_473 ( .A(_abc_40319_new_n3065_), .Y(_abc_40319_new_n3066_));
INVX1 INVX1_474 ( .A(_abc_40319_new_n3083_), .Y(_abc_40319_new_n3084_));
INVX1 INVX1_475 ( .A(_abc_40319_new_n3086_), .Y(_abc_40319_new_n3087_));
INVX1 INVX1_476 ( .A(_abc_40319_new_n3091_), .Y(_abc_40319_new_n3092_));
INVX1 INVX1_477 ( .A(_abc_40319_new_n3095_), .Y(_abc_40319_new_n3096_));
INVX1 INVX1_478 ( .A(_abc_40319_new_n3099_), .Y(_abc_40319_new_n3100_));
INVX1 INVX1_479 ( .A(_abc_40319_new_n3101_), .Y(_abc_40319_new_n3102_));
INVX1 INVX1_48 ( .A(_abc_40319_new_n661_), .Y(n1341));
INVX1 INVX1_480 ( .A(_abc_40319_new_n3106_), .Y(_abc_40319_new_n3107_));
INVX1 INVX1_481 ( .A(_abc_40319_new_n3113_), .Y(_abc_40319_new_n3114_));
INVX1 INVX1_482 ( .A(_abc_40319_new_n3115_), .Y(_abc_40319_new_n3116_));
INVX1 INVX1_483 ( .A(_abc_40319_new_n3118_), .Y(_abc_40319_new_n3119_));
INVX1 INVX1_484 ( .A(_abc_40319_new_n3123_), .Y(_abc_40319_new_n3124_));
INVX1 INVX1_485 ( .A(_abc_40319_new_n3127_), .Y(_abc_40319_new_n3128_));
INVX1 INVX1_486 ( .A(_abc_40319_new_n3133_), .Y(_abc_40319_new_n3134_));
INVX1 INVX1_487 ( .A(_abc_40319_new_n3137_), .Y(_abc_40319_new_n3138_));
INVX1 INVX1_488 ( .A(_abc_40319_new_n3142_), .Y(_abc_40319_new_n3143_));
INVX1 INVX1_489 ( .A(_abc_40319_new_n3146_), .Y(_abc_40319_new_n3147_));
INVX1 INVX1_49 ( .A(_abc_40319_new_n598_), .Y(_abc_40319_new_n663_));
INVX1 INVX1_490 ( .A(_abc_40319_new_n3153_), .Y(_abc_40319_new_n3154_));
INVX1 INVX1_491 ( .A(_abc_40319_new_n3157_), .Y(_abc_40319_new_n3158_));
INVX1 INVX1_492 ( .A(_abc_40319_new_n2560_), .Y(_abc_40319_new_n3159_));
INVX1 INVX1_493 ( .A(_abc_40319_new_n3160_), .Y(_abc_40319_new_n3161_));
INVX1 INVX1_494 ( .A(_abc_40319_new_n2553_), .Y(_abc_40319_new_n3162_));
INVX1 INVX1_495 ( .A(_abc_40319_new_n3163_), .Y(_abc_40319_new_n3164_));
INVX1 INVX1_496 ( .A(_abc_40319_new_n3075_), .Y(_abc_40319_new_n3166_));
INVX1 INVX1_497 ( .A(_abc_40319_new_n3167_), .Y(_abc_40319_new_n3168_));
INVX1 INVX1_498 ( .A(_abc_40319_new_n3069_), .Y(_abc_40319_new_n3169_));
INVX1 INVX1_499 ( .A(_abc_40319_new_n3170_), .Y(_abc_40319_new_n3171_));
INVX1 INVX1_5 ( .A(IR_REG_2_), .Y(_abc_40319_new_n528_));
INVX1 INVX1_50 ( .A(_abc_40319_new_n664_), .Y(_abc_40319_new_n665_));
INVX1 INVX1_500 ( .A(_abc_40319_new_n3176_), .Y(_abc_40319_new_n3177_));
INVX1 INVX1_501 ( .A(_abc_40319_new_n3185_), .Y(_abc_40319_new_n3186_));
INVX1 INVX1_502 ( .A(_abc_40319_new_n3189_), .Y(_abc_40319_new_n3190_));
INVX1 INVX1_503 ( .A(_abc_40319_new_n3195_), .Y(_abc_40319_new_n3196_));
INVX1 INVX1_504 ( .A(_abc_40319_new_n3199_), .Y(_abc_40319_new_n3200_));
INVX1 INVX1_505 ( .A(_abc_40319_new_n3203_), .Y(_abc_40319_new_n3204_));
INVX1 INVX1_506 ( .A(_abc_40319_new_n3207_), .Y(_abc_40319_new_n3208_));
INVX1 INVX1_507 ( .A(_abc_40319_new_n3211_), .Y(_abc_40319_new_n3212_));
INVX1 INVX1_508 ( .A(_abc_40319_new_n3215_), .Y(_abc_40319_new_n3216_));
INVX1 INVX1_509 ( .A(_abc_40319_new_n784_), .Y(_abc_40319_new_n3218_));
INVX1 INVX1_51 ( .A(_abc_40319_new_n650_), .Y(_abc_40319_new_n666_));
INVX1 INVX1_510 ( .A(_abc_40319_new_n795_), .Y(_abc_40319_new_n3220_));
INVX1 INVX1_511 ( .A(_abc_40319_new_n3222_), .Y(_abc_40319_new_n3223_));
INVX1 INVX1_512 ( .A(_abc_40319_new_n3226_), .Y(_abc_40319_new_n3227_));
INVX1 INVX1_513 ( .A(_abc_40319_new_n3231_), .Y(_abc_40319_new_n3232_));
INVX1 INVX1_514 ( .A(_abc_40319_new_n3235_), .Y(_abc_40319_new_n3236_));
INVX1 INVX1_515 ( .A(_abc_40319_new_n3249_), .Y(_abc_40319_new_n3250_));
INVX1 INVX1_516 ( .A(_abc_40319_new_n3253_), .Y(_abc_40319_new_n3254_));
INVX1 INVX1_517 ( .A(_abc_40319_new_n3257_), .Y(_abc_40319_new_n3258_));
INVX1 INVX1_518 ( .A(_abc_40319_new_n3261_), .Y(_abc_40319_new_n3262_));
INVX1 INVX1_519 ( .A(_abc_40319_new_n3247_), .Y(_abc_40319_new_n3268_));
INVX1 INVX1_52 ( .A(_abc_40319_new_n670_), .Y(_abc_40319_new_n671_));
INVX1 INVX1_520 ( .A(_abc_40319_new_n3251_), .Y(_abc_40319_new_n3270_));
INVX1 INVX1_521 ( .A(_abc_40319_new_n3273_), .Y(_abc_40319_new_n3274_));
INVX1 INVX1_522 ( .A(_abc_40319_new_n3193_), .Y(_abc_40319_new_n3275_));
INVX1 INVX1_523 ( .A(_abc_40319_new_n3259_), .Y(_abc_40319_new_n3276_));
INVX1 INVX1_524 ( .A(_abc_40319_new_n3278_), .Y(_abc_40319_new_n3279_));
INVX1 INVX1_525 ( .A(_abc_40319_new_n3283_), .Y(_abc_40319_new_n3284_));
INVX1 INVX1_526 ( .A(_abc_40319_new_n3201_), .Y(_abc_40319_new_n3286_));
INVX1 INVX1_527 ( .A(_abc_40319_new_n3287_), .Y(_abc_40319_new_n3288_));
INVX1 INVX1_528 ( .A(_abc_40319_new_n3229_), .Y(_abc_40319_new_n3290_));
INVX1 INVX1_529 ( .A(_abc_40319_new_n3151_), .Y(_abc_40319_new_n3291_));
INVX1 INVX1_53 ( .A(_abc_40319_new_n531_), .Y(_abc_40319_new_n674_));
INVX1 INVX1_530 ( .A(_abc_40319_new_n3187_), .Y(_abc_40319_new_n3292_));
INVX1 INVX1_531 ( .A(_abc_40319_new_n3293_), .Y(_abc_40319_new_n3294_));
INVX1 INVX1_532 ( .A(_abc_40319_new_n3152_), .Y(_abc_40319_new_n3295_));
INVX1 INVX1_533 ( .A(_abc_40319_new_n3297_), .Y(_abc_40319_new_n3298_));
INVX1 INVX1_534 ( .A(_abc_40319_new_n3233_), .Y(_abc_40319_new_n3303_));
INVX1 INVX1_535 ( .A(_abc_40319_new_n3140_), .Y(_abc_40319_new_n3304_));
INVX1 INVX1_536 ( .A(_abc_40319_new_n3111_), .Y(_abc_40319_new_n3307_));
INVX1 INVX1_537 ( .A(_abc_40319_new_n3144_), .Y(_abc_40319_new_n3308_));
INVX1 INVX1_538 ( .A(_abc_40319_new_n3205_), .Y(_abc_40319_new_n3312_));
INVX1 INVX1_539 ( .A(_abc_40319_new_n3224_), .Y(_abc_40319_new_n3313_));
INVX1 INVX1_54 ( .A(_abc_40319_new_n675_), .Y(_abc_40319_new_n676_));
INVX1 INVX1_540 ( .A(_abc_40319_new_n3209_), .Y(_abc_40319_new_n3316_));
INVX1 INVX1_541 ( .A(_abc_40319_new_n3155_), .Y(_abc_40319_new_n3317_));
INVX1 INVX1_542 ( .A(_abc_40319_new_n3174_), .Y(_abc_40319_new_n3318_));
INVX1 INVX1_543 ( .A(_abc_40319_new_n3325_), .Y(_abc_40319_new_n3326_));
INVX1 INVX1_544 ( .A(_abc_40319_new_n3213_), .Y(_abc_40319_new_n3328_));
INVX1 INVX1_545 ( .A(_abc_40319_new_n3121_), .Y(_abc_40319_new_n3332_));
INVX1 INVX1_546 ( .A(_abc_40319_new_n3219_), .Y(_abc_40319_new_n3335_));
INVX1 INVX1_547 ( .A(_abc_40319_new_n3132_), .Y(_abc_40319_new_n3336_));
INVX1 INVX1_548 ( .A(_abc_40319_new_n3125_), .Y(_abc_40319_new_n3337_));
INVX1 INVX1_549 ( .A(_abc_40319_new_n3344_), .Y(_abc_40319_new_n3345_));
INVX1 INVX1_55 ( .A(_abc_40319_new_n677_), .Y(_abc_40319_new_n678_));
INVX1 INVX1_550 ( .A(_abc_40319_new_n3197_), .Y(_abc_40319_new_n3349_));
INVX1 INVX1_551 ( .A(_abc_40319_new_n3353_), .Y(_abc_40319_new_n3354_));
INVX1 INVX1_552 ( .A(_abc_40319_new_n3364_), .Y(_abc_40319_new_n3365_));
INVX1 INVX1_553 ( .A(_abc_40319_new_n3373_), .Y(_abc_40319_new_n3374_));
INVX1 INVX1_554 ( .A(_abc_40319_new_n3376_), .Y(_abc_40319_new_n3377_));
INVX1 INVX1_555 ( .A(_abc_40319_new_n3105_), .Y(_abc_40319_new_n3378_));
INVX1 INVX1_556 ( .A(_abc_40319_new_n3256_), .Y(_abc_40319_new_n3379_));
INVX1 INVX1_557 ( .A(_abc_40319_new_n3384_), .Y(_abc_40319_new_n3385_));
INVX1 INVX1_558 ( .A(_abc_40319_new_n3388_), .Y(_abc_40319_new_n3389_));
INVX1 INVX1_559 ( .A(_abc_40319_new_n3202_), .Y(_abc_40319_new_n3398_));
INVX1 INVX1_56 ( .A(_abc_40319_new_n680_), .Y(_abc_40319_new_n681_));
INVX1 INVX1_560 ( .A(_abc_40319_new_n3198_), .Y(_abc_40319_new_n3399_));
INVX1 INVX1_561 ( .A(_abc_40319_new_n3289_), .Y(_abc_40319_new_n3401_));
INVX1 INVX1_562 ( .A(_abc_40319_new_n3184_), .Y(_abc_40319_new_n3402_));
INVX1 INVX1_563 ( .A(_abc_40319_new_n3407_), .Y(_abc_40319_new_n3408_));
INVX1 INVX1_564 ( .A(_abc_40319_new_n3439_), .Y(_abc_40319_new_n3440_));
INVX1 INVX1_565 ( .A(_abc_40319_new_n3441_), .Y(_abc_40319_new_n3442_));
INVX1 INVX1_566 ( .A(_abc_40319_new_n3397_), .Y(_abc_40319_new_n3465_));
INVX1 INVX1_567 ( .A(_abc_40319_new_n3104_), .Y(_abc_40319_new_n3466_));
INVX1 INVX1_568 ( .A(_abc_40319_new_n3467_), .Y(_abc_40319_new_n3468_));
INVX1 INVX1_569 ( .A(_abc_40319_new_n3470_), .Y(_abc_40319_new_n3471_));
INVX1 INVX1_57 ( .A(_abc_40319_new_n684_), .Y(_abc_40319_new_n685_));
INVX1 INVX1_570 ( .A(_abc_40319_new_n3188_), .Y(_abc_40319_new_n3472_));
INVX1 INVX1_571 ( .A(_abc_40319_new_n3366_), .Y(_abc_40319_new_n3473_));
INVX1 INVX1_572 ( .A(_abc_40319_new_n3474_), .Y(_abc_40319_new_n3475_));
INVX1 INVX1_573 ( .A(_abc_40319_new_n3145_), .Y(_abc_40319_new_n3476_));
INVX1 INVX1_574 ( .A(_abc_40319_new_n3230_), .Y(_abc_40319_new_n3477_));
INVX1 INVX1_575 ( .A(_abc_40319_new_n3112_), .Y(_abc_40319_new_n3478_));
INVX1 INVX1_576 ( .A(_abc_40319_new_n3480_), .Y(_abc_40319_new_n3481_));
INVX1 INVX1_577 ( .A(_abc_40319_new_n3225_), .Y(_abc_40319_new_n3483_));
INVX1 INVX1_578 ( .A(_abc_40319_new_n3206_), .Y(_abc_40319_new_n3484_));
INVX1 INVX1_579 ( .A(_abc_40319_new_n3486_), .Y(_abc_40319_new_n3487_));
INVX1 INVX1_58 ( .A(_abc_40319_new_n686_), .Y(_abc_40319_new_n687_));
INVX1 INVX1_580 ( .A(_abc_40319_new_n3221_), .Y(_abc_40319_new_n3496_));
INVX1 INVX1_581 ( .A(_abc_40319_new_n3497_), .Y(_abc_40319_new_n3498_));
INVX1 INVX1_582 ( .A(_abc_40319_new_n3499_), .Y(_abc_40319_new_n3500_));
INVX1 INVX1_583 ( .A(_abc_40319_new_n3156_), .Y(_abc_40319_new_n3510_));
INVX1 INVX1_584 ( .A(_abc_40319_new_n3511_), .Y(_abc_40319_new_n3512_));
INVX1 INVX1_585 ( .A(_abc_40319_new_n3520_), .Y(_abc_40319_new_n3521_));
INVX1 INVX1_586 ( .A(_abc_40319_new_n3524_), .Y(_abc_40319_new_n3525_));
INVX1 INVX1_587 ( .A(_abc_40319_new_n3526_), .Y(_abc_40319_new_n3527_));
INVX1 INVX1_588 ( .A(_abc_40319_new_n3533_), .Y(_abc_40319_new_n3534_));
INVX1 INVX1_589 ( .A(_abc_40319_new_n3541_), .Y(_abc_40319_new_n3542_));
INVX1 INVX1_59 ( .A(_abc_40319_new_n691_), .Y(_abc_40319_new_n692_));
INVX1 INVX1_590 ( .A(_abc_40319_new_n3266_), .Y(_abc_40319_new_n3544_));
INVX1 INVX1_591 ( .A(_abc_40319_new_n3556_), .Y(_abc_40319_new_n3557_));
INVX1 INVX1_592 ( .A(_abc_40319_new_n3567_), .Y(_abc_40319_new_n3568_));
INVX1 INVX1_593 ( .A(_abc_40319_new_n3573_), .Y(_abc_40319_new_n3574_));
INVX1 INVX1_594 ( .A(_abc_40319_new_n3584_), .Y(_abc_40319_new_n3585_));
INVX1 INVX1_595 ( .A(REG2_REG_1_), .Y(_abc_40319_new_n3589_));
INVX1 INVX1_596 ( .A(_abc_40319_new_n3590_), .Y(_abc_40319_new_n3591_));
INVX1 INVX1_597 ( .A(_abc_40319_new_n3592_), .Y(_abc_40319_new_n3593_));
INVX1 INVX1_598 ( .A(_abc_40319_new_n886_), .Y(_abc_40319_new_n3596_));
INVX1 INVX1_599 ( .A(_abc_40319_new_n3594_), .Y(_abc_40319_new_n3597_));
INVX1 INVX1_6 ( .A(_abc_40319_new_n529_), .Y(_abc_40319_new_n530_));
INVX1 INVX1_60 ( .A(_abc_40319_new_n649_), .Y(_abc_40319_new_n693_));
INVX1 INVX1_600 ( .A(_abc_40319_new_n3601_), .Y(_abc_40319_new_n3602_));
INVX1 INVX1_601 ( .A(REG1_REG_1_), .Y(_abc_40319_new_n3603_));
INVX1 INVX1_602 ( .A(_abc_40319_new_n3604_), .Y(_abc_40319_new_n3605_));
INVX1 INVX1_603 ( .A(_abc_40319_new_n3606_), .Y(_abc_40319_new_n3608_));
INVX1 INVX1_604 ( .A(_abc_40319_new_n843_), .Y(_abc_40319_new_n3625_));
INVX1 INVX1_605 ( .A(_abc_40319_new_n3626_), .Y(_abc_40319_new_n3627_));
INVX1 INVX1_606 ( .A(_abc_40319_new_n3628_), .Y(_abc_40319_new_n3629_));
INVX1 INVX1_607 ( .A(_abc_40319_new_n3630_), .Y(_abc_40319_new_n3631_));
INVX1 INVX1_608 ( .A(_abc_40319_new_n3633_), .Y(_abc_40319_new_n3635_));
INVX1 INVX1_609 ( .A(_abc_40319_new_n3639_), .Y(_abc_40319_new_n3640_));
INVX1 INVX1_61 ( .A(_abc_40319_new_n697_), .Y(_abc_40319_new_n698_));
INVX1 INVX1_610 ( .A(_abc_40319_new_n3641_), .Y(_abc_40319_new_n3642_));
INVX1 INVX1_611 ( .A(_abc_40319_new_n3643_), .Y(_abc_40319_new_n3644_));
INVX1 INVX1_612 ( .A(_abc_40319_new_n3646_), .Y(_abc_40319_new_n3647_));
INVX1 INVX1_613 ( .A(REG2_REG_3_), .Y(_abc_40319_new_n3663_));
INVX1 INVX1_614 ( .A(_abc_40319_new_n3664_), .Y(_abc_40319_new_n3665_));
INVX1 INVX1_615 ( .A(_abc_40319_new_n3666_), .Y(_abc_40319_new_n3667_));
INVX1 INVX1_616 ( .A(_abc_40319_new_n3660_), .Y(_abc_40319_new_n3669_));
INVX1 INVX1_617 ( .A(REG1_REG_3_), .Y(_abc_40319_new_n3674_));
INVX1 INVX1_618 ( .A(_abc_40319_new_n3676_), .Y(_abc_40319_new_n3677_));
INVX1 INVX1_619 ( .A(_abc_40319_new_n3678_), .Y(_abc_40319_new_n3679_));
INVX1 INVX1_62 ( .A(_abc_40319_new_n700_), .Y(_abc_40319_new_n701_));
INVX1 INVX1_620 ( .A(_abc_40319_new_n3680_), .Y(_abc_40319_new_n3681_));
INVX1 INVX1_621 ( .A(_abc_40319_new_n3682_), .Y(_abc_40319_new_n3683_));
INVX1 INVX1_622 ( .A(_abc_40319_new_n3696_), .Y(_abc_40319_new_n3697_));
INVX1 INVX1_623 ( .A(REG2_REG_4_), .Y(_abc_40319_new_n3698_));
INVX1 INVX1_624 ( .A(_abc_40319_new_n3699_), .Y(_abc_40319_new_n3700_));
INVX1 INVX1_625 ( .A(_abc_40319_new_n3702_), .Y(_abc_40319_new_n3703_));
INVX1 INVX1_626 ( .A(_abc_40319_new_n3705_), .Y(_abc_40319_new_n3706_));
INVX1 INVX1_627 ( .A(REG1_REG_4_), .Y(_abc_40319_new_n3713_));
INVX1 INVX1_628 ( .A(_abc_40319_new_n3712_), .Y(_abc_40319_new_n3717_));
INVX1 INVX1_629 ( .A(_abc_40319_new_n3710_), .Y(_abc_40319_new_n3718_));
INVX1 INVX1_63 ( .A(_abc_40319_new_n704_), .Y(_abc_40319_new_n705_));
INVX1 INVX1_630 ( .A(_abc_40319_new_n3714_), .Y(_abc_40319_new_n3719_));
INVX1 INVX1_631 ( .A(_abc_40319_new_n3733_), .Y(_abc_40319_new_n3734_));
INVX1 INVX1_632 ( .A(_abc_40319_new_n3735_), .Y(_abc_40319_new_n3736_));
INVX1 INVX1_633 ( .A(REG1_REG_5_), .Y(_abc_40319_new_n3737_));
INVX1 INVX1_634 ( .A(_abc_40319_new_n3738_), .Y(_abc_40319_new_n3739_));
INVX1 INVX1_635 ( .A(_abc_40319_new_n3740_), .Y(_abc_40319_new_n3741_));
INVX1 INVX1_636 ( .A(REG2_REG_5_), .Y(_abc_40319_new_n3747_));
INVX1 INVX1_637 ( .A(_abc_40319_new_n3748_), .Y(_abc_40319_new_n3749_));
INVX1 INVX1_638 ( .A(_abc_40319_new_n3750_), .Y(_abc_40319_new_n3751_));
INVX1 INVX1_639 ( .A(_abc_40319_new_n3746_), .Y(_abc_40319_new_n3754_));
INVX1 INVX1_64 ( .A(IR_REG_30_), .Y(_abc_40319_new_n706_));
INVX1 INVX1_640 ( .A(_abc_40319_new_n3752_), .Y(_abc_40319_new_n3755_));
INVX1 INVX1_641 ( .A(_abc_40319_new_n3768_), .Y(_abc_40319_new_n3769_));
INVX1 INVX1_642 ( .A(_abc_40319_new_n3771_), .Y(_abc_40319_new_n3772_));
INVX1 INVX1_643 ( .A(_abc_40319_new_n3766_), .Y(_abc_40319_new_n3774_));
INVX1 INVX1_644 ( .A(_abc_40319_new_n3782_), .Y(_abc_40319_new_n3783_));
INVX1 INVX1_645 ( .A(_abc_40319_new_n3781_), .Y(_abc_40319_new_n3786_));
INVX1 INVX1_646 ( .A(_abc_40319_new_n3779_), .Y(_abc_40319_new_n3787_));
INVX1 INVX1_647 ( .A(_abc_40319_new_n3800_), .Y(_abc_40319_new_n3801_));
INVX1 INVX1_648 ( .A(_abc_40319_new_n3803_), .Y(_abc_40319_new_n3804_));
INVX1 INVX1_649 ( .A(_abc_40319_new_n3799_), .Y(_abc_40319_new_n3806_));
INVX1 INVX1_65 ( .A(IR_REG_29_), .Y(_abc_40319_new_n708_));
INVX1 INVX1_650 ( .A(_abc_40319_new_n3813_), .Y(_abc_40319_new_n3814_));
INVX1 INVX1_651 ( .A(_abc_40319_new_n3812_), .Y(_abc_40319_new_n3817_));
INVX1 INVX1_652 ( .A(_abc_40319_new_n3811_), .Y(_abc_40319_new_n3818_));
INVX1 INVX1_653 ( .A(_abc_40319_new_n3832_), .Y(_abc_40319_new_n3833_));
INVX1 INVX1_654 ( .A(_abc_40319_new_n3835_), .Y(_abc_40319_new_n3836_));
INVX1 INVX1_655 ( .A(_abc_40319_new_n3831_), .Y(_abc_40319_new_n3838_));
INVX1 INVX1_656 ( .A(REG1_REG_8_), .Y(_abc_40319_new_n3843_));
INVX1 INVX1_657 ( .A(_abc_40319_new_n3846_), .Y(_abc_40319_new_n3847_));
INVX1 INVX1_658 ( .A(_abc_40319_new_n3845_), .Y(_abc_40319_new_n3850_));
INVX1 INVX1_659 ( .A(_abc_40319_new_n3865_), .Y(_abc_40319_new_n3866_));
INVX1 INVX1_66 ( .A(_abc_40319_new_n710_), .Y(_abc_40319_new_n712_));
INVX1 INVX1_660 ( .A(_abc_40319_new_n3868_), .Y(_abc_40319_new_n3869_));
INVX1 INVX1_661 ( .A(_abc_40319_new_n3870_), .Y(_abc_40319_new_n3871_));
INVX1 INVX1_662 ( .A(_abc_40319_new_n3876_), .Y(_abc_40319_new_n3877_));
INVX1 INVX1_663 ( .A(_abc_40319_new_n3879_), .Y(_abc_40319_new_n3882_));
INVX1 INVX1_664 ( .A(_abc_40319_new_n3880_), .Y(_abc_40319_new_n3883_));
INVX1 INVX1_665 ( .A(_abc_40319_new_n1754_), .Y(_abc_40319_new_n3897_));
INVX1 INVX1_666 ( .A(_abc_40319_new_n3878_), .Y(_abc_40319_new_n3899_));
INVX1 INVX1_667 ( .A(_abc_40319_new_n3901_), .Y(_abc_40319_new_n3902_));
INVX1 INVX1_668 ( .A(_abc_40319_new_n3903_), .Y(_abc_40319_new_n3904_));
INVX1 INVX1_669 ( .A(REG1_REG_10_), .Y(_abc_40319_new_n3905_));
INVX1 INVX1_67 ( .A(_abc_40319_new_n707_), .Y(_abc_40319_new_n724_));
INVX1 INVX1_670 ( .A(_abc_40319_new_n3906_), .Y(_abc_40319_new_n3907_));
INVX1 INVX1_671 ( .A(_abc_40319_new_n3908_), .Y(_abc_40319_new_n3909_));
INVX1 INVX1_672 ( .A(_abc_40319_new_n3922_), .Y(_abc_40319_new_n3923_));
INVX1 INVX1_673 ( .A(_abc_40319_new_n3925_), .Y(_abc_40319_new_n3929_));
INVX1 INVX1_674 ( .A(_abc_40319_new_n3927_), .Y(_abc_40319_new_n3930_));
INVX1 INVX1_675 ( .A(_abc_40319_new_n1720_), .Y(_abc_40319_new_n3940_));
INVX1 INVX1_676 ( .A(_abc_40319_new_n3941_), .Y(_abc_40319_new_n3942_));
INVX1 INVX1_677 ( .A(_abc_40319_new_n3944_), .Y(_abc_40319_new_n3945_));
INVX1 INVX1_678 ( .A(_abc_40319_new_n3947_), .Y(_abc_40319_new_n3948_));
INVX1 INVX1_679 ( .A(_abc_40319_new_n3955_), .Y(_abc_40319_new_n3956_));
INVX1 INVX1_68 ( .A(_abc_40319_new_n711_), .Y(_abc_40319_new_n725_));
INVX1 INVX1_680 ( .A(_abc_40319_new_n3958_), .Y(_abc_40319_new_n3959_));
INVX1 INVX1_681 ( .A(_abc_40319_new_n3961_), .Y(_abc_40319_new_n3963_));
INVX1 INVX1_682 ( .A(_abc_40319_new_n1686_), .Y(_abc_40319_new_n3976_));
INVX1 INVX1_683 ( .A(_abc_40319_new_n3977_), .Y(_abc_40319_new_n3978_));
INVX1 INVX1_684 ( .A(_abc_40319_new_n3980_), .Y(_abc_40319_new_n3981_));
INVX1 INVX1_685 ( .A(_abc_40319_new_n3943_), .Y(_abc_40319_new_n3982_));
INVX1 INVX1_686 ( .A(_abc_40319_new_n3984_), .Y(_abc_40319_new_n3985_));
INVX1 INVX1_687 ( .A(_abc_40319_new_n3990_), .Y(_abc_40319_new_n3991_));
INVX1 INVX1_688 ( .A(_abc_40319_new_n3993_), .Y(_abc_40319_new_n3994_));
INVX1 INVX1_689 ( .A(_abc_40319_new_n3996_), .Y(_abc_40319_new_n3998_));
INVX1 INVX1_69 ( .A(_abc_40319_new_n719_), .Y(_abc_40319_new_n730_));
INVX1 INVX1_690 ( .A(_abc_40319_new_n1651_), .Y(_abc_40319_new_n4011_));
INVX1 INVX1_691 ( .A(REG1_REG_13_), .Y(_abc_40319_new_n4012_));
INVX1 INVX1_692 ( .A(_abc_40319_new_n3979_), .Y(_abc_40319_new_n4013_));
INVX1 INVX1_693 ( .A(_abc_40319_new_n4016_), .Y(_abc_40319_new_n4017_));
INVX1 INVX1_694 ( .A(_abc_40319_new_n4015_), .Y(_abc_40319_new_n4018_));
INVX1 INVX1_695 ( .A(_abc_40319_new_n4019_), .Y(_abc_40319_new_n4020_));
INVX1 INVX1_696 ( .A(_abc_40319_new_n4021_), .Y(_abc_40319_new_n4022_));
INVX1 INVX1_697 ( .A(_abc_40319_new_n4027_), .Y(_abc_40319_new_n4028_));
INVX1 INVX1_698 ( .A(_abc_40319_new_n4030_), .Y(_abc_40319_new_n4034_));
INVX1 INVX1_699 ( .A(_abc_40319_new_n4032_), .Y(_abc_40319_new_n4035_));
INVX1 INVX1_7 ( .A(IR_REG_3_), .Y(_abc_40319_new_n532_));
INVX1 INVX1_70 ( .A(_abc_40319_new_n720_), .Y(_abc_40319_new_n731_));
INVX1 INVX1_700 ( .A(REG1_REG_14_), .Y(_abc_40319_new_n4048_));
INVX1 INVX1_701 ( .A(_abc_40319_new_n4052_), .Y(_abc_40319_new_n4053_));
INVX1 INVX1_702 ( .A(_abc_40319_new_n4051_), .Y(_abc_40319_new_n4056_));
INVX1 INVX1_703 ( .A(_abc_40319_new_n4061_), .Y(_abc_40319_new_n4062_));
INVX1 INVX1_704 ( .A(_abc_40319_new_n4064_), .Y(_abc_40319_new_n4065_));
INVX1 INVX1_705 ( .A(_abc_40319_new_n4067_), .Y(_abc_40319_new_n4068_));
INVX1 INVX1_706 ( .A(REG1_REG_15_), .Y(_abc_40319_new_n4084_));
INVX1 INVX1_707 ( .A(_abc_40319_new_n4086_), .Y(_abc_40319_new_n4087_));
INVX1 INVX1_708 ( .A(_abc_40319_new_n4085_), .Y(_abc_40319_new_n4088_));
INVX1 INVX1_709 ( .A(_abc_40319_new_n4089_), .Y(_abc_40319_new_n4090_));
INVX1 INVX1_71 ( .A(_abc_40319_new_n740_), .Y(_abc_40319_new_n741_));
INVX1 INVX1_710 ( .A(_abc_40319_new_n4091_), .Y(_abc_40319_new_n4093_));
INVX1 INVX1_711 ( .A(_abc_40319_new_n4098_), .Y(_abc_40319_new_n4099_));
INVX1 INVX1_712 ( .A(_abc_40319_new_n4101_), .Y(_abc_40319_new_n4102_));
INVX1 INVX1_713 ( .A(_abc_40319_new_n4104_), .Y(_abc_40319_new_n4105_));
INVX1 INVX1_714 ( .A(_abc_40319_new_n1394_), .Y(_abc_40319_new_n4120_));
INVX1 INVX1_715 ( .A(_abc_40319_new_n4121_), .Y(_abc_40319_new_n4122_));
INVX1 INVX1_716 ( .A(_abc_40319_new_n4124_), .Y(_abc_40319_new_n4125_));
INVX1 INVX1_717 ( .A(_abc_40319_new_n4127_), .Y(_abc_40319_new_n4128_));
INVX1 INVX1_718 ( .A(_abc_40319_new_n4133_), .Y(_abc_40319_new_n4134_));
INVX1 INVX1_719 ( .A(_abc_40319_new_n4136_), .Y(_abc_40319_new_n4137_));
INVX1 INVX1_72 ( .A(_abc_40319_new_n653_), .Y(_abc_40319_new_n749_));
INVX1 INVX1_720 ( .A(_abc_40319_new_n4139_), .Y(_abc_40319_new_n4140_));
INVX1 INVX1_721 ( .A(_abc_40319_new_n4156_), .Y(_abc_40319_new_n4157_));
INVX1 INVX1_722 ( .A(_abc_40319_new_n4159_), .Y(_abc_40319_new_n4160_));
INVX1 INVX1_723 ( .A(_abc_40319_new_n4162_), .Y(_abc_40319_new_n4164_));
INVX1 INVX1_724 ( .A(_abc_40319_new_n4169_), .Y(_abc_40319_new_n4170_));
INVX1 INVX1_725 ( .A(_abc_40319_new_n4172_), .Y(_abc_40319_new_n4173_));
INVX1 INVX1_726 ( .A(_abc_40319_new_n4175_), .Y(_abc_40319_new_n4176_));
INVX1 INVX1_727 ( .A(REG1_REG_18_), .Y(_abc_40319_new_n4191_));
INVX1 INVX1_728 ( .A(_abc_40319_new_n4192_), .Y(_abc_40319_new_n4193_));
INVX1 INVX1_729 ( .A(_abc_40319_new_n4194_), .Y(_abc_40319_new_n4195_));
INVX1 INVX1_73 ( .A(_abc_40319_new_n654_), .Y(_abc_40319_new_n750_));
INVX1 INVX1_730 ( .A(_abc_40319_new_n4196_), .Y(_abc_40319_new_n4197_));
INVX1 INVX1_731 ( .A(_abc_40319_new_n4199_), .Y(_abc_40319_new_n4201_));
INVX1 INVX1_732 ( .A(REG2_REG_18_), .Y(_abc_40319_new_n4205_));
INVX1 INVX1_733 ( .A(_abc_40319_new_n4206_), .Y(_abc_40319_new_n4207_));
INVX1 INVX1_734 ( .A(_abc_40319_new_n4208_), .Y(_abc_40319_new_n4209_));
INVX1 INVX1_735 ( .A(_abc_40319_new_n4210_), .Y(_abc_40319_new_n4214_));
INVX1 INVX1_736 ( .A(_abc_40319_new_n4212_), .Y(_abc_40319_new_n4215_));
INVX1 INVX1_737 ( .A(_abc_40319_new_n4231_), .Y(_abc_40319_new_n4232_));
INVX1 INVX1_738 ( .A(_abc_40319_new_n4234_), .Y(_abc_40319_new_n4235_));
INVX1 INVX1_739 ( .A(_abc_40319_new_n4236_), .Y(_abc_40319_new_n4237_));
INVX1 INVX1_74 ( .A(_abc_40319_new_n760_), .Y(_abc_40319_new_n761_));
INVX1 INVX1_740 ( .A(_abc_40319_new_n4243_), .Y(_abc_40319_new_n4244_));
INVX1 INVX1_741 ( .A(_abc_40319_new_n4245_), .Y(_abc_40319_new_n4246_));
INVX1 INVX1_742 ( .A(_abc_40319_new_n4248_), .Y(_abc_40319_new_n4250_));
INVX1 INVX1_743 ( .A(_abc_40319_new_n1112_), .Y(_abc_40319_new_n4265_));
INVX1 INVX1_744 ( .A(_abc_40319_new_n1159_), .Y(_abc_40319_new_n4267_));
INVX1 INVX1_745 ( .A(_abc_40319_new_n891_), .Y(_abc_40319_new_n4273_));
INVX1 INVX1_746 ( .A(_abc_40319_new_n4303_), .Y(_abc_40319_new_n4304_));
INVX1 INVX1_747 ( .A(_abc_40319_new_n4271_), .Y(_abc_40319_new_n4309_));
INVX1 INVX1_748 ( .A(_abc_40319_new_n4331_), .Y(_abc_40319_new_n4332_));
INVX1 INVX1_749 ( .A(_abc_40319_new_n4333_), .Y(_abc_40319_new_n4334_));
INVX1 INVX1_75 ( .A(_abc_40319_new_n757_), .Y(_abc_40319_new_n768_));
INVX1 INVX1_750 ( .A(_abc_40319_new_n4335_), .Y(_abc_40319_new_n4336_));
INVX1 INVX1_751 ( .A(_abc_40319_new_n4337_), .Y(_abc_40319_new_n4338_));
INVX1 INVX1_752 ( .A(_abc_40319_new_n4341_), .Y(_abc_40319_new_n4342_));
INVX1 INVX1_753 ( .A(_abc_40319_new_n4344_), .Y(_abc_40319_new_n4345_));
INVX1 INVX1_754 ( .A(_abc_40319_new_n4347_), .Y(_abc_40319_new_n4348_));
INVX1 INVX1_755 ( .A(_abc_40319_new_n4349_), .Y(_abc_40319_new_n4350_));
INVX1 INVX1_756 ( .A(_abc_40319_new_n4352_), .Y(_abc_40319_new_n4353_));
INVX1 INVX1_757 ( .A(_abc_40319_new_n3108_), .Y(_abc_40319_new_n4354_));
INVX1 INVX1_758 ( .A(_abc_40319_new_n4365_), .Y(_abc_40319_new_n4366_));
INVX1 INVX1_759 ( .A(_abc_40319_new_n4368_), .Y(_abc_40319_new_n4369_));
INVX1 INVX1_76 ( .A(_abc_40319_new_n766_), .Y(_abc_40319_new_n769_));
INVX1 INVX1_760 ( .A(_abc_40319_new_n4372_), .Y(_abc_40319_new_n4373_));
INVX1 INVX1_761 ( .A(_abc_40319_new_n4374_), .Y(_abc_40319_new_n4375_));
INVX1 INVX1_762 ( .A(_abc_40319_new_n4377_), .Y(_abc_40319_new_n4378_));
INVX1 INVX1_763 ( .A(_abc_40319_new_n4379_), .Y(_abc_40319_new_n4380_));
INVX1 INVX1_764 ( .A(_abc_40319_new_n4382_), .Y(_abc_40319_new_n4383_));
INVX1 INVX1_765 ( .A(_abc_40319_new_n4385_), .Y(_abc_40319_new_n4386_));
INVX1 INVX1_766 ( .A(_abc_40319_new_n4388_), .Y(_abc_40319_new_n4389_));
INVX1 INVX1_767 ( .A(_abc_40319_new_n4397_), .Y(_abc_40319_new_n4398_));
INVX1 INVX1_768 ( .A(_abc_40319_new_n4399_), .Y(_abc_40319_new_n4400_));
INVX1 INVX1_769 ( .A(_abc_40319_new_n4401_), .Y(_abc_40319_new_n4402_));
INVX1 INVX1_77 ( .A(_abc_40319_new_n775_), .Y(_abc_40319_new_n776_));
INVX1 INVX1_770 ( .A(_abc_40319_new_n4410_), .Y(_abc_40319_new_n4411_));
INVX1 INVX1_771 ( .A(_abc_40319_new_n4412_), .Y(_abc_40319_new_n4413_));
INVX1 INVX1_772 ( .A(_abc_40319_new_n4416_), .Y(_abc_40319_new_n4417_));
INVX1 INVX1_773 ( .A(_abc_40319_new_n4418_), .Y(_abc_40319_new_n4419_));
INVX1 INVX1_774 ( .A(_abc_40319_new_n4421_), .Y(_abc_40319_new_n4422_));
INVX1 INVX1_775 ( .A(_abc_40319_new_n4424_), .Y(_abc_40319_new_n4425_));
INVX1 INVX1_776 ( .A(_abc_40319_new_n4426_), .Y(_abc_40319_new_n4427_));
INVX1 INVX1_777 ( .A(_abc_40319_new_n4428_), .Y(_abc_40319_new_n4429_));
INVX1 INVX1_778 ( .A(_abc_40319_new_n4431_), .Y(_abc_40319_new_n4432_));
INVX1 INVX1_779 ( .A(_abc_40319_new_n4433_), .Y(_abc_40319_new_n4434_));
INVX1 INVX1_78 ( .A(_abc_40319_new_n779_), .Y(_abc_40319_new_n780_));
INVX1 INVX1_780 ( .A(_abc_40319_new_n4459_), .Y(_abc_40319_new_n4460_));
INVX1 INVX1_781 ( .A(_abc_40319_new_n4467_), .Y(_abc_40319_new_n4468_));
INVX1 INVX1_782 ( .A(_abc_40319_new_n4469_), .Y(_abc_40319_new_n4470_));
INVX1 INVX1_783 ( .A(_abc_40319_new_n4487_), .Y(_abc_40319_new_n4488_));
INVX1 INVX1_784 ( .A(_abc_40319_new_n4489_), .Y(_abc_40319_new_n4490_));
INVX1 INVX1_785 ( .A(_abc_40319_new_n3537_), .Y(_abc_40319_new_n4501_));
INVX1 INVX1_786 ( .A(_abc_40319_new_n4502_), .Y(_abc_40319_new_n4503_));
INVX1 INVX1_787 ( .A(_abc_40319_new_n4301_), .Y(_abc_40319_new_n4514_));
INVX1 INVX1_788 ( .A(_abc_40319_new_n4476_), .Y(_abc_40319_new_n4531_));
INVX1 INVX1_789 ( .A(_abc_40319_new_n4533_), .Y(_abc_40319_new_n4535_));
INVX1 INVX1_79 ( .A(_abc_40319_new_n781_), .Y(_abc_40319_new_n782_));
INVX1 INVX1_790 ( .A(_abc_40319_new_n3536_), .Y(_abc_40319_new_n4540_));
INVX1 INVX1_791 ( .A(_abc_40319_new_n4541_), .Y(_abc_40319_new_n4542_));
INVX1 INVX1_792 ( .A(_abc_40319_new_n4300_), .Y(_abc_40319_new_n4551_));
INVX1 INVX1_793 ( .A(_abc_40319_new_n4480_), .Y(_abc_40319_new_n4572_));
INVX1 INVX1_794 ( .A(_abc_40319_new_n4568_), .Y(_abc_40319_new_n4573_));
INVX1 INVX1_795 ( .A(_abc_40319_new_n4339_), .Y(_abc_40319_new_n4575_));
INVX1 INVX1_796 ( .A(_abc_40319_new_n4299_), .Y(_abc_40319_new_n4590_));
INVX1 INVX1_797 ( .A(_abc_40319_new_n4611_), .Y(_abc_40319_new_n4613_));
INVX1 INVX1_798 ( .A(_abc_40319_new_n4298_), .Y(_abc_40319_new_n4621_));
INVX1 INVX1_799 ( .A(_abc_40319_new_n4642_), .Y(_abc_40319_new_n4643_));
INVX1 INVX1_8 ( .A(IR_REG_5_), .Y(_abc_40319_new_n533_));
INVX1 INVX1_80 ( .A(_abc_40319_new_n739_), .Y(_abc_40319_new_n790_));
INVX1 INVX1_800 ( .A(_abc_40319_new_n4650_), .Y(_abc_40319_new_n4651_));
INVX1 INVX1_801 ( .A(_abc_40319_new_n4657_), .Y(_abc_40319_new_n4658_));
INVX1 INVX1_802 ( .A(_abc_40319_new_n4297_), .Y(_abc_40319_new_n4667_));
INVX1 INVX1_803 ( .A(_abc_40319_new_n4684_), .Y(_abc_40319_new_n4685_));
INVX1 INVX1_804 ( .A(_abc_40319_new_n4474_), .Y(_abc_40319_new_n4700_));
INVX1 INVX1_805 ( .A(_abc_40319_new_n4296_), .Y(_abc_40319_new_n4709_));
INVX1 INVX1_806 ( .A(_abc_40319_new_n4687_), .Y(_abc_40319_new_n4726_));
INVX1 INVX1_807 ( .A(_abc_40319_new_n4472_), .Y(_abc_40319_new_n4731_));
INVX1 INVX1_808 ( .A(_abc_40319_new_n4295_), .Y(_abc_40319_new_n4740_));
INVX1 INVX1_809 ( .A(_abc_40319_new_n4464_), .Y(_abc_40319_new_n4756_));
INVX1 INVX1_81 ( .A(_abc_40319_new_n800_), .Y(_abc_40319_new_n802_));
INVX1 INVX1_810 ( .A(_abc_40319_new_n4762_), .Y(_abc_40319_new_n4764_));
INVX1 INVX1_811 ( .A(_abc_40319_new_n4294_), .Y(_abc_40319_new_n4777_));
INVX1 INVX1_812 ( .A(_abc_40319_new_n4794_), .Y(_abc_40319_new_n4795_));
INVX1 INVX1_813 ( .A(_abc_40319_new_n3110_), .Y(_abc_40319_new_n4797_));
INVX1 INVX1_814 ( .A(_abc_40319_new_n4803_), .Y(_abc_40319_new_n4805_));
INVX1 INVX1_815 ( .A(_abc_40319_new_n4293_), .Y(_abc_40319_new_n4813_));
INVX1 INVX1_816 ( .A(_abc_40319_new_n4760_), .Y(_abc_40319_new_n4830_));
INVX1 INVX1_817 ( .A(_abc_40319_new_n4645_), .Y(_abc_40319_new_n4835_));
INVX1 INVX1_818 ( .A(_abc_40319_new_n4292_), .Y(_abc_40319_new_n4844_));
INVX1 INVX1_819 ( .A(_abc_40319_new_n4758_), .Y(_abc_40319_new_n4860_));
INVX1 INVX1_82 ( .A(_abc_40319_new_n804_), .Y(_abc_40319_new_n805_));
INVX1 INVX1_820 ( .A(_abc_40319_new_n4866_), .Y(_abc_40319_new_n4867_));
INVX1 INVX1_821 ( .A(_abc_40319_new_n4291_), .Y(_abc_40319_new_n4876_));
INVX1 INVX1_822 ( .A(_abc_40319_new_n4466_), .Y(_abc_40319_new_n4892_));
INVX1 INVX1_823 ( .A(_abc_40319_new_n4894_), .Y(_abc_40319_new_n4896_));
INVX1 INVX1_824 ( .A(_abc_40319_new_n4901_), .Y(_abc_40319_new_n4902_));
INVX1 INVX1_825 ( .A(_abc_40319_new_n4290_), .Y(_abc_40319_new_n4911_));
INVX1 INVX1_826 ( .A(_abc_40319_new_n3518_), .Y(_abc_40319_new_n4928_));
INVX1 INVX1_827 ( .A(_abc_40319_new_n4932_), .Y(_abc_40319_new_n4934_));
INVX1 INVX1_828 ( .A(_abc_40319_new_n4289_), .Y(_abc_40319_new_n4947_));
INVX1 INVX1_829 ( .A(_abc_40319_new_n4930_), .Y(_abc_40319_new_n4965_));
INVX1 INVX1_83 ( .A(_abc_40319_new_n809_), .Y(_abc_40319_new_n810_));
INVX1 INVX1_830 ( .A(_abc_40319_new_n4462_), .Y(_abc_40319_new_n4970_));
INVX1 INVX1_831 ( .A(_abc_40319_new_n4288_), .Y(_abc_40319_new_n4979_));
INVX1 INVX1_832 ( .A(_abc_40319_new_n4287_), .Y(_abc_40319_new_n5008_));
INVX1 INVX1_833 ( .A(_abc_40319_new_n3516_), .Y(_abc_40319_new_n5024_));
INVX1 INVX1_834 ( .A(_abc_40319_new_n5032_), .Y(_abc_40319_new_n5034_));
INVX1 INVX1_835 ( .A(_abc_40319_new_n4286_), .Y(_abc_40319_new_n5042_));
INVX1 INVX1_836 ( .A(_abc_40319_new_n3514_), .Y(_abc_40319_new_n5058_));
INVX1 INVX1_837 ( .A(_abc_40319_new_n5030_), .Y(_abc_40319_new_n5065_));
INVX1 INVX1_838 ( .A(_abc_40319_new_n4285_), .Y(_abc_40319_new_n5073_));
INVX1 INVX1_839 ( .A(_abc_40319_new_n3509_), .Y(_abc_40319_new_n5089_));
INVX1 INVX1_84 ( .A(_abc_40319_new_n813_), .Y(_abc_40319_new_n814_));
INVX1 INVX1_840 ( .A(_abc_40319_new_n5093_), .Y(_abc_40319_new_n5095_));
INVX1 INVX1_841 ( .A(_abc_40319_new_n4456_), .Y(_abc_40319_new_n5101_));
INVX1 INVX1_842 ( .A(_abc_40319_new_n4284_), .Y(_abc_40319_new_n5109_));
INVX1 INVX1_843 ( .A(_abc_40319_new_n5091_), .Y(_abc_40319_new_n5126_));
INVX1 INVX1_844 ( .A(_abc_40319_new_n5133_), .Y(_abc_40319_new_n5135_));
INVX1 INVX1_845 ( .A(_abc_40319_new_n4283_), .Y(_abc_40319_new_n5143_));
INVX1 INVX1_846 ( .A(_abc_40319_new_n5131_), .Y(_abc_40319_new_n5166_));
INVX1 INVX1_847 ( .A(_abc_40319_new_n4282_), .Y(_abc_40319_new_n5174_));
INVX1 INVX1_848 ( .A(_abc_40319_new_n5190_), .Y(_abc_40319_new_n5191_));
INVX1 INVX1_849 ( .A(_abc_40319_new_n4452_), .Y(_abc_40319_new_n5198_));
INVX1 INVX1_85 ( .A(DATAI_3_), .Y(_abc_40319_new_n816_));
INVX1 INVX1_850 ( .A(_abc_40319_new_n4281_), .Y(_abc_40319_new_n5206_));
INVX1 INVX1_851 ( .A(_abc_40319_new_n3505_), .Y(_abc_40319_new_n5222_));
INVX1 INVX1_852 ( .A(_abc_40319_new_n4450_), .Y(_abc_40319_new_n5229_));
INVX1 INVX1_853 ( .A(_abc_40319_new_n4280_), .Y(_abc_40319_new_n5237_));
INVX1 INVX1_854 ( .A(_abc_40319_new_n3495_), .Y(_abc_40319_new_n5253_));
INVX1 INVX1_855 ( .A(_abc_40319_new_n5255_), .Y(_abc_40319_new_n5256_));
INVX1 INVX1_856 ( .A(_abc_40319_new_n5258_), .Y(_abc_40319_new_n5259_));
INVX1 INVX1_857 ( .A(_abc_40319_new_n4448_), .Y(_abc_40319_new_n5266_));
INVX1 INVX1_858 ( .A(_abc_40319_new_n4279_), .Y(_abc_40319_new_n5274_));
INVX1 INVX1_859 ( .A(_abc_40319_new_n4439_), .Y(_abc_40319_new_n5295_));
INVX1 INVX1_86 ( .A(_abc_40319_new_n819_), .Y(_abc_40319_new_n820_));
INVX1 INVX1_860 ( .A(_abc_40319_new_n5296_), .Y(_abc_40319_new_n5297_));
INVX1 INVX1_861 ( .A(_abc_40319_new_n5299_), .Y(_abc_40319_new_n5300_));
INVX1 INVX1_862 ( .A(_abc_40319_new_n4277_), .Y(_abc_40319_new_n5315_));
INVX1 INVX1_863 ( .A(_abc_40319_new_n5331_), .Y(_abc_40319_new_n5332_));
INVX1 INVX1_864 ( .A(_abc_40319_new_n4278_), .Y(_abc_40319_new_n5345_));
INVX1 INVX1_865 ( .A(_abc_40319_new_n3493_), .Y(_abc_40319_new_n5357_));
INVX1 INVX1_866 ( .A(_abc_40319_new_n5362_), .Y(_abc_40319_new_n5363_));
INVX1 INVX1_867 ( .A(_abc_40319_new_n4276_), .Y(_abc_40319_new_n5376_));
INVX1 INVX1_868 ( .A(_abc_40319_new_n3491_), .Y(_abc_40319_new_n5392_));
INVX1 INVX1_869 ( .A(_abc_40319_new_n4275_), .Y(_abc_40319_new_n5404_));
INVX1 INVX1_87 ( .A(REG3_REG_3_), .Y(_abc_40319_new_n826_));
INVX1 INVX1_870 ( .A(_abc_40319_new_n3136_), .Y(_abc_40319_new_n5418_));
INVX1 INVX1_871 ( .A(_abc_40319_new_n4274_), .Y(_abc_40319_new_n5430_));
INVX1 INVX1_872 ( .A(_abc_40319_new_n5468_), .Y(_abc_40319_new_n5469_));
INVX1 INVX1_873 ( .A(_abc_40319_new_n643_), .Y(_abc_40319_new_n5547_));
INVX1 INVX1_874 ( .A(_abc_40319_new_n1392_), .Y(_abc_40319_new_n5584_));
INVX1 INVX1_875 ( .A(_abc_40319_new_n1649_), .Y(_abc_40319_new_n5603_));
INVX1 INVX1_876 ( .A(_abc_40319_new_n1684_), .Y(_abc_40319_new_n5610_));
INVX1 INVX1_877 ( .A(_abc_40319_new_n1718_), .Y(_abc_40319_new_n5617_));
INVX1 INVX1_878 ( .A(_abc_40319_new_n1752_), .Y(_abc_40319_new_n5624_));
INVX1 INVX1_879 ( .A(_abc_40319_new_n3103_), .Y(_abc_40319_new_n5691_));
INVX1 INVX1_88 ( .A(_abc_40319_new_n831_), .Y(_abc_40319_new_n832_));
INVX1 INVX1_880 ( .A(_abc_40319_new_n3539_), .Y(_abc_40319_new_n5692_));
INVX1 INVX1_881 ( .A(_abc_40319_new_n5697_), .Y(_abc_40319_new_n5698_));
INVX1 INVX1_882 ( .A(_abc_40319_new_n5700_), .Y(_abc_40319_new_n5702_));
INVX1 INVX1_883 ( .A(_abc_40319_new_n4302_), .Y(_abc_40319_new_n5716_));
INVX1 INVX1_884 ( .A(_abc_40319_new_n1076_), .Y(_abc_40319_new_n5740_));
INVX1 INVX1_885 ( .A(_abc_40319_new_n1168_), .Y(_abc_40319_new_n5741_));
INVX1 INVX1_886 ( .A(_abc_40319_new_n5744_), .Y(_abc_40319_new_n5753_));
INVX1 INVX1_887 ( .A(_abc_40319_new_n6057_), .Y(_abc_40319_new_n6059_));
INVX1 INVX1_888 ( .A(_abc_40319_new_n615_), .Y(_abc_40319_new_n6188_));
INVX1 INVX1_89 ( .A(_abc_40319_new_n841_), .Y(_abc_40319_new_n842_));
INVX1 INVX1_9 ( .A(IR_REG_4_), .Y(_abc_40319_new_n534_));
INVX1 INVX1_90 ( .A(DATAI_2_), .Y(_abc_40319_new_n845_));
INVX1 INVX1_91 ( .A(_abc_40319_new_n847_), .Y(_abc_40319_new_n848_));
INVX1 INVX1_92 ( .A(REG3_REG_2_), .Y(_abc_40319_new_n850_));
INVX1 INVX1_93 ( .A(REG1_REG_2_), .Y(_abc_40319_new_n853_));
INVX1 INVX1_94 ( .A(REG0_REG_2_), .Y(_abc_40319_new_n857_));
INVX1 INVX1_95 ( .A(REG2_REG_2_), .Y(_abc_40319_new_n860_));
INVX1 INVX1_96 ( .A(_abc_40319_new_n864_), .Y(_abc_40319_new_n865_));
INVX1 INVX1_97 ( .A(_abc_40319_new_n868_), .Y(_abc_40319_new_n872_));
INVX1 INVX1_98 ( .A(_abc_40319_new_n869_), .Y(_abc_40319_new_n873_));
INVX1 INVX1_99 ( .A(_abc_40319_new_n882_), .Y(_abc_40319_new_n883_));
OR2X2 OR2X2_1 ( .A(IR_REG_0_), .B(IR_REG_1_), .Y(_abc_40319_new_n529_));
OR2X2 OR2X2_10 ( .A(_abc_40319_new_n603_), .B(_abc_40319_new_n604_), .Y(_abc_40319_new_n605_));
OR2X2 OR2X2_100 ( .A(_abc_40319_new_n922_), .B(_abc_40319_new_n921_), .Y(_abc_40319_new_n923_));
OR2X2 OR2X2_1000 ( .A(_abc_40319_new_n3758_), .B(_abc_40319_new_n3759_), .Y(_abc_40319_new_n3760_));
OR2X2 OR2X2_1001 ( .A(_abc_40319_new_n3760_), .B(_abc_40319_new_n3745_), .Y(_abc_40319_new_n3761_));
OR2X2 OR2X2_1002 ( .A(_abc_40319_new_n3763_), .B(_abc_40319_new_n2276_), .Y(_abc_40319_new_n3764_));
OR2X2 OR2X2_1003 ( .A(_abc_40319_new_n3762_), .B(_abc_40319_new_n3764_), .Y(n1034));
OR2X2 OR2X2_1004 ( .A(_abc_40319_new_n3767_), .B(_abc_40319_new_n3748_), .Y(_abc_40319_new_n3768_));
OR2X2 OR2X2_1005 ( .A(_abc_40319_new_n993_), .B(REG2_REG_6_), .Y(_abc_40319_new_n3770_));
OR2X2 OR2X2_1006 ( .A(_abc_40319_new_n3772_), .B(_abc_40319_new_n3766_), .Y(_abc_40319_new_n3773_));
OR2X2 OR2X2_1007 ( .A(_abc_40319_new_n3769_), .B(_abc_40319_new_n3775_), .Y(_abc_40319_new_n3776_));
OR2X2 OR2X2_1008 ( .A(_abc_40319_new_n3738_), .B(_abc_40319_new_n685_), .Y(_abc_40319_new_n3780_));
OR2X2 OR2X2_1009 ( .A(_abc_40319_new_n993_), .B(REG1_REG_6_), .Y(_abc_40319_new_n3782_));
OR2X2 OR2X2_101 ( .A(_abc_40319_new_n920_), .B(_abc_40319_new_n923_), .Y(_abc_40319_new_n924_));
OR2X2 OR2X2_1010 ( .A(_abc_40319_new_n3781_), .B(_abc_40319_new_n3783_), .Y(_abc_40319_new_n3784_));
OR2X2 OR2X2_1011 ( .A(_abc_40319_new_n3784_), .B(_abc_40319_new_n3779_), .Y(_abc_40319_new_n3785_));
OR2X2 OR2X2_1012 ( .A(_abc_40319_new_n3786_), .B(_abc_40319_new_n3788_), .Y(_abc_40319_new_n3789_));
OR2X2 OR2X2_1013 ( .A(_abc_40319_new_n3791_), .B(_abc_40319_new_n3792_), .Y(_abc_40319_new_n3793_));
OR2X2 OR2X2_1014 ( .A(_abc_40319_new_n3778_), .B(_abc_40319_new_n3793_), .Y(_abc_40319_new_n3794_));
OR2X2 OR2X2_1015 ( .A(_abc_40319_new_n3796_), .B(_abc_40319_new_n2503_), .Y(_abc_40319_new_n3797_));
OR2X2 OR2X2_1016 ( .A(_abc_40319_new_n3795_), .B(_abc_40319_new_n3797_), .Y(n1030));
OR2X2 OR2X2_1017 ( .A(_abc_40319_new_n1029_), .B(REG2_REG_7_), .Y(_abc_40319_new_n3802_));
OR2X2 OR2X2_1018 ( .A(_abc_40319_new_n3804_), .B(_abc_40319_new_n3799_), .Y(_abc_40319_new_n3805_));
OR2X2 OR2X2_1019 ( .A(_abc_40319_new_n3801_), .B(_abc_40319_new_n3807_), .Y(_abc_40319_new_n3808_));
OR2X2 OR2X2_102 ( .A(_abc_40319_new_n817_), .B(IR_REG_0_), .Y(_abc_40319_new_n926_));
OR2X2 OR2X2_1020 ( .A(_abc_40319_new_n1029_), .B(REG1_REG_7_), .Y(_abc_40319_new_n3813_));
OR2X2 OR2X2_1021 ( .A(_abc_40319_new_n3812_), .B(_abc_40319_new_n3814_), .Y(_abc_40319_new_n3815_));
OR2X2 OR2X2_1022 ( .A(_abc_40319_new_n3815_), .B(_abc_40319_new_n3811_), .Y(_abc_40319_new_n3816_));
OR2X2 OR2X2_1023 ( .A(_abc_40319_new_n3817_), .B(_abc_40319_new_n3819_), .Y(_abc_40319_new_n3820_));
OR2X2 OR2X2_1024 ( .A(_abc_40319_new_n3822_), .B(_abc_40319_new_n3823_), .Y(_abc_40319_new_n3824_));
OR2X2 OR2X2_1025 ( .A(_abc_40319_new_n3810_), .B(_abc_40319_new_n3824_), .Y(_abc_40319_new_n3825_));
OR2X2 OR2X2_1026 ( .A(_abc_40319_new_n3827_), .B(_abc_40319_new_n1175_), .Y(_abc_40319_new_n3828_));
OR2X2 OR2X2_1027 ( .A(_abc_40319_new_n3826_), .B(_abc_40319_new_n3828_), .Y(n1026));
OR2X2 OR2X2_1028 ( .A(_abc_40319_new_n1567_), .B(REG2_REG_8_), .Y(_abc_40319_new_n3834_));
OR2X2 OR2X2_1029 ( .A(_abc_40319_new_n3836_), .B(_abc_40319_new_n3831_), .Y(_abc_40319_new_n3837_));
OR2X2 OR2X2_103 ( .A(_abc_40319_new_n931_), .B(_abc_40319_new_n932_), .Y(_abc_40319_new_n933_));
OR2X2 OR2X2_1030 ( .A(_abc_40319_new_n3833_), .B(_abc_40319_new_n3839_), .Y(_abc_40319_new_n3840_));
OR2X2 OR2X2_1031 ( .A(_abc_40319_new_n3844_), .B(_abc_40319_new_n3843_), .Y(_abc_40319_new_n3846_));
OR2X2 OR2X2_1032 ( .A(_abc_40319_new_n3847_), .B(_abc_40319_new_n3845_), .Y(_abc_40319_new_n3848_));
OR2X2 OR2X2_1033 ( .A(_abc_40319_new_n3849_), .B(_abc_40319_new_n3852_), .Y(_abc_40319_new_n3853_));
OR2X2 OR2X2_1034 ( .A(_abc_40319_new_n3842_), .B(_abc_40319_new_n3854_), .Y(_abc_40319_new_n3855_));
OR2X2 OR2X2_1035 ( .A(_abc_40319_new_n3855_), .B(_abc_40319_new_n3830_), .Y(_abc_40319_new_n3856_));
OR2X2 OR2X2_1036 ( .A(_abc_40319_new_n3860_), .B(_abc_40319_new_n2152_), .Y(_abc_40319_new_n3861_));
OR2X2 OR2X2_1037 ( .A(_abc_40319_new_n3861_), .B(_abc_40319_new_n3859_), .Y(_abc_40319_new_n3862_));
OR2X2 OR2X2_1038 ( .A(_abc_40319_new_n3858_), .B(_abc_40319_new_n3862_), .Y(_abc_40319_new_n3863_));
OR2X2 OR2X2_1039 ( .A(_abc_40319_new_n3863_), .B(_abc_40319_new_n3857_), .Y(n1022));
OR2X2 OR2X2_104 ( .A(_abc_40319_new_n933_), .B(_abc_40319_new_n925_), .Y(_abc_40319_new_n934_));
OR2X2 OR2X2_1040 ( .A(_abc_40319_new_n1609_), .B(REG2_REG_9_), .Y(_abc_40319_new_n3867_));
OR2X2 OR2X2_1041 ( .A(_abc_40319_new_n3872_), .B(_abc_40319_new_n3873_), .Y(_abc_40319_new_n3874_));
OR2X2 OR2X2_1042 ( .A(_abc_40319_new_n1609_), .B(REG1_REG_9_), .Y(_abc_40319_new_n3878_));
OR2X2 OR2X2_1043 ( .A(_abc_40319_new_n3851_), .B(_abc_40319_new_n3845_), .Y(_abc_40319_new_n3880_));
OR2X2 OR2X2_1044 ( .A(_abc_40319_new_n3884_), .B(_abc_40319_new_n3881_), .Y(_abc_40319_new_n3885_));
OR2X2 OR2X2_1045 ( .A(_abc_40319_new_n3875_), .B(_abc_40319_new_n3886_), .Y(_abc_40319_new_n3887_));
OR2X2 OR2X2_1046 ( .A(_abc_40319_new_n3889_), .B(_abc_40319_new_n3891_), .Y(_abc_40319_new_n3892_));
OR2X2 OR2X2_1047 ( .A(_abc_40319_new_n3893_), .B(_abc_40319_new_n2352_), .Y(_abc_40319_new_n3894_));
OR2X2 OR2X2_1048 ( .A(_abc_40319_new_n3892_), .B(_abc_40319_new_n3894_), .Y(_abc_40319_new_n3895_));
OR2X2 OR2X2_1049 ( .A(_abc_40319_new_n3888_), .B(_abc_40319_new_n3895_), .Y(n1018));
OR2X2 OR2X2_105 ( .A(_abc_40319_new_n934_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n935_));
OR2X2 OR2X2_1050 ( .A(_abc_40319_new_n3880_), .B(_abc_40319_new_n3899_), .Y(_abc_40319_new_n3900_));
OR2X2 OR2X2_1051 ( .A(_abc_40319_new_n3909_), .B(_abc_40319_new_n1754_), .Y(_abc_40319_new_n3910_));
OR2X2 OR2X2_1052 ( .A(_abc_40319_new_n3908_), .B(_abc_40319_new_n3897_), .Y(_abc_40319_new_n3911_));
OR2X2 OR2X2_1053 ( .A(_abc_40319_new_n3913_), .B(_abc_40319_new_n3898_), .Y(_abc_40319_new_n3914_));
OR2X2 OR2X2_1054 ( .A(_abc_40319_new_n3919_), .B(_abc_40319_new_n2042_), .Y(_abc_40319_new_n3920_));
OR2X2 OR2X2_1055 ( .A(_abc_40319_new_n3920_), .B(_abc_40319_new_n3918_), .Y(_abc_40319_new_n3921_));
OR2X2 OR2X2_1056 ( .A(_abc_40319_new_n3897_), .B(REG2_REG_10_), .Y(_abc_40319_new_n3924_));
OR2X2 OR2X2_1057 ( .A(_abc_40319_new_n3926_), .B(_abc_40319_new_n3865_), .Y(_abc_40319_new_n3927_));
OR2X2 OR2X2_1058 ( .A(_abc_40319_new_n3927_), .B(_abc_40319_new_n3925_), .Y(_abc_40319_new_n3928_));
OR2X2 OR2X2_1059 ( .A(_abc_40319_new_n3930_), .B(_abc_40319_new_n3929_), .Y(_abc_40319_new_n3931_));
OR2X2 OR2X2_106 ( .A(_abc_40319_new_n760_), .B(_abc_40319_new_n598_), .Y(_abc_40319_new_n938_));
OR2X2 OR2X2_1060 ( .A(_abc_40319_new_n3932_), .B(_abc_40319_new_n3933_), .Y(_abc_40319_new_n3934_));
OR2X2 OR2X2_1061 ( .A(_abc_40319_new_n3936_), .B(_abc_40319_new_n3921_), .Y(_abc_40319_new_n3937_));
OR2X2 OR2X2_1062 ( .A(_abc_40319_new_n3937_), .B(_abc_40319_new_n3917_), .Y(_abc_40319_new_n3938_));
OR2X2 OR2X2_1063 ( .A(_abc_40319_new_n3938_), .B(_abc_40319_new_n3915_), .Y(n1014));
OR2X2 OR2X2_1064 ( .A(_abc_40319_new_n3940_), .B(REG1_REG_11_), .Y(_abc_40319_new_n3943_));
OR2X2 OR2X2_1065 ( .A(_abc_40319_new_n3906_), .B(_abc_40319_new_n1754_), .Y(_abc_40319_new_n3946_));
OR2X2 OR2X2_1066 ( .A(_abc_40319_new_n3949_), .B(_abc_40319_new_n3950_), .Y(_abc_40319_new_n3951_));
OR2X2 OR2X2_1067 ( .A(_abc_40319_new_n3916_), .B(_abc_40319_new_n3952_), .Y(_abc_40319_new_n3953_));
OR2X2 OR2X2_1068 ( .A(_abc_40319_new_n3940_), .B(REG2_REG_11_), .Y(_abc_40319_new_n3957_));
OR2X2 OR2X2_1069 ( .A(_abc_40319_new_n3960_), .B(_abc_40319_new_n3922_), .Y(_abc_40319_new_n3961_));
OR2X2 OR2X2_107 ( .A(_abc_40319_new_n941_), .B(_abc_40319_new_n928_), .Y(_abc_40319_new_n942_));
OR2X2 OR2X2_1070 ( .A(_abc_40319_new_n3964_), .B(_abc_40319_new_n3962_), .Y(_abc_40319_new_n3965_));
OR2X2 OR2X2_1071 ( .A(_abc_40319_new_n3967_), .B(_abc_40319_new_n2448_), .Y(_abc_40319_new_n3968_));
OR2X2 OR2X2_1072 ( .A(_abc_40319_new_n3970_), .B(_abc_40319_new_n3971_), .Y(_abc_40319_new_n3972_));
OR2X2 OR2X2_1073 ( .A(_abc_40319_new_n3968_), .B(_abc_40319_new_n3972_), .Y(_abc_40319_new_n3973_));
OR2X2 OR2X2_1074 ( .A(_abc_40319_new_n3966_), .B(_abc_40319_new_n3973_), .Y(_abc_40319_new_n3974_));
OR2X2 OR2X2_1075 ( .A(_abc_40319_new_n3974_), .B(_abc_40319_new_n3954_), .Y(n1010));
OR2X2 OR2X2_1076 ( .A(_abc_40319_new_n3976_), .B(REG1_REG_12_), .Y(_abc_40319_new_n3979_));
OR2X2 OR2X2_1077 ( .A(_abc_40319_new_n3947_), .B(_abc_40319_new_n3982_), .Y(_abc_40319_new_n3983_));
OR2X2 OR2X2_1078 ( .A(_abc_40319_new_n3986_), .B(_abc_40319_new_n3987_), .Y(_abc_40319_new_n3988_));
OR2X2 OR2X2_1079 ( .A(_abc_40319_new_n3976_), .B(REG2_REG_12_), .Y(_abc_40319_new_n3992_));
OR2X2 OR2X2_108 ( .A(_abc_40319_new_n942_), .B(_abc_40319_new_n939_), .Y(_abc_40319_new_n943_));
OR2X2 OR2X2_1080 ( .A(_abc_40319_new_n3995_), .B(_abc_40319_new_n3955_), .Y(_abc_40319_new_n3996_));
OR2X2 OR2X2_1081 ( .A(_abc_40319_new_n3999_), .B(_abc_40319_new_n3997_), .Y(_abc_40319_new_n4000_));
OR2X2 OR2X2_1082 ( .A(_abc_40319_new_n4002_), .B(_abc_40319_new_n2220_), .Y(_abc_40319_new_n4003_));
OR2X2 OR2X2_1083 ( .A(_abc_40319_new_n4005_), .B(_abc_40319_new_n4006_), .Y(_abc_40319_new_n4007_));
OR2X2 OR2X2_1084 ( .A(_abc_40319_new_n4003_), .B(_abc_40319_new_n4007_), .Y(_abc_40319_new_n4008_));
OR2X2 OR2X2_1085 ( .A(_abc_40319_new_n4001_), .B(_abc_40319_new_n4008_), .Y(_abc_40319_new_n4009_));
OR2X2 OR2X2_1086 ( .A(_abc_40319_new_n4009_), .B(_abc_40319_new_n3989_), .Y(n1006));
OR2X2 OR2X2_1087 ( .A(_abc_40319_new_n3984_), .B(_abc_40319_new_n4013_), .Y(_abc_40319_new_n4014_));
OR2X2 OR2X2_1088 ( .A(_abc_40319_new_n4023_), .B(_abc_40319_new_n4024_), .Y(_abc_40319_new_n4025_));
OR2X2 OR2X2_1089 ( .A(_abc_40319_new_n4011_), .B(REG2_REG_13_), .Y(_abc_40319_new_n4029_));
OR2X2 OR2X2_109 ( .A(_abc_40319_new_n861_), .B(_abc_40319_new_n944_), .Y(_abc_40319_new_n945_));
OR2X2 OR2X2_1090 ( .A(_abc_40319_new_n4031_), .B(_abc_40319_new_n3990_), .Y(_abc_40319_new_n4032_));
OR2X2 OR2X2_1091 ( .A(_abc_40319_new_n4032_), .B(_abc_40319_new_n4030_), .Y(_abc_40319_new_n4033_));
OR2X2 OR2X2_1092 ( .A(_abc_40319_new_n4035_), .B(_abc_40319_new_n4034_), .Y(_abc_40319_new_n4036_));
OR2X2 OR2X2_1093 ( .A(_abc_40319_new_n4039_), .B(_abc_40319_new_n4041_), .Y(_abc_40319_new_n4042_));
OR2X2 OR2X2_1094 ( .A(_abc_40319_new_n4043_), .B(_abc_40319_new_n2412_), .Y(_abc_40319_new_n4044_));
OR2X2 OR2X2_1095 ( .A(_abc_40319_new_n4042_), .B(_abc_40319_new_n4044_), .Y(_abc_40319_new_n4045_));
OR2X2 OR2X2_1096 ( .A(_abc_40319_new_n4038_), .B(_abc_40319_new_n4045_), .Y(_abc_40319_new_n4046_));
OR2X2 OR2X2_1097 ( .A(_abc_40319_new_n4046_), .B(_abc_40319_new_n4026_), .Y(n1002));
OR2X2 OR2X2_1098 ( .A(_abc_40319_new_n4016_), .B(_abc_40319_new_n1651_), .Y(_abc_40319_new_n4049_));
OR2X2 OR2X2_1099 ( .A(_abc_40319_new_n4050_), .B(_abc_40319_new_n4048_), .Y(_abc_40319_new_n4052_));
OR2X2 OR2X2_11 ( .A(_abc_40319_new_n602_), .B(_abc_40319_new_n605_), .Y(_abc_40319_new_n606_));
OR2X2 OR2X2_110 ( .A(_abc_40319_new_n858_), .B(_abc_40319_new_n946_), .Y(_abc_40319_new_n947_));
OR2X2 OR2X2_1100 ( .A(_abc_40319_new_n4053_), .B(_abc_40319_new_n4051_), .Y(_abc_40319_new_n4054_));
OR2X2 OR2X2_1101 ( .A(_abc_40319_new_n4055_), .B(_abc_40319_new_n4058_), .Y(_abc_40319_new_n4059_));
OR2X2 OR2X2_1102 ( .A(_abc_40319_new_n1501_), .B(REG2_REG_14_), .Y(_abc_40319_new_n4063_));
OR2X2 OR2X2_1103 ( .A(_abc_40319_new_n4066_), .B(_abc_40319_new_n4027_), .Y(_abc_40319_new_n4067_));
OR2X2 OR2X2_1104 ( .A(_abc_40319_new_n4068_), .B(_abc_40319_new_n4065_), .Y(_abc_40319_new_n4069_));
OR2X2 OR2X2_1105 ( .A(_abc_40319_new_n4067_), .B(_abc_40319_new_n4064_), .Y(_abc_40319_new_n4070_));
OR2X2 OR2X2_1106 ( .A(_abc_40319_new_n4075_), .B(_abc_40319_new_n2005_), .Y(_abc_40319_new_n4076_));
OR2X2 OR2X2_1107 ( .A(_abc_40319_new_n4076_), .B(_abc_40319_new_n4073_), .Y(_abc_40319_new_n4077_));
OR2X2 OR2X2_1108 ( .A(_abc_40319_new_n4072_), .B(_abc_40319_new_n4077_), .Y(_abc_40319_new_n4078_));
OR2X2 OR2X2_1109 ( .A(_abc_40319_new_n4079_), .B(_abc_40319_new_n4074_), .Y(_abc_40319_new_n4080_));
OR2X2 OR2X2_111 ( .A(_abc_40319_new_n851_), .B(_abc_40319_new_n949_), .Y(_abc_40319_new_n950_));
OR2X2 OR2X2_1110 ( .A(_abc_40319_new_n4081_), .B(_abc_40319_new_n4078_), .Y(_abc_40319_new_n4082_));
OR2X2 OR2X2_1111 ( .A(_abc_40319_new_n4082_), .B(_abc_40319_new_n4060_), .Y(n998));
OR2X2 OR2X2_1112 ( .A(_abc_40319_new_n4057_), .B(_abc_40319_new_n4051_), .Y(_abc_40319_new_n4085_));
OR2X2 OR2X2_1113 ( .A(_abc_40319_new_n4091_), .B(_abc_40319_new_n1466_), .Y(_abc_40319_new_n4092_));
OR2X2 OR2X2_1114 ( .A(_abc_40319_new_n4093_), .B(_abc_40319_new_n1467_), .Y(_abc_40319_new_n4094_));
OR2X2 OR2X2_1115 ( .A(_abc_40319_new_n1466_), .B(REG2_REG_15_), .Y(_abc_40319_new_n4100_));
OR2X2 OR2X2_1116 ( .A(_abc_40319_new_n4103_), .B(_abc_40319_new_n4061_), .Y(_abc_40319_new_n4104_));
OR2X2 OR2X2_1117 ( .A(_abc_40319_new_n4105_), .B(_abc_40319_new_n4102_), .Y(_abc_40319_new_n4106_));
OR2X2 OR2X2_1118 ( .A(_abc_40319_new_n4104_), .B(_abc_40319_new_n4101_), .Y(_abc_40319_new_n4107_));
OR2X2 OR2X2_1119 ( .A(_abc_40319_new_n4109_), .B(_abc_40319_new_n4097_), .Y(_abc_40319_new_n4110_));
OR2X2 OR2X2_112 ( .A(_abc_40319_new_n854_), .B(_abc_40319_new_n951_), .Y(_abc_40319_new_n952_));
OR2X2 OR2X2_1120 ( .A(_abc_40319_new_n4114_), .B(_abc_40319_new_n2543_), .Y(_abc_40319_new_n4115_));
OR2X2 OR2X2_1121 ( .A(_abc_40319_new_n4115_), .B(_abc_40319_new_n4113_), .Y(_abc_40319_new_n4116_));
OR2X2 OR2X2_1122 ( .A(_abc_40319_new_n4112_), .B(_abc_40319_new_n4116_), .Y(_abc_40319_new_n4117_));
OR2X2 OR2X2_1123 ( .A(_abc_40319_new_n4111_), .B(_abc_40319_new_n4117_), .Y(_abc_40319_new_n4118_));
OR2X2 OR2X2_1124 ( .A(_abc_40319_new_n4118_), .B(_abc_40319_new_n4096_), .Y(n994));
OR2X2 OR2X2_1125 ( .A(_abc_40319_new_n4120_), .B(REG1_REG_16_), .Y(_abc_40319_new_n4123_));
OR2X2 OR2X2_1126 ( .A(_abc_40319_new_n4086_), .B(_abc_40319_new_n1467_), .Y(_abc_40319_new_n4126_));
OR2X2 OR2X2_1127 ( .A(_abc_40319_new_n4129_), .B(_abc_40319_new_n4130_), .Y(_abc_40319_new_n4131_));
OR2X2 OR2X2_1128 ( .A(_abc_40319_new_n4120_), .B(REG2_REG_16_), .Y(_abc_40319_new_n4135_));
OR2X2 OR2X2_1129 ( .A(_abc_40319_new_n4138_), .B(_abc_40319_new_n4098_), .Y(_abc_40319_new_n4139_));
OR2X2 OR2X2_113 ( .A(_abc_40319_new_n954_), .B(_abc_40319_new_n909_), .Y(_abc_40319_new_n955_));
OR2X2 OR2X2_1130 ( .A(_abc_40319_new_n4140_), .B(_abc_40319_new_n4137_), .Y(_abc_40319_new_n4141_));
OR2X2 OR2X2_1131 ( .A(_abc_40319_new_n4139_), .B(_abc_40319_new_n4136_), .Y(_abc_40319_new_n4142_));
OR2X2 OR2X2_1132 ( .A(_abc_40319_new_n4147_), .B(_abc_40319_new_n4146_), .Y(_abc_40319_new_n4148_));
OR2X2 OR2X2_1133 ( .A(_abc_40319_new_n4148_), .B(_abc_40319_new_n2258_), .Y(_abc_40319_new_n4149_));
OR2X2 OR2X2_1134 ( .A(_abc_40319_new_n4144_), .B(_abc_40319_new_n4149_), .Y(_abc_40319_new_n4150_));
OR2X2 OR2X2_1135 ( .A(_abc_40319_new_n4151_), .B(_abc_40319_new_n4145_), .Y(_abc_40319_new_n4152_));
OR2X2 OR2X2_1136 ( .A(_abc_40319_new_n4153_), .B(_abc_40319_new_n4150_), .Y(_abc_40319_new_n4154_));
OR2X2 OR2X2_1137 ( .A(_abc_40319_new_n4154_), .B(_abc_40319_new_n4132_), .Y(n990));
OR2X2 OR2X2_1138 ( .A(_abc_40319_new_n1428_), .B(REG1_REG_17_), .Y(_abc_40319_new_n4158_));
OR2X2 OR2X2_1139 ( .A(_abc_40319_new_n4161_), .B(_abc_40319_new_n4121_), .Y(_abc_40319_new_n4162_));
OR2X2 OR2X2_114 ( .A(_abc_40319_new_n956_), .B(_abc_40319_new_n768_), .Y(_abc_40319_new_n957_));
OR2X2 OR2X2_1140 ( .A(_abc_40319_new_n4165_), .B(_abc_40319_new_n4163_), .Y(_abc_40319_new_n4166_));
OR2X2 OR2X2_1141 ( .A(_abc_40319_new_n1428_), .B(REG2_REG_17_), .Y(_abc_40319_new_n4171_));
OR2X2 OR2X2_1142 ( .A(_abc_40319_new_n4174_), .B(_abc_40319_new_n4133_), .Y(_abc_40319_new_n4175_));
OR2X2 OR2X2_1143 ( .A(_abc_40319_new_n4176_), .B(_abc_40319_new_n4173_), .Y(_abc_40319_new_n4177_));
OR2X2 OR2X2_1144 ( .A(_abc_40319_new_n4175_), .B(_abc_40319_new_n4172_), .Y(_abc_40319_new_n4178_));
OR2X2 OR2X2_1145 ( .A(_abc_40319_new_n4180_), .B(_abc_40319_new_n4168_), .Y(_abc_40319_new_n4181_));
OR2X2 OR2X2_1146 ( .A(_abc_40319_new_n4185_), .B(_abc_40319_new_n2297_), .Y(_abc_40319_new_n4186_));
OR2X2 OR2X2_1147 ( .A(_abc_40319_new_n4186_), .B(_abc_40319_new_n4184_), .Y(_abc_40319_new_n4187_));
OR2X2 OR2X2_1148 ( .A(_abc_40319_new_n4183_), .B(_abc_40319_new_n4187_), .Y(_abc_40319_new_n4188_));
OR2X2 OR2X2_1149 ( .A(_abc_40319_new_n4182_), .B(_abc_40319_new_n4188_), .Y(_abc_40319_new_n4189_));
OR2X2 OR2X2_115 ( .A(_abc_40319_new_n958_), .B(_abc_40319_new_n959_), .Y(_abc_40319_new_n960_));
OR2X2 OR2X2_1150 ( .A(_abc_40319_new_n4189_), .B(_abc_40319_new_n4167_), .Y(n986));
OR2X2 OR2X2_1151 ( .A(_abc_40319_new_n4198_), .B(_abc_40319_new_n4156_), .Y(_abc_40319_new_n4199_));
OR2X2 OR2X2_1152 ( .A(_abc_40319_new_n4202_), .B(_abc_40319_new_n4200_), .Y(_abc_40319_new_n4203_));
OR2X2 OR2X2_1153 ( .A(_abc_40319_new_n4211_), .B(_abc_40319_new_n4169_), .Y(_abc_40319_new_n4212_));
OR2X2 OR2X2_1154 ( .A(_abc_40319_new_n4212_), .B(_abc_40319_new_n4210_), .Y(_abc_40319_new_n4213_));
OR2X2 OR2X2_1155 ( .A(_abc_40319_new_n4215_), .B(_abc_40319_new_n4214_), .Y(_abc_40319_new_n4216_));
OR2X2 OR2X2_1156 ( .A(_abc_40319_new_n4204_), .B(_abc_40319_new_n4218_), .Y(_abc_40319_new_n4219_));
OR2X2 OR2X2_1157 ( .A(_abc_40319_new_n4222_), .B(_abc_40319_new_n2485_), .Y(_abc_40319_new_n4223_));
OR2X2 OR2X2_1158 ( .A(_abc_40319_new_n4224_), .B(_abc_40319_new_n4225_), .Y(_abc_40319_new_n4226_));
OR2X2 OR2X2_1159 ( .A(_abc_40319_new_n4226_), .B(_abc_40319_new_n4223_), .Y(_abc_40319_new_n4227_));
OR2X2 OR2X2_116 ( .A(_abc_40319_new_n757_), .B(_abc_40319_new_n961_), .Y(_abc_40319_new_n962_));
OR2X2 OR2X2_1160 ( .A(_abc_40319_new_n4220_), .B(_abc_40319_new_n4227_), .Y(n982));
OR2X2 OR2X2_1161 ( .A(_abc_40319_new_n4230_), .B(_abc_40319_new_n4208_), .Y(_abc_40319_new_n4231_));
OR2X2 OR2X2_1162 ( .A(_abc_40319_new_n698_), .B(REG2_REG_19_), .Y(_abc_40319_new_n4234_));
OR2X2 OR2X2_1163 ( .A(_abc_40319_new_n4235_), .B(_abc_40319_new_n4233_), .Y(_abc_40319_new_n4236_));
OR2X2 OR2X2_1164 ( .A(_abc_40319_new_n4232_), .B(_abc_40319_new_n4237_), .Y(_abc_40319_new_n4238_));
OR2X2 OR2X2_1165 ( .A(_abc_40319_new_n4231_), .B(_abc_40319_new_n4236_), .Y(_abc_40319_new_n4239_));
OR2X2 OR2X2_1166 ( .A(_abc_40319_new_n698_), .B(REG1_REG_19_), .Y(_abc_40319_new_n4243_));
OR2X2 OR2X2_1167 ( .A(_abc_40319_new_n4244_), .B(_abc_40319_new_n4242_), .Y(_abc_40319_new_n4245_));
OR2X2 OR2X2_1168 ( .A(_abc_40319_new_n4247_), .B(_abc_40319_new_n4194_), .Y(_abc_40319_new_n4248_));
OR2X2 OR2X2_1169 ( .A(_abc_40319_new_n4251_), .B(_abc_40319_new_n4249_), .Y(_abc_40319_new_n4252_));
OR2X2 OR2X2_117 ( .A(_abc_40319_new_n960_), .B(_abc_40319_new_n962_), .Y(_abc_40319_new_n963_));
OR2X2 OR2X2_1170 ( .A(_abc_40319_new_n4253_), .B(_abc_40319_new_n4241_), .Y(_abc_40319_new_n4254_));
OR2X2 OR2X2_1171 ( .A(_abc_40319_new_n4254_), .B(_abc_40319_new_n4229_), .Y(_abc_40319_new_n4255_));
OR2X2 OR2X2_1172 ( .A(_abc_40319_new_n4259_), .B(_abc_40319_new_n2083_), .Y(_abc_40319_new_n4260_));
OR2X2 OR2X2_1173 ( .A(_abc_40319_new_n4260_), .B(_abc_40319_new_n4258_), .Y(_abc_40319_new_n4261_));
OR2X2 OR2X2_1174 ( .A(_abc_40319_new_n4257_), .B(_abc_40319_new_n4261_), .Y(_abc_40319_new_n4262_));
OR2X2 OR2X2_1175 ( .A(_abc_40319_new_n4256_), .B(_abc_40319_new_n4262_), .Y(n978));
OR2X2 OR2X2_1176 ( .A(_abc_40319_new_n4270_), .B(_abc_40319_new_n1169_), .Y(_abc_40319_new_n4271_));
OR2X2 OR2X2_1177 ( .A(_abc_40319_new_n4305_), .B(_abc_40319_new_n4306_), .Y(_abc_40319_new_n4307_));
OR2X2 OR2X2_1178 ( .A(_abc_40319_new_n629_), .B(_abc_40319_new_n1069_), .Y(_abc_40319_new_n4311_));
OR2X2 OR2X2_1179 ( .A(_abc_40319_new_n4309_), .B(_abc_40319_new_n4313_), .Y(_abc_40319_new_n4314_));
OR2X2 OR2X2_118 ( .A(_abc_40319_new_n964_), .B(_abc_40319_new_n936_), .Y(_abc_40319_new_n965_));
OR2X2 OR2X2_1180 ( .A(_abc_40319_new_n4271_), .B(REG2_REG_31_), .Y(_abc_40319_new_n4315_));
OR2X2 OR2X2_1181 ( .A(_abc_40319_new_n4316_), .B(_abc_40319_new_n4318_), .Y(_abc_40319_new_n4319_));
OR2X2 OR2X2_1182 ( .A(_abc_40319_new_n4319_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n4320_));
OR2X2 OR2X2_1183 ( .A(_abc_40319_new_n4308_), .B(_abc_40319_new_n4320_), .Y(n973));
OR2X2 OR2X2_1184 ( .A(_abc_40319_new_n4302_), .B(_abc_40319_new_n3169_), .Y(_abc_40319_new_n4322_));
OR2X2 OR2X2_1185 ( .A(_abc_40319_new_n4271_), .B(REG2_REG_30_), .Y(_abc_40319_new_n4325_));
OR2X2 OR2X2_1186 ( .A(_abc_40319_new_n4326_), .B(_abc_40319_new_n4327_), .Y(_abc_40319_new_n4328_));
OR2X2 OR2X2_1187 ( .A(_abc_40319_new_n4328_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n4329_));
OR2X2 OR2X2_1188 ( .A(_abc_40319_new_n4324_), .B(_abc_40319_new_n4329_), .Y(n968));
OR2X2 OR2X2_1189 ( .A(_abc_40319_new_n3109_), .B(_abc_40319_new_n4359_), .Y(_abc_40319_new_n4360_));
OR2X2 OR2X2_119 ( .A(_abc_40319_new_n966_), .B(_abc_40319_new_n917_), .Y(_abc_40319_new_n967_));
OR2X2 OR2X2_1190 ( .A(_abc_40319_new_n4361_), .B(_abc_40319_new_n4358_), .Y(_abc_40319_new_n4362_));
OR2X2 OR2X2_1191 ( .A(_abc_40319_new_n4357_), .B(_abc_40319_new_n4362_), .Y(_abc_40319_new_n4363_));
OR2X2 OR2X2_1192 ( .A(_abc_40319_new_n4370_), .B(_abc_40319_new_n2858_), .Y(_abc_40319_new_n4371_));
OR2X2 OR2X2_1193 ( .A(_abc_40319_new_n4364_), .B(_abc_40319_new_n4376_), .Y(_abc_40319_new_n4377_));
OR2X2 OR2X2_1194 ( .A(_abc_40319_new_n4392_), .B(_abc_40319_new_n4393_), .Y(_abc_40319_new_n4394_));
OR2X2 OR2X2_1195 ( .A(_abc_40319_new_n4391_), .B(_abc_40319_new_n4394_), .Y(_abc_40319_new_n4395_));
OR2X2 OR2X2_1196 ( .A(_abc_40319_new_n4406_), .B(_abc_40319_new_n4407_), .Y(_abc_40319_new_n4408_));
OR2X2 OR2X2_1197 ( .A(_abc_40319_new_n4405_), .B(_abc_40319_new_n4408_), .Y(_abc_40319_new_n4409_));
OR2X2 OR2X2_1198 ( .A(_abc_40319_new_n4422_), .B(_abc_40319_new_n4420_), .Y(_abc_40319_new_n4423_));
OR2X2 OR2X2_1199 ( .A(_abc_40319_new_n4440_), .B(_abc_40319_new_n4438_), .Y(_abc_40319_new_n4441_));
OR2X2 OR2X2_12 ( .A(_abc_40319_new_n572_), .B(_abc_40319_new_n524_), .Y(_abc_40319_new_n611_));
OR2X2 OR2X2_120 ( .A(_abc_40319_new_n870_), .B(_abc_40319_new_n768_), .Y(_abc_40319_new_n973_));
OR2X2 OR2X2_1200 ( .A(_abc_40319_new_n4445_), .B(_abc_40319_new_n4443_), .Y(_abc_40319_new_n4446_));
OR2X2 OR2X2_1201 ( .A(_abc_40319_new_n4442_), .B(_abc_40319_new_n4446_), .Y(_abc_40319_new_n4447_));
OR2X2 OR2X2_1202 ( .A(_abc_40319_new_n4447_), .B(_abc_40319_new_n4437_), .Y(_abc_40319_new_n4448_));
OR2X2 OR2X2_1203 ( .A(_abc_40319_new_n4449_), .B(_abc_40319_new_n4415_), .Y(_abc_40319_new_n4450_));
OR2X2 OR2X2_1204 ( .A(_abc_40319_new_n4450_), .B(_abc_40319_new_n4414_), .Y(_abc_40319_new_n4451_));
OR2X2 OR2X2_1205 ( .A(_abc_40319_new_n4454_), .B(_abc_40319_new_n4409_), .Y(_abc_40319_new_n4455_));
OR2X2 OR2X2_1206 ( .A(_abc_40319_new_n4458_), .B(_abc_40319_new_n4396_), .Y(_abc_40319_new_n4459_));
OR2X2 OR2X2_1207 ( .A(_abc_40319_new_n4460_), .B(_abc_40319_new_n4384_), .Y(_abc_40319_new_n4461_));
OR2X2 OR2X2_1208 ( .A(_abc_40319_new_n4462_), .B(_abc_40319_new_n4381_), .Y(_abc_40319_new_n4463_));
OR2X2 OR2X2_1209 ( .A(_abc_40319_new_n4465_), .B(_abc_40319_new_n4466_), .Y(_abc_40319_new_n4467_));
OR2X2 OR2X2_121 ( .A(_abc_40319_new_n874_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n974_));
OR2X2 OR2X2_1210 ( .A(_abc_40319_new_n4464_), .B(_abc_40319_new_n4470_), .Y(_abc_40319_new_n4471_));
OR2X2 OR2X2_1211 ( .A(_abc_40319_new_n4473_), .B(_abc_40319_new_n4346_), .Y(_abc_40319_new_n4474_));
OR2X2 OR2X2_1212 ( .A(_abc_40319_new_n4475_), .B(_abc_40319_new_n4343_), .Y(_abc_40319_new_n4476_));
OR2X2 OR2X2_1213 ( .A(_abc_40319_new_n4476_), .B(_abc_40319_new_n4342_), .Y(_abc_40319_new_n4477_));
OR2X2 OR2X2_1214 ( .A(_abc_40319_new_n4479_), .B(_abc_40319_new_n4480_), .Y(_abc_40319_new_n4481_));
OR2X2 OR2X2_1215 ( .A(_abc_40319_new_n4484_), .B(_abc_40319_new_n4482_), .Y(_abc_40319_new_n4485_));
OR2X2 OR2X2_1216 ( .A(_abc_40319_new_n4486_), .B(_abc_40319_new_n4478_), .Y(_abc_40319_new_n4487_));
OR2X2 OR2X2_1217 ( .A(_abc_40319_new_n4491_), .B(_abc_40319_new_n4492_), .Y(_abc_40319_new_n4493_));
OR2X2 OR2X2_1218 ( .A(_abc_40319_new_n672_), .B(_abc_40319_new_n646_), .Y(_abc_40319_new_n4494_));
OR2X2 OR2X2_1219 ( .A(_abc_40319_new_n1115_), .B(_abc_40319_new_n670_), .Y(_abc_40319_new_n4495_));
OR2X2 OR2X2_122 ( .A(_abc_40319_new_n971_), .B(_abc_40319_new_n976_), .Y(_abc_40319_new_n977_));
OR2X2 OR2X2_1220 ( .A(_abc_40319_new_n4501_), .B(_abc_40319_new_n3252_), .Y(_abc_40319_new_n4502_));
OR2X2 OR2X2_1221 ( .A(_abc_40319_new_n4504_), .B(_abc_40319_new_n4505_), .Y(_abc_40319_new_n4506_));
OR2X2 OR2X2_1222 ( .A(_abc_40319_new_n754_), .B(_abc_40319_new_n3452_), .Y(_abc_40319_new_n4507_));
OR2X2 OR2X2_1223 ( .A(_abc_40319_new_n4508_), .B(_abc_40319_new_n4500_), .Y(_abc_40319_new_n4509_));
OR2X2 OR2X2_1224 ( .A(_abc_40319_new_n4509_), .B(_abc_40319_new_n4498_), .Y(_abc_40319_new_n4510_));
OR2X2 OR2X2_1225 ( .A(_abc_40319_new_n4300_), .B(_abc_40319_new_n3042_), .Y(_abc_40319_new_n4515_));
OR2X2 OR2X2_1226 ( .A(_abc_40319_new_n4271_), .B(REG2_REG_28_), .Y(_abc_40319_new_n4521_));
OR2X2 OR2X2_1227 ( .A(_abc_40319_new_n4309_), .B(_abc_40319_new_n4522_), .Y(_abc_40319_new_n4523_));
OR2X2 OR2X2_1228 ( .A(_abc_40319_new_n4524_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n4525_));
OR2X2 OR2X2_1229 ( .A(_abc_40319_new_n4520_), .B(_abc_40319_new_n4525_), .Y(_abc_40319_new_n4526_));
OR2X2 OR2X2_123 ( .A(_abc_40319_new_n979_), .B(_abc_40319_new_n881_), .Y(_abc_40319_new_n980_));
OR2X2 OR2X2_1230 ( .A(_abc_40319_new_n4526_), .B(_abc_40319_new_n4519_), .Y(_abc_40319_new_n4527_));
OR2X2 OR2X2_1231 ( .A(_abc_40319_new_n4517_), .B(_abc_40319_new_n4527_), .Y(_abc_40319_new_n4528_));
OR2X2 OR2X2_1232 ( .A(_abc_40319_new_n4513_), .B(_abc_40319_new_n4528_), .Y(_abc_40319_new_n4529_));
OR2X2 OR2X2_1233 ( .A(_abc_40319_new_n4511_), .B(_abc_40319_new_n4529_), .Y(n958));
OR2X2 OR2X2_1234 ( .A(_abc_40319_new_n4532_), .B(_abc_40319_new_n4485_), .Y(_abc_40319_new_n4533_));
OR2X2 OR2X2_1235 ( .A(_abc_40319_new_n4533_), .B(_abc_40319_new_n3253_), .Y(_abc_40319_new_n4534_));
OR2X2 OR2X2_1236 ( .A(_abc_40319_new_n4535_), .B(_abc_40319_new_n3254_), .Y(_abc_40319_new_n4536_));
OR2X2 OR2X2_1237 ( .A(_abc_40319_new_n4542_), .B(_abc_40319_new_n3254_), .Y(_abc_40319_new_n4543_));
OR2X2 OR2X2_1238 ( .A(_abc_40319_new_n4541_), .B(_abc_40319_new_n3253_), .Y(_abc_40319_new_n4544_));
OR2X2 OR2X2_1239 ( .A(_abc_40319_new_n4546_), .B(_abc_40319_new_n4539_), .Y(_abc_40319_new_n4547_));
OR2X2 OR2X2_124 ( .A(_abc_40319_new_n981_), .B(_abc_40319_new_n806_), .Y(_abc_40319_new_n982_));
OR2X2 OR2X2_1240 ( .A(_abc_40319_new_n4538_), .B(_abc_40319_new_n4547_), .Y(_abc_40319_new_n4548_));
OR2X2 OR2X2_1241 ( .A(_abc_40319_new_n4299_), .B(_abc_40319_new_n3025_), .Y(_abc_40319_new_n4552_));
OR2X2 OR2X2_1242 ( .A(_abc_40319_new_n4271_), .B(REG2_REG_27_), .Y(_abc_40319_new_n4557_));
OR2X2 OR2X2_1243 ( .A(_abc_40319_new_n4309_), .B(_abc_40319_new_n4558_), .Y(_abc_40319_new_n4559_));
OR2X2 OR2X2_1244 ( .A(_abc_40319_new_n4560_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n4561_));
OR2X2 OR2X2_1245 ( .A(_abc_40319_new_n4561_), .B(_abc_40319_new_n4556_), .Y(_abc_40319_new_n4562_));
OR2X2 OR2X2_1246 ( .A(_abc_40319_new_n4555_), .B(_abc_40319_new_n4562_), .Y(_abc_40319_new_n4563_));
OR2X2 OR2X2_1247 ( .A(_abc_40319_new_n4554_), .B(_abc_40319_new_n4563_), .Y(_abc_40319_new_n4564_));
OR2X2 OR2X2_1248 ( .A(_abc_40319_new_n4550_), .B(_abc_40319_new_n4564_), .Y(_abc_40319_new_n4565_));
OR2X2 OR2X2_1249 ( .A(_abc_40319_new_n4549_), .B(_abc_40319_new_n4565_), .Y(n953));
OR2X2 OR2X2_125 ( .A(_abc_40319_new_n983_), .B(_abc_40319_new_n772_), .Y(_abc_40319_new_n984_));
OR2X2 OR2X2_1250 ( .A(_abc_40319_new_n4567_), .B(_abc_40319_new_n4483_), .Y(_abc_40319_new_n4568_));
OR2X2 OR2X2_1251 ( .A(_abc_40319_new_n4569_), .B(_abc_40319_new_n4480_), .Y(_abc_40319_new_n4570_));
OR2X2 OR2X2_1252 ( .A(_abc_40319_new_n4570_), .B(_abc_40319_new_n3106_), .Y(_abc_40319_new_n4571_));
OR2X2 OR2X2_1253 ( .A(_abc_40319_new_n4575_), .B(_abc_40319_new_n4479_), .Y(_abc_40319_new_n4576_));
OR2X2 OR2X2_1254 ( .A(_abc_40319_new_n4574_), .B(_abc_40319_new_n4576_), .Y(_abc_40319_new_n4577_));
OR2X2 OR2X2_1255 ( .A(_abc_40319_new_n4540_), .B(_abc_40319_new_n3104_), .Y(_abc_40319_new_n4581_));
OR2X2 OR2X2_1256 ( .A(_abc_40319_new_n4582_), .B(_abc_40319_new_n3107_), .Y(_abc_40319_new_n4583_));
OR2X2 OR2X2_1257 ( .A(_abc_40319_new_n4585_), .B(_abc_40319_new_n4580_), .Y(_abc_40319_new_n4586_));
OR2X2 OR2X2_1258 ( .A(_abc_40319_new_n4579_), .B(_abc_40319_new_n4586_), .Y(_abc_40319_new_n4587_));
OR2X2 OR2X2_1259 ( .A(_abc_40319_new_n4298_), .B(_abc_40319_new_n3009_), .Y(_abc_40319_new_n4591_));
OR2X2 OR2X2_126 ( .A(_abc_40319_new_n988_), .B(_abc_40319_new_n986_), .Y(_abc_40319_new_n989_));
OR2X2 OR2X2_1260 ( .A(_abc_40319_new_n4271_), .B(REG2_REG_26_), .Y(_abc_40319_new_n4596_));
OR2X2 OR2X2_1261 ( .A(_abc_40319_new_n4309_), .B(_abc_40319_new_n4597_), .Y(_abc_40319_new_n4598_));
OR2X2 OR2X2_1262 ( .A(_abc_40319_new_n4599_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n4600_));
OR2X2 OR2X2_1263 ( .A(_abc_40319_new_n4600_), .B(_abc_40319_new_n4595_), .Y(_abc_40319_new_n4601_));
OR2X2 OR2X2_1264 ( .A(_abc_40319_new_n4601_), .B(_abc_40319_new_n4594_), .Y(_abc_40319_new_n4602_));
OR2X2 OR2X2_1265 ( .A(_abc_40319_new_n4593_), .B(_abc_40319_new_n4602_), .Y(_abc_40319_new_n4603_));
OR2X2 OR2X2_1266 ( .A(_abc_40319_new_n4589_), .B(_abc_40319_new_n4603_), .Y(_abc_40319_new_n4604_));
OR2X2 OR2X2_1267 ( .A(_abc_40319_new_n4588_), .B(_abc_40319_new_n4604_), .Y(n948));
OR2X2 OR2X2_1268 ( .A(_abc_40319_new_n4607_), .B(_abc_40319_new_n4606_), .Y(_abc_40319_new_n4608_));
OR2X2 OR2X2_1269 ( .A(_abc_40319_new_n3534_), .B(_abc_40319_new_n3194_), .Y(_abc_40319_new_n4611_));
OR2X2 OR2X2_127 ( .A(_abc_40319_new_n991_), .B(_abc_40319_new_n992_), .Y(_abc_40319_new_n993_));
OR2X2 OR2X2_1270 ( .A(_abc_40319_new_n4611_), .B(_abc_40319_new_n3258_), .Y(_abc_40319_new_n4612_));
OR2X2 OR2X2_1271 ( .A(_abc_40319_new_n4613_), .B(_abc_40319_new_n3257_), .Y(_abc_40319_new_n4614_));
OR2X2 OR2X2_1272 ( .A(_abc_40319_new_n4616_), .B(_abc_40319_new_n4610_), .Y(_abc_40319_new_n4617_));
OR2X2 OR2X2_1273 ( .A(_abc_40319_new_n4609_), .B(_abc_40319_new_n4617_), .Y(_abc_40319_new_n4618_));
OR2X2 OR2X2_1274 ( .A(_abc_40319_new_n4297_), .B(_abc_40319_new_n2992_), .Y(_abc_40319_new_n4622_));
OR2X2 OR2X2_1275 ( .A(_abc_40319_new_n4271_), .B(REG2_REG_25_), .Y(_abc_40319_new_n4627_));
OR2X2 OR2X2_1276 ( .A(_abc_40319_new_n4309_), .B(_abc_40319_new_n4628_), .Y(_abc_40319_new_n4629_));
OR2X2 OR2X2_1277 ( .A(_abc_40319_new_n4630_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n4631_));
OR2X2 OR2X2_1278 ( .A(_abc_40319_new_n4631_), .B(_abc_40319_new_n4626_), .Y(_abc_40319_new_n4632_));
OR2X2 OR2X2_1279 ( .A(_abc_40319_new_n4632_), .B(_abc_40319_new_n4625_), .Y(_abc_40319_new_n4633_));
OR2X2 OR2X2_128 ( .A(_abc_40319_new_n640_), .B(DATAI_6_), .Y(_abc_40319_new_n997_));
OR2X2 OR2X2_1280 ( .A(_abc_40319_new_n4624_), .B(_abc_40319_new_n4633_), .Y(_abc_40319_new_n4634_));
OR2X2 OR2X2_1281 ( .A(_abc_40319_new_n4620_), .B(_abc_40319_new_n4634_), .Y(_abc_40319_new_n4635_));
OR2X2 OR2X2_1282 ( .A(_abc_40319_new_n4619_), .B(_abc_40319_new_n4635_), .Y(n943));
OR2X2 OR2X2_1283 ( .A(_abc_40319_new_n4637_), .B(_abc_40319_new_n4638_), .Y(_abc_40319_new_n4639_));
OR2X2 OR2X2_1284 ( .A(_abc_40319_new_n4644_), .B(_abc_40319_new_n3151_), .Y(_abc_40319_new_n4645_));
OR2X2 OR2X2_1285 ( .A(_abc_40319_new_n4649_), .B(_abc_40319_new_n3366_), .Y(_abc_40319_new_n4650_));
OR2X2 OR2X2_1286 ( .A(_abc_40319_new_n4653_), .B(_abc_40319_new_n3469_), .Y(_abc_40319_new_n4654_));
OR2X2 OR2X2_1287 ( .A(_abc_40319_new_n4652_), .B(_abc_40319_new_n4654_), .Y(_abc_40319_new_n4655_));
OR2X2 OR2X2_1288 ( .A(_abc_40319_new_n4648_), .B(_abc_40319_new_n4656_), .Y(_abc_40319_new_n4657_));
OR2X2 OR2X2_1289 ( .A(_abc_40319_new_n4658_), .B(_abc_40319_new_n3195_), .Y(_abc_40319_new_n4659_));
OR2X2 OR2X2_129 ( .A(_abc_40319_new_n740_), .B(REG3_REG_6_), .Y(_abc_40319_new_n1002_));
OR2X2 OR2X2_1290 ( .A(_abc_40319_new_n4657_), .B(_abc_40319_new_n3196_), .Y(_abc_40319_new_n4660_));
OR2X2 OR2X2_1291 ( .A(_abc_40319_new_n4662_), .B(_abc_40319_new_n4641_), .Y(_abc_40319_new_n4663_));
OR2X2 OR2X2_1292 ( .A(_abc_40319_new_n4640_), .B(_abc_40319_new_n4663_), .Y(_abc_40319_new_n4664_));
OR2X2 OR2X2_1293 ( .A(_abc_40319_new_n4296_), .B(_abc_40319_new_n2976_), .Y(_abc_40319_new_n4668_));
OR2X2 OR2X2_1294 ( .A(_abc_40319_new_n4271_), .B(REG2_REG_24_), .Y(_abc_40319_new_n4673_));
OR2X2 OR2X2_1295 ( .A(_abc_40319_new_n4309_), .B(_abc_40319_new_n4674_), .Y(_abc_40319_new_n4675_));
OR2X2 OR2X2_1296 ( .A(_abc_40319_new_n4676_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n4677_));
OR2X2 OR2X2_1297 ( .A(_abc_40319_new_n4677_), .B(_abc_40319_new_n4672_), .Y(_abc_40319_new_n4678_));
OR2X2 OR2X2_1298 ( .A(_abc_40319_new_n4678_), .B(_abc_40319_new_n4671_), .Y(_abc_40319_new_n4679_));
OR2X2 OR2X2_1299 ( .A(_abc_40319_new_n4670_), .B(_abc_40319_new_n4679_), .Y(_abc_40319_new_n4680_));
OR2X2 OR2X2_13 ( .A(_abc_40319_new_n610_), .B(_abc_40319_new_n611_), .Y(_abc_40319_new_n612_));
OR2X2 OR2X2_130 ( .A(_abc_40319_new_n1005_), .B(_abc_40319_new_n1004_), .Y(_abc_40319_new_n1006_));
OR2X2 OR2X2_1300 ( .A(_abc_40319_new_n4666_), .B(_abc_40319_new_n4680_), .Y(_abc_40319_new_n4681_));
OR2X2 OR2X2_1301 ( .A(_abc_40319_new_n4665_), .B(_abc_40319_new_n4681_), .Y(n938));
OR2X2 OR2X2_1302 ( .A(_abc_40319_new_n4683_), .B(_abc_40319_new_n4651_), .Y(_abc_40319_new_n4684_));
OR2X2 OR2X2_1303 ( .A(_abc_40319_new_n4686_), .B(_abc_40319_new_n3202_), .Y(_abc_40319_new_n4687_));
OR2X2 OR2X2_1304 ( .A(_abc_40319_new_n4653_), .B(_abc_40319_new_n3197_), .Y(_abc_40319_new_n4692_));
OR2X2 OR2X2_1305 ( .A(_abc_40319_new_n4693_), .B(_abc_40319_new_n4694_), .Y(_abc_40319_new_n4695_));
OR2X2 OR2X2_1306 ( .A(_abc_40319_new_n4691_), .B(_abc_40319_new_n4695_), .Y(_abc_40319_new_n4696_));
OR2X2 OR2X2_1307 ( .A(_abc_40319_new_n4689_), .B(_abc_40319_new_n4696_), .Y(_abc_40319_new_n4697_));
OR2X2 OR2X2_1308 ( .A(_abc_40319_new_n4701_), .B(_abc_40319_new_n4702_), .Y(_abc_40319_new_n4703_));
OR2X2 OR2X2_1309 ( .A(_abc_40319_new_n4704_), .B(_abc_40319_new_n4699_), .Y(_abc_40319_new_n4705_));
OR2X2 OR2X2_131 ( .A(_abc_40319_new_n1007_), .B(_abc_40319_new_n1008_), .Y(_abc_40319_new_n1009_));
OR2X2 OR2X2_1310 ( .A(_abc_40319_new_n4705_), .B(_abc_40319_new_n4698_), .Y(_abc_40319_new_n4706_));
OR2X2 OR2X2_1311 ( .A(_abc_40319_new_n4295_), .B(_abc_40319_new_n2959_), .Y(_abc_40319_new_n4710_));
OR2X2 OR2X2_1312 ( .A(_abc_40319_new_n4271_), .B(REG2_REG_23_), .Y(_abc_40319_new_n4715_));
OR2X2 OR2X2_1313 ( .A(_abc_40319_new_n4309_), .B(_abc_40319_new_n4716_), .Y(_abc_40319_new_n4717_));
OR2X2 OR2X2_1314 ( .A(_abc_40319_new_n4718_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n4719_));
OR2X2 OR2X2_1315 ( .A(_abc_40319_new_n4719_), .B(_abc_40319_new_n4714_), .Y(_abc_40319_new_n4720_));
OR2X2 OR2X2_1316 ( .A(_abc_40319_new_n4720_), .B(_abc_40319_new_n4713_), .Y(_abc_40319_new_n4721_));
OR2X2 OR2X2_1317 ( .A(_abc_40319_new_n4712_), .B(_abc_40319_new_n4721_), .Y(_abc_40319_new_n4722_));
OR2X2 OR2X2_1318 ( .A(_abc_40319_new_n4708_), .B(_abc_40319_new_n4722_), .Y(_abc_40319_new_n4723_));
OR2X2 OR2X2_1319 ( .A(_abc_40319_new_n4707_), .B(_abc_40319_new_n4723_), .Y(n933));
OR2X2 OR2X2_132 ( .A(_abc_40319_new_n1006_), .B(_abc_40319_new_n1009_), .Y(_abc_40319_new_n1010_));
OR2X2 OR2X2_1320 ( .A(_abc_40319_new_n4727_), .B(_abc_40319_new_n4725_), .Y(_abc_40319_new_n4728_));
OR2X2 OR2X2_1321 ( .A(_abc_40319_new_n4732_), .B(_abc_40319_new_n4733_), .Y(_abc_40319_new_n4734_));
OR2X2 OR2X2_1322 ( .A(_abc_40319_new_n4735_), .B(_abc_40319_new_n4730_), .Y(_abc_40319_new_n4736_));
OR2X2 OR2X2_1323 ( .A(_abc_40319_new_n4729_), .B(_abc_40319_new_n4736_), .Y(_abc_40319_new_n4737_));
OR2X2 OR2X2_1324 ( .A(_abc_40319_new_n4294_), .B(_abc_40319_new_n2943_), .Y(_abc_40319_new_n4741_));
OR2X2 OR2X2_1325 ( .A(_abc_40319_new_n4271_), .B(REG2_REG_22_), .Y(_abc_40319_new_n4745_));
OR2X2 OR2X2_1326 ( .A(_abc_40319_new_n4309_), .B(_abc_40319_new_n4746_), .Y(_abc_40319_new_n4747_));
OR2X2 OR2X2_1327 ( .A(_abc_40319_new_n4749_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n4750_));
OR2X2 OR2X2_1328 ( .A(_abc_40319_new_n4748_), .B(_abc_40319_new_n4750_), .Y(_abc_40319_new_n4751_));
OR2X2 OR2X2_1329 ( .A(_abc_40319_new_n4751_), .B(_abc_40319_new_n4744_), .Y(_abc_40319_new_n4752_));
OR2X2 OR2X2_133 ( .A(_abc_40319_new_n1011_), .B(_abc_40319_new_n999_), .Y(_abc_40319_new_n1012_));
OR2X2 OR2X2_1330 ( .A(_abc_40319_new_n4743_), .B(_abc_40319_new_n4752_), .Y(_abc_40319_new_n4753_));
OR2X2 OR2X2_1331 ( .A(_abc_40319_new_n4739_), .B(_abc_40319_new_n4753_), .Y(_abc_40319_new_n4754_));
OR2X2 OR2X2_1332 ( .A(_abc_40319_new_n4738_), .B(_abc_40319_new_n4754_), .Y(n928));
OR2X2 OR2X2_1333 ( .A(_abc_40319_new_n4757_), .B(_abc_40319_new_n4375_), .Y(_abc_40319_new_n4758_));
OR2X2 OR2X2_1334 ( .A(_abc_40319_new_n4759_), .B(_abc_40319_new_n4351_), .Y(_abc_40319_new_n4760_));
OR2X2 OR2X2_1335 ( .A(_abc_40319_new_n4761_), .B(_abc_40319_new_n4361_), .Y(_abc_40319_new_n4762_));
OR2X2 OR2X2_1336 ( .A(_abc_40319_new_n4762_), .B(_abc_40319_new_n3203_), .Y(_abc_40319_new_n4763_));
OR2X2 OR2X2_1337 ( .A(_abc_40319_new_n4764_), .B(_abc_40319_new_n3204_), .Y(_abc_40319_new_n4765_));
OR2X2 OR2X2_1338 ( .A(_abc_40319_new_n4685_), .B(_abc_40319_new_n3203_), .Y(_abc_40319_new_n4769_));
OR2X2 OR2X2_1339 ( .A(_abc_40319_new_n4684_), .B(_abc_40319_new_n3204_), .Y(_abc_40319_new_n4770_));
OR2X2 OR2X2_134 ( .A(_abc_40319_new_n1014_), .B(_abc_40319_new_n1015_), .Y(_abc_40319_new_n1016_));
OR2X2 OR2X2_1340 ( .A(_abc_40319_new_n4772_), .B(_abc_40319_new_n4768_), .Y(_abc_40319_new_n4773_));
OR2X2 OR2X2_1341 ( .A(_abc_40319_new_n4767_), .B(_abc_40319_new_n4773_), .Y(_abc_40319_new_n4774_));
OR2X2 OR2X2_1342 ( .A(_abc_40319_new_n4293_), .B(_abc_40319_new_n2926_), .Y(_abc_40319_new_n4778_));
OR2X2 OR2X2_1343 ( .A(_abc_40319_new_n4782_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n4783_));
OR2X2 OR2X2_1344 ( .A(_abc_40319_new_n4784_), .B(_abc_40319_new_n4786_), .Y(_abc_40319_new_n4787_));
OR2X2 OR2X2_1345 ( .A(_abc_40319_new_n4787_), .B(_abc_40319_new_n4783_), .Y(_abc_40319_new_n4788_));
OR2X2 OR2X2_1346 ( .A(_abc_40319_new_n4788_), .B(_abc_40319_new_n4781_), .Y(_abc_40319_new_n4789_));
OR2X2 OR2X2_1347 ( .A(_abc_40319_new_n4780_), .B(_abc_40319_new_n4789_), .Y(_abc_40319_new_n4790_));
OR2X2 OR2X2_1348 ( .A(_abc_40319_new_n4776_), .B(_abc_40319_new_n4790_), .Y(_abc_40319_new_n4791_));
OR2X2 OR2X2_1349 ( .A(_abc_40319_new_n4775_), .B(_abc_40319_new_n4791_), .Y(n923));
OR2X2 OR2X2_135 ( .A(_abc_40319_new_n1016_), .B(_abc_40319_new_n768_), .Y(_abc_40319_new_n1017_));
OR2X2 OR2X2_1350 ( .A(_abc_40319_new_n4793_), .B(_abc_40319_new_n4359_), .Y(_abc_40319_new_n4794_));
OR2X2 OR2X2_1351 ( .A(_abc_40319_new_n4795_), .B(_abc_40319_new_n3110_), .Y(_abc_40319_new_n4796_));
OR2X2 OR2X2_1352 ( .A(_abc_40319_new_n4794_), .B(_abc_40319_new_n4797_), .Y(_abc_40319_new_n4798_));
OR2X2 OR2X2_1353 ( .A(_abc_40319_new_n4802_), .B(_abc_40319_new_n3187_), .Y(_abc_40319_new_n4803_));
OR2X2 OR2X2_1354 ( .A(_abc_40319_new_n4803_), .B(_abc_40319_new_n3110_), .Y(_abc_40319_new_n4804_));
OR2X2 OR2X2_1355 ( .A(_abc_40319_new_n4805_), .B(_abc_40319_new_n4797_), .Y(_abc_40319_new_n4806_));
OR2X2 OR2X2_1356 ( .A(_abc_40319_new_n4808_), .B(_abc_40319_new_n4801_), .Y(_abc_40319_new_n4809_));
OR2X2 OR2X2_1357 ( .A(_abc_40319_new_n4800_), .B(_abc_40319_new_n4809_), .Y(_abc_40319_new_n4810_));
OR2X2 OR2X2_1358 ( .A(_abc_40319_new_n4292_), .B(_abc_40319_new_n2910_), .Y(_abc_40319_new_n4814_));
OR2X2 OR2X2_1359 ( .A(_abc_40319_new_n4821_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n4822_));
OR2X2 OR2X2_136 ( .A(_abc_40319_new_n1018_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1019_));
OR2X2 OR2X2_1360 ( .A(_abc_40319_new_n4820_), .B(_abc_40319_new_n4822_), .Y(_abc_40319_new_n4823_));
OR2X2 OR2X2_1361 ( .A(_abc_40319_new_n4823_), .B(_abc_40319_new_n4819_), .Y(_abc_40319_new_n4824_));
OR2X2 OR2X2_1362 ( .A(_abc_40319_new_n4824_), .B(_abc_40319_new_n4817_), .Y(_abc_40319_new_n4825_));
OR2X2 OR2X2_1363 ( .A(_abc_40319_new_n4816_), .B(_abc_40319_new_n4825_), .Y(_abc_40319_new_n4826_));
OR2X2 OR2X2_1364 ( .A(_abc_40319_new_n4812_), .B(_abc_40319_new_n4826_), .Y(_abc_40319_new_n4827_));
OR2X2 OR2X2_1365 ( .A(_abc_40319_new_n4811_), .B(_abc_40319_new_n4827_), .Y(n918));
OR2X2 OR2X2_1366 ( .A(_abc_40319_new_n4831_), .B(_abc_40319_new_n4829_), .Y(_abc_40319_new_n4832_));
OR2X2 OR2X2_1367 ( .A(_abc_40319_new_n4835_), .B(_abc_40319_new_n3189_), .Y(_abc_40319_new_n4836_));
OR2X2 OR2X2_1368 ( .A(_abc_40319_new_n4645_), .B(_abc_40319_new_n3190_), .Y(_abc_40319_new_n4837_));
OR2X2 OR2X2_1369 ( .A(_abc_40319_new_n4839_), .B(_abc_40319_new_n4834_), .Y(_abc_40319_new_n4840_));
OR2X2 OR2X2_137 ( .A(_abc_40319_new_n1020_), .B(_abc_40319_new_n1013_), .Y(_abc_40319_new_n1021_));
OR2X2 OR2X2_1370 ( .A(_abc_40319_new_n4833_), .B(_abc_40319_new_n4840_), .Y(_abc_40319_new_n4841_));
OR2X2 OR2X2_1371 ( .A(_abc_40319_new_n4291_), .B(_abc_40319_new_n2893_), .Y(_abc_40319_new_n4845_));
OR2X2 OR2X2_1372 ( .A(_abc_40319_new_n4852_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n4853_));
OR2X2 OR2X2_1373 ( .A(_abc_40319_new_n4851_), .B(_abc_40319_new_n4853_), .Y(_abc_40319_new_n4854_));
OR2X2 OR2X2_1374 ( .A(_abc_40319_new_n4854_), .B(_abc_40319_new_n4849_), .Y(_abc_40319_new_n4855_));
OR2X2 OR2X2_1375 ( .A(_abc_40319_new_n4855_), .B(_abc_40319_new_n4848_), .Y(_abc_40319_new_n4856_));
OR2X2 OR2X2_1376 ( .A(_abc_40319_new_n4847_), .B(_abc_40319_new_n4856_), .Y(_abc_40319_new_n4857_));
OR2X2 OR2X2_1377 ( .A(_abc_40319_new_n4843_), .B(_abc_40319_new_n4857_), .Y(_abc_40319_new_n4858_));
OR2X2 OR2X2_1378 ( .A(_abc_40319_new_n4842_), .B(_abc_40319_new_n4858_), .Y(n913));
OR2X2 OR2X2_1379 ( .A(_abc_40319_new_n4861_), .B(_abc_40319_new_n4862_), .Y(_abc_40319_new_n4863_));
OR2X2 OR2X2_138 ( .A(_abc_40319_new_n986_), .B(_abc_40319_new_n548_), .Y(_abc_40319_new_n1025_));
OR2X2 OR2X2_1380 ( .A(_abc_40319_new_n4867_), .B(_abc_40319_new_n3153_), .Y(_abc_40319_new_n4868_));
OR2X2 OR2X2_1381 ( .A(_abc_40319_new_n4866_), .B(_abc_40319_new_n3154_), .Y(_abc_40319_new_n4869_));
OR2X2 OR2X2_1382 ( .A(_abc_40319_new_n4871_), .B(_abc_40319_new_n4865_), .Y(_abc_40319_new_n4872_));
OR2X2 OR2X2_1383 ( .A(_abc_40319_new_n4864_), .B(_abc_40319_new_n4872_), .Y(_abc_40319_new_n4873_));
OR2X2 OR2X2_1384 ( .A(_abc_40319_new_n4290_), .B(_abc_40319_new_n2877_), .Y(_abc_40319_new_n4877_));
OR2X2 OR2X2_1385 ( .A(_abc_40319_new_n4884_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n4885_));
OR2X2 OR2X2_1386 ( .A(_abc_40319_new_n4883_), .B(_abc_40319_new_n4885_), .Y(_abc_40319_new_n4886_));
OR2X2 OR2X2_1387 ( .A(_abc_40319_new_n4886_), .B(_abc_40319_new_n4881_), .Y(_abc_40319_new_n4887_));
OR2X2 OR2X2_1388 ( .A(_abc_40319_new_n4887_), .B(_abc_40319_new_n4880_), .Y(_abc_40319_new_n4888_));
OR2X2 OR2X2_1389 ( .A(_abc_40319_new_n4879_), .B(_abc_40319_new_n4888_), .Y(_abc_40319_new_n4889_));
OR2X2 OR2X2_139 ( .A(_abc_40319_new_n1027_), .B(_abc_40319_new_n1028_), .Y(_abc_40319_new_n1029_));
OR2X2 OR2X2_1390 ( .A(_abc_40319_new_n4875_), .B(_abc_40319_new_n4889_), .Y(_abc_40319_new_n4890_));
OR2X2 OR2X2_1391 ( .A(_abc_40319_new_n4874_), .B(_abc_40319_new_n4890_), .Y(n908));
OR2X2 OR2X2_1392 ( .A(_abc_40319_new_n4893_), .B(_abc_40319_new_n4368_), .Y(_abc_40319_new_n4894_));
OR2X2 OR2X2_1393 ( .A(_abc_40319_new_n4894_), .B(_abc_40319_new_n3185_), .Y(_abc_40319_new_n4895_));
OR2X2 OR2X2_1394 ( .A(_abc_40319_new_n4896_), .B(_abc_40319_new_n3186_), .Y(_abc_40319_new_n4897_));
OR2X2 OR2X2_1395 ( .A(_abc_40319_new_n4902_), .B(_abc_40319_new_n3186_), .Y(_abc_40319_new_n4903_));
OR2X2 OR2X2_1396 ( .A(_abc_40319_new_n4901_), .B(_abc_40319_new_n3185_), .Y(_abc_40319_new_n4904_));
OR2X2 OR2X2_1397 ( .A(_abc_40319_new_n4906_), .B(_abc_40319_new_n4900_), .Y(_abc_40319_new_n4907_));
OR2X2 OR2X2_1398 ( .A(_abc_40319_new_n4899_), .B(_abc_40319_new_n4907_), .Y(_abc_40319_new_n4908_));
OR2X2 OR2X2_1399 ( .A(_abc_40319_new_n4289_), .B(_abc_40319_new_n2860_), .Y(_abc_40319_new_n4912_));
OR2X2 OR2X2_14 ( .A(_abc_40319_new_n619_), .B(_abc_40319_new_n623_), .Y(_abc_40319_new_n624_));
OR2X2 OR2X2_140 ( .A(_abc_40319_new_n640_), .B(DATAI_7_), .Y(_abc_40319_new_n1033_));
OR2X2 OR2X2_1400 ( .A(_abc_40319_new_n4920_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n4921_));
OR2X2 OR2X2_1401 ( .A(_abc_40319_new_n4919_), .B(_abc_40319_new_n4921_), .Y(_abc_40319_new_n4922_));
OR2X2 OR2X2_1402 ( .A(_abc_40319_new_n4922_), .B(_abc_40319_new_n4918_), .Y(_abc_40319_new_n4923_));
OR2X2 OR2X2_1403 ( .A(_abc_40319_new_n4923_), .B(_abc_40319_new_n4916_), .Y(_abc_40319_new_n4924_));
OR2X2 OR2X2_1404 ( .A(_abc_40319_new_n4914_), .B(_abc_40319_new_n4924_), .Y(_abc_40319_new_n4925_));
OR2X2 OR2X2_1405 ( .A(_abc_40319_new_n4910_), .B(_abc_40319_new_n4925_), .Y(_abc_40319_new_n4926_));
OR2X2 OR2X2_1406 ( .A(_abc_40319_new_n4909_), .B(_abc_40319_new_n4926_), .Y(n903));
OR2X2 OR2X2_1407 ( .A(_abc_40319_new_n4929_), .B(_abc_40319_new_n3144_), .Y(_abc_40319_new_n4930_));
OR2X2 OR2X2_1408 ( .A(_abc_40319_new_n4931_), .B(_abc_40319_new_n3111_), .Y(_abc_40319_new_n4932_));
OR2X2 OR2X2_1409 ( .A(_abc_40319_new_n4935_), .B(_abc_40319_new_n4933_), .Y(_abc_40319_new_n4936_));
OR2X2 OR2X2_141 ( .A(_abc_40319_new_n1036_), .B(_abc_40319_new_n1037_), .Y(_abc_40319_new_n1038_));
OR2X2 OR2X2_1410 ( .A(_abc_40319_new_n4939_), .B(_abc_40319_new_n4940_), .Y(_abc_40319_new_n4941_));
OR2X2 OR2X2_1411 ( .A(_abc_40319_new_n4942_), .B(_abc_40319_new_n4938_), .Y(_abc_40319_new_n4943_));
OR2X2 OR2X2_1412 ( .A(_abc_40319_new_n4943_), .B(_abc_40319_new_n4937_), .Y(_abc_40319_new_n4944_));
OR2X2 OR2X2_1413 ( .A(_abc_40319_new_n4288_), .B(_abc_40319_new_n2844_), .Y(_abc_40319_new_n4948_));
OR2X2 OR2X2_1414 ( .A(_abc_40319_new_n4953_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n4954_));
OR2X2 OR2X2_1415 ( .A(_abc_40319_new_n4952_), .B(_abc_40319_new_n4954_), .Y(_abc_40319_new_n4955_));
OR2X2 OR2X2_1416 ( .A(_abc_40319_new_n4958_), .B(_abc_40319_new_n4957_), .Y(_abc_40319_new_n4959_));
OR2X2 OR2X2_1417 ( .A(_abc_40319_new_n4959_), .B(_abc_40319_new_n4955_), .Y(_abc_40319_new_n4960_));
OR2X2 OR2X2_1418 ( .A(_abc_40319_new_n4950_), .B(_abc_40319_new_n4960_), .Y(_abc_40319_new_n4961_));
OR2X2 OR2X2_1419 ( .A(_abc_40319_new_n4946_), .B(_abc_40319_new_n4961_), .Y(_abc_40319_new_n4962_));
OR2X2 OR2X2_142 ( .A(_abc_40319_new_n1000_), .B(REG3_REG_7_), .Y(_abc_40319_new_n1041_));
OR2X2 OR2X2_1420 ( .A(_abc_40319_new_n4945_), .B(_abc_40319_new_n4962_), .Y(n898));
OR2X2 OR2X2_1421 ( .A(_abc_40319_new_n4966_), .B(_abc_40319_new_n4964_), .Y(_abc_40319_new_n4967_));
OR2X2 OR2X2_1422 ( .A(_abc_40319_new_n4971_), .B(_abc_40319_new_n4972_), .Y(_abc_40319_new_n4973_));
OR2X2 OR2X2_1423 ( .A(_abc_40319_new_n4974_), .B(_abc_40319_new_n4969_), .Y(_abc_40319_new_n4975_));
OR2X2 OR2X2_1424 ( .A(_abc_40319_new_n4975_), .B(_abc_40319_new_n4968_), .Y(_abc_40319_new_n4976_));
OR2X2 OR2X2_1425 ( .A(_abc_40319_new_n4287_), .B(_abc_40319_new_n2827_), .Y(_abc_40319_new_n4980_));
OR2X2 OR2X2_1426 ( .A(_abc_40319_new_n4271_), .B(REG2_REG_15_), .Y(_abc_40319_new_n4983_));
OR2X2 OR2X2_1427 ( .A(_abc_40319_new_n4309_), .B(_abc_40319_new_n4985_), .Y(_abc_40319_new_n4986_));
OR2X2 OR2X2_1428 ( .A(_abc_40319_new_n4986_), .B(_abc_40319_new_n4984_), .Y(_abc_40319_new_n4987_));
OR2X2 OR2X2_1429 ( .A(_abc_40319_new_n4989_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n4990_));
OR2X2 OR2X2_143 ( .A(_abc_40319_new_n1044_), .B(_abc_40319_new_n1043_), .Y(_abc_40319_new_n1045_));
OR2X2 OR2X2_1430 ( .A(_abc_40319_new_n4988_), .B(_abc_40319_new_n4990_), .Y(_abc_40319_new_n4991_));
OR2X2 OR2X2_1431 ( .A(_abc_40319_new_n4982_), .B(_abc_40319_new_n4991_), .Y(_abc_40319_new_n4992_));
OR2X2 OR2X2_1432 ( .A(_abc_40319_new_n4978_), .B(_abc_40319_new_n4992_), .Y(_abc_40319_new_n4993_));
OR2X2 OR2X2_1433 ( .A(_abc_40319_new_n4977_), .B(_abc_40319_new_n4993_), .Y(n893));
OR2X2 OR2X2_1434 ( .A(_abc_40319_new_n4928_), .B(_abc_40319_new_n3147_), .Y(_abc_40319_new_n4995_));
OR2X2 OR2X2_1435 ( .A(_abc_40319_new_n3518_), .B(_abc_40319_new_n3146_), .Y(_abc_40319_new_n4996_));
OR2X2 OR2X2_1436 ( .A(_abc_40319_new_n5001_), .B(_abc_40319_new_n5000_), .Y(_abc_40319_new_n5002_));
OR2X2 OR2X2_1437 ( .A(_abc_40319_new_n5003_), .B(_abc_40319_new_n4999_), .Y(_abc_40319_new_n5004_));
OR2X2 OR2X2_1438 ( .A(_abc_40319_new_n5004_), .B(_abc_40319_new_n4998_), .Y(_abc_40319_new_n5005_));
OR2X2 OR2X2_1439 ( .A(_abc_40319_new_n4286_), .B(_abc_40319_new_n2809_), .Y(_abc_40319_new_n5009_));
OR2X2 OR2X2_144 ( .A(_abc_40319_new_n1038_), .B(_abc_40319_new_n1045_), .Y(_abc_40319_new_n1046_));
OR2X2 OR2X2_1440 ( .A(_abc_40319_new_n5012_), .B(_abc_40319_new_n5013_), .Y(_abc_40319_new_n5014_));
OR2X2 OR2X2_1441 ( .A(_abc_40319_new_n5017_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5018_));
OR2X2 OR2X2_1442 ( .A(_abc_40319_new_n5016_), .B(_abc_40319_new_n5018_), .Y(_abc_40319_new_n5019_));
OR2X2 OR2X2_1443 ( .A(_abc_40319_new_n5019_), .B(_abc_40319_new_n5015_), .Y(_abc_40319_new_n5020_));
OR2X2 OR2X2_1444 ( .A(_abc_40319_new_n5011_), .B(_abc_40319_new_n5020_), .Y(_abc_40319_new_n5021_));
OR2X2 OR2X2_1445 ( .A(_abc_40319_new_n5007_), .B(_abc_40319_new_n5021_), .Y(_abc_40319_new_n5022_));
OR2X2 OR2X2_1446 ( .A(_abc_40319_new_n5006_), .B(_abc_40319_new_n5022_), .Y(n888));
OR2X2 OR2X2_1447 ( .A(_abc_40319_new_n5025_), .B(_abc_40319_new_n5026_), .Y(_abc_40319_new_n5027_));
OR2X2 OR2X2_1448 ( .A(_abc_40319_new_n4457_), .B(_abc_40319_new_n4387_), .Y(_abc_40319_new_n5030_));
OR2X2 OR2X2_1449 ( .A(_abc_40319_new_n5031_), .B(_abc_40319_new_n4392_), .Y(_abc_40319_new_n5032_));
OR2X2 OR2X2_145 ( .A(_abc_40319_new_n1047_), .B(_abc_40319_new_n1035_), .Y(_abc_40319_new_n1048_));
OR2X2 OR2X2_1450 ( .A(_abc_40319_new_n5032_), .B(_abc_40319_new_n3142_), .Y(_abc_40319_new_n5033_));
OR2X2 OR2X2_1451 ( .A(_abc_40319_new_n5034_), .B(_abc_40319_new_n3143_), .Y(_abc_40319_new_n5035_));
OR2X2 OR2X2_1452 ( .A(_abc_40319_new_n5037_), .B(_abc_40319_new_n5029_), .Y(_abc_40319_new_n5038_));
OR2X2 OR2X2_1453 ( .A(_abc_40319_new_n5038_), .B(_abc_40319_new_n5028_), .Y(_abc_40319_new_n5039_));
OR2X2 OR2X2_1454 ( .A(_abc_40319_new_n4285_), .B(_abc_40319_new_n2755_), .Y(_abc_40319_new_n5043_));
OR2X2 OR2X2_1455 ( .A(_abc_40319_new_n4271_), .B(REG2_REG_13_), .Y(_abc_40319_new_n5046_));
OR2X2 OR2X2_1456 ( .A(_abc_40319_new_n4309_), .B(_abc_40319_new_n5048_), .Y(_abc_40319_new_n5049_));
OR2X2 OR2X2_1457 ( .A(_abc_40319_new_n5049_), .B(_abc_40319_new_n5047_), .Y(_abc_40319_new_n5050_));
OR2X2 OR2X2_1458 ( .A(_abc_40319_new_n5052_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5053_));
OR2X2 OR2X2_1459 ( .A(_abc_40319_new_n5051_), .B(_abc_40319_new_n5053_), .Y(_abc_40319_new_n5054_));
OR2X2 OR2X2_146 ( .A(_abc_40319_new_n1050_), .B(_abc_40319_new_n1051_), .Y(_abc_40319_new_n1052_));
OR2X2 OR2X2_1460 ( .A(_abc_40319_new_n5045_), .B(_abc_40319_new_n5054_), .Y(_abc_40319_new_n5055_));
OR2X2 OR2X2_1461 ( .A(_abc_40319_new_n5041_), .B(_abc_40319_new_n5055_), .Y(_abc_40319_new_n5056_));
OR2X2 OR2X2_1462 ( .A(_abc_40319_new_n5040_), .B(_abc_40319_new_n5056_), .Y(n883));
OR2X2 OR2X2_1463 ( .A(_abc_40319_new_n5059_), .B(_abc_40319_new_n5060_), .Y(_abc_40319_new_n5061_));
OR2X2 OR2X2_1464 ( .A(_abc_40319_new_n5066_), .B(_abc_40319_new_n5064_), .Y(_abc_40319_new_n5067_));
OR2X2 OR2X2_1465 ( .A(_abc_40319_new_n5068_), .B(_abc_40319_new_n5063_), .Y(_abc_40319_new_n5069_));
OR2X2 OR2X2_1466 ( .A(_abc_40319_new_n5069_), .B(_abc_40319_new_n5062_), .Y(_abc_40319_new_n5070_));
OR2X2 OR2X2_1467 ( .A(_abc_40319_new_n4284_), .B(_abc_40319_new_n2762_), .Y(_abc_40319_new_n5074_));
OR2X2 OR2X2_1468 ( .A(_abc_40319_new_n4271_), .B(REG2_REG_12_), .Y(_abc_40319_new_n5077_));
OR2X2 OR2X2_1469 ( .A(_abc_40319_new_n4309_), .B(_abc_40319_new_n5079_), .Y(_abc_40319_new_n5080_));
OR2X2 OR2X2_147 ( .A(_abc_40319_new_n1052_), .B(_abc_40319_new_n768_), .Y(_abc_40319_new_n1053_));
OR2X2 OR2X2_1470 ( .A(_abc_40319_new_n5080_), .B(_abc_40319_new_n5078_), .Y(_abc_40319_new_n5081_));
OR2X2 OR2X2_1471 ( .A(_abc_40319_new_n5083_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5084_));
OR2X2 OR2X2_1472 ( .A(_abc_40319_new_n5082_), .B(_abc_40319_new_n5084_), .Y(_abc_40319_new_n5085_));
OR2X2 OR2X2_1473 ( .A(_abc_40319_new_n5076_), .B(_abc_40319_new_n5085_), .Y(_abc_40319_new_n5086_));
OR2X2 OR2X2_1474 ( .A(_abc_40319_new_n5072_), .B(_abc_40319_new_n5086_), .Y(_abc_40319_new_n5087_));
OR2X2 OR2X2_1475 ( .A(_abc_40319_new_n5071_), .B(_abc_40319_new_n5087_), .Y(n878));
OR2X2 OR2X2_1476 ( .A(_abc_40319_new_n5090_), .B(_abc_40319_new_n3155_), .Y(_abc_40319_new_n5091_));
OR2X2 OR2X2_1477 ( .A(_abc_40319_new_n5092_), .B(_abc_40319_new_n3205_), .Y(_abc_40319_new_n5093_));
OR2X2 OR2X2_1478 ( .A(_abc_40319_new_n5096_), .B(_abc_40319_new_n5094_), .Y(_abc_40319_new_n5097_));
OR2X2 OR2X2_1479 ( .A(_abc_40319_new_n4456_), .B(_abc_40319_new_n3226_), .Y(_abc_40319_new_n5100_));
OR2X2 OR2X2_148 ( .A(_abc_40319_new_n1054_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1055_));
OR2X2 OR2X2_1480 ( .A(_abc_40319_new_n5101_), .B(_abc_40319_new_n3227_), .Y(_abc_40319_new_n5102_));
OR2X2 OR2X2_1481 ( .A(_abc_40319_new_n5104_), .B(_abc_40319_new_n5099_), .Y(_abc_40319_new_n5105_));
OR2X2 OR2X2_1482 ( .A(_abc_40319_new_n5098_), .B(_abc_40319_new_n5105_), .Y(_abc_40319_new_n5106_));
OR2X2 OR2X2_1483 ( .A(_abc_40319_new_n4283_), .B(_abc_40319_new_n2784_), .Y(_abc_40319_new_n5110_));
OR2X2 OR2X2_1484 ( .A(_abc_40319_new_n5113_), .B(_abc_40319_new_n5114_), .Y(_abc_40319_new_n5115_));
OR2X2 OR2X2_1485 ( .A(_abc_40319_new_n5118_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5119_));
OR2X2 OR2X2_1486 ( .A(_abc_40319_new_n5117_), .B(_abc_40319_new_n5119_), .Y(_abc_40319_new_n5120_));
OR2X2 OR2X2_1487 ( .A(_abc_40319_new_n5120_), .B(_abc_40319_new_n5116_), .Y(_abc_40319_new_n5121_));
OR2X2 OR2X2_1488 ( .A(_abc_40319_new_n5112_), .B(_abc_40319_new_n5121_), .Y(_abc_40319_new_n5122_));
OR2X2 OR2X2_1489 ( .A(_abc_40319_new_n5108_), .B(_abc_40319_new_n5122_), .Y(_abc_40319_new_n5123_));
OR2X2 OR2X2_149 ( .A(_abc_40319_new_n1056_), .B(_abc_40319_new_n1049_), .Y(_abc_40319_new_n1057_));
OR2X2 OR2X2_1490 ( .A(_abc_40319_new_n5107_), .B(_abc_40319_new_n5123_), .Y(n873));
OR2X2 OR2X2_1491 ( .A(_abc_40319_new_n5127_), .B(_abc_40319_new_n5125_), .Y(_abc_40319_new_n5128_));
OR2X2 OR2X2_1492 ( .A(_abc_40319_new_n4453_), .B(_abc_40319_new_n4403_), .Y(_abc_40319_new_n5131_));
OR2X2 OR2X2_1493 ( .A(_abc_40319_new_n5131_), .B(_abc_40319_new_n4406_), .Y(_abc_40319_new_n5132_));
OR2X2 OR2X2_1494 ( .A(_abc_40319_new_n5133_), .B(_abc_40319_new_n3207_), .Y(_abc_40319_new_n5134_));
OR2X2 OR2X2_1495 ( .A(_abc_40319_new_n5135_), .B(_abc_40319_new_n3208_), .Y(_abc_40319_new_n5136_));
OR2X2 OR2X2_1496 ( .A(_abc_40319_new_n5138_), .B(_abc_40319_new_n5130_), .Y(_abc_40319_new_n5139_));
OR2X2 OR2X2_1497 ( .A(_abc_40319_new_n5139_), .B(_abc_40319_new_n5129_), .Y(_abc_40319_new_n5140_));
OR2X2 OR2X2_1498 ( .A(_abc_40319_new_n4282_), .B(_abc_40319_new_n2703_), .Y(_abc_40319_new_n5144_));
OR2X2 OR2X2_1499 ( .A(_abc_40319_new_n5148_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5149_));
OR2X2 OR2X2_15 ( .A(_abc_40319_new_n626_), .B(_abc_40319_new_n627_), .Y(_abc_40319_new_n628_));
OR2X2 OR2X2_150 ( .A(_abc_40319_new_n1059_), .B(_abc_40319_new_n1060_), .Y(_abc_40319_new_n1061_));
OR2X2 OR2X2_1500 ( .A(_abc_40319_new_n5147_), .B(_abc_40319_new_n5149_), .Y(_abc_40319_new_n5150_));
OR2X2 OR2X2_1501 ( .A(_abc_40319_new_n5152_), .B(_abc_40319_new_n5154_), .Y(_abc_40319_new_n5155_));
OR2X2 OR2X2_1502 ( .A(_abc_40319_new_n5150_), .B(_abc_40319_new_n5155_), .Y(_abc_40319_new_n5156_));
OR2X2 OR2X2_1503 ( .A(_abc_40319_new_n5146_), .B(_abc_40319_new_n5156_), .Y(_abc_40319_new_n5157_));
OR2X2 OR2X2_1504 ( .A(_abc_40319_new_n5142_), .B(_abc_40319_new_n5157_), .Y(_abc_40319_new_n5158_));
OR2X2 OR2X2_1505 ( .A(_abc_40319_new_n5141_), .B(_abc_40319_new_n5158_), .Y(n868));
OR2X2 OR2X2_1506 ( .A(_abc_40319_new_n3509_), .B(_abc_40319_new_n3157_), .Y(_abc_40319_new_n5160_));
OR2X2 OR2X2_1507 ( .A(_abc_40319_new_n5089_), .B(_abc_40319_new_n3158_), .Y(_abc_40319_new_n5161_));
OR2X2 OR2X2_1508 ( .A(_abc_40319_new_n5167_), .B(_abc_40319_new_n5165_), .Y(_abc_40319_new_n5168_));
OR2X2 OR2X2_1509 ( .A(_abc_40319_new_n5169_), .B(_abc_40319_new_n5164_), .Y(_abc_40319_new_n5170_));
OR2X2 OR2X2_151 ( .A(_abc_40319_new_n1061_), .B(_abc_40319_new_n1058_), .Y(_abc_40319_new_n1062_));
OR2X2 OR2X2_1510 ( .A(_abc_40319_new_n5170_), .B(_abc_40319_new_n5163_), .Y(_abc_40319_new_n5171_));
OR2X2 OR2X2_1511 ( .A(_abc_40319_new_n4281_), .B(_abc_40319_new_n2714_), .Y(_abc_40319_new_n5175_));
OR2X2 OR2X2_1512 ( .A(_abc_40319_new_n5178_), .B(_abc_40319_new_n5179_), .Y(_abc_40319_new_n5180_));
OR2X2 OR2X2_1513 ( .A(_abc_40319_new_n5183_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5184_));
OR2X2 OR2X2_1514 ( .A(_abc_40319_new_n5182_), .B(_abc_40319_new_n5184_), .Y(_abc_40319_new_n5185_));
OR2X2 OR2X2_1515 ( .A(_abc_40319_new_n5185_), .B(_abc_40319_new_n5181_), .Y(_abc_40319_new_n5186_));
OR2X2 OR2X2_1516 ( .A(_abc_40319_new_n5177_), .B(_abc_40319_new_n5186_), .Y(_abc_40319_new_n5187_));
OR2X2 OR2X2_1517 ( .A(_abc_40319_new_n5173_), .B(_abc_40319_new_n5187_), .Y(_abc_40319_new_n5188_));
OR2X2 OR2X2_1518 ( .A(_abc_40319_new_n5172_), .B(_abc_40319_new_n5188_), .Y(n863));
OR2X2 OR2X2_1519 ( .A(_abc_40319_new_n5192_), .B(_abc_40319_new_n5193_), .Y(_abc_40319_new_n5194_));
OR2X2 OR2X2_152 ( .A(_abc_40319_new_n1022_), .B(_abc_40319_new_n1062_), .Y(_abc_40319_new_n1063_));
OR2X2 OR2X2_1520 ( .A(_abc_40319_new_n4452_), .B(_abc_40319_new_n3176_), .Y(_abc_40319_new_n5197_));
OR2X2 OR2X2_1521 ( .A(_abc_40319_new_n5198_), .B(_abc_40319_new_n3177_), .Y(_abc_40319_new_n5199_));
OR2X2 OR2X2_1522 ( .A(_abc_40319_new_n5201_), .B(_abc_40319_new_n5196_), .Y(_abc_40319_new_n5202_));
OR2X2 OR2X2_1523 ( .A(_abc_40319_new_n5202_), .B(_abc_40319_new_n5195_), .Y(_abc_40319_new_n5203_));
OR2X2 OR2X2_1524 ( .A(_abc_40319_new_n4280_), .B(_abc_40319_new_n2730_), .Y(_abc_40319_new_n5207_));
OR2X2 OR2X2_1525 ( .A(_abc_40319_new_n5210_), .B(_abc_40319_new_n5211_), .Y(_abc_40319_new_n5212_));
OR2X2 OR2X2_1526 ( .A(_abc_40319_new_n5215_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5216_));
OR2X2 OR2X2_1527 ( .A(_abc_40319_new_n5214_), .B(_abc_40319_new_n5216_), .Y(_abc_40319_new_n5217_));
OR2X2 OR2X2_1528 ( .A(_abc_40319_new_n5217_), .B(_abc_40319_new_n5213_), .Y(_abc_40319_new_n5218_));
OR2X2 OR2X2_1529 ( .A(_abc_40319_new_n5209_), .B(_abc_40319_new_n5218_), .Y(_abc_40319_new_n5219_));
OR2X2 OR2X2_153 ( .A(_abc_40319_new_n1068_), .B(_abc_40319_new_n1070_), .Y(_abc_40319_new_n1071_));
OR2X2 OR2X2_1530 ( .A(_abc_40319_new_n5205_), .B(_abc_40319_new_n5219_), .Y(_abc_40319_new_n5220_));
OR2X2 OR2X2_1531 ( .A(_abc_40319_new_n5204_), .B(_abc_40319_new_n5220_), .Y(n858));
OR2X2 OR2X2_1532 ( .A(_abc_40319_new_n5223_), .B(_abc_40319_new_n5224_), .Y(_abc_40319_new_n5225_));
OR2X2 OR2X2_1533 ( .A(_abc_40319_new_n5230_), .B(_abc_40319_new_n5228_), .Y(_abc_40319_new_n5231_));
OR2X2 OR2X2_1534 ( .A(_abc_40319_new_n5232_), .B(_abc_40319_new_n5227_), .Y(_abc_40319_new_n5233_));
OR2X2 OR2X2_1535 ( .A(_abc_40319_new_n5233_), .B(_abc_40319_new_n5226_), .Y(_abc_40319_new_n5234_));
OR2X2 OR2X2_1536 ( .A(_abc_40319_new_n4279_), .B(_abc_40319_new_n2578_), .Y(_abc_40319_new_n5238_));
OR2X2 OR2X2_1537 ( .A(_abc_40319_new_n4271_), .B(REG2_REG_7_), .Y(_abc_40319_new_n5241_));
OR2X2 OR2X2_1538 ( .A(_abc_40319_new_n5242_), .B(_abc_40319_new_n5243_), .Y(_abc_40319_new_n5244_));
OR2X2 OR2X2_1539 ( .A(_abc_40319_new_n4309_), .B(_abc_40319_new_n5244_), .Y(_abc_40319_new_n5245_));
OR2X2 OR2X2_154 ( .A(_abc_40319_new_n1071_), .B(_abc_40319_new_n1067_), .Y(_abc_40319_new_n1072_));
OR2X2 OR2X2_1540 ( .A(_abc_40319_new_n5247_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5248_));
OR2X2 OR2X2_1541 ( .A(_abc_40319_new_n5246_), .B(_abc_40319_new_n5248_), .Y(_abc_40319_new_n5249_));
OR2X2 OR2X2_1542 ( .A(_abc_40319_new_n5240_), .B(_abc_40319_new_n5249_), .Y(_abc_40319_new_n5250_));
OR2X2 OR2X2_1543 ( .A(_abc_40319_new_n5236_), .B(_abc_40319_new_n5250_), .Y(_abc_40319_new_n5251_));
OR2X2 OR2X2_1544 ( .A(_abc_40319_new_n5235_), .B(_abc_40319_new_n5251_), .Y(n853));
OR2X2 OR2X2_1545 ( .A(_abc_40319_new_n5254_), .B(_abc_40319_new_n3219_), .Y(_abc_40319_new_n5255_));
OR2X2 OR2X2_1546 ( .A(_abc_40319_new_n5257_), .B(_abc_40319_new_n3122_), .Y(_abc_40319_new_n5258_));
OR2X2 OR2X2_1547 ( .A(_abc_40319_new_n5260_), .B(_abc_40319_new_n5261_), .Y(_abc_40319_new_n5262_));
OR2X2 OR2X2_1548 ( .A(_abc_40319_new_n5267_), .B(_abc_40319_new_n5265_), .Y(_abc_40319_new_n5268_));
OR2X2 OR2X2_1549 ( .A(_abc_40319_new_n5269_), .B(_abc_40319_new_n5264_), .Y(_abc_40319_new_n5270_));
OR2X2 OR2X2_155 ( .A(_abc_40319_new_n1072_), .B(D_REG_1_), .Y(_abc_40319_new_n1073_));
OR2X2 OR2X2_1550 ( .A(_abc_40319_new_n5263_), .B(_abc_40319_new_n5270_), .Y(_abc_40319_new_n5271_));
OR2X2 OR2X2_1551 ( .A(_abc_40319_new_n4278_), .B(_abc_40319_new_n2585_), .Y(_abc_40319_new_n5275_));
OR2X2 OR2X2_1552 ( .A(_abc_40319_new_n4271_), .B(REG2_REG_6_), .Y(_abc_40319_new_n5278_));
OR2X2 OR2X2_1553 ( .A(_abc_40319_new_n5280_), .B(_abc_40319_new_n5279_), .Y(_abc_40319_new_n5281_));
OR2X2 OR2X2_1554 ( .A(_abc_40319_new_n4309_), .B(_abc_40319_new_n5281_), .Y(_abc_40319_new_n5282_));
OR2X2 OR2X2_1555 ( .A(_abc_40319_new_n5284_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5285_));
OR2X2 OR2X2_1556 ( .A(_abc_40319_new_n5283_), .B(_abc_40319_new_n5285_), .Y(_abc_40319_new_n5286_));
OR2X2 OR2X2_1557 ( .A(_abc_40319_new_n5277_), .B(_abc_40319_new_n5286_), .Y(_abc_40319_new_n5287_));
OR2X2 OR2X2_1558 ( .A(_abc_40319_new_n5273_), .B(_abc_40319_new_n5287_), .Y(_abc_40319_new_n5288_));
OR2X2 OR2X2_1559 ( .A(_abc_40319_new_n5272_), .B(_abc_40319_new_n5288_), .Y(n848));
OR2X2 OR2X2_156 ( .A(D_REG_15_), .B(D_REG_14_), .Y(_abc_40319_new_n1078_));
OR2X2 OR2X2_1560 ( .A(_abc_40319_new_n5290_), .B(_abc_40319_new_n5291_), .Y(_abc_40319_new_n5292_));
OR2X2 OR2X2_1561 ( .A(_abc_40319_new_n5298_), .B(_abc_40319_new_n4438_), .Y(_abc_40319_new_n5299_));
OR2X2 OR2X2_1562 ( .A(_abc_40319_new_n5300_), .B(_abc_40319_new_n3223_), .Y(_abc_40319_new_n5301_));
OR2X2 OR2X2_1563 ( .A(_abc_40319_new_n5299_), .B(_abc_40319_new_n3222_), .Y(_abc_40319_new_n5302_));
OR2X2 OR2X2_1564 ( .A(_abc_40319_new_n5304_), .B(_abc_40319_new_n5294_), .Y(_abc_40319_new_n5305_));
OR2X2 OR2X2_1565 ( .A(_abc_40319_new_n5305_), .B(_abc_40319_new_n5293_), .Y(_abc_40319_new_n5306_));
OR2X2 OR2X2_1566 ( .A(_abc_40319_new_n4271_), .B(REG2_REG_4_), .Y(_abc_40319_new_n5309_));
OR2X2 OR2X2_1567 ( .A(_abc_40319_new_n5310_), .B(_abc_40319_new_n5311_), .Y(_abc_40319_new_n5312_));
OR2X2 OR2X2_1568 ( .A(_abc_40319_new_n4309_), .B(_abc_40319_new_n5312_), .Y(_abc_40319_new_n5313_));
OR2X2 OR2X2_1569 ( .A(_abc_40319_new_n4276_), .B(_abc_40319_new_n3218_), .Y(_abc_40319_new_n5316_));
OR2X2 OR2X2_157 ( .A(D_REG_12_), .B(D_REG_17_), .Y(_abc_40319_new_n1079_));
OR2X2 OR2X2_1570 ( .A(_abc_40319_new_n5319_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5320_));
OR2X2 OR2X2_1571 ( .A(_abc_40319_new_n5318_), .B(_abc_40319_new_n5320_), .Y(_abc_40319_new_n5321_));
OR2X2 OR2X2_1572 ( .A(_abc_40319_new_n5321_), .B(_abc_40319_new_n5314_), .Y(_abc_40319_new_n5322_));
OR2X2 OR2X2_1573 ( .A(_abc_40319_new_n5308_), .B(_abc_40319_new_n5322_), .Y(_abc_40319_new_n5323_));
OR2X2 OR2X2_1574 ( .A(_abc_40319_new_n5307_), .B(_abc_40319_new_n5323_), .Y(n838));
OR2X2 OR2X2_1575 ( .A(_abc_40319_new_n5256_), .B(_abc_40319_new_n3123_), .Y(_abc_40319_new_n5325_));
OR2X2 OR2X2_1576 ( .A(_abc_40319_new_n5255_), .B(_abc_40319_new_n3124_), .Y(_abc_40319_new_n5326_));
OR2X2 OR2X2_1577 ( .A(_abc_40319_new_n5330_), .B(_abc_40319_new_n4444_), .Y(_abc_40319_new_n5331_));
OR2X2 OR2X2_1578 ( .A(_abc_40319_new_n5333_), .B(_abc_40319_new_n5334_), .Y(_abc_40319_new_n5335_));
OR2X2 OR2X2_1579 ( .A(_abc_40319_new_n5336_), .B(_abc_40319_new_n5329_), .Y(_abc_40319_new_n5337_));
OR2X2 OR2X2_158 ( .A(_abc_40319_new_n1078_), .B(_abc_40319_new_n1079_), .Y(_abc_40319_new_n1080_));
OR2X2 OR2X2_1580 ( .A(_abc_40319_new_n5337_), .B(_abc_40319_new_n5328_), .Y(_abc_40319_new_n5338_));
OR2X2 OR2X2_1581 ( .A(_abc_40319_new_n5339_), .B(_abc_40319_new_n5340_), .Y(_abc_40319_new_n5341_));
OR2X2 OR2X2_1582 ( .A(_abc_40319_new_n5338_), .B(_abc_40319_new_n5341_), .Y(_abc_40319_new_n5342_));
OR2X2 OR2X2_1583 ( .A(_abc_40319_new_n4277_), .B(_abc_40319_new_n2605_), .Y(_abc_40319_new_n5346_));
OR2X2 OR2X2_1584 ( .A(_abc_40319_new_n5350_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5351_));
OR2X2 OR2X2_1585 ( .A(_abc_40319_new_n5349_), .B(_abc_40319_new_n5351_), .Y(_abc_40319_new_n5352_));
OR2X2 OR2X2_1586 ( .A(_abc_40319_new_n5348_), .B(_abc_40319_new_n5352_), .Y(_abc_40319_new_n5353_));
OR2X2 OR2X2_1587 ( .A(_abc_40319_new_n5344_), .B(_abc_40319_new_n5353_), .Y(_abc_40319_new_n5354_));
OR2X2 OR2X2_1588 ( .A(_abc_40319_new_n5343_), .B(_abc_40319_new_n5354_), .Y(n843));
OR2X2 OR2X2_1589 ( .A(_abc_40319_new_n3493_), .B(_abc_40319_new_n3133_), .Y(_abc_40319_new_n5356_));
OR2X2 OR2X2_159 ( .A(D_REG_5_), .B(D_REG_11_), .Y(_abc_40319_new_n1081_));
OR2X2 OR2X2_1590 ( .A(_abc_40319_new_n5357_), .B(_abc_40319_new_n3134_), .Y(_abc_40319_new_n5358_));
OR2X2 OR2X2_1591 ( .A(_abc_40319_new_n5363_), .B(_abc_40319_new_n3134_), .Y(_abc_40319_new_n5364_));
OR2X2 OR2X2_1592 ( .A(_abc_40319_new_n5362_), .B(_abc_40319_new_n3133_), .Y(_abc_40319_new_n5365_));
OR2X2 OR2X2_1593 ( .A(_abc_40319_new_n5367_), .B(_abc_40319_new_n5361_), .Y(_abc_40319_new_n5368_));
OR2X2 OR2X2_1594 ( .A(_abc_40319_new_n5368_), .B(_abc_40319_new_n5360_), .Y(_abc_40319_new_n5369_));
OR2X2 OR2X2_1595 ( .A(_abc_40319_new_n5370_), .B(_abc_40319_new_n5371_), .Y(_abc_40319_new_n5372_));
OR2X2 OR2X2_1596 ( .A(_abc_40319_new_n5369_), .B(_abc_40319_new_n5372_), .Y(_abc_40319_new_n5373_));
OR2X2 OR2X2_1597 ( .A(_abc_40319_new_n4275_), .B(_abc_40319_new_n819_), .Y(_abc_40319_new_n5377_));
OR2X2 OR2X2_1598 ( .A(_abc_40319_new_n5381_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5382_));
OR2X2 OR2X2_1599 ( .A(_abc_40319_new_n5380_), .B(_abc_40319_new_n5382_), .Y(_abc_40319_new_n5383_));
OR2X2 OR2X2_16 ( .A(_abc_40319_new_n623_), .B(_abc_40319_new_n630_), .Y(_abc_40319_new_n635_));
OR2X2 OR2X2_160 ( .A(D_REG_10_), .B(D_REG_13_), .Y(_abc_40319_new_n1082_));
OR2X2 OR2X2_1600 ( .A(_abc_40319_new_n5383_), .B(_abc_40319_new_n5379_), .Y(_abc_40319_new_n5384_));
OR2X2 OR2X2_1601 ( .A(_abc_40319_new_n5375_), .B(_abc_40319_new_n5384_), .Y(_abc_40319_new_n5385_));
OR2X2 OR2X2_1602 ( .A(_abc_40319_new_n5374_), .B(_abc_40319_new_n5385_), .Y(n833));
OR2X2 OR2X2_1603 ( .A(_abc_40319_new_n4271_), .B(REG2_REG_2_), .Y(_abc_40319_new_n5387_));
OR2X2 OR2X2_1604 ( .A(_abc_40319_new_n5388_), .B(_abc_40319_new_n5389_), .Y(_abc_40319_new_n5390_));
OR2X2 OR2X2_1605 ( .A(_abc_40319_new_n5392_), .B(_abc_40319_new_n3128_), .Y(_abc_40319_new_n5393_));
OR2X2 OR2X2_1606 ( .A(_abc_40319_new_n3491_), .B(_abc_40319_new_n3127_), .Y(_abc_40319_new_n5394_));
OR2X2 OR2X2_1607 ( .A(_abc_40319_new_n5398_), .B(_abc_40319_new_n5399_), .Y(_abc_40319_new_n5400_));
OR2X2 OR2X2_1608 ( .A(_abc_40319_new_n5400_), .B(_abc_40319_new_n5397_), .Y(_abc_40319_new_n5401_));
OR2X2 OR2X2_1609 ( .A(_abc_40319_new_n5396_), .B(_abc_40319_new_n5401_), .Y(_abc_40319_new_n5402_));
OR2X2 OR2X2_161 ( .A(_abc_40319_new_n1081_), .B(_abc_40319_new_n1082_), .Y(_abc_40319_new_n1083_));
OR2X2 OR2X2_1610 ( .A(_abc_40319_new_n5402_), .B(_abc_40319_new_n5391_), .Y(_abc_40319_new_n5403_));
OR2X2 OR2X2_1611 ( .A(_abc_40319_new_n4274_), .B(_abc_40319_new_n847_), .Y(_abc_40319_new_n5406_));
OR2X2 OR2X2_1612 ( .A(_abc_40319_new_n5409_), .B(_abc_40319_new_n4309_), .Y(_abc_40319_new_n5410_));
OR2X2 OR2X2_1613 ( .A(_abc_40319_new_n5403_), .B(_abc_40319_new_n5410_), .Y(_abc_40319_new_n5411_));
OR2X2 OR2X2_1614 ( .A(_abc_40319_new_n5414_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5415_));
OR2X2 OR2X2_1615 ( .A(_abc_40319_new_n5413_), .B(_abc_40319_new_n5415_), .Y(_abc_40319_new_n5416_));
OR2X2 OR2X2_1616 ( .A(_abc_40319_new_n5412_), .B(_abc_40319_new_n5416_), .Y(n828));
OR2X2 OR2X2_1617 ( .A(_abc_40319_new_n3119_), .B(_abc_40319_new_n5418_), .Y(_abc_40319_new_n5419_));
OR2X2 OR2X2_1618 ( .A(_abc_40319_new_n3490_), .B(_abc_40319_new_n3116_), .Y(_abc_40319_new_n5420_));
OR2X2 OR2X2_1619 ( .A(_abc_40319_new_n5425_), .B(_abc_40319_new_n5424_), .Y(_abc_40319_new_n5426_));
OR2X2 OR2X2_162 ( .A(_abc_40319_new_n1080_), .B(_abc_40319_new_n1083_), .Y(_abc_40319_new_n1084_));
OR2X2 OR2X2_1620 ( .A(_abc_40319_new_n5427_), .B(_abc_40319_new_n5423_), .Y(_abc_40319_new_n5428_));
OR2X2 OR2X2_1621 ( .A(_abc_40319_new_n5428_), .B(_abc_40319_new_n5422_), .Y(_abc_40319_new_n5429_));
OR2X2 OR2X2_1622 ( .A(_abc_40319_new_n4273_), .B(_abc_40319_new_n942_), .Y(_abc_40319_new_n5431_));
OR2X2 OR2X2_1623 ( .A(_abc_40319_new_n5435_), .B(_abc_40319_new_n5436_), .Y(_abc_40319_new_n5437_));
OR2X2 OR2X2_1624 ( .A(_abc_40319_new_n5434_), .B(_abc_40319_new_n5437_), .Y(_abc_40319_new_n5438_));
OR2X2 OR2X2_1625 ( .A(_abc_40319_new_n5429_), .B(_abc_40319_new_n5438_), .Y(_abc_40319_new_n5439_));
OR2X2 OR2X2_1626 ( .A(_abc_40319_new_n5443_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5444_));
OR2X2 OR2X2_1627 ( .A(_abc_40319_new_n5442_), .B(_abc_40319_new_n5444_), .Y(_abc_40319_new_n5445_));
OR2X2 OR2X2_1628 ( .A(_abc_40319_new_n5441_), .B(_abc_40319_new_n5445_), .Y(_abc_40319_new_n5446_));
OR2X2 OR2X2_1629 ( .A(_abc_40319_new_n5440_), .B(_abc_40319_new_n5446_), .Y(n823));
OR2X2 OR2X2_163 ( .A(D_REG_19_), .B(D_REG_18_), .Y(_abc_40319_new_n1085_));
OR2X2 OR2X2_1630 ( .A(_abc_40319_new_n4497_), .B(_abc_40319_new_n4507_), .Y(_abc_40319_new_n5448_));
OR2X2 OR2X2_1631 ( .A(_abc_40319_new_n5449_), .B(_abc_40319_new_n5450_), .Y(_abc_40319_new_n5451_));
OR2X2 OR2X2_1632 ( .A(_abc_40319_new_n4264_), .B(_abc_40319_new_n1152_), .Y(_abc_40319_new_n5452_));
OR2X2 OR2X2_1633 ( .A(_abc_40319_new_n4309_), .B(_abc_40319_new_n5453_), .Y(_abc_40319_new_n5454_));
OR2X2 OR2X2_1634 ( .A(_abc_40319_new_n5454_), .B(_abc_40319_new_n5451_), .Y(_abc_40319_new_n5455_));
OR2X2 OR2X2_1635 ( .A(_abc_40319_new_n4271_), .B(REG2_REG_0_), .Y(_abc_40319_new_n5456_));
OR2X2 OR2X2_1636 ( .A(_abc_40319_new_n5459_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5460_));
OR2X2 OR2X2_1637 ( .A(_abc_40319_new_n5458_), .B(_abc_40319_new_n5460_), .Y(_abc_40319_new_n5461_));
OR2X2 OR2X2_1638 ( .A(_abc_40319_new_n5457_), .B(_abc_40319_new_n5461_), .Y(n818));
OR2X2 OR2X2_1639 ( .A(_abc_40319_new_n5465_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5466_));
OR2X2 OR2X2_164 ( .A(D_REG_21_), .B(D_REG_20_), .Y(_abc_40319_new_n1086_));
OR2X2 OR2X2_1640 ( .A(_abc_40319_new_n5464_), .B(_abc_40319_new_n5466_), .Y(n333));
OR2X2 OR2X2_1641 ( .A(_abc_40319_new_n5504_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5505_));
OR2X2 OR2X2_1642 ( .A(_abc_40319_new_n5505_), .B(_abc_40319_new_n5503_), .Y(_abc_40319_new_n5506_));
OR2X2 OR2X2_1643 ( .A(_abc_40319_new_n5501_), .B(_abc_40319_new_n5506_), .Y(n328));
OR2X2 OR2X2_1644 ( .A(_abc_40319_new_n5510_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5511_));
OR2X2 OR2X2_1645 ( .A(_abc_40319_new_n5511_), .B(_abc_40319_new_n5509_), .Y(_abc_40319_new_n5512_));
OR2X2 OR2X2_1646 ( .A(_abc_40319_new_n5508_), .B(_abc_40319_new_n5512_), .Y(n323));
OR2X2 OR2X2_1647 ( .A(_abc_40319_new_n5516_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5517_));
OR2X2 OR2X2_1648 ( .A(_abc_40319_new_n5517_), .B(_abc_40319_new_n5515_), .Y(_abc_40319_new_n5518_));
OR2X2 OR2X2_1649 ( .A(_abc_40319_new_n5514_), .B(_abc_40319_new_n5518_), .Y(n318));
OR2X2 OR2X2_165 ( .A(_abc_40319_new_n1085_), .B(_abc_40319_new_n1086_), .Y(_abc_40319_new_n1087_));
OR2X2 OR2X2_1650 ( .A(_abc_40319_new_n5522_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5523_));
OR2X2 OR2X2_1651 ( .A(_abc_40319_new_n5523_), .B(_abc_40319_new_n5521_), .Y(_abc_40319_new_n5524_));
OR2X2 OR2X2_1652 ( .A(_abc_40319_new_n5520_), .B(_abc_40319_new_n5524_), .Y(n313));
OR2X2 OR2X2_1653 ( .A(_abc_40319_new_n5528_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5529_));
OR2X2 OR2X2_1654 ( .A(_abc_40319_new_n5529_), .B(_abc_40319_new_n5527_), .Y(_abc_40319_new_n5530_));
OR2X2 OR2X2_1655 ( .A(_abc_40319_new_n5526_), .B(_abc_40319_new_n5530_), .Y(n308));
OR2X2 OR2X2_1656 ( .A(_abc_40319_new_n5534_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5535_));
OR2X2 OR2X2_1657 ( .A(_abc_40319_new_n5535_), .B(_abc_40319_new_n5533_), .Y(_abc_40319_new_n5536_));
OR2X2 OR2X2_1658 ( .A(_abc_40319_new_n5532_), .B(_abc_40319_new_n5536_), .Y(n303));
OR2X2 OR2X2_1659 ( .A(_abc_40319_new_n5540_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5541_));
OR2X2 OR2X2_166 ( .A(D_REG_16_), .B(D_REG_24_), .Y(_abc_40319_new_n1088_));
OR2X2 OR2X2_1660 ( .A(_abc_40319_new_n5541_), .B(_abc_40319_new_n5539_), .Y(_abc_40319_new_n5542_));
OR2X2 OR2X2_1661 ( .A(_abc_40319_new_n5538_), .B(_abc_40319_new_n5542_), .Y(n298));
OR2X2 OR2X2_1662 ( .A(_abc_40319_new_n5544_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5545_));
OR2X2 OR2X2_1663 ( .A(_abc_40319_new_n2550_), .B(_abc_40319_new_n5545_), .Y(n293));
OR2X2 OR2X2_1664 ( .A(_abc_40319_new_n5550_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5551_));
OR2X2 OR2X2_1665 ( .A(_abc_40319_new_n5551_), .B(_abc_40319_new_n5549_), .Y(_abc_40319_new_n5552_));
OR2X2 OR2X2_1666 ( .A(_abc_40319_new_n5548_), .B(_abc_40319_new_n5552_), .Y(n288));
OR2X2 OR2X2_1667 ( .A(_abc_40319_new_n5556_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5557_));
OR2X2 OR2X2_1668 ( .A(_abc_40319_new_n5557_), .B(_abc_40319_new_n5555_), .Y(_abc_40319_new_n5558_));
OR2X2 OR2X2_1669 ( .A(_abc_40319_new_n5554_), .B(_abc_40319_new_n5558_), .Y(n283));
OR2X2 OR2X2_167 ( .A(D_REG_23_), .B(D_REG_22_), .Y(_abc_40319_new_n1089_));
OR2X2 OR2X2_1670 ( .A(_abc_40319_new_n5562_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5563_));
OR2X2 OR2X2_1671 ( .A(_abc_40319_new_n5563_), .B(_abc_40319_new_n5561_), .Y(_abc_40319_new_n5564_));
OR2X2 OR2X2_1672 ( .A(_abc_40319_new_n5560_), .B(_abc_40319_new_n5564_), .Y(n278));
OR2X2 OR2X2_1673 ( .A(_abc_40319_new_n5568_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5569_));
OR2X2 OR2X2_1674 ( .A(_abc_40319_new_n5569_), .B(_abc_40319_new_n5567_), .Y(_abc_40319_new_n5570_));
OR2X2 OR2X2_1675 ( .A(_abc_40319_new_n5566_), .B(_abc_40319_new_n5570_), .Y(n273));
OR2X2 OR2X2_1676 ( .A(_abc_40319_new_n5574_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5575_));
OR2X2 OR2X2_1677 ( .A(_abc_40319_new_n5575_), .B(_abc_40319_new_n5573_), .Y(_abc_40319_new_n5576_));
OR2X2 OR2X2_1678 ( .A(_abc_40319_new_n5572_), .B(_abc_40319_new_n5576_), .Y(n268));
OR2X2 OR2X2_1679 ( .A(_abc_40319_new_n5580_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5581_));
OR2X2 OR2X2_168 ( .A(_abc_40319_new_n1088_), .B(_abc_40319_new_n1089_), .Y(_abc_40319_new_n1090_));
OR2X2 OR2X2_1680 ( .A(_abc_40319_new_n5581_), .B(_abc_40319_new_n5579_), .Y(_abc_40319_new_n5582_));
OR2X2 OR2X2_1681 ( .A(_abc_40319_new_n5578_), .B(_abc_40319_new_n5582_), .Y(n263));
OR2X2 OR2X2_1682 ( .A(_abc_40319_new_n5587_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5588_));
OR2X2 OR2X2_1683 ( .A(_abc_40319_new_n5588_), .B(_abc_40319_new_n5586_), .Y(_abc_40319_new_n5589_));
OR2X2 OR2X2_1684 ( .A(_abc_40319_new_n5585_), .B(_abc_40319_new_n5589_), .Y(n258));
OR2X2 OR2X2_1685 ( .A(_abc_40319_new_n5593_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5594_));
OR2X2 OR2X2_1686 ( .A(_abc_40319_new_n5594_), .B(_abc_40319_new_n5592_), .Y(_abc_40319_new_n5595_));
OR2X2 OR2X2_1687 ( .A(_abc_40319_new_n5591_), .B(_abc_40319_new_n5595_), .Y(n253));
OR2X2 OR2X2_1688 ( .A(_abc_40319_new_n5599_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5600_));
OR2X2 OR2X2_1689 ( .A(_abc_40319_new_n5600_), .B(_abc_40319_new_n5598_), .Y(_abc_40319_new_n5601_));
OR2X2 OR2X2_169 ( .A(_abc_40319_new_n1087_), .B(_abc_40319_new_n1090_), .Y(_abc_40319_new_n1091_));
OR2X2 OR2X2_1690 ( .A(_abc_40319_new_n5597_), .B(_abc_40319_new_n5601_), .Y(n248));
OR2X2 OR2X2_1691 ( .A(_abc_40319_new_n5606_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5607_));
OR2X2 OR2X2_1692 ( .A(_abc_40319_new_n5607_), .B(_abc_40319_new_n5605_), .Y(_abc_40319_new_n5608_));
OR2X2 OR2X2_1693 ( .A(_abc_40319_new_n5604_), .B(_abc_40319_new_n5608_), .Y(n243));
OR2X2 OR2X2_1694 ( .A(_abc_40319_new_n5613_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5614_));
OR2X2 OR2X2_1695 ( .A(_abc_40319_new_n5614_), .B(_abc_40319_new_n5612_), .Y(_abc_40319_new_n5615_));
OR2X2 OR2X2_1696 ( .A(_abc_40319_new_n5611_), .B(_abc_40319_new_n5615_), .Y(n238));
OR2X2 OR2X2_1697 ( .A(_abc_40319_new_n5620_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5621_));
OR2X2 OR2X2_1698 ( .A(_abc_40319_new_n5621_), .B(_abc_40319_new_n5619_), .Y(_abc_40319_new_n5622_));
OR2X2 OR2X2_1699 ( .A(_abc_40319_new_n5618_), .B(_abc_40319_new_n5622_), .Y(n233));
OR2X2 OR2X2_17 ( .A(_abc_40319_new_n636_), .B(_abc_40319_new_n524_), .Y(_abc_40319_new_n637_));
OR2X2 OR2X2_170 ( .A(_abc_40319_new_n1084_), .B(_abc_40319_new_n1091_), .Y(_abc_40319_new_n1092_));
OR2X2 OR2X2_1700 ( .A(_abc_40319_new_n5627_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5628_));
OR2X2 OR2X2_1701 ( .A(_abc_40319_new_n5628_), .B(_abc_40319_new_n5626_), .Y(_abc_40319_new_n5629_));
OR2X2 OR2X2_1702 ( .A(_abc_40319_new_n5625_), .B(_abc_40319_new_n5629_), .Y(n228));
OR2X2 OR2X2_1703 ( .A(_abc_40319_new_n5633_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5634_));
OR2X2 OR2X2_1704 ( .A(_abc_40319_new_n5634_), .B(_abc_40319_new_n5632_), .Y(_abc_40319_new_n5635_));
OR2X2 OR2X2_1705 ( .A(_abc_40319_new_n5631_), .B(_abc_40319_new_n5635_), .Y(n223));
OR2X2 OR2X2_1706 ( .A(_abc_40319_new_n5639_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5640_));
OR2X2 OR2X2_1707 ( .A(_abc_40319_new_n5640_), .B(_abc_40319_new_n5638_), .Y(_abc_40319_new_n5641_));
OR2X2 OR2X2_1708 ( .A(_abc_40319_new_n5637_), .B(_abc_40319_new_n5641_), .Y(n218));
OR2X2 OR2X2_1709 ( .A(_abc_40319_new_n5645_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5646_));
OR2X2 OR2X2_171 ( .A(D_REG_26_), .B(D_REG_25_), .Y(_abc_40319_new_n1093_));
OR2X2 OR2X2_1710 ( .A(_abc_40319_new_n5646_), .B(_abc_40319_new_n5644_), .Y(_abc_40319_new_n5647_));
OR2X2 OR2X2_1711 ( .A(_abc_40319_new_n5643_), .B(_abc_40319_new_n5647_), .Y(n213));
OR2X2 OR2X2_1712 ( .A(_abc_40319_new_n5651_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5652_));
OR2X2 OR2X2_1713 ( .A(_abc_40319_new_n5652_), .B(_abc_40319_new_n5650_), .Y(_abc_40319_new_n5653_));
OR2X2 OR2X2_1714 ( .A(_abc_40319_new_n5649_), .B(_abc_40319_new_n5653_), .Y(n208));
OR2X2 OR2X2_1715 ( .A(_abc_40319_new_n5657_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5658_));
OR2X2 OR2X2_1716 ( .A(_abc_40319_new_n5658_), .B(_abc_40319_new_n5656_), .Y(_abc_40319_new_n5659_));
OR2X2 OR2X2_1717 ( .A(_abc_40319_new_n5655_), .B(_abc_40319_new_n5659_), .Y(n203));
OR2X2 OR2X2_1718 ( .A(_abc_40319_new_n5663_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5664_));
OR2X2 OR2X2_1719 ( .A(_abc_40319_new_n5664_), .B(_abc_40319_new_n5662_), .Y(_abc_40319_new_n5665_));
OR2X2 OR2X2_172 ( .A(D_REG_2_), .B(D_REG_29_), .Y(_abc_40319_new_n1094_));
OR2X2 OR2X2_1720 ( .A(_abc_40319_new_n5661_), .B(_abc_40319_new_n5665_), .Y(n198));
OR2X2 OR2X2_1721 ( .A(_abc_40319_new_n5669_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5670_));
OR2X2 OR2X2_1722 ( .A(_abc_40319_new_n5670_), .B(_abc_40319_new_n5668_), .Y(_abc_40319_new_n5671_));
OR2X2 OR2X2_1723 ( .A(_abc_40319_new_n5667_), .B(_abc_40319_new_n5671_), .Y(n193));
OR2X2 OR2X2_1724 ( .A(_abc_40319_new_n530_), .B(_abc_40319_new_n528_), .Y(_abc_40319_new_n5673_));
OR2X2 OR2X2_1725 ( .A(_abc_40319_new_n5677_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5678_));
OR2X2 OR2X2_1726 ( .A(_abc_40319_new_n5678_), .B(_abc_40319_new_n5676_), .Y(_abc_40319_new_n5679_));
OR2X2 OR2X2_1727 ( .A(_abc_40319_new_n5675_), .B(_abc_40319_new_n5679_), .Y(n188));
OR2X2 OR2X2_1728 ( .A(_abc_40319_new_n5682_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5683_));
OR2X2 OR2X2_1729 ( .A(_abc_40319_new_n5681_), .B(_abc_40319_new_n5683_), .Y(n183));
OR2X2 OR2X2_173 ( .A(D_REG_28_), .B(D_REG_27_), .Y(_abc_40319_new_n1095_));
OR2X2 OR2X2_1730 ( .A(_abc_40319_new_n5686_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5687_));
OR2X2 OR2X2_1731 ( .A(_abc_40319_new_n5685_), .B(_abc_40319_new_n5687_), .Y(n178));
OR2X2 OR2X2_1732 ( .A(_abc_40319_new_n3539_), .B(_abc_40319_new_n3103_), .Y(_abc_40319_new_n5690_));
OR2X2 OR2X2_1733 ( .A(_abc_40319_new_n5692_), .B(_abc_40319_new_n5691_), .Y(_abc_40319_new_n5693_));
OR2X2 OR2X2_1734 ( .A(_abc_40319_new_n5699_), .B(_abc_40319_new_n5696_), .Y(_abc_40319_new_n5700_));
OR2X2 OR2X2_1735 ( .A(_abc_40319_new_n5700_), .B(_abc_40319_new_n3103_), .Y(_abc_40319_new_n5701_));
OR2X2 OR2X2_1736 ( .A(_abc_40319_new_n5702_), .B(_abc_40319_new_n5691_), .Y(_abc_40319_new_n5703_));
OR2X2 OR2X2_1737 ( .A(_abc_40319_new_n3453_), .B(_abc_40319_new_n754_), .Y(_abc_40319_new_n5706_));
OR2X2 OR2X2_1738 ( .A(_abc_40319_new_n5709_), .B(_abc_40319_new_n5708_), .Y(_abc_40319_new_n5710_));
OR2X2 OR2X2_1739 ( .A(_abc_40319_new_n5707_), .B(_abc_40319_new_n5710_), .Y(_abc_40319_new_n5711_));
OR2X2 OR2X2_174 ( .A(_abc_40319_new_n1094_), .B(_abc_40319_new_n1095_), .Y(_abc_40319_new_n1096_));
OR2X2 OR2X2_1740 ( .A(_abc_40319_new_n5705_), .B(_abc_40319_new_n5711_), .Y(_abc_40319_new_n5712_));
OR2X2 OR2X2_1741 ( .A(_abc_40319_new_n5712_), .B(_abc_40319_new_n5695_), .Y(_abc_40319_new_n5713_));
OR2X2 OR2X2_1742 ( .A(_abc_40319_new_n4301_), .B(_abc_40319_new_n3059_), .Y(_abc_40319_new_n5717_));
OR2X2 OR2X2_1743 ( .A(_abc_40319_new_n5723_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5724_));
OR2X2 OR2X2_1744 ( .A(_abc_40319_new_n5724_), .B(_abc_40319_new_n5722_), .Y(_abc_40319_new_n5725_));
OR2X2 OR2X2_1745 ( .A(_abc_40319_new_n5720_), .B(_abc_40319_new_n5725_), .Y(_abc_40319_new_n5726_));
OR2X2 OR2X2_1746 ( .A(_abc_40319_new_n5719_), .B(_abc_40319_new_n5726_), .Y(_abc_40319_new_n5727_));
OR2X2 OR2X2_1747 ( .A(_abc_40319_new_n5715_), .B(_abc_40319_new_n5727_), .Y(_abc_40319_new_n5728_));
OR2X2 OR2X2_1748 ( .A(_abc_40319_new_n5714_), .B(_abc_40319_new_n5728_), .Y(n963));
OR2X2 OR2X2_1749 ( .A(_abc_40319_new_n5730_), .B(_abc_40319_new_n596_), .Y(_abc_40319_new_n5731_));
OR2X2 OR2X2_175 ( .A(_abc_40319_new_n1096_), .B(_abc_40319_new_n1093_), .Y(_abc_40319_new_n1097_));
OR2X2 OR2X2_1750 ( .A(_abc_40319_new_n5733_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5734_));
OR2X2 OR2X2_1751 ( .A(_abc_40319_new_n5734_), .B(_abc_40319_new_n5732_), .Y(n338));
OR2X2 OR2X2_1752 ( .A(_abc_40319_new_n5737_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5738_));
OR2X2 OR2X2_1753 ( .A(_abc_40319_new_n5738_), .B(_abc_40319_new_n5736_), .Y(n343));
OR2X2 OR2X2_1754 ( .A(_abc_40319_new_n5747_), .B(_abc_40319_new_n4818_), .Y(_abc_40319_new_n5748_));
OR2X2 OR2X2_1755 ( .A(_abc_40319_new_n5746_), .B(_abc_40319_new_n5748_), .Y(_abc_40319_new_n5749_));
OR2X2 OR2X2_1756 ( .A(_abc_40319_new_n5745_), .B(_abc_40319_new_n5749_), .Y(_abc_40319_new_n5750_));
OR2X2 OR2X2_1757 ( .A(_abc_40319_new_n4810_), .B(_abc_40319_new_n5750_), .Y(_abc_40319_new_n5751_));
OR2X2 OR2X2_1758 ( .A(_abc_40319_new_n5754_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5755_));
OR2X2 OR2X2_1759 ( .A(_abc_40319_new_n5752_), .B(_abc_40319_new_n5755_), .Y(n598));
OR2X2 OR2X2_176 ( .A(D_REG_4_), .B(D_REG_3_), .Y(_abc_40319_new_n1098_));
OR2X2 OR2X2_1760 ( .A(_abc_40319_new_n5757_), .B(_abc_40319_new_n5758_), .Y(_abc_40319_new_n5759_));
OR2X2 OR2X2_1761 ( .A(_abc_40319_new_n5451_), .B(_abc_40319_new_n5759_), .Y(_abc_40319_new_n5760_));
OR2X2 OR2X2_1762 ( .A(_abc_40319_new_n5762_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5763_));
OR2X2 OR2X2_1763 ( .A(_abc_40319_new_n5761_), .B(_abc_40319_new_n5763_), .Y(n498));
OR2X2 OR2X2_1764 ( .A(_abc_40319_new_n5433_), .B(_abc_40319_new_n5437_), .Y(_abc_40319_new_n5766_));
OR2X2 OR2X2_1765 ( .A(_abc_40319_new_n5765_), .B(_abc_40319_new_n5766_), .Y(_abc_40319_new_n5767_));
OR2X2 OR2X2_1766 ( .A(_abc_40319_new_n5429_), .B(_abc_40319_new_n5767_), .Y(_abc_40319_new_n5768_));
OR2X2 OR2X2_1767 ( .A(_abc_40319_new_n5770_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5771_));
OR2X2 OR2X2_1768 ( .A(_abc_40319_new_n5769_), .B(_abc_40319_new_n5771_), .Y(n503));
OR2X2 OR2X2_1769 ( .A(_abc_40319_new_n5773_), .B(_abc_40319_new_n5408_), .Y(_abc_40319_new_n5774_));
OR2X2 OR2X2_177 ( .A(D_REG_7_), .B(D_REG_6_), .Y(_abc_40319_new_n1099_));
OR2X2 OR2X2_1770 ( .A(_abc_40319_new_n5403_), .B(_abc_40319_new_n5774_), .Y(_abc_40319_new_n5775_));
OR2X2 OR2X2_1771 ( .A(_abc_40319_new_n5777_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5778_));
OR2X2 OR2X2_1772 ( .A(_abc_40319_new_n5776_), .B(_abc_40319_new_n5778_), .Y(n508));
OR2X2 OR2X2_1773 ( .A(_abc_40319_new_n5781_), .B(_abc_40319_new_n5372_), .Y(_abc_40319_new_n5782_));
OR2X2 OR2X2_1774 ( .A(_abc_40319_new_n5780_), .B(_abc_40319_new_n5782_), .Y(_abc_40319_new_n5783_));
OR2X2 OR2X2_1775 ( .A(_abc_40319_new_n5369_), .B(_abc_40319_new_n5783_), .Y(_abc_40319_new_n5784_));
OR2X2 OR2X2_1776 ( .A(_abc_40319_new_n5786_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5787_));
OR2X2 OR2X2_1777 ( .A(_abc_40319_new_n5785_), .B(_abc_40319_new_n5787_), .Y(n513));
OR2X2 OR2X2_1778 ( .A(_abc_40319_new_n5790_), .B(_abc_40319_new_n5312_), .Y(_abc_40319_new_n5791_));
OR2X2 OR2X2_1779 ( .A(_abc_40319_new_n5789_), .B(_abc_40319_new_n5791_), .Y(_abc_40319_new_n5792_));
OR2X2 OR2X2_178 ( .A(_abc_40319_new_n1098_), .B(_abc_40319_new_n1099_), .Y(_abc_40319_new_n1100_));
OR2X2 OR2X2_1780 ( .A(_abc_40319_new_n5306_), .B(_abc_40319_new_n5792_), .Y(_abc_40319_new_n5793_));
OR2X2 OR2X2_1781 ( .A(_abc_40319_new_n5795_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5796_));
OR2X2 OR2X2_1782 ( .A(_abc_40319_new_n5794_), .B(_abc_40319_new_n5796_), .Y(n518));
OR2X2 OR2X2_1783 ( .A(_abc_40319_new_n5799_), .B(_abc_40319_new_n5341_), .Y(_abc_40319_new_n5800_));
OR2X2 OR2X2_1784 ( .A(_abc_40319_new_n5798_), .B(_abc_40319_new_n5800_), .Y(_abc_40319_new_n5801_));
OR2X2 OR2X2_1785 ( .A(_abc_40319_new_n5338_), .B(_abc_40319_new_n5801_), .Y(_abc_40319_new_n5802_));
OR2X2 OR2X2_1786 ( .A(_abc_40319_new_n5804_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5805_));
OR2X2 OR2X2_1787 ( .A(_abc_40319_new_n5803_), .B(_abc_40319_new_n5805_), .Y(n523));
OR2X2 OR2X2_1788 ( .A(_abc_40319_new_n5807_), .B(_abc_40319_new_n5281_), .Y(_abc_40319_new_n5808_));
OR2X2 OR2X2_1789 ( .A(_abc_40319_new_n5809_), .B(_abc_40319_new_n5808_), .Y(_abc_40319_new_n5810_));
OR2X2 OR2X2_179 ( .A(D_REG_9_), .B(D_REG_8_), .Y(_abc_40319_new_n1101_));
OR2X2 OR2X2_1790 ( .A(_abc_40319_new_n5271_), .B(_abc_40319_new_n5810_), .Y(_abc_40319_new_n5811_));
OR2X2 OR2X2_1791 ( .A(_abc_40319_new_n5813_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5814_));
OR2X2 OR2X2_1792 ( .A(_abc_40319_new_n5812_), .B(_abc_40319_new_n5814_), .Y(n528));
OR2X2 OR2X2_1793 ( .A(_abc_40319_new_n5817_), .B(_abc_40319_new_n5244_), .Y(_abc_40319_new_n5818_));
OR2X2 OR2X2_1794 ( .A(_abc_40319_new_n5816_), .B(_abc_40319_new_n5818_), .Y(_abc_40319_new_n5819_));
OR2X2 OR2X2_1795 ( .A(_abc_40319_new_n5234_), .B(_abc_40319_new_n5819_), .Y(_abc_40319_new_n5820_));
OR2X2 OR2X2_1796 ( .A(_abc_40319_new_n5822_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5823_));
OR2X2 OR2X2_1797 ( .A(_abc_40319_new_n5821_), .B(_abc_40319_new_n5823_), .Y(n533));
OR2X2 OR2X2_1798 ( .A(_abc_40319_new_n5826_), .B(_abc_40319_new_n5212_), .Y(_abc_40319_new_n5827_));
OR2X2 OR2X2_1799 ( .A(_abc_40319_new_n5825_), .B(_abc_40319_new_n5827_), .Y(_abc_40319_new_n5828_));
OR2X2 OR2X2_18 ( .A(_abc_40319_new_n608_), .B(_abc_40319_new_n642_), .Y(_abc_40319_new_n643_));
OR2X2 OR2X2_180 ( .A(D_REG_31_), .B(D_REG_30_), .Y(_abc_40319_new_n1102_));
OR2X2 OR2X2_1800 ( .A(_abc_40319_new_n5203_), .B(_abc_40319_new_n5828_), .Y(_abc_40319_new_n5829_));
OR2X2 OR2X2_1801 ( .A(_abc_40319_new_n5831_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5832_));
OR2X2 OR2X2_1802 ( .A(_abc_40319_new_n5830_), .B(_abc_40319_new_n5832_), .Y(n538));
OR2X2 OR2X2_1803 ( .A(_abc_40319_new_n5835_), .B(_abc_40319_new_n5180_), .Y(_abc_40319_new_n5836_));
OR2X2 OR2X2_1804 ( .A(_abc_40319_new_n5834_), .B(_abc_40319_new_n5836_), .Y(_abc_40319_new_n5837_));
OR2X2 OR2X2_1805 ( .A(_abc_40319_new_n5171_), .B(_abc_40319_new_n5837_), .Y(_abc_40319_new_n5838_));
OR2X2 OR2X2_1806 ( .A(_abc_40319_new_n5840_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5841_));
OR2X2 OR2X2_1807 ( .A(_abc_40319_new_n5839_), .B(_abc_40319_new_n5841_), .Y(n543));
OR2X2 OR2X2_1808 ( .A(_abc_40319_new_n5151_), .B(_abc_40319_new_n5153_), .Y(_abc_40319_new_n5845_));
OR2X2 OR2X2_1809 ( .A(_abc_40319_new_n5844_), .B(_abc_40319_new_n5845_), .Y(_abc_40319_new_n5846_));
OR2X2 OR2X2_181 ( .A(_abc_40319_new_n1101_), .B(_abc_40319_new_n1102_), .Y(_abc_40319_new_n1103_));
OR2X2 OR2X2_1810 ( .A(_abc_40319_new_n5843_), .B(_abc_40319_new_n5846_), .Y(_abc_40319_new_n5847_));
OR2X2 OR2X2_1811 ( .A(_abc_40319_new_n5140_), .B(_abc_40319_new_n5847_), .Y(_abc_40319_new_n5848_));
OR2X2 OR2X2_1812 ( .A(_abc_40319_new_n5850_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5851_));
OR2X2 OR2X2_1813 ( .A(_abc_40319_new_n5849_), .B(_abc_40319_new_n5851_), .Y(n548));
OR2X2 OR2X2_1814 ( .A(_abc_40319_new_n5854_), .B(_abc_40319_new_n5115_), .Y(_abc_40319_new_n5855_));
OR2X2 OR2X2_1815 ( .A(_abc_40319_new_n5853_), .B(_abc_40319_new_n5855_), .Y(_abc_40319_new_n5856_));
OR2X2 OR2X2_1816 ( .A(_abc_40319_new_n5106_), .B(_abc_40319_new_n5856_), .Y(_abc_40319_new_n5857_));
OR2X2 OR2X2_1817 ( .A(_abc_40319_new_n5859_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5860_));
OR2X2 OR2X2_1818 ( .A(_abc_40319_new_n5858_), .B(_abc_40319_new_n5860_), .Y(n553));
OR2X2 OR2X2_1819 ( .A(_abc_40319_new_n5079_), .B(_abc_40319_new_n5078_), .Y(_abc_40319_new_n5864_));
OR2X2 OR2X2_182 ( .A(_abc_40319_new_n1100_), .B(_abc_40319_new_n1103_), .Y(_abc_40319_new_n1104_));
OR2X2 OR2X2_1820 ( .A(_abc_40319_new_n5863_), .B(_abc_40319_new_n5864_), .Y(_abc_40319_new_n5865_));
OR2X2 OR2X2_1821 ( .A(_abc_40319_new_n5862_), .B(_abc_40319_new_n5865_), .Y(_abc_40319_new_n5866_));
OR2X2 OR2X2_1822 ( .A(_abc_40319_new_n5070_), .B(_abc_40319_new_n5866_), .Y(_abc_40319_new_n5867_));
OR2X2 OR2X2_1823 ( .A(_abc_40319_new_n5869_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5870_));
OR2X2 OR2X2_1824 ( .A(_abc_40319_new_n5868_), .B(_abc_40319_new_n5870_), .Y(n558));
OR2X2 OR2X2_1825 ( .A(_abc_40319_new_n5048_), .B(_abc_40319_new_n5047_), .Y(_abc_40319_new_n5874_));
OR2X2 OR2X2_1826 ( .A(_abc_40319_new_n5873_), .B(_abc_40319_new_n5874_), .Y(_abc_40319_new_n5875_));
OR2X2 OR2X2_1827 ( .A(_abc_40319_new_n5872_), .B(_abc_40319_new_n5875_), .Y(_abc_40319_new_n5876_));
OR2X2 OR2X2_1828 ( .A(_abc_40319_new_n5039_), .B(_abc_40319_new_n5876_), .Y(_abc_40319_new_n5877_));
OR2X2 OR2X2_1829 ( .A(_abc_40319_new_n5879_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5880_));
OR2X2 OR2X2_183 ( .A(_abc_40319_new_n1104_), .B(_abc_40319_new_n1097_), .Y(_abc_40319_new_n1105_));
OR2X2 OR2X2_1830 ( .A(_abc_40319_new_n5878_), .B(_abc_40319_new_n5880_), .Y(n563));
OR2X2 OR2X2_1831 ( .A(_abc_40319_new_n5882_), .B(_abc_40319_new_n5014_), .Y(_abc_40319_new_n5883_));
OR2X2 OR2X2_1832 ( .A(_abc_40319_new_n5884_), .B(_abc_40319_new_n5883_), .Y(_abc_40319_new_n5885_));
OR2X2 OR2X2_1833 ( .A(_abc_40319_new_n5005_), .B(_abc_40319_new_n5885_), .Y(_abc_40319_new_n5886_));
OR2X2 OR2X2_1834 ( .A(_abc_40319_new_n5888_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5889_));
OR2X2 OR2X2_1835 ( .A(_abc_40319_new_n5887_), .B(_abc_40319_new_n5889_), .Y(n568));
OR2X2 OR2X2_1836 ( .A(_abc_40319_new_n4985_), .B(_abc_40319_new_n4984_), .Y(_abc_40319_new_n5893_));
OR2X2 OR2X2_1837 ( .A(_abc_40319_new_n5892_), .B(_abc_40319_new_n5893_), .Y(_abc_40319_new_n5894_));
OR2X2 OR2X2_1838 ( .A(_abc_40319_new_n5891_), .B(_abc_40319_new_n5894_), .Y(_abc_40319_new_n5895_));
OR2X2 OR2X2_1839 ( .A(_abc_40319_new_n4976_), .B(_abc_40319_new_n5895_), .Y(_abc_40319_new_n5896_));
OR2X2 OR2X2_184 ( .A(_abc_40319_new_n1092_), .B(_abc_40319_new_n1105_), .Y(_abc_40319_new_n1106_));
OR2X2 OR2X2_1840 ( .A(_abc_40319_new_n5898_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5899_));
OR2X2 OR2X2_1841 ( .A(_abc_40319_new_n5897_), .B(_abc_40319_new_n5899_), .Y(n573));
OR2X2 OR2X2_1842 ( .A(_abc_40319_new_n4956_), .B(_abc_40319_new_n4951_), .Y(_abc_40319_new_n5903_));
OR2X2 OR2X2_1843 ( .A(_abc_40319_new_n5902_), .B(_abc_40319_new_n5903_), .Y(_abc_40319_new_n5904_));
OR2X2 OR2X2_1844 ( .A(_abc_40319_new_n5901_), .B(_abc_40319_new_n5904_), .Y(_abc_40319_new_n5905_));
OR2X2 OR2X2_1845 ( .A(_abc_40319_new_n4944_), .B(_abc_40319_new_n5905_), .Y(_abc_40319_new_n5906_));
OR2X2 OR2X2_1846 ( .A(_abc_40319_new_n5908_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5909_));
OR2X2 OR2X2_1847 ( .A(_abc_40319_new_n5907_), .B(_abc_40319_new_n5909_), .Y(n578));
OR2X2 OR2X2_1848 ( .A(_abc_40319_new_n4915_), .B(_abc_40319_new_n4917_), .Y(_abc_40319_new_n5912_));
OR2X2 OR2X2_1849 ( .A(_abc_40319_new_n5911_), .B(_abc_40319_new_n5912_), .Y(_abc_40319_new_n5913_));
OR2X2 OR2X2_185 ( .A(_abc_40319_new_n1072_), .B(D_REG_0_), .Y(_abc_40319_new_n1109_));
OR2X2 OR2X2_1850 ( .A(_abc_40319_new_n5914_), .B(_abc_40319_new_n5913_), .Y(_abc_40319_new_n5915_));
OR2X2 OR2X2_1851 ( .A(_abc_40319_new_n4908_), .B(_abc_40319_new_n5915_), .Y(_abc_40319_new_n5916_));
OR2X2 OR2X2_1852 ( .A(_abc_40319_new_n5918_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5919_));
OR2X2 OR2X2_1853 ( .A(_abc_40319_new_n5917_), .B(_abc_40319_new_n5919_), .Y(n583));
OR2X2 OR2X2_1854 ( .A(_abc_40319_new_n5923_), .B(_abc_40319_new_n4882_), .Y(_abc_40319_new_n5924_));
OR2X2 OR2X2_1855 ( .A(_abc_40319_new_n5922_), .B(_abc_40319_new_n5924_), .Y(_abc_40319_new_n5925_));
OR2X2 OR2X2_1856 ( .A(_abc_40319_new_n5921_), .B(_abc_40319_new_n5925_), .Y(_abc_40319_new_n5926_));
OR2X2 OR2X2_1857 ( .A(_abc_40319_new_n5926_), .B(_abc_40319_new_n4873_), .Y(_abc_40319_new_n5927_));
OR2X2 OR2X2_1858 ( .A(_abc_40319_new_n5929_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5930_));
OR2X2 OR2X2_1859 ( .A(_abc_40319_new_n5928_), .B(_abc_40319_new_n5930_), .Y(n588));
OR2X2 OR2X2_186 ( .A(_abc_40319_new_n759_), .B(_abc_40319_new_n1116_), .Y(_abc_40319_new_n1117_));
OR2X2 OR2X2_1860 ( .A(_abc_40319_new_n5934_), .B(_abc_40319_new_n4850_), .Y(_abc_40319_new_n5935_));
OR2X2 OR2X2_1861 ( .A(_abc_40319_new_n5933_), .B(_abc_40319_new_n5935_), .Y(_abc_40319_new_n5936_));
OR2X2 OR2X2_1862 ( .A(_abc_40319_new_n5932_), .B(_abc_40319_new_n5936_), .Y(_abc_40319_new_n5937_));
OR2X2 OR2X2_1863 ( .A(_abc_40319_new_n5937_), .B(_abc_40319_new_n4841_), .Y(_abc_40319_new_n5938_));
OR2X2 OR2X2_1864 ( .A(_abc_40319_new_n5940_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5941_));
OR2X2 OR2X2_1865 ( .A(_abc_40319_new_n5939_), .B(_abc_40319_new_n5941_), .Y(n593));
OR2X2 OR2X2_1866 ( .A(_abc_40319_new_n5944_), .B(_abc_40319_new_n4785_), .Y(_abc_40319_new_n5945_));
OR2X2 OR2X2_1867 ( .A(_abc_40319_new_n5943_), .B(_abc_40319_new_n5945_), .Y(_abc_40319_new_n5946_));
OR2X2 OR2X2_1868 ( .A(_abc_40319_new_n5947_), .B(_abc_40319_new_n5946_), .Y(_abc_40319_new_n5948_));
OR2X2 OR2X2_1869 ( .A(_abc_40319_new_n4774_), .B(_abc_40319_new_n5948_), .Y(_abc_40319_new_n5949_));
OR2X2 OR2X2_187 ( .A(_abc_40319_new_n1127_), .B(_abc_40319_new_n1125_), .Y(_abc_40319_new_n1128_));
OR2X2 OR2X2_1870 ( .A(_abc_40319_new_n5951_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5952_));
OR2X2 OR2X2_1871 ( .A(_abc_40319_new_n5950_), .B(_abc_40319_new_n5952_), .Y(n603));
OR2X2 OR2X2_1872 ( .A(_abc_40319_new_n5956_), .B(_abc_40319_new_n4746_), .Y(_abc_40319_new_n5957_));
OR2X2 OR2X2_1873 ( .A(_abc_40319_new_n5955_), .B(_abc_40319_new_n5957_), .Y(_abc_40319_new_n5958_));
OR2X2 OR2X2_1874 ( .A(_abc_40319_new_n5954_), .B(_abc_40319_new_n5958_), .Y(_abc_40319_new_n5959_));
OR2X2 OR2X2_1875 ( .A(_abc_40319_new_n4737_), .B(_abc_40319_new_n5959_), .Y(_abc_40319_new_n5960_));
OR2X2 OR2X2_1876 ( .A(_abc_40319_new_n5962_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5963_));
OR2X2 OR2X2_1877 ( .A(_abc_40319_new_n5961_), .B(_abc_40319_new_n5963_), .Y(n608));
OR2X2 OR2X2_1878 ( .A(_abc_40319_new_n5967_), .B(_abc_40319_new_n4716_), .Y(_abc_40319_new_n5968_));
OR2X2 OR2X2_1879 ( .A(_abc_40319_new_n5966_), .B(_abc_40319_new_n5968_), .Y(_abc_40319_new_n5969_));
OR2X2 OR2X2_188 ( .A(_abc_40319_new_n1124_), .B(_abc_40319_new_n1128_), .Y(_abc_40319_new_n1129_));
OR2X2 OR2X2_1880 ( .A(_abc_40319_new_n5965_), .B(_abc_40319_new_n5969_), .Y(_abc_40319_new_n5970_));
OR2X2 OR2X2_1881 ( .A(_abc_40319_new_n4706_), .B(_abc_40319_new_n5970_), .Y(_abc_40319_new_n5971_));
OR2X2 OR2X2_1882 ( .A(_abc_40319_new_n5973_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5974_));
OR2X2 OR2X2_1883 ( .A(_abc_40319_new_n5972_), .B(_abc_40319_new_n5974_), .Y(n613));
OR2X2 OR2X2_1884 ( .A(_abc_40319_new_n5978_), .B(_abc_40319_new_n4674_), .Y(_abc_40319_new_n5979_));
OR2X2 OR2X2_1885 ( .A(_abc_40319_new_n5977_), .B(_abc_40319_new_n5979_), .Y(_abc_40319_new_n5980_));
OR2X2 OR2X2_1886 ( .A(_abc_40319_new_n5976_), .B(_abc_40319_new_n5980_), .Y(_abc_40319_new_n5981_));
OR2X2 OR2X2_1887 ( .A(_abc_40319_new_n5981_), .B(_abc_40319_new_n4664_), .Y(_abc_40319_new_n5982_));
OR2X2 OR2X2_1888 ( .A(_abc_40319_new_n5984_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5985_));
OR2X2 OR2X2_1889 ( .A(_abc_40319_new_n5983_), .B(_abc_40319_new_n5985_), .Y(n618));
OR2X2 OR2X2_189 ( .A(_abc_40319_new_n1039_), .B(REG3_REG_8_), .Y(_abc_40319_new_n1136_));
OR2X2 OR2X2_1890 ( .A(_abc_40319_new_n5989_), .B(_abc_40319_new_n4628_), .Y(_abc_40319_new_n5990_));
OR2X2 OR2X2_1891 ( .A(_abc_40319_new_n5988_), .B(_abc_40319_new_n5990_), .Y(_abc_40319_new_n5991_));
OR2X2 OR2X2_1892 ( .A(_abc_40319_new_n5987_), .B(_abc_40319_new_n5991_), .Y(_abc_40319_new_n5992_));
OR2X2 OR2X2_1893 ( .A(_abc_40319_new_n5992_), .B(_abc_40319_new_n4618_), .Y(_abc_40319_new_n5993_));
OR2X2 OR2X2_1894 ( .A(_abc_40319_new_n5995_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n5996_));
OR2X2 OR2X2_1895 ( .A(_abc_40319_new_n5994_), .B(_abc_40319_new_n5996_), .Y(n623));
OR2X2 OR2X2_1896 ( .A(_abc_40319_new_n6000_), .B(_abc_40319_new_n4597_), .Y(_abc_40319_new_n6001_));
OR2X2 OR2X2_1897 ( .A(_abc_40319_new_n5999_), .B(_abc_40319_new_n6001_), .Y(_abc_40319_new_n6002_));
OR2X2 OR2X2_1898 ( .A(_abc_40319_new_n5998_), .B(_abc_40319_new_n6002_), .Y(_abc_40319_new_n6003_));
OR2X2 OR2X2_1899 ( .A(_abc_40319_new_n6003_), .B(_abc_40319_new_n4587_), .Y(_abc_40319_new_n6004_));
OR2X2 OR2X2_19 ( .A(_abc_40319_new_n644_), .B(_abc_40319_new_n641_), .Y(_abc_40319_new_n645_));
OR2X2 OR2X2_190 ( .A(_abc_40319_new_n1141_), .B(_abc_40319_new_n1140_), .Y(_abc_40319_new_n1142_));
OR2X2 OR2X2_1900 ( .A(_abc_40319_new_n6006_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6007_));
OR2X2 OR2X2_1901 ( .A(_abc_40319_new_n6005_), .B(_abc_40319_new_n6007_), .Y(n628));
OR2X2 OR2X2_1902 ( .A(_abc_40319_new_n6011_), .B(_abc_40319_new_n4558_), .Y(_abc_40319_new_n6012_));
OR2X2 OR2X2_1903 ( .A(_abc_40319_new_n6010_), .B(_abc_40319_new_n6012_), .Y(_abc_40319_new_n6013_));
OR2X2 OR2X2_1904 ( .A(_abc_40319_new_n6009_), .B(_abc_40319_new_n6013_), .Y(_abc_40319_new_n6014_));
OR2X2 OR2X2_1905 ( .A(_abc_40319_new_n6014_), .B(_abc_40319_new_n4548_), .Y(_abc_40319_new_n6015_));
OR2X2 OR2X2_1906 ( .A(_abc_40319_new_n6017_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6018_));
OR2X2 OR2X2_1907 ( .A(_abc_40319_new_n6016_), .B(_abc_40319_new_n6018_), .Y(n633));
OR2X2 OR2X2_1908 ( .A(_abc_40319_new_n6022_), .B(_abc_40319_new_n4522_), .Y(_abc_40319_new_n6023_));
OR2X2 OR2X2_1909 ( .A(_abc_40319_new_n6021_), .B(_abc_40319_new_n6023_), .Y(_abc_40319_new_n6024_));
OR2X2 OR2X2_191 ( .A(_abc_40319_new_n1143_), .B(_abc_40319_new_n1144_), .Y(_abc_40319_new_n1145_));
OR2X2 OR2X2_1910 ( .A(_abc_40319_new_n6020_), .B(_abc_40319_new_n6024_), .Y(_abc_40319_new_n6025_));
OR2X2 OR2X2_1911 ( .A(_abc_40319_new_n4510_), .B(_abc_40319_new_n6025_), .Y(_abc_40319_new_n6026_));
OR2X2 OR2X2_1912 ( .A(_abc_40319_new_n6028_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6029_));
OR2X2 OR2X2_1913 ( .A(_abc_40319_new_n6027_), .B(_abc_40319_new_n6029_), .Y(n638));
OR2X2 OR2X2_1914 ( .A(_abc_40319_new_n6032_), .B(_abc_40319_new_n5721_), .Y(_abc_40319_new_n6033_));
OR2X2 OR2X2_1915 ( .A(_abc_40319_new_n5695_), .B(_abc_40319_new_n6033_), .Y(_abc_40319_new_n6034_));
OR2X2 OR2X2_1916 ( .A(_abc_40319_new_n6031_), .B(_abc_40319_new_n6034_), .Y(_abc_40319_new_n6035_));
OR2X2 OR2X2_1917 ( .A(_abc_40319_new_n5712_), .B(_abc_40319_new_n6035_), .Y(_abc_40319_new_n6036_));
OR2X2 OR2X2_1918 ( .A(_abc_40319_new_n6038_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6039_));
OR2X2 OR2X2_1919 ( .A(_abc_40319_new_n6037_), .B(_abc_40319_new_n6039_), .Y(n643));
OR2X2 OR2X2_192 ( .A(_abc_40319_new_n1142_), .B(_abc_40319_new_n1145_), .Y(_abc_40319_new_n1146_));
OR2X2 OR2X2_1920 ( .A(_abc_40319_new_n4313_), .B(_abc_40319_new_n6042_), .Y(_abc_40319_new_n6043_));
OR2X2 OR2X2_1921 ( .A(_abc_40319_new_n6041_), .B(_abc_40319_new_n6043_), .Y(_abc_40319_new_n6044_));
OR2X2 OR2X2_1922 ( .A(_abc_40319_new_n6046_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6047_));
OR2X2 OR2X2_1923 ( .A(_abc_40319_new_n6045_), .B(_abc_40319_new_n6047_), .Y(n648));
OR2X2 OR2X2_1924 ( .A(_abc_40319_new_n4313_), .B(_abc_40319_new_n6050_), .Y(_abc_40319_new_n6051_));
OR2X2 OR2X2_1925 ( .A(_abc_40319_new_n6049_), .B(_abc_40319_new_n6051_), .Y(_abc_40319_new_n6052_));
OR2X2 OR2X2_1926 ( .A(_abc_40319_new_n6054_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6055_));
OR2X2 OR2X2_1927 ( .A(_abc_40319_new_n6053_), .B(_abc_40319_new_n6055_), .Y(n653));
OR2X2 OR2X2_1928 ( .A(_abc_40319_new_n6060_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6061_));
OR2X2 OR2X2_1929 ( .A(_abc_40319_new_n6058_), .B(_abc_40319_new_n6061_), .Y(n658));
OR2X2 OR2X2_193 ( .A(_abc_40319_new_n1135_), .B(_abc_40319_new_n1148_), .Y(_abc_40319_new_n1149_));
OR2X2 OR2X2_1930 ( .A(_abc_40319_new_n6064_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6065_));
OR2X2 OR2X2_1931 ( .A(_abc_40319_new_n6063_), .B(_abc_40319_new_n6065_), .Y(n663));
OR2X2 OR2X2_1932 ( .A(_abc_40319_new_n6068_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6069_));
OR2X2 OR2X2_1933 ( .A(_abc_40319_new_n6067_), .B(_abc_40319_new_n6069_), .Y(n668));
OR2X2 OR2X2_1934 ( .A(_abc_40319_new_n6072_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6073_));
OR2X2 OR2X2_1935 ( .A(_abc_40319_new_n6071_), .B(_abc_40319_new_n6073_), .Y(n673));
OR2X2 OR2X2_1936 ( .A(_abc_40319_new_n6076_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6077_));
OR2X2 OR2X2_1937 ( .A(_abc_40319_new_n6075_), .B(_abc_40319_new_n6077_), .Y(n678));
OR2X2 OR2X2_1938 ( .A(_abc_40319_new_n6080_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6081_));
OR2X2 OR2X2_1939 ( .A(_abc_40319_new_n6079_), .B(_abc_40319_new_n6081_), .Y(n683));
OR2X2 OR2X2_194 ( .A(_abc_40319_new_n1153_), .B(_abc_40319_new_n1154_), .Y(_abc_40319_new_n1155_));
OR2X2 OR2X2_1940 ( .A(_abc_40319_new_n6084_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6085_));
OR2X2 OR2X2_1941 ( .A(_abc_40319_new_n6083_), .B(_abc_40319_new_n6085_), .Y(n688));
OR2X2 OR2X2_1942 ( .A(_abc_40319_new_n6088_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6089_));
OR2X2 OR2X2_1943 ( .A(_abc_40319_new_n6087_), .B(_abc_40319_new_n6089_), .Y(n693));
OR2X2 OR2X2_1944 ( .A(_abc_40319_new_n6092_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6093_));
OR2X2 OR2X2_1945 ( .A(_abc_40319_new_n6091_), .B(_abc_40319_new_n6093_), .Y(n698));
OR2X2 OR2X2_1946 ( .A(_abc_40319_new_n6096_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6097_));
OR2X2 OR2X2_1947 ( .A(_abc_40319_new_n6095_), .B(_abc_40319_new_n6097_), .Y(n703));
OR2X2 OR2X2_1948 ( .A(_abc_40319_new_n6100_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6101_));
OR2X2 OR2X2_1949 ( .A(_abc_40319_new_n6099_), .B(_abc_40319_new_n6101_), .Y(n708));
OR2X2 OR2X2_195 ( .A(_abc_40319_new_n1157_), .B(_abc_40319_new_n1159_), .Y(_abc_40319_new_n1160_));
OR2X2 OR2X2_1950 ( .A(_abc_40319_new_n6104_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6105_));
OR2X2 OR2X2_1951 ( .A(_abc_40319_new_n6103_), .B(_abc_40319_new_n6105_), .Y(n713));
OR2X2 OR2X2_1952 ( .A(_abc_40319_new_n6108_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6109_));
OR2X2 OR2X2_1953 ( .A(_abc_40319_new_n6107_), .B(_abc_40319_new_n6109_), .Y(n718));
OR2X2 OR2X2_1954 ( .A(_abc_40319_new_n6112_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6113_));
OR2X2 OR2X2_1955 ( .A(_abc_40319_new_n6111_), .B(_abc_40319_new_n6113_), .Y(n723));
OR2X2 OR2X2_1956 ( .A(_abc_40319_new_n6116_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6117_));
OR2X2 OR2X2_1957 ( .A(_abc_40319_new_n6115_), .B(_abc_40319_new_n6117_), .Y(n728));
OR2X2 OR2X2_1958 ( .A(_abc_40319_new_n6120_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6121_));
OR2X2 OR2X2_1959 ( .A(_abc_40319_new_n6119_), .B(_abc_40319_new_n6121_), .Y(n733));
OR2X2 OR2X2_196 ( .A(_abc_40319_new_n1156_), .B(_abc_40319_new_n1161_), .Y(_abc_40319_new_n1162_));
OR2X2 OR2X2_1960 ( .A(_abc_40319_new_n6124_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6125_));
OR2X2 OR2X2_1961 ( .A(_abc_40319_new_n6123_), .B(_abc_40319_new_n6125_), .Y(n738));
OR2X2 OR2X2_1962 ( .A(_abc_40319_new_n6128_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6129_));
OR2X2 OR2X2_1963 ( .A(_abc_40319_new_n6127_), .B(_abc_40319_new_n6129_), .Y(n743));
OR2X2 OR2X2_1964 ( .A(_abc_40319_new_n6132_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6133_));
OR2X2 OR2X2_1965 ( .A(_abc_40319_new_n6131_), .B(_abc_40319_new_n6133_), .Y(n748));
OR2X2 OR2X2_1966 ( .A(_abc_40319_new_n6136_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6137_));
OR2X2 OR2X2_1967 ( .A(_abc_40319_new_n6135_), .B(_abc_40319_new_n6137_), .Y(n753));
OR2X2 OR2X2_1968 ( .A(_abc_40319_new_n6140_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6141_));
OR2X2 OR2X2_1969 ( .A(_abc_40319_new_n6139_), .B(_abc_40319_new_n6141_), .Y(n758));
OR2X2 OR2X2_197 ( .A(_abc_40319_new_n1162_), .B(_abc_40319_new_n1163_), .Y(_abc_40319_new_n1164_));
OR2X2 OR2X2_1970 ( .A(_abc_40319_new_n6144_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6145_));
OR2X2 OR2X2_1971 ( .A(_abc_40319_new_n6143_), .B(_abc_40319_new_n6145_), .Y(n763));
OR2X2 OR2X2_1972 ( .A(_abc_40319_new_n6148_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6149_));
OR2X2 OR2X2_1973 ( .A(_abc_40319_new_n6147_), .B(_abc_40319_new_n6149_), .Y(n768));
OR2X2 OR2X2_1974 ( .A(_abc_40319_new_n6152_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6153_));
OR2X2 OR2X2_1975 ( .A(_abc_40319_new_n6151_), .B(_abc_40319_new_n6153_), .Y(n773));
OR2X2 OR2X2_1976 ( .A(_abc_40319_new_n6156_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6157_));
OR2X2 OR2X2_1977 ( .A(_abc_40319_new_n6155_), .B(_abc_40319_new_n6157_), .Y(n778));
OR2X2 OR2X2_1978 ( .A(_abc_40319_new_n6160_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6161_));
OR2X2 OR2X2_1979 ( .A(_abc_40319_new_n6159_), .B(_abc_40319_new_n6161_), .Y(n783));
OR2X2 OR2X2_198 ( .A(_abc_40319_new_n1170_), .B(_abc_40319_new_n1169_), .Y(_abc_40319_new_n1171_));
OR2X2 OR2X2_1980 ( .A(_abc_40319_new_n6164_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6165_));
OR2X2 OR2X2_1981 ( .A(_abc_40319_new_n6163_), .B(_abc_40319_new_n6165_), .Y(n788));
OR2X2 OR2X2_1982 ( .A(_abc_40319_new_n6168_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6169_));
OR2X2 OR2X2_1983 ( .A(_abc_40319_new_n6167_), .B(_abc_40319_new_n6169_), .Y(n793));
OR2X2 OR2X2_1984 ( .A(_abc_40319_new_n6172_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6173_));
OR2X2 OR2X2_1985 ( .A(_abc_40319_new_n6171_), .B(_abc_40319_new_n6173_), .Y(n798));
OR2X2 OR2X2_1986 ( .A(_abc_40319_new_n6176_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6177_));
OR2X2 OR2X2_1987 ( .A(_abc_40319_new_n6175_), .B(_abc_40319_new_n6177_), .Y(n803));
OR2X2 OR2X2_1988 ( .A(_abc_40319_new_n6180_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6181_));
OR2X2 OR2X2_1989 ( .A(_abc_40319_new_n6179_), .B(_abc_40319_new_n6181_), .Y(n808));
OR2X2 OR2X2_199 ( .A(_abc_40319_new_n1174_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n1175_));
OR2X2 OR2X2_1990 ( .A(_abc_40319_new_n6184_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6185_));
OR2X2 OR2X2_1991 ( .A(_abc_40319_new_n6183_), .B(_abc_40319_new_n6185_), .Y(n813));
OR2X2 OR2X2_1992 ( .A(_abc_40319_new_n6189_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6190_));
OR2X2 OR2X2_1993 ( .A(_abc_40319_new_n6187_), .B(_abc_40319_new_n6190_), .Y(n1058));
OR2X2 OR2X2_1994 ( .A(_abc_40319_new_n6193_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6194_));
OR2X2 OR2X2_1995 ( .A(_abc_40319_new_n6192_), .B(_abc_40319_new_n6194_), .Y(n1062));
OR2X2 OR2X2_1996 ( .A(_abc_40319_new_n6197_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6198_));
OR2X2 OR2X2_1997 ( .A(_abc_40319_new_n6196_), .B(_abc_40319_new_n6198_), .Y(n1066));
OR2X2 OR2X2_1998 ( .A(_abc_40319_new_n6201_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6202_));
OR2X2 OR2X2_1999 ( .A(_abc_40319_new_n6200_), .B(_abc_40319_new_n6202_), .Y(n1070));
OR2X2 OR2X2_2 ( .A(IR_REG_23_), .B(IR_REG_18_), .Y(_abc_40319_new_n567_));
OR2X2 OR2X2_20 ( .A(_abc_40319_new_n650_), .B(_abc_40319_new_n564_), .Y(_abc_40319_new_n651_));
OR2X2 OR2X2_200 ( .A(_abc_40319_new_n1172_), .B(_abc_40319_new_n1175_), .Y(_abc_40319_new_n1176_));
OR2X2 OR2X2_2000 ( .A(_abc_40319_new_n6205_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6206_));
OR2X2 OR2X2_2001 ( .A(_abc_40319_new_n6204_), .B(_abc_40319_new_n6206_), .Y(n1074));
OR2X2 OR2X2_2002 ( .A(_abc_40319_new_n6209_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6210_));
OR2X2 OR2X2_2003 ( .A(_abc_40319_new_n6208_), .B(_abc_40319_new_n6210_), .Y(n1078));
OR2X2 OR2X2_2004 ( .A(_abc_40319_new_n6213_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6214_));
OR2X2 OR2X2_2005 ( .A(_abc_40319_new_n6212_), .B(_abc_40319_new_n6214_), .Y(n1082));
OR2X2 OR2X2_2006 ( .A(_abc_40319_new_n6217_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6218_));
OR2X2 OR2X2_2007 ( .A(_abc_40319_new_n6216_), .B(_abc_40319_new_n6218_), .Y(n1086));
OR2X2 OR2X2_2008 ( .A(_abc_40319_new_n6221_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6222_));
OR2X2 OR2X2_2009 ( .A(_abc_40319_new_n6220_), .B(_abc_40319_new_n6222_), .Y(n1090));
OR2X2 OR2X2_201 ( .A(_abc_40319_new_n1165_), .B(_abc_40319_new_n1176_), .Y(_abc_40319_new_n1177_));
OR2X2 OR2X2_2010 ( .A(_abc_40319_new_n6225_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6226_));
OR2X2 OR2X2_2011 ( .A(_abc_40319_new_n6224_), .B(_abc_40319_new_n6226_), .Y(n1094));
OR2X2 OR2X2_2012 ( .A(_abc_40319_new_n6229_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6230_));
OR2X2 OR2X2_2013 ( .A(_abc_40319_new_n6228_), .B(_abc_40319_new_n6230_), .Y(n1098));
OR2X2 OR2X2_2014 ( .A(_abc_40319_new_n6233_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6234_));
OR2X2 OR2X2_2015 ( .A(_abc_40319_new_n6232_), .B(_abc_40319_new_n6234_), .Y(n1102));
OR2X2 OR2X2_2016 ( .A(_abc_40319_new_n6237_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6238_));
OR2X2 OR2X2_2017 ( .A(_abc_40319_new_n6236_), .B(_abc_40319_new_n6238_), .Y(n1106));
OR2X2 OR2X2_2018 ( .A(_abc_40319_new_n6241_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6242_));
OR2X2 OR2X2_2019 ( .A(_abc_40319_new_n6240_), .B(_abc_40319_new_n6242_), .Y(n1110));
OR2X2 OR2X2_202 ( .A(_abc_40319_new_n1177_), .B(_abc_40319_new_n1150_), .Y(_abc_40319_new_n1178_));
OR2X2 OR2X2_2020 ( .A(_abc_40319_new_n6245_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6246_));
OR2X2 OR2X2_2021 ( .A(_abc_40319_new_n6244_), .B(_abc_40319_new_n6246_), .Y(n1114));
OR2X2 OR2X2_2022 ( .A(_abc_40319_new_n6249_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6250_));
OR2X2 OR2X2_2023 ( .A(_abc_40319_new_n6248_), .B(_abc_40319_new_n6250_), .Y(n1118));
OR2X2 OR2X2_2024 ( .A(_abc_40319_new_n6253_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6254_));
OR2X2 OR2X2_2025 ( .A(_abc_40319_new_n6252_), .B(_abc_40319_new_n6254_), .Y(n1122));
OR2X2 OR2X2_2026 ( .A(_abc_40319_new_n6257_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6258_));
OR2X2 OR2X2_2027 ( .A(_abc_40319_new_n6256_), .B(_abc_40319_new_n6258_), .Y(n1126));
OR2X2 OR2X2_2028 ( .A(_abc_40319_new_n6261_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6262_));
OR2X2 OR2X2_2029 ( .A(_abc_40319_new_n6260_), .B(_abc_40319_new_n6262_), .Y(n1130));
OR2X2 OR2X2_203 ( .A(_abc_40319_new_n1131_), .B(_abc_40319_new_n1178_), .Y(n1331));
OR2X2 OR2X2_2030 ( .A(_abc_40319_new_n6265_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6266_));
OR2X2 OR2X2_2031 ( .A(_abc_40319_new_n6264_), .B(_abc_40319_new_n6266_), .Y(n1134));
OR2X2 OR2X2_2032 ( .A(_abc_40319_new_n6269_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6270_));
OR2X2 OR2X2_2033 ( .A(_abc_40319_new_n6268_), .B(_abc_40319_new_n6270_), .Y(n1138));
OR2X2 OR2X2_2034 ( .A(_abc_40319_new_n6273_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6274_));
OR2X2 OR2X2_2035 ( .A(_abc_40319_new_n6272_), .B(_abc_40319_new_n6274_), .Y(n1142));
OR2X2 OR2X2_2036 ( .A(_abc_40319_new_n6277_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6278_));
OR2X2 OR2X2_2037 ( .A(_abc_40319_new_n6276_), .B(_abc_40319_new_n6278_), .Y(n1146));
OR2X2 OR2X2_2038 ( .A(_abc_40319_new_n6281_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6282_));
OR2X2 OR2X2_2039 ( .A(_abc_40319_new_n6280_), .B(_abc_40319_new_n6282_), .Y(n1150));
OR2X2 OR2X2_204 ( .A(_abc_40319_new_n1199_), .B(REG3_REG_27_), .Y(_abc_40319_new_n1200_));
OR2X2 OR2X2_2040 ( .A(_abc_40319_new_n6285_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6286_));
OR2X2 OR2X2_2041 ( .A(_abc_40319_new_n6284_), .B(_abc_40319_new_n6286_), .Y(n1154));
OR2X2 OR2X2_2042 ( .A(_abc_40319_new_n6289_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6290_));
OR2X2 OR2X2_2043 ( .A(_abc_40319_new_n6288_), .B(_abc_40319_new_n6290_), .Y(n1158));
OR2X2 OR2X2_2044 ( .A(_abc_40319_new_n6293_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6294_));
OR2X2 OR2X2_2045 ( .A(_abc_40319_new_n6292_), .B(_abc_40319_new_n6294_), .Y(n1162));
OR2X2 OR2X2_2046 ( .A(_abc_40319_new_n6297_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6298_));
OR2X2 OR2X2_2047 ( .A(_abc_40319_new_n6296_), .B(_abc_40319_new_n6298_), .Y(n1166));
OR2X2 OR2X2_2048 ( .A(_abc_40319_new_n6301_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6302_));
OR2X2 OR2X2_2049 ( .A(_abc_40319_new_n6300_), .B(_abc_40319_new_n6302_), .Y(n1170));
OR2X2 OR2X2_205 ( .A(_abc_40319_new_n1206_), .B(_abc_40319_new_n1207_), .Y(_abc_40319_new_n1208_));
OR2X2 OR2X2_2050 ( .A(_abc_40319_new_n6305_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6306_));
OR2X2 OR2X2_2051 ( .A(_abc_40319_new_n6304_), .B(_abc_40319_new_n6306_), .Y(n1174));
OR2X2 OR2X2_2052 ( .A(_abc_40319_new_n6309_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6310_));
OR2X2 OR2X2_2053 ( .A(_abc_40319_new_n6308_), .B(_abc_40319_new_n6310_), .Y(n1178));
OR2X2 OR2X2_2054 ( .A(_abc_40319_new_n6313_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n6314_));
OR2X2 OR2X2_2055 ( .A(_abc_40319_new_n6312_), .B(_abc_40319_new_n6314_), .Y(n1182));
OR2X2 OR2X2_206 ( .A(_abc_40319_new_n1208_), .B(_abc_40319_new_n1205_), .Y(_abc_40319_new_n1209_));
OR2X2 OR2X2_207 ( .A(_abc_40319_new_n1204_), .B(_abc_40319_new_n1209_), .Y(_abc_40319_new_n1210_));
OR2X2 OR2X2_208 ( .A(_abc_40319_new_n1211_), .B(_abc_40319_new_n1181_), .Y(_abc_40319_new_n1212_));
OR2X2 OR2X2_209 ( .A(_abc_40319_new_n1214_), .B(_abc_40319_new_n1213_), .Y(_abc_40319_new_n1215_));
OR2X2 OR2X2_21 ( .A(_abc_40319_new_n653_), .B(_abc_40319_new_n654_), .Y(_abc_40319_new_n655_));
OR2X2 OR2X2_210 ( .A(_abc_40319_new_n1217_), .B(_abc_40319_new_n1218_), .Y(_abc_40319_new_n1219_));
OR2X2 OR2X2_211 ( .A(_abc_40319_new_n1219_), .B(_abc_40319_new_n1212_), .Y(_abc_40319_new_n1222_));
OR2X2 OR2X2_212 ( .A(_abc_40319_new_n1198_), .B(REG3_REG_26_), .Y(_abc_40319_new_n1227_));
OR2X2 OR2X2_213 ( .A(_abc_40319_new_n1231_), .B(_abc_40319_new_n1232_), .Y(_abc_40319_new_n1233_));
OR2X2 OR2X2_214 ( .A(_abc_40319_new_n1233_), .B(_abc_40319_new_n1230_), .Y(_abc_40319_new_n1234_));
OR2X2 OR2X2_215 ( .A(_abc_40319_new_n1229_), .B(_abc_40319_new_n1234_), .Y(_abc_40319_new_n1235_));
OR2X2 OR2X2_216 ( .A(_abc_40319_new_n1236_), .B(_abc_40319_new_n1225_), .Y(_abc_40319_new_n1237_));
OR2X2 OR2X2_217 ( .A(_abc_40319_new_n1240_), .B(_abc_40319_new_n1239_), .Y(_abc_40319_new_n1241_));
OR2X2 OR2X2_218 ( .A(_abc_40319_new_n1243_), .B(_abc_40319_new_n1244_), .Y(_abc_40319_new_n1245_));
OR2X2 OR2X2_219 ( .A(_abc_40319_new_n1197_), .B(REG3_REG_25_), .Y(_abc_40319_new_n1252_));
OR2X2 OR2X2_22 ( .A(_abc_40319_new_n656_), .B(_abc_40319_new_n598_), .Y(_abc_40319_new_n657_));
OR2X2 OR2X2_220 ( .A(_abc_40319_new_n1256_), .B(_abc_40319_new_n1257_), .Y(_abc_40319_new_n1258_));
OR2X2 OR2X2_221 ( .A(_abc_40319_new_n1258_), .B(_abc_40319_new_n1255_), .Y(_abc_40319_new_n1259_));
OR2X2 OR2X2_222 ( .A(_abc_40319_new_n1254_), .B(_abc_40319_new_n1259_), .Y(_abc_40319_new_n1260_));
OR2X2 OR2X2_223 ( .A(_abc_40319_new_n1261_), .B(_abc_40319_new_n1250_), .Y(_abc_40319_new_n1262_));
OR2X2 OR2X2_224 ( .A(_abc_40319_new_n1265_), .B(_abc_40319_new_n1264_), .Y(_abc_40319_new_n1266_));
OR2X2 OR2X2_225 ( .A(_abc_40319_new_n1268_), .B(_abc_40319_new_n1269_), .Y(_abc_40319_new_n1270_));
OR2X2 OR2X2_226 ( .A(_abc_40319_new_n1196_), .B(REG3_REG_24_), .Y(_abc_40319_new_n1277_));
OR2X2 OR2X2_227 ( .A(_abc_40319_new_n1281_), .B(_abc_40319_new_n1282_), .Y(_abc_40319_new_n1283_));
OR2X2 OR2X2_228 ( .A(_abc_40319_new_n1283_), .B(_abc_40319_new_n1280_), .Y(_abc_40319_new_n1284_));
OR2X2 OR2X2_229 ( .A(_abc_40319_new_n1279_), .B(_abc_40319_new_n1284_), .Y(_abc_40319_new_n1285_));
OR2X2 OR2X2_23 ( .A(_abc_40319_new_n658_), .B(_abc_40319_new_n640_), .Y(_abc_40319_new_n659_));
OR2X2 OR2X2_230 ( .A(_abc_40319_new_n1286_), .B(_abc_40319_new_n1275_), .Y(_abc_40319_new_n1287_));
OR2X2 OR2X2_231 ( .A(_abc_40319_new_n1289_), .B(_abc_40319_new_n1288_), .Y(_abc_40319_new_n1290_));
OR2X2 OR2X2_232 ( .A(_abc_40319_new_n1292_), .B(_abc_40319_new_n1293_), .Y(_abc_40319_new_n1294_));
OR2X2 OR2X2_233 ( .A(_abc_40319_new_n1270_), .B(_abc_40319_new_n1263_), .Y(_abc_40319_new_n1301_));
OR2X2 OR2X2_234 ( .A(_abc_40319_new_n1303_), .B(_abc_40319_new_n1247_), .Y(_abc_40319_new_n1304_));
OR2X2 OR2X2_235 ( .A(_abc_40319_new_n1195_), .B(REG3_REG_23_), .Y(_abc_40319_new_n1309_));
OR2X2 OR2X2_236 ( .A(_abc_40319_new_n1313_), .B(_abc_40319_new_n1314_), .Y(_abc_40319_new_n1315_));
OR2X2 OR2X2_237 ( .A(_abc_40319_new_n1315_), .B(_abc_40319_new_n1312_), .Y(_abc_40319_new_n1316_));
OR2X2 OR2X2_238 ( .A(_abc_40319_new_n1311_), .B(_abc_40319_new_n1316_), .Y(_abc_40319_new_n1317_));
OR2X2 OR2X2_239 ( .A(_abc_40319_new_n1318_), .B(_abc_40319_new_n1307_), .Y(_abc_40319_new_n1319_));
OR2X2 OR2X2_24 ( .A(_abc_40319_new_n649_), .B(_abc_40319_new_n563_), .Y(_abc_40319_new_n667_));
OR2X2 OR2X2_240 ( .A(_abc_40319_new_n1321_), .B(_abc_40319_new_n1320_), .Y(_abc_40319_new_n1322_));
OR2X2 OR2X2_241 ( .A(_abc_40319_new_n1322_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1323_));
OR2X2 OR2X2_242 ( .A(_abc_40319_new_n1324_), .B(_abc_40319_new_n768_), .Y(_abc_40319_new_n1325_));
OR2X2 OR2X2_243 ( .A(_abc_40319_new_n1326_), .B(_abc_40319_new_n1319_), .Y(_abc_40319_new_n1328_));
OR2X2 OR2X2_244 ( .A(_abc_40319_new_n1194_), .B(REG3_REG_22_), .Y(_abc_40319_new_n1332_));
OR2X2 OR2X2_245 ( .A(_abc_40319_new_n1336_), .B(_abc_40319_new_n1337_), .Y(_abc_40319_new_n1338_));
OR2X2 OR2X2_246 ( .A(_abc_40319_new_n1338_), .B(_abc_40319_new_n1335_), .Y(_abc_40319_new_n1339_));
OR2X2 OR2X2_247 ( .A(_abc_40319_new_n1334_), .B(_abc_40319_new_n1339_), .Y(_abc_40319_new_n1340_));
OR2X2 OR2X2_248 ( .A(_abc_40319_new_n1341_), .B(_abc_40319_new_n1330_), .Y(_abc_40319_new_n1342_));
OR2X2 OR2X2_249 ( .A(_abc_40319_new_n1344_), .B(_abc_40319_new_n1343_), .Y(_abc_40319_new_n1345_));
OR2X2 OR2X2_25 ( .A(_abc_40319_new_n668_), .B(_abc_40319_new_n524_), .Y(_abc_40319_new_n669_));
OR2X2 OR2X2_250 ( .A(_abc_40319_new_n1347_), .B(_abc_40319_new_n1348_), .Y(_abc_40319_new_n1349_));
OR2X2 OR2X2_251 ( .A(_abc_40319_new_n1350_), .B(_abc_40319_new_n1342_), .Y(_abc_40319_new_n1352_));
OR2X2 OR2X2_252 ( .A(_abc_40319_new_n1353_), .B(_abc_40319_new_n648_), .Y(_abc_40319_new_n1354_));
OR2X2 OR2X2_253 ( .A(_abc_40319_new_n1356_), .B(_abc_40319_new_n1357_), .Y(_abc_40319_new_n1358_));
OR2X2 OR2X2_254 ( .A(_abc_40319_new_n640_), .B(DATAI_18_), .Y(_abc_40319_new_n1362_));
OR2X2 OR2X2_255 ( .A(_abc_40319_new_n1190_), .B(REG3_REG_18_), .Y(_abc_40319_new_n1367_));
OR2X2 OR2X2_256 ( .A(_abc_40319_new_n1371_), .B(_abc_40319_new_n1370_), .Y(_abc_40319_new_n1372_));
OR2X2 OR2X2_257 ( .A(_abc_40319_new_n1372_), .B(_abc_40319_new_n1369_), .Y(_abc_40319_new_n1373_));
OR2X2 OR2X2_258 ( .A(_abc_40319_new_n1373_), .B(_abc_40319_new_n1365_), .Y(_abc_40319_new_n1374_));
OR2X2 OR2X2_259 ( .A(_abc_40319_new_n1375_), .B(_abc_40319_new_n1364_), .Y(_abc_40319_new_n1376_));
OR2X2 OR2X2_26 ( .A(_abc_40319_new_n674_), .B(IR_REG_3_), .Y(_abc_40319_new_n675_));
OR2X2 OR2X2_260 ( .A(_abc_40319_new_n1378_), .B(_abc_40319_new_n1377_), .Y(_abc_40319_new_n1379_));
OR2X2 OR2X2_261 ( .A(_abc_40319_new_n1381_), .B(_abc_40319_new_n1382_), .Y(_abc_40319_new_n1383_));
OR2X2 OR2X2_262 ( .A(_abc_40319_new_n1384_), .B(_abc_40319_new_n1376_), .Y(_abc_40319_new_n1386_));
OR2X2 OR2X2_263 ( .A(_abc_40319_new_n1391_), .B(_abc_40319_new_n1388_), .Y(_abc_40319_new_n1392_));
OR2X2 OR2X2_264 ( .A(_abc_40319_new_n1393_), .B(_abc_40319_new_n1387_), .Y(_abc_40319_new_n1394_));
OR2X2 OR2X2_265 ( .A(_abc_40319_new_n640_), .B(DATAI_16_), .Y(_abc_40319_new_n1397_));
OR2X2 OR2X2_266 ( .A(_abc_40319_new_n1400_), .B(_abc_40319_new_n1401_), .Y(_abc_40319_new_n1402_));
OR2X2 OR2X2_267 ( .A(_abc_40319_new_n1188_), .B(REG3_REG_16_), .Y(_abc_40319_new_n1403_));
OR2X2 OR2X2_268 ( .A(_abc_40319_new_n1408_), .B(_abc_40319_new_n1407_), .Y(_abc_40319_new_n1409_));
OR2X2 OR2X2_269 ( .A(_abc_40319_new_n1402_), .B(_abc_40319_new_n1409_), .Y(_abc_40319_new_n1410_));
OR2X2 OR2X2_27 ( .A(_abc_40319_new_n679_), .B(_abc_40319_new_n537_), .Y(_abc_40319_new_n680_));
OR2X2 OR2X2_270 ( .A(_abc_40319_new_n1411_), .B(_abc_40319_new_n1399_), .Y(_abc_40319_new_n1412_));
OR2X2 OR2X2_271 ( .A(_abc_40319_new_n1414_), .B(_abc_40319_new_n1415_), .Y(_abc_40319_new_n1416_));
OR2X2 OR2X2_272 ( .A(_abc_40319_new_n1416_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1417_));
OR2X2 OR2X2_273 ( .A(_abc_40319_new_n1418_), .B(_abc_40319_new_n768_), .Y(_abc_40319_new_n1419_));
OR2X2 OR2X2_274 ( .A(_abc_40319_new_n1388_), .B(_abc_40319_new_n555_), .Y(_abc_40319_new_n1424_));
OR2X2 OR2X2_275 ( .A(_abc_40319_new_n1426_), .B(_abc_40319_new_n1427_), .Y(_abc_40319_new_n1428_));
OR2X2 OR2X2_276 ( .A(_abc_40319_new_n640_), .B(DATAI_17_), .Y(_abc_40319_new_n1432_));
OR2X2 OR2X2_277 ( .A(_abc_40319_new_n1435_), .B(_abc_40319_new_n1436_), .Y(_abc_40319_new_n1437_));
OR2X2 OR2X2_278 ( .A(_abc_40319_new_n1404_), .B(REG3_REG_17_), .Y(_abc_40319_new_n1439_));
OR2X2 OR2X2_279 ( .A(_abc_40319_new_n1442_), .B(_abc_40319_new_n1441_), .Y(_abc_40319_new_n1443_));
OR2X2 OR2X2_28 ( .A(_abc_40319_new_n682_), .B(_abc_40319_new_n683_), .Y(_abc_40319_new_n684_));
OR2X2 OR2X2_280 ( .A(_abc_40319_new_n1437_), .B(_abc_40319_new_n1443_), .Y(_abc_40319_new_n1444_));
OR2X2 OR2X2_281 ( .A(_abc_40319_new_n1445_), .B(_abc_40319_new_n1434_), .Y(_abc_40319_new_n1446_));
OR2X2 OR2X2_282 ( .A(_abc_40319_new_n1448_), .B(_abc_40319_new_n1449_), .Y(_abc_40319_new_n1450_));
OR2X2 OR2X2_283 ( .A(_abc_40319_new_n1450_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1451_));
OR2X2 OR2X2_284 ( .A(_abc_40319_new_n1452_), .B(_abc_40319_new_n768_), .Y(_abc_40319_new_n1453_));
OR2X2 OR2X2_285 ( .A(_abc_40319_new_n1461_), .B(_abc_40319_new_n1389_), .Y(_abc_40319_new_n1462_));
OR2X2 OR2X2_286 ( .A(_abc_40319_new_n1464_), .B(_abc_40319_new_n1465_), .Y(_abc_40319_new_n1466_));
OR2X2 OR2X2_287 ( .A(_abc_40319_new_n640_), .B(DATAI_15_), .Y(_abc_40319_new_n1470_));
OR2X2 OR2X2_288 ( .A(_abc_40319_new_n1473_), .B(_abc_40319_new_n1474_), .Y(_abc_40319_new_n1475_));
OR2X2 OR2X2_289 ( .A(_abc_40319_new_n1478_), .B(REG3_REG_15_), .Y(_abc_40319_new_n1479_));
OR2X2 OR2X2_29 ( .A(_abc_40319_new_n640_), .B(DATAI_5_), .Y(_abc_40319_new_n688_));
OR2X2 OR2X2_290 ( .A(_abc_40319_new_n1476_), .B(_abc_40319_new_n1481_), .Y(_abc_40319_new_n1482_));
OR2X2 OR2X2_291 ( .A(_abc_40319_new_n1475_), .B(_abc_40319_new_n1482_), .Y(_abc_40319_new_n1483_));
OR2X2 OR2X2_292 ( .A(_abc_40319_new_n1484_), .B(_abc_40319_new_n1472_), .Y(_abc_40319_new_n1485_));
OR2X2 OR2X2_293 ( .A(_abc_40319_new_n1486_), .B(_abc_40319_new_n1487_), .Y(_abc_40319_new_n1488_));
OR2X2 OR2X2_294 ( .A(_abc_40319_new_n1488_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1489_));
OR2X2 OR2X2_295 ( .A(_abc_40319_new_n1490_), .B(_abc_40319_new_n768_), .Y(_abc_40319_new_n1491_));
OR2X2 OR2X2_296 ( .A(_abc_40319_new_n1492_), .B(_abc_40319_new_n1485_), .Y(_abc_40319_new_n1494_));
OR2X2 OR2X2_297 ( .A(_abc_40319_new_n1496_), .B(_abc_40319_new_n1459_), .Y(_abc_40319_new_n1497_));
OR2X2 OR2X2_298 ( .A(_abc_40319_new_n1499_), .B(_abc_40319_new_n1500_), .Y(_abc_40319_new_n1501_));
OR2X2 OR2X2_299 ( .A(_abc_40319_new_n640_), .B(DATAI_14_), .Y(_abc_40319_new_n1505_));
OR2X2 OR2X2_3 ( .A(_abc_40319_new_n576_), .B(_abc_40319_new_n525_), .Y(_abc_40319_new_n577_));
OR2X2 OR2X2_30 ( .A(_abc_40319_new_n648_), .B(_abc_40319_new_n562_), .Y(_abc_40319_new_n694_));
OR2X2 OR2X2_300 ( .A(_abc_40319_new_n1508_), .B(_abc_40319_new_n1509_), .Y(_abc_40319_new_n1510_));
OR2X2 OR2X2_301 ( .A(_abc_40319_new_n1186_), .B(REG3_REG_14_), .Y(_abc_40319_new_n1512_));
OR2X2 OR2X2_302 ( .A(_abc_40319_new_n1515_), .B(_abc_40319_new_n1514_), .Y(_abc_40319_new_n1516_));
OR2X2 OR2X2_303 ( .A(_abc_40319_new_n1510_), .B(_abc_40319_new_n1516_), .Y(_abc_40319_new_n1517_));
OR2X2 OR2X2_304 ( .A(_abc_40319_new_n1518_), .B(_abc_40319_new_n1507_), .Y(_abc_40319_new_n1519_));
OR2X2 OR2X2_305 ( .A(_abc_40319_new_n1520_), .B(_abc_40319_new_n1521_), .Y(_abc_40319_new_n1522_));
OR2X2 OR2X2_306 ( .A(_abc_40319_new_n1522_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1523_));
OR2X2 OR2X2_307 ( .A(_abc_40319_new_n1524_), .B(_abc_40319_new_n768_), .Y(_abc_40319_new_n1525_));
OR2X2 OR2X2_308 ( .A(_abc_40319_new_n1526_), .B(_abc_40319_new_n1519_), .Y(_abc_40319_new_n1528_));
OR2X2 OR2X2_309 ( .A(_abc_40319_new_n975_), .B(_abc_40319_new_n972_), .Y(_abc_40319_new_n1531_));
OR2X2 OR2X2_31 ( .A(_abc_40319_new_n695_), .B(_abc_40319_new_n524_), .Y(_abc_40319_new_n696_));
OR2X2 OR2X2_310 ( .A(_abc_40319_new_n1532_), .B(_abc_40319_new_n969_), .Y(_abc_40319_new_n1533_));
OR2X2 OR2X2_311 ( .A(_abc_40319_new_n912_), .B(_abc_40319_new_n768_), .Y(_abc_40319_new_n1538_));
OR2X2 OR2X2_312 ( .A(_abc_40319_new_n911_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1539_));
OR2X2 OR2X2_313 ( .A(_abc_40319_new_n942_), .B(_abc_40319_new_n909_), .Y(_abc_40319_new_n1544_));
OR2X2 OR2X2_314 ( .A(_abc_40319_new_n956_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1549_));
OR2X2 OR2X2_315 ( .A(_abc_40319_new_n960_), .B(_abc_40319_new_n1550_), .Y(_abc_40319_new_n1551_));
OR2X2 OR2X2_316 ( .A(_abc_40319_new_n1552_), .B(_abc_40319_new_n1548_), .Y(_abc_40319_new_n1553_));
OR2X2 OR2X2_317 ( .A(_abc_40319_new_n1554_), .B(_abc_40319_new_n1541_), .Y(_abc_40319_new_n1555_));
OR2X2 OR2X2_318 ( .A(_abc_40319_new_n1556_), .B(_abc_40319_new_n977_), .Y(_abc_40319_new_n1557_));
OR2X2 OR2X2_319 ( .A(_abc_40319_new_n1558_), .B(_abc_40319_new_n1530_), .Y(_abc_40319_new_n1559_));
OR2X2 OR2X2_32 ( .A(_abc_40319_new_n699_), .B(_abc_40319_new_n670_), .Y(_abc_40319_new_n700_));
OR2X2 OR2X2_320 ( .A(_abc_40319_new_n1562_), .B(_abc_40319_new_n1561_), .Y(_abc_40319_new_n1563_));
OR2X2 OR2X2_321 ( .A(_abc_40319_new_n1565_), .B(_abc_40319_new_n1566_), .Y(_abc_40319_new_n1567_));
OR2X2 OR2X2_322 ( .A(_abc_40319_new_n640_), .B(DATAI_8_), .Y(_abc_40319_new_n1571_));
OR2X2 OR2X2_323 ( .A(_abc_40319_new_n1574_), .B(_abc_40319_new_n1573_), .Y(_abc_40319_new_n1575_));
OR2X2 OR2X2_324 ( .A(_abc_40319_new_n1577_), .B(_abc_40319_new_n1578_), .Y(_abc_40319_new_n1579_));
OR2X2 OR2X2_325 ( .A(_abc_40319_new_n1579_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1580_));
OR2X2 OR2X2_326 ( .A(_abc_40319_new_n1581_), .B(_abc_40319_new_n768_), .Y(_abc_40319_new_n1582_));
OR2X2 OR2X2_327 ( .A(_abc_40319_new_n1560_), .B(_abc_40319_new_n1590_), .Y(_abc_40319_new_n1591_));
OR2X2 OR2X2_328 ( .A(_abc_40319_new_n1061_), .B(_abc_40319_new_n1594_), .Y(_abc_40319_new_n1595_));
OR2X2 OR2X2_329 ( .A(_abc_40319_new_n1596_), .B(_abc_40319_new_n1060_), .Y(_abc_40319_new_n1597_));
OR2X2 OR2X2_33 ( .A(_abc_40319_new_n655_), .B(_abc_40319_new_n698_), .Y(_abc_40319_new_n702_));
OR2X2 OR2X2_330 ( .A(_abc_40319_new_n1599_), .B(_abc_40319_new_n1585_), .Y(_abc_40319_new_n1600_));
OR2X2 OR2X2_331 ( .A(_abc_40319_new_n1561_), .B(_abc_40319_new_n545_), .Y(_abc_40319_new_n1606_));
OR2X2 OR2X2_332 ( .A(_abc_40319_new_n1607_), .B(_abc_40319_new_n524_), .Y(_abc_40319_new_n1608_));
OR2X2 OR2X2_333 ( .A(_abc_40319_new_n640_), .B(DATAI_9_), .Y(_abc_40319_new_n1613_));
OR2X2 OR2X2_334 ( .A(_abc_40319_new_n1137_), .B(REG3_REG_9_), .Y(_abc_40319_new_n1617_));
OR2X2 OR2X2_335 ( .A(_abc_40319_new_n1620_), .B(_abc_40319_new_n1619_), .Y(_abc_40319_new_n1621_));
OR2X2 OR2X2_336 ( .A(_abc_40319_new_n1622_), .B(_abc_40319_new_n1623_), .Y(_abc_40319_new_n1624_));
OR2X2 OR2X2_337 ( .A(_abc_40319_new_n1621_), .B(_abc_40319_new_n1624_), .Y(_abc_40319_new_n1625_));
OR2X2 OR2X2_338 ( .A(_abc_40319_new_n1615_), .B(_abc_40319_new_n1626_), .Y(_abc_40319_new_n1627_));
OR2X2 OR2X2_339 ( .A(_abc_40319_new_n1627_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1628_));
OR2X2 OR2X2_34 ( .A(_abc_40319_new_n703_), .B(_abc_40319_new_n598_), .Y(_abc_40319_new_n704_));
OR2X2 OR2X2_340 ( .A(_abc_40319_new_n1629_), .B(_abc_40319_new_n768_), .Y(_abc_40319_new_n1630_));
OR2X2 OR2X2_341 ( .A(_abc_40319_new_n1635_), .B(_abc_40319_new_n1636_), .Y(_abc_40319_new_n1637_));
OR2X2 OR2X2_342 ( .A(_abc_40319_new_n1640_), .B(_abc_40319_new_n1639_), .Y(_abc_40319_new_n1641_));
OR2X2 OR2X2_343 ( .A(_abc_40319_new_n1638_), .B(_abc_40319_new_n1641_), .Y(_abc_40319_new_n1642_));
OR2X2 OR2X2_344 ( .A(_abc_40319_new_n1648_), .B(_abc_40319_new_n553_), .Y(_abc_40319_new_n1649_));
OR2X2 OR2X2_345 ( .A(_abc_40319_new_n1650_), .B(_abc_40319_new_n1644_), .Y(_abc_40319_new_n1651_));
OR2X2 OR2X2_346 ( .A(_abc_40319_new_n640_), .B(DATAI_13_), .Y(_abc_40319_new_n1654_));
OR2X2 OR2X2_347 ( .A(_abc_40319_new_n1658_), .B(REG3_REG_13_), .Y(_abc_40319_new_n1659_));
OR2X2 OR2X2_348 ( .A(_abc_40319_new_n1662_), .B(_abc_40319_new_n1661_), .Y(_abc_40319_new_n1663_));
OR2X2 OR2X2_349 ( .A(_abc_40319_new_n1664_), .B(_abc_40319_new_n1665_), .Y(_abc_40319_new_n1666_));
OR2X2 OR2X2_35 ( .A(_abc_40319_new_n713_), .B(_abc_40319_new_n711_), .Y(_abc_40319_new_n714_));
OR2X2 OR2X2_350 ( .A(_abc_40319_new_n1663_), .B(_abc_40319_new_n1666_), .Y(_abc_40319_new_n1667_));
OR2X2 OR2X2_351 ( .A(_abc_40319_new_n1668_), .B(_abc_40319_new_n1656_), .Y(_abc_40319_new_n1669_));
OR2X2 OR2X2_352 ( .A(_abc_40319_new_n1671_), .B(_abc_40319_new_n1672_), .Y(_abc_40319_new_n1673_));
OR2X2 OR2X2_353 ( .A(_abc_40319_new_n1673_), .B(_abc_40319_new_n768_), .Y(_abc_40319_new_n1674_));
OR2X2 OR2X2_354 ( .A(_abc_40319_new_n1675_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1676_));
OR2X2 OR2X2_355 ( .A(_abc_40319_new_n1683_), .B(_abc_40319_new_n1646_), .Y(_abc_40319_new_n1684_));
OR2X2 OR2X2_356 ( .A(_abc_40319_new_n1685_), .B(_abc_40319_new_n1680_), .Y(_abc_40319_new_n1686_));
OR2X2 OR2X2_357 ( .A(_abc_40319_new_n640_), .B(DATAI_12_), .Y(_abc_40319_new_n1689_));
OR2X2 OR2X2_358 ( .A(_abc_40319_new_n1692_), .B(_abc_40319_new_n1693_), .Y(_abc_40319_new_n1694_));
OR2X2 OR2X2_359 ( .A(_abc_40319_new_n1184_), .B(REG3_REG_12_), .Y(_abc_40319_new_n1697_));
OR2X2 OR2X2_36 ( .A(_abc_40319_new_n715_), .B(_abc_40319_new_n707_), .Y(_abc_40319_new_n716_));
OR2X2 OR2X2_360 ( .A(_abc_40319_new_n1695_), .B(_abc_40319_new_n1699_), .Y(_abc_40319_new_n1700_));
OR2X2 OR2X2_361 ( .A(_abc_40319_new_n1694_), .B(_abc_40319_new_n1700_), .Y(_abc_40319_new_n1701_));
OR2X2 OR2X2_362 ( .A(_abc_40319_new_n1702_), .B(_abc_40319_new_n1691_), .Y(_abc_40319_new_n1703_));
OR2X2 OR2X2_363 ( .A(_abc_40319_new_n1705_), .B(_abc_40319_new_n1706_), .Y(_abc_40319_new_n1707_));
OR2X2 OR2X2_364 ( .A(_abc_40319_new_n1707_), .B(_abc_40319_new_n768_), .Y(_abc_40319_new_n1708_));
OR2X2 OR2X2_365 ( .A(_abc_40319_new_n1709_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1710_));
OR2X2 OR2X2_366 ( .A(_abc_40319_new_n1717_), .B(_abc_40319_new_n1681_), .Y(_abc_40319_new_n1718_));
OR2X2 OR2X2_367 ( .A(_abc_40319_new_n1719_), .B(_abc_40319_new_n1715_), .Y(_abc_40319_new_n1720_));
OR2X2 OR2X2_368 ( .A(_abc_40319_new_n640_), .B(DATAI_11_), .Y(_abc_40319_new_n1723_));
OR2X2 OR2X2_369 ( .A(_abc_40319_new_n1726_), .B(_abc_40319_new_n1727_), .Y(_abc_40319_new_n1728_));
OR2X2 OR2X2_37 ( .A(_abc_40319_new_n633_), .B(_abc_40319_new_n708_), .Y(_abc_40319_new_n717_));
OR2X2 OR2X2_370 ( .A(_abc_40319_new_n1183_), .B(REG3_REG_11_), .Y(_abc_40319_new_n1731_));
OR2X2 OR2X2_371 ( .A(_abc_40319_new_n1729_), .B(_abc_40319_new_n1733_), .Y(_abc_40319_new_n1734_));
OR2X2 OR2X2_372 ( .A(_abc_40319_new_n1728_), .B(_abc_40319_new_n1734_), .Y(_abc_40319_new_n1735_));
OR2X2 OR2X2_373 ( .A(_abc_40319_new_n1736_), .B(_abc_40319_new_n1725_), .Y(_abc_40319_new_n1737_));
OR2X2 OR2X2_374 ( .A(_abc_40319_new_n1739_), .B(_abc_40319_new_n1740_), .Y(_abc_40319_new_n1741_));
OR2X2 OR2X2_375 ( .A(_abc_40319_new_n1741_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1742_));
OR2X2 OR2X2_376 ( .A(_abc_40319_new_n1743_), .B(_abc_40319_new_n768_), .Y(_abc_40319_new_n1744_));
OR2X2 OR2X2_377 ( .A(_abc_40319_new_n1751_), .B(_abc_40319_new_n1645_), .Y(_abc_40319_new_n1752_));
OR2X2 OR2X2_378 ( .A(_abc_40319_new_n1753_), .B(_abc_40319_new_n1750_), .Y(_abc_40319_new_n1754_));
OR2X2 OR2X2_379 ( .A(_abc_40319_new_n640_), .B(DATAI_10_), .Y(_abc_40319_new_n1757_));
OR2X2 OR2X2_38 ( .A(_abc_40319_new_n719_), .B(_abc_40319_new_n720_), .Y(_abc_40319_new_n721_));
OR2X2 OR2X2_380 ( .A(_abc_40319_new_n1760_), .B(_abc_40319_new_n1761_), .Y(_abc_40319_new_n1762_));
OR2X2 OR2X2_381 ( .A(_abc_40319_new_n1182_), .B(REG3_REG_10_), .Y(_abc_40319_new_n1765_));
OR2X2 OR2X2_382 ( .A(_abc_40319_new_n1763_), .B(_abc_40319_new_n1767_), .Y(_abc_40319_new_n1768_));
OR2X2 OR2X2_383 ( .A(_abc_40319_new_n1762_), .B(_abc_40319_new_n1768_), .Y(_abc_40319_new_n1769_));
OR2X2 OR2X2_384 ( .A(_abc_40319_new_n1770_), .B(_abc_40319_new_n1759_), .Y(_abc_40319_new_n1771_));
OR2X2 OR2X2_385 ( .A(_abc_40319_new_n1773_), .B(_abc_40319_new_n1774_), .Y(_abc_40319_new_n1775_));
OR2X2 OR2X2_386 ( .A(_abc_40319_new_n1775_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n1776_));
OR2X2 OR2X2_387 ( .A(_abc_40319_new_n1777_), .B(_abc_40319_new_n768_), .Y(_abc_40319_new_n1778_));
OR2X2 OR2X2_388 ( .A(_abc_40319_new_n1711_), .B(_abc_40319_new_n1704_), .Y(_abc_40319_new_n1791_));
OR2X2 OR2X2_389 ( .A(_abc_40319_new_n1677_), .B(_abc_40319_new_n1670_), .Y(_abc_40319_new_n1792_));
OR2X2 OR2X2_39 ( .A(_abc_40319_new_n710_), .B(_abc_40319_new_n706_), .Y(_abc_40319_new_n726_));
OR2X2 OR2X2_390 ( .A(_abc_40319_new_n1794_), .B(_abc_40319_new_n1678_), .Y(_abc_40319_new_n1795_));
OR2X2 OR2X2_391 ( .A(_abc_40319_new_n1784_), .B(_abc_40319_new_n1797_), .Y(_abc_40319_new_n1798_));
OR2X2 OR2X2_392 ( .A(_abc_40319_new_n1799_), .B(_abc_40319_new_n1527_), .Y(_abc_40319_new_n1800_));
OR2X2 OR2X2_393 ( .A(_abc_40319_new_n1801_), .B(_abc_40319_new_n1493_), .Y(_abc_40319_new_n1802_));
OR2X2 OR2X2_394 ( .A(_abc_40319_new_n1808_), .B(_abc_40319_new_n1456_), .Y(_abc_40319_new_n1809_));
OR2X2 OR2X2_395 ( .A(_abc_40319_new_n1803_), .B(_abc_40319_new_n1810_), .Y(_abc_40319_new_n1811_));
OR2X2 OR2X2_396 ( .A(_abc_40319_new_n1812_), .B(_abc_40319_new_n1385_), .Y(_abc_40319_new_n1813_));
OR2X2 OR2X2_397 ( .A(_abc_40319_new_n640_), .B(DATAI_19_), .Y(_abc_40319_new_n1816_));
OR2X2 OR2X2_398 ( .A(_abc_40319_new_n1191_), .B(REG3_REG_19_), .Y(_abc_40319_new_n1821_));
OR2X2 OR2X2_399 ( .A(_abc_40319_new_n1825_), .B(_abc_40319_new_n1824_), .Y(_abc_40319_new_n1826_));
OR2X2 OR2X2_4 ( .A(_abc_40319_new_n580_), .B(_abc_40319_new_n524_), .Y(_abc_40319_new_n581_));
OR2X2 OR2X2_40 ( .A(_abc_40319_new_n727_), .B(_abc_40319_new_n524_), .Y(_abc_40319_new_n728_));
OR2X2 OR2X2_400 ( .A(_abc_40319_new_n1826_), .B(_abc_40319_new_n1823_), .Y(_abc_40319_new_n1827_));
OR2X2 OR2X2_401 ( .A(_abc_40319_new_n1827_), .B(_abc_40319_new_n1819_), .Y(_abc_40319_new_n1828_));
OR2X2 OR2X2_402 ( .A(_abc_40319_new_n1829_), .B(_abc_40319_new_n1818_), .Y(_abc_40319_new_n1830_));
OR2X2 OR2X2_403 ( .A(_abc_40319_new_n1833_), .B(_abc_40319_new_n1832_), .Y(_abc_40319_new_n1834_));
OR2X2 OR2X2_404 ( .A(_abc_40319_new_n1836_), .B(_abc_40319_new_n1837_), .Y(_abc_40319_new_n1838_));
OR2X2 OR2X2_405 ( .A(_abc_40319_new_n1192_), .B(REG3_REG_20_), .Y(_abc_40319_new_n1845_));
OR2X2 OR2X2_406 ( .A(_abc_40319_new_n1849_), .B(_abc_40319_new_n1848_), .Y(_abc_40319_new_n1850_));
OR2X2 OR2X2_407 ( .A(_abc_40319_new_n1850_), .B(_abc_40319_new_n1847_), .Y(_abc_40319_new_n1851_));
OR2X2 OR2X2_408 ( .A(_abc_40319_new_n1851_), .B(_abc_40319_new_n1843_), .Y(_abc_40319_new_n1852_));
OR2X2 OR2X2_409 ( .A(_abc_40319_new_n1853_), .B(_abc_40319_new_n1842_), .Y(_abc_40319_new_n1854_));
OR2X2 OR2X2_41 ( .A(_abc_40319_new_n723_), .B(_abc_40319_new_n734_), .Y(_abc_40319_new_n735_));
OR2X2 OR2X2_410 ( .A(_abc_40319_new_n1857_), .B(_abc_40319_new_n1856_), .Y(_abc_40319_new_n1858_));
OR2X2 OR2X2_411 ( .A(_abc_40319_new_n1860_), .B(_abc_40319_new_n1861_), .Y(_abc_40319_new_n1862_));
OR2X2 OR2X2_412 ( .A(_abc_40319_new_n1193_), .B(REG3_REG_21_), .Y(_abc_40319_new_n1868_));
OR2X2 OR2X2_413 ( .A(_abc_40319_new_n1872_), .B(_abc_40319_new_n1873_), .Y(_abc_40319_new_n1874_));
OR2X2 OR2X2_414 ( .A(_abc_40319_new_n1874_), .B(_abc_40319_new_n1871_), .Y(_abc_40319_new_n1875_));
OR2X2 OR2X2_415 ( .A(_abc_40319_new_n1875_), .B(_abc_40319_new_n1870_), .Y(_abc_40319_new_n1876_));
OR2X2 OR2X2_416 ( .A(_abc_40319_new_n1877_), .B(_abc_40319_new_n1866_), .Y(_abc_40319_new_n1878_));
OR2X2 OR2X2_417 ( .A(_abc_40319_new_n1881_), .B(_abc_40319_new_n1880_), .Y(_abc_40319_new_n1882_));
OR2X2 OR2X2_418 ( .A(_abc_40319_new_n1884_), .B(_abc_40319_new_n1885_), .Y(_abc_40319_new_n1886_));
OR2X2 OR2X2_419 ( .A(_abc_40319_new_n1838_), .B(_abc_40319_new_n1831_), .Y(_abc_40319_new_n1893_));
OR2X2 OR2X2_42 ( .A(_abc_40319_new_n739_), .B(REG3_REG_5_), .Y(_abc_40319_new_n742_));
OR2X2 OR2X2_420 ( .A(_abc_40319_new_n1862_), .B(_abc_40319_new_n1855_), .Y(_abc_40319_new_n1899_));
OR2X2 OR2X2_421 ( .A(_abc_40319_new_n1901_), .B(_abc_40319_new_n1888_), .Y(_abc_40319_new_n1902_));
OR2X2 OR2X2_422 ( .A(_abc_40319_new_n1892_), .B(_abc_40319_new_n1903_), .Y(_abc_40319_new_n1904_));
OR2X2 OR2X2_423 ( .A(_abc_40319_new_n1905_), .B(_abc_40319_new_n1351_), .Y(_abc_40319_new_n1906_));
OR2X2 OR2X2_424 ( .A(_abc_40319_new_n1907_), .B(_abc_40319_new_n1327_), .Y(_abc_40319_new_n1908_));
OR2X2 OR2X2_425 ( .A(_abc_40319_new_n1295_), .B(_abc_40319_new_n1287_), .Y(_abc_40319_new_n1909_));
OR2X2 OR2X2_426 ( .A(_abc_40319_new_n1911_), .B(_abc_40319_new_n1305_), .Y(_abc_40319_new_n1912_));
OR2X2 OR2X2_427 ( .A(_abc_40319_new_n1912_), .B(_abc_40319_new_n1223_), .Y(_abc_40319_new_n1913_));
OR2X2 OR2X2_428 ( .A(_abc_40319_new_n1633_), .B(_abc_40319_new_n1927_), .Y(_abc_40319_new_n1928_));
OR2X2 OR2X2_429 ( .A(_abc_40319_new_n1929_), .B(_abc_40319_new_n1930_), .Y(_abc_40319_new_n1931_));
OR2X2 OR2X2_43 ( .A(_abc_40319_new_n737_), .B(_abc_40319_new_n744_), .Y(_abc_40319_new_n745_));
OR2X2 OR2X2_430 ( .A(_abc_40319_new_n1932_), .B(_abc_40319_new_n1925_), .Y(_abc_40319_new_n1933_));
OR2X2 OR2X2_431 ( .A(_abc_40319_new_n1934_), .B(_abc_40319_new_n1923_), .Y(_abc_40319_new_n1935_));
OR2X2 OR2X2_432 ( .A(_abc_40319_new_n1936_), .B(_abc_40319_new_n1921_), .Y(_abc_40319_new_n1937_));
OR2X2 OR2X2_433 ( .A(_abc_40319_new_n1938_), .B(_abc_40319_new_n1920_), .Y(_abc_40319_new_n1939_));
OR2X2 OR2X2_434 ( .A(_abc_40319_new_n1940_), .B(_abc_40319_new_n1941_), .Y(_abc_40319_new_n1942_));
OR2X2 OR2X2_435 ( .A(_abc_40319_new_n1943_), .B(_abc_40319_new_n1918_), .Y(_abc_40319_new_n1944_));
OR2X2 OR2X2_436 ( .A(_abc_40319_new_n1945_), .B(_abc_40319_new_n1916_), .Y(_abc_40319_new_n1946_));
OR2X2 OR2X2_437 ( .A(_abc_40319_new_n1947_), .B(_abc_40319_new_n1948_), .Y(_abc_40319_new_n1949_));
OR2X2 OR2X2_438 ( .A(_abc_40319_new_n1950_), .B(_abc_40319_new_n1914_), .Y(_abc_40319_new_n1951_));
OR2X2 OR2X2_439 ( .A(_abc_40319_new_n1969_), .B(REG3_REG_28_), .Y(_abc_40319_new_n1972_));
OR2X2 OR2X2_44 ( .A(_abc_40319_new_n735_), .B(_abc_40319_new_n745_), .Y(_abc_40319_new_n746_));
OR2X2 OR2X2_440 ( .A(_abc_40319_new_n1976_), .B(_abc_40319_new_n1977_), .Y(_abc_40319_new_n1978_));
OR2X2 OR2X2_441 ( .A(_abc_40319_new_n1978_), .B(_abc_40319_new_n1975_), .Y(_abc_40319_new_n1979_));
OR2X2 OR2X2_442 ( .A(_abc_40319_new_n1974_), .B(_abc_40319_new_n1979_), .Y(_abc_40319_new_n1980_));
OR2X2 OR2X2_443 ( .A(_abc_40319_new_n1981_), .B(_abc_40319_new_n1954_), .Y(_abc_40319_new_n1982_));
OR2X2 OR2X2_444 ( .A(_abc_40319_new_n1986_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n1987_));
OR2X2 OR2X2_445 ( .A(_abc_40319_new_n1985_), .B(_abc_40319_new_n1987_), .Y(_abc_40319_new_n1988_));
OR2X2 OR2X2_446 ( .A(_abc_40319_new_n1984_), .B(_abc_40319_new_n1988_), .Y(_abc_40319_new_n1989_));
OR2X2 OR2X2_447 ( .A(_abc_40319_new_n1983_), .B(_abc_40319_new_n1989_), .Y(_abc_40319_new_n1990_));
OR2X2 OR2X2_448 ( .A(_abc_40319_new_n1953_), .B(_abc_40319_new_n1990_), .Y(n1326));
OR2X2 OR2X2_449 ( .A(_abc_40319_new_n1932_), .B(_abc_40319_new_n1993_), .Y(_abc_40319_new_n1994_));
OR2X2 OR2X2_45 ( .A(_abc_40319_new_n747_), .B(_abc_40319_new_n690_), .Y(_abc_40319_new_n748_));
OR2X2 OR2X2_450 ( .A(_abc_40319_new_n1798_), .B(_abc_40319_new_n1992_), .Y(_abc_40319_new_n1995_));
OR2X2 OR2X2_451 ( .A(_abc_40319_new_n1998_), .B(_abc_40319_new_n1999_), .Y(_abc_40319_new_n2000_));
OR2X2 OR2X2_452 ( .A(_abc_40319_new_n2004_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n2005_));
OR2X2 OR2X2_453 ( .A(_abc_40319_new_n2003_), .B(_abc_40319_new_n2005_), .Y(_abc_40319_new_n2006_));
OR2X2 OR2X2_454 ( .A(_abc_40319_new_n2002_), .B(_abc_40319_new_n2006_), .Y(_abc_40319_new_n2007_));
OR2X2 OR2X2_455 ( .A(_abc_40319_new_n2007_), .B(_abc_40319_new_n2001_), .Y(_abc_40319_new_n2008_));
OR2X2 OR2X2_456 ( .A(_abc_40319_new_n1997_), .B(_abc_40319_new_n2008_), .Y(n1321));
OR2X2 OR2X2_457 ( .A(_abc_40319_new_n1945_), .B(_abc_40319_new_n2011_), .Y(_abc_40319_new_n2012_));
OR2X2 OR2X2_458 ( .A(_abc_40319_new_n1906_), .B(_abc_40319_new_n2010_), .Y(_abc_40319_new_n2013_));
OR2X2 OR2X2_459 ( .A(_abc_40319_new_n2017_), .B(_abc_40319_new_n2016_), .Y(_abc_40319_new_n2018_));
OR2X2 OR2X2_46 ( .A(_abc_40319_new_n753_), .B(_abc_40319_new_n754_), .Y(_abc_40319_new_n755_));
OR2X2 OR2X2_460 ( .A(_abc_40319_new_n2022_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n2023_));
OR2X2 OR2X2_461 ( .A(_abc_40319_new_n2021_), .B(_abc_40319_new_n2023_), .Y(_abc_40319_new_n2024_));
OR2X2 OR2X2_462 ( .A(_abc_40319_new_n2020_), .B(_abc_40319_new_n2024_), .Y(_abc_40319_new_n2025_));
OR2X2 OR2X2_463 ( .A(_abc_40319_new_n2025_), .B(_abc_40319_new_n2019_), .Y(_abc_40319_new_n2026_));
OR2X2 OR2X2_464 ( .A(_abc_40319_new_n2015_), .B(_abc_40319_new_n2026_), .Y(n1316));
OR2X2 OR2X2_465 ( .A(_abc_40319_new_n1929_), .B(_abc_40319_new_n2030_), .Y(_abc_40319_new_n2031_));
OR2X2 OR2X2_466 ( .A(_abc_40319_new_n1643_), .B(_abc_40319_new_n2029_), .Y(_abc_40319_new_n2032_));
OR2X2 OR2X2_467 ( .A(_abc_40319_new_n2035_), .B(_abc_40319_new_n2036_), .Y(_abc_40319_new_n2037_));
OR2X2 OR2X2_468 ( .A(_abc_40319_new_n2041_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n2042_));
OR2X2 OR2X2_469 ( .A(_abc_40319_new_n2040_), .B(_abc_40319_new_n2042_), .Y(_abc_40319_new_n2043_));
OR2X2 OR2X2_47 ( .A(_abc_40319_new_n755_), .B(_abc_40319_new_n752_), .Y(_abc_40319_new_n756_));
OR2X2 OR2X2_470 ( .A(_abc_40319_new_n2039_), .B(_abc_40319_new_n2043_), .Y(_abc_40319_new_n2044_));
OR2X2 OR2X2_471 ( .A(_abc_40319_new_n2044_), .B(_abc_40319_new_n2038_), .Y(_abc_40319_new_n2045_));
OR2X2 OR2X2_472 ( .A(_abc_40319_new_n2034_), .B(_abc_40319_new_n2045_), .Y(n1311));
OR2X2 OR2X2_473 ( .A(_abc_40319_new_n971_), .B(_abc_40319_new_n2047_), .Y(_abc_40319_new_n2048_));
OR2X2 OR2X2_474 ( .A(_abc_40319_new_n2050_), .B(_abc_40319_new_n877_), .Y(_abc_40319_new_n2051_));
OR2X2 OR2X2_475 ( .A(_abc_40319_new_n2052_), .B(_abc_40319_new_n2048_), .Y(_abc_40319_new_n2053_));
OR2X2 OR2X2_476 ( .A(_abc_40319_new_n2051_), .B(_abc_40319_new_n2054_), .Y(_abc_40319_new_n2055_));
OR2X2 OR2X2_477 ( .A(_abc_40319_new_n2058_), .B(_abc_40319_new_n2059_), .Y(_abc_40319_new_n2060_));
OR2X2 OR2X2_478 ( .A(_abc_40319_new_n2063_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n2064_));
OR2X2 OR2X2_479 ( .A(_abc_40319_new_n2062_), .B(_abc_40319_new_n2064_), .Y(_abc_40319_new_n2065_));
OR2X2 OR2X2_48 ( .A(_abc_40319_new_n655_), .B(_abc_40319_new_n646_), .Y(_abc_40319_new_n759_));
OR2X2 OR2X2_480 ( .A(_abc_40319_new_n2066_), .B(_abc_40319_new_n2065_), .Y(_abc_40319_new_n2067_));
OR2X2 OR2X2_481 ( .A(_abc_40319_new_n2067_), .B(_abc_40319_new_n2061_), .Y(_abc_40319_new_n2068_));
OR2X2 OR2X2_482 ( .A(_abc_40319_new_n2057_), .B(_abc_40319_new_n2068_), .Y(n1306));
OR2X2 OR2X2_483 ( .A(_abc_40319_new_n1940_), .B(_abc_40319_new_n2071_), .Y(_abc_40319_new_n2072_));
OR2X2 OR2X2_484 ( .A(_abc_40319_new_n1813_), .B(_abc_40319_new_n2070_), .Y(_abc_40319_new_n2073_));
OR2X2 OR2X2_485 ( .A(_abc_40319_new_n2076_), .B(_abc_40319_new_n2077_), .Y(_abc_40319_new_n2078_));
OR2X2 OR2X2_486 ( .A(_abc_40319_new_n2082_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n2083_));
OR2X2 OR2X2_487 ( .A(_abc_40319_new_n2081_), .B(_abc_40319_new_n2083_), .Y(_abc_40319_new_n2084_));
OR2X2 OR2X2_488 ( .A(_abc_40319_new_n2080_), .B(_abc_40319_new_n2084_), .Y(_abc_40319_new_n2085_));
OR2X2 OR2X2_489 ( .A(_abc_40319_new_n2085_), .B(_abc_40319_new_n2079_), .Y(_abc_40319_new_n2086_));
OR2X2 OR2X2_49 ( .A(_abc_40319_new_n762_), .B(_abc_40319_new_n758_), .Y(_abc_40319_new_n763_));
OR2X2 OR2X2_490 ( .A(_abc_40319_new_n2075_), .B(_abc_40319_new_n2086_), .Y(n1301));
OR2X2 OR2X2_491 ( .A(_abc_40319_new_n1912_), .B(_abc_40319_new_n1220_), .Y(_abc_40319_new_n2088_));
OR2X2 OR2X2_492 ( .A(_abc_40319_new_n2091_), .B(_abc_40319_new_n2090_), .Y(_abc_40319_new_n2092_));
OR2X2 OR2X2_493 ( .A(_abc_40319_new_n2094_), .B(_abc_40319_new_n2093_), .Y(_abc_40319_new_n2095_));
OR2X2 OR2X2_494 ( .A(_abc_40319_new_n2097_), .B(_abc_40319_new_n2098_), .Y(_abc_40319_new_n2099_));
OR2X2 OR2X2_495 ( .A(_abc_40319_new_n2099_), .B(_abc_40319_new_n2092_), .Y(_abc_40319_new_n2100_));
OR2X2 OR2X2_496 ( .A(_abc_40319_new_n2102_), .B(_abc_40319_new_n2101_), .Y(_abc_40319_new_n2103_));
OR2X2 OR2X2_497 ( .A(_abc_40319_new_n1950_), .B(_abc_40319_new_n2108_), .Y(_abc_40319_new_n2109_));
OR2X2 OR2X2_498 ( .A(_abc_40319_new_n2107_), .B(_abc_40319_new_n2111_), .Y(_abc_40319_new_n2112_));
OR2X2 OR2X2_499 ( .A(_abc_40319_new_n2120_), .B(_abc_40319_new_n2117_), .Y(_abc_40319_new_n2121_));
OR2X2 OR2X2_5 ( .A(_abc_40319_new_n584_), .B(_abc_40319_new_n574_), .Y(_abc_40319_new_n585_));
OR2X2 OR2X2_50 ( .A(_abc_40319_new_n764_), .B(_abc_40319_new_n765_), .Y(_abc_40319_new_n766_));
OR2X2 OR2X2_500 ( .A(_abc_40319_new_n2121_), .B(_abc_40319_new_n2116_), .Y(_abc_40319_new_n2122_));
OR2X2 OR2X2_501 ( .A(_abc_40319_new_n2122_), .B(_abc_40319_new_n2115_), .Y(_abc_40319_new_n2123_));
OR2X2 OR2X2_502 ( .A(_abc_40319_new_n2124_), .B(_abc_40319_new_n2114_), .Y(_abc_40319_new_n2125_));
OR2X2 OR2X2_503 ( .A(_abc_40319_new_n2129_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n2130_));
OR2X2 OR2X2_504 ( .A(_abc_40319_new_n2128_), .B(_abc_40319_new_n2130_), .Y(_abc_40319_new_n2131_));
OR2X2 OR2X2_505 ( .A(_abc_40319_new_n2127_), .B(_abc_40319_new_n2131_), .Y(_abc_40319_new_n2132_));
OR2X2 OR2X2_506 ( .A(_abc_40319_new_n2132_), .B(_abc_40319_new_n2126_), .Y(_abc_40319_new_n2133_));
OR2X2 OR2X2_507 ( .A(_abc_40319_new_n2113_), .B(_abc_40319_new_n2133_), .Y(n1296));
OR2X2 OR2X2_508 ( .A(_abc_40319_new_n2139_), .B(_abc_40319_new_n2135_), .Y(_abc_40319_new_n2140_));
OR2X2 OR2X2_509 ( .A(_abc_40319_new_n2138_), .B(_abc_40319_new_n2141_), .Y(_abc_40319_new_n2142_));
OR2X2 OR2X2_51 ( .A(_abc_40319_new_n766_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n767_));
OR2X2 OR2X2_510 ( .A(_abc_40319_new_n2145_), .B(_abc_40319_new_n2146_), .Y(_abc_40319_new_n2147_));
OR2X2 OR2X2_511 ( .A(_abc_40319_new_n2151_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n2152_));
OR2X2 OR2X2_512 ( .A(_abc_40319_new_n2150_), .B(_abc_40319_new_n2152_), .Y(_abc_40319_new_n2153_));
OR2X2 OR2X2_513 ( .A(_abc_40319_new_n2149_), .B(_abc_40319_new_n2153_), .Y(_abc_40319_new_n2154_));
OR2X2 OR2X2_514 ( .A(_abc_40319_new_n2154_), .B(_abc_40319_new_n2148_), .Y(_abc_40319_new_n2155_));
OR2X2 OR2X2_515 ( .A(_abc_40319_new_n2144_), .B(_abc_40319_new_n2155_), .Y(n1291));
OR2X2 OR2X2_516 ( .A(_abc_40319_new_n1555_), .B(_abc_40319_new_n917_), .Y(_abc_40319_new_n2157_));
OR2X2 OR2X2_517 ( .A(_abc_40319_new_n2158_), .B(_abc_40319_new_n966_), .Y(_abc_40319_new_n2159_));
OR2X2 OR2X2_518 ( .A(_abc_40319_new_n2162_), .B(_abc_40319_new_n2163_), .Y(_abc_40319_new_n2164_));
OR2X2 OR2X2_519 ( .A(_abc_40319_new_n2167_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n2168_));
OR2X2 OR2X2_52 ( .A(_abc_40319_new_n769_), .B(_abc_40319_new_n768_), .Y(_abc_40319_new_n770_));
OR2X2 OR2X2_520 ( .A(_abc_40319_new_n2166_), .B(_abc_40319_new_n2168_), .Y(_abc_40319_new_n2169_));
OR2X2 OR2X2_521 ( .A(_abc_40319_new_n2170_), .B(_abc_40319_new_n2169_), .Y(_abc_40319_new_n2171_));
OR2X2 OR2X2_522 ( .A(_abc_40319_new_n2171_), .B(_abc_40319_new_n2165_), .Y(_abc_40319_new_n2172_));
OR2X2 OR2X2_523 ( .A(_abc_40319_new_n2161_), .B(_abc_40319_new_n2172_), .Y(n1286));
OR2X2 OR2X2_524 ( .A(_abc_40319_new_n2174_), .B(_abc_40319_new_n1894_), .Y(_abc_40319_new_n2175_));
OR2X2 OR2X2_525 ( .A(_abc_40319_new_n2178_), .B(_abc_40319_new_n1897_), .Y(_abc_40319_new_n2179_));
OR2X2 OR2X2_526 ( .A(_abc_40319_new_n2177_), .B(_abc_40319_new_n2179_), .Y(_abc_40319_new_n2180_));
OR2X2 OR2X2_527 ( .A(_abc_40319_new_n2183_), .B(_abc_40319_new_n2182_), .Y(_abc_40319_new_n2184_));
OR2X2 OR2X2_528 ( .A(_abc_40319_new_n2181_), .B(_abc_40319_new_n2184_), .Y(_abc_40319_new_n2185_));
OR2X2 OR2X2_529 ( .A(_abc_40319_new_n2189_), .B(_abc_40319_new_n2190_), .Y(_abc_40319_new_n2191_));
OR2X2 OR2X2_53 ( .A(_abc_40319_new_n771_), .B(_abc_40319_new_n748_), .Y(_abc_40319_new_n773_));
OR2X2 OR2X2_530 ( .A(_abc_40319_new_n2191_), .B(_abc_40319_new_n2188_), .Y(_abc_40319_new_n2192_));
OR2X2 OR2X2_531 ( .A(_abc_40319_new_n2196_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n2197_));
OR2X2 OR2X2_532 ( .A(_abc_40319_new_n2195_), .B(_abc_40319_new_n2197_), .Y(_abc_40319_new_n2198_));
OR2X2 OR2X2_533 ( .A(_abc_40319_new_n2198_), .B(_abc_40319_new_n2194_), .Y(_abc_40319_new_n2199_));
OR2X2 OR2X2_534 ( .A(_abc_40319_new_n2199_), .B(_abc_40319_new_n2193_), .Y(_abc_40319_new_n2200_));
OR2X2 OR2X2_535 ( .A(_abc_40319_new_n2187_), .B(_abc_40319_new_n2200_), .Y(n1281));
OR2X2 OR2X2_536 ( .A(_abc_40319_new_n2203_), .B(_abc_40319_new_n1785_), .Y(_abc_40319_new_n2204_));
OR2X2 OR2X2_537 ( .A(_abc_40319_new_n2205_), .B(_abc_40319_new_n1788_), .Y(_abc_40319_new_n2206_));
OR2X2 OR2X2_538 ( .A(_abc_40319_new_n2206_), .B(_abc_40319_new_n2202_), .Y(_abc_40319_new_n2207_));
OR2X2 OR2X2_539 ( .A(_abc_40319_new_n2209_), .B(_abc_40319_new_n2208_), .Y(_abc_40319_new_n2210_));
OR2X2 OR2X2_54 ( .A(_abc_40319_new_n677_), .B(_abc_40319_new_n774_), .Y(_abc_40319_new_n775_));
OR2X2 OR2X2_540 ( .A(_abc_40319_new_n2213_), .B(_abc_40319_new_n2214_), .Y(_abc_40319_new_n2215_));
OR2X2 OR2X2_541 ( .A(_abc_40319_new_n2219_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n2220_));
OR2X2 OR2X2_542 ( .A(_abc_40319_new_n2218_), .B(_abc_40319_new_n2220_), .Y(_abc_40319_new_n2221_));
OR2X2 OR2X2_543 ( .A(_abc_40319_new_n2217_), .B(_abc_40319_new_n2221_), .Y(_abc_40319_new_n2222_));
OR2X2 OR2X2_544 ( .A(_abc_40319_new_n2222_), .B(_abc_40319_new_n2216_), .Y(_abc_40319_new_n2223_));
OR2X2 OR2X2_545 ( .A(_abc_40319_new_n2212_), .B(_abc_40319_new_n2223_), .Y(n1276));
OR2X2 OR2X2_546 ( .A(_abc_40319_new_n2226_), .B(_abc_40319_new_n1296_), .Y(_abc_40319_new_n2227_));
OR2X2 OR2X2_547 ( .A(_abc_40319_new_n2227_), .B(_abc_40319_new_n2225_), .Y(_abc_40319_new_n2228_));
OR2X2 OR2X2_548 ( .A(_abc_40319_new_n2230_), .B(_abc_40319_new_n2229_), .Y(_abc_40319_new_n2231_));
OR2X2 OR2X2_549 ( .A(_abc_40319_new_n2235_), .B(_abc_40319_new_n2234_), .Y(_abc_40319_new_n2236_));
OR2X2 OR2X2_55 ( .A(_abc_40319_new_n777_), .B(_abc_40319_new_n778_), .Y(_abc_40319_new_n779_));
OR2X2 OR2X2_550 ( .A(_abc_40319_new_n2240_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n2241_));
OR2X2 OR2X2_551 ( .A(_abc_40319_new_n2239_), .B(_abc_40319_new_n2241_), .Y(_abc_40319_new_n2242_));
OR2X2 OR2X2_552 ( .A(_abc_40319_new_n2238_), .B(_abc_40319_new_n2242_), .Y(_abc_40319_new_n2243_));
OR2X2 OR2X2_553 ( .A(_abc_40319_new_n2237_), .B(_abc_40319_new_n2243_), .Y(_abc_40319_new_n2244_));
OR2X2 OR2X2_554 ( .A(_abc_40319_new_n2233_), .B(_abc_40319_new_n2244_), .Y(n1271));
OR2X2 OR2X2_555 ( .A(_abc_40319_new_n1936_), .B(_abc_40319_new_n2247_), .Y(_abc_40319_new_n2248_));
OR2X2 OR2X2_556 ( .A(_abc_40319_new_n1802_), .B(_abc_40319_new_n2246_), .Y(_abc_40319_new_n2249_));
OR2X2 OR2X2_557 ( .A(_abc_40319_new_n2252_), .B(_abc_40319_new_n2253_), .Y(_abc_40319_new_n2254_));
OR2X2 OR2X2_558 ( .A(_abc_40319_new_n2257_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n2258_));
OR2X2 OR2X2_559 ( .A(_abc_40319_new_n2256_), .B(_abc_40319_new_n2258_), .Y(_abc_40319_new_n2259_));
OR2X2 OR2X2_56 ( .A(_abc_40319_new_n640_), .B(DATAI_4_), .Y(_abc_40319_new_n783_));
OR2X2 OR2X2_560 ( .A(_abc_40319_new_n2260_), .B(_abc_40319_new_n2259_), .Y(_abc_40319_new_n2261_));
OR2X2 OR2X2_561 ( .A(_abc_40319_new_n2261_), .B(_abc_40319_new_n2255_), .Y(_abc_40319_new_n2262_));
OR2X2 OR2X2_562 ( .A(_abc_40319_new_n2251_), .B(_abc_40319_new_n2262_), .Y(n1266));
OR2X2 OR2X2_563 ( .A(_abc_40319_new_n1560_), .B(_abc_40319_new_n2265_), .Y(_abc_40319_new_n2266_));
OR2X2 OR2X2_564 ( .A(_abc_40319_new_n982_), .B(_abc_40319_new_n2264_), .Y(_abc_40319_new_n2267_));
OR2X2 OR2X2_565 ( .A(_abc_40319_new_n2270_), .B(_abc_40319_new_n2271_), .Y(_abc_40319_new_n2272_));
OR2X2 OR2X2_566 ( .A(_abc_40319_new_n2275_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n2276_));
OR2X2 OR2X2_567 ( .A(_abc_40319_new_n2274_), .B(_abc_40319_new_n2276_), .Y(_abc_40319_new_n2277_));
OR2X2 OR2X2_568 ( .A(_abc_40319_new_n2278_), .B(_abc_40319_new_n2277_), .Y(_abc_40319_new_n2279_));
OR2X2 OR2X2_569 ( .A(_abc_40319_new_n2279_), .B(_abc_40319_new_n2273_), .Y(_abc_40319_new_n2280_));
OR2X2 OR2X2_57 ( .A(_abc_40319_new_n786_), .B(_abc_40319_new_n787_), .Y(_abc_40319_new_n788_));
OR2X2 OR2X2_570 ( .A(_abc_40319_new_n2269_), .B(_abc_40319_new_n2280_), .Y(n1261));
OR2X2 OR2X2_571 ( .A(_abc_40319_new_n2283_), .B(_abc_40319_new_n1804_), .Y(_abc_40319_new_n2284_));
OR2X2 OR2X2_572 ( .A(_abc_40319_new_n2282_), .B(_abc_40319_new_n2284_), .Y(_abc_40319_new_n2285_));
OR2X2 OR2X2_573 ( .A(_abc_40319_new_n1921_), .B(_abc_40319_new_n1806_), .Y(_abc_40319_new_n2287_));
OR2X2 OR2X2_574 ( .A(_abc_40319_new_n2286_), .B(_abc_40319_new_n2287_), .Y(_abc_40319_new_n2288_));
OR2X2 OR2X2_575 ( .A(_abc_40319_new_n2291_), .B(_abc_40319_new_n2292_), .Y(_abc_40319_new_n2293_));
OR2X2 OR2X2_576 ( .A(_abc_40319_new_n2296_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n2297_));
OR2X2 OR2X2_577 ( .A(_abc_40319_new_n2295_), .B(_abc_40319_new_n2297_), .Y(_abc_40319_new_n2298_));
OR2X2 OR2X2_578 ( .A(_abc_40319_new_n2299_), .B(_abc_40319_new_n2298_), .Y(_abc_40319_new_n2300_));
OR2X2 OR2X2_579 ( .A(_abc_40319_new_n2300_), .B(_abc_40319_new_n2294_), .Y(_abc_40319_new_n2301_));
OR2X2 OR2X2_58 ( .A(REG3_REG_3_), .B(REG3_REG_4_), .Y(_abc_40319_new_n791_));
OR2X2 OR2X2_580 ( .A(_abc_40319_new_n2290_), .B(_abc_40319_new_n2301_), .Y(n1256));
OR2X2 OR2X2_581 ( .A(_abc_40319_new_n1947_), .B(_abc_40319_new_n2305_), .Y(_abc_40319_new_n2306_));
OR2X2 OR2X2_582 ( .A(_abc_40319_new_n1908_), .B(_abc_40319_new_n2304_), .Y(_abc_40319_new_n2307_));
OR2X2 OR2X2_583 ( .A(_abc_40319_new_n2311_), .B(_abc_40319_new_n2310_), .Y(_abc_40319_new_n2312_));
OR2X2 OR2X2_584 ( .A(_abc_40319_new_n2316_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n2317_));
OR2X2 OR2X2_585 ( .A(_abc_40319_new_n2315_), .B(_abc_40319_new_n2317_), .Y(_abc_40319_new_n2318_));
OR2X2 OR2X2_586 ( .A(_abc_40319_new_n2314_), .B(_abc_40319_new_n2318_), .Y(_abc_40319_new_n2319_));
OR2X2 OR2X2_587 ( .A(_abc_40319_new_n2313_), .B(_abc_40319_new_n2319_), .Y(_abc_40319_new_n2320_));
OR2X2 OR2X2_588 ( .A(_abc_40319_new_n2309_), .B(_abc_40319_new_n2320_), .Y(n1251));
OR2X2 OR2X2_589 ( .A(_abc_40319_new_n1558_), .B(_abc_40319_new_n2323_), .Y(_abc_40319_new_n2324_));
OR2X2 OR2X2_59 ( .A(_abc_40319_new_n789_), .B(_abc_40319_new_n793_), .Y(_abc_40319_new_n794_));
OR2X2 OR2X2_590 ( .A(_abc_40319_new_n980_), .B(_abc_40319_new_n2322_), .Y(_abc_40319_new_n2325_));
OR2X2 OR2X2_591 ( .A(_abc_40319_new_n2328_), .B(_abc_40319_new_n2329_), .Y(_abc_40319_new_n2330_));
OR2X2 OR2X2_592 ( .A(_abc_40319_new_n2333_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n2334_));
OR2X2 OR2X2_593 ( .A(_abc_40319_new_n2332_), .B(_abc_40319_new_n2334_), .Y(_abc_40319_new_n2335_));
OR2X2 OR2X2_594 ( .A(_abc_40319_new_n2336_), .B(_abc_40319_new_n2335_), .Y(_abc_40319_new_n2337_));
OR2X2 OR2X2_595 ( .A(_abc_40319_new_n2337_), .B(_abc_40319_new_n2331_), .Y(_abc_40319_new_n2338_));
OR2X2 OR2X2_596 ( .A(_abc_40319_new_n2327_), .B(_abc_40319_new_n2338_), .Y(n1246));
OR2X2 OR2X2_597 ( .A(_abc_40319_new_n1928_), .B(_abc_40319_new_n1638_), .Y(_abc_40319_new_n2340_));
OR2X2 OR2X2_598 ( .A(_abc_40319_new_n2341_), .B(_abc_40319_new_n1641_), .Y(_abc_40319_new_n2342_));
OR2X2 OR2X2_599 ( .A(_abc_40319_new_n2345_), .B(_abc_40319_new_n2346_), .Y(_abc_40319_new_n2347_));
OR2X2 OR2X2_6 ( .A(_abc_40319_new_n587_), .B(_abc_40319_new_n588_), .Y(_abc_40319_new_n589_));
OR2X2 OR2X2_60 ( .A(_abc_40319_new_n788_), .B(_abc_40319_new_n794_), .Y(_abc_40319_new_n795_));
OR2X2 OR2X2_600 ( .A(_abc_40319_new_n2351_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n2352_));
OR2X2 OR2X2_601 ( .A(_abc_40319_new_n2350_), .B(_abc_40319_new_n2352_), .Y(_abc_40319_new_n2353_));
OR2X2 OR2X2_602 ( .A(_abc_40319_new_n2349_), .B(_abc_40319_new_n2353_), .Y(_abc_40319_new_n2354_));
OR2X2 OR2X2_603 ( .A(_abc_40319_new_n2354_), .B(_abc_40319_new_n2348_), .Y(_abc_40319_new_n2355_));
OR2X2 OR2X2_604 ( .A(_abc_40319_new_n2344_), .B(_abc_40319_new_n2355_), .Y(n1241));
OR2X2 OR2X2_605 ( .A(_abc_40319_new_n2358_), .B(_abc_40319_new_n1552_), .Y(_abc_40319_new_n2359_));
OR2X2 OR2X2_606 ( .A(_abc_40319_new_n2357_), .B(_abc_40319_new_n964_), .Y(_abc_40319_new_n2360_));
OR2X2 OR2X2_607 ( .A(_abc_40319_new_n2362_), .B(_abc_40319_new_n2363_), .Y(_abc_40319_new_n2364_));
OR2X2 OR2X2_608 ( .A(_abc_40319_new_n2365_), .B(_abc_40319_new_n2367_), .Y(_abc_40319_new_n2368_));
OR2X2 OR2X2_609 ( .A(_abc_40319_new_n2369_), .B(_abc_40319_new_n2368_), .Y(_abc_40319_new_n2370_));
OR2X2 OR2X2_61 ( .A(_abc_40319_new_n796_), .B(_abc_40319_new_n785_), .Y(_abc_40319_new_n797_));
OR2X2 OR2X2_610 ( .A(_abc_40319_new_n2370_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n2371_));
OR2X2 OR2X2_611 ( .A(_abc_40319_new_n2364_), .B(_abc_40319_new_n2371_), .Y(n1236));
OR2X2 OR2X2_612 ( .A(_abc_40319_new_n2176_), .B(_abc_40319_new_n2374_), .Y(_abc_40319_new_n2375_));
OR2X2 OR2X2_613 ( .A(_abc_40319_new_n2175_), .B(_abc_40319_new_n2373_), .Y(_abc_40319_new_n2376_));
OR2X2 OR2X2_614 ( .A(_abc_40319_new_n2379_), .B(_abc_40319_new_n2380_), .Y(_abc_40319_new_n2381_));
OR2X2 OR2X2_615 ( .A(_abc_40319_new_n2384_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n2385_));
OR2X2 OR2X2_616 ( .A(_abc_40319_new_n2383_), .B(_abc_40319_new_n2385_), .Y(_abc_40319_new_n2386_));
OR2X2 OR2X2_617 ( .A(_abc_40319_new_n2387_), .B(_abc_40319_new_n2386_), .Y(_abc_40319_new_n2388_));
OR2X2 OR2X2_618 ( .A(_abc_40319_new_n2388_), .B(_abc_40319_new_n2382_), .Y(_abc_40319_new_n2389_));
OR2X2 OR2X2_619 ( .A(_abc_40319_new_n2378_), .B(_abc_40319_new_n2389_), .Y(n1231));
OR2X2 OR2X2_62 ( .A(_abc_40319_new_n798_), .B(_abc_40319_new_n799_), .Y(_abc_40319_new_n800_));
OR2X2 OR2X2_620 ( .A(_abc_40319_new_n2392_), .B(_abc_40319_new_n2393_), .Y(_abc_40319_new_n2394_));
OR2X2 OR2X2_621 ( .A(_abc_40319_new_n2391_), .B(_abc_40319_new_n2394_), .Y(_abc_40319_new_n2395_));
OR2X2 OR2X2_622 ( .A(_abc_40319_new_n2398_), .B(_abc_40319_new_n2397_), .Y(_abc_40319_new_n2399_));
OR2X2 OR2X2_623 ( .A(_abc_40319_new_n2396_), .B(_abc_40319_new_n2399_), .Y(_abc_40319_new_n2400_));
OR2X2 OR2X2_624 ( .A(_abc_40319_new_n2404_), .B(_abc_40319_new_n2405_), .Y(_abc_40319_new_n2406_));
OR2X2 OR2X2_625 ( .A(_abc_40319_new_n2406_), .B(_abc_40319_new_n2403_), .Y(_abc_40319_new_n2407_));
OR2X2 OR2X2_626 ( .A(_abc_40319_new_n2411_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n2412_));
OR2X2 OR2X2_627 ( .A(_abc_40319_new_n2410_), .B(_abc_40319_new_n2412_), .Y(_abc_40319_new_n2413_));
OR2X2 OR2X2_628 ( .A(_abc_40319_new_n2413_), .B(_abc_40319_new_n2409_), .Y(_abc_40319_new_n2414_));
OR2X2 OR2X2_629 ( .A(_abc_40319_new_n2414_), .B(_abc_40319_new_n2408_), .Y(_abc_40319_new_n2415_));
OR2X2 OR2X2_63 ( .A(_abc_40319_new_n800_), .B(_abc_40319_new_n768_), .Y(_abc_40319_new_n801_));
OR2X2 OR2X2_630 ( .A(_abc_40319_new_n2402_), .B(_abc_40319_new_n2415_), .Y(n1226));
OR2X2 OR2X2_631 ( .A(_abc_40319_new_n1904_), .B(_abc_40319_new_n2417_), .Y(_abc_40319_new_n2418_));
OR2X2 OR2X2_632 ( .A(_abc_40319_new_n1943_), .B(_abc_40319_new_n2419_), .Y(_abc_40319_new_n2420_));
OR2X2 OR2X2_633 ( .A(_abc_40319_new_n2424_), .B(_abc_40319_new_n2423_), .Y(_abc_40319_new_n2425_));
OR2X2 OR2X2_634 ( .A(_abc_40319_new_n2429_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n2430_));
OR2X2 OR2X2_635 ( .A(_abc_40319_new_n2428_), .B(_abc_40319_new_n2430_), .Y(_abc_40319_new_n2431_));
OR2X2 OR2X2_636 ( .A(_abc_40319_new_n2427_), .B(_abc_40319_new_n2431_), .Y(_abc_40319_new_n2432_));
OR2X2 OR2X2_637 ( .A(_abc_40319_new_n2432_), .B(_abc_40319_new_n2426_), .Y(_abc_40319_new_n2433_));
OR2X2 OR2X2_638 ( .A(_abc_40319_new_n2422_), .B(_abc_40319_new_n2433_), .Y(n1221));
OR2X2 OR2X2_639 ( .A(_abc_40319_new_n1747_), .B(_abc_40319_new_n1788_), .Y(_abc_40319_new_n2436_));
OR2X2 OR2X2_64 ( .A(_abc_40319_new_n802_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n803_));
OR2X2 OR2X2_640 ( .A(_abc_40319_new_n2435_), .B(_abc_40319_new_n2436_), .Y(_abc_40319_new_n2437_));
OR2X2 OR2X2_641 ( .A(_abc_40319_new_n2204_), .B(_abc_40319_new_n2438_), .Y(_abc_40319_new_n2439_));
OR2X2 OR2X2_642 ( .A(_abc_40319_new_n2442_), .B(_abc_40319_new_n2443_), .Y(_abc_40319_new_n2444_));
OR2X2 OR2X2_643 ( .A(_abc_40319_new_n2447_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n2448_));
OR2X2 OR2X2_644 ( .A(_abc_40319_new_n2446_), .B(_abc_40319_new_n2448_), .Y(_abc_40319_new_n2449_));
OR2X2 OR2X2_645 ( .A(_abc_40319_new_n2450_), .B(_abc_40319_new_n2449_), .Y(_abc_40319_new_n2451_));
OR2X2 OR2X2_646 ( .A(_abc_40319_new_n2451_), .B(_abc_40319_new_n2445_), .Y(_abc_40319_new_n2452_));
OR2X2 OR2X2_647 ( .A(_abc_40319_new_n2441_), .B(_abc_40319_new_n2452_), .Y(n1216));
OR2X2 OR2X2_648 ( .A(_abc_40319_new_n1556_), .B(_abc_40319_new_n2455_), .Y(_abc_40319_new_n2456_));
OR2X2 OR2X2_649 ( .A(_abc_40319_new_n968_), .B(_abc_40319_new_n2454_), .Y(_abc_40319_new_n2457_));
OR2X2 OR2X2_65 ( .A(_abc_40319_new_n805_), .B(_abc_40319_new_n797_), .Y(_abc_40319_new_n807_));
OR2X2 OR2X2_650 ( .A(_abc_40319_new_n2460_), .B(_abc_40319_new_n2461_), .Y(_abc_40319_new_n2462_));
OR2X2 OR2X2_651 ( .A(_abc_40319_new_n2466_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n2467_));
OR2X2 OR2X2_652 ( .A(_abc_40319_new_n2465_), .B(_abc_40319_new_n2467_), .Y(_abc_40319_new_n2468_));
OR2X2 OR2X2_653 ( .A(_abc_40319_new_n2464_), .B(_abc_40319_new_n2468_), .Y(_abc_40319_new_n2469_));
OR2X2 OR2X2_654 ( .A(_abc_40319_new_n2469_), .B(_abc_40319_new_n2463_), .Y(_abc_40319_new_n2470_));
OR2X2 OR2X2_655 ( .A(_abc_40319_new_n2459_), .B(_abc_40319_new_n2470_), .Y(n1211));
OR2X2 OR2X2_656 ( .A(_abc_40319_new_n1811_), .B(_abc_40319_new_n2472_), .Y(_abc_40319_new_n2473_));
OR2X2 OR2X2_657 ( .A(_abc_40319_new_n1938_), .B(_abc_40319_new_n2474_), .Y(_abc_40319_new_n2475_));
OR2X2 OR2X2_658 ( .A(_abc_40319_new_n2478_), .B(_abc_40319_new_n2479_), .Y(_abc_40319_new_n2480_));
OR2X2 OR2X2_659 ( .A(_abc_40319_new_n2484_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n2485_));
OR2X2 OR2X2_66 ( .A(_abc_40319_new_n676_), .B(_abc_40319_new_n808_), .Y(_abc_40319_new_n809_));
OR2X2 OR2X2_660 ( .A(_abc_40319_new_n2483_), .B(_abc_40319_new_n2485_), .Y(_abc_40319_new_n2486_));
OR2X2 OR2X2_661 ( .A(_abc_40319_new_n2482_), .B(_abc_40319_new_n2486_), .Y(_abc_40319_new_n2487_));
OR2X2 OR2X2_662 ( .A(_abc_40319_new_n2487_), .B(_abc_40319_new_n2481_), .Y(_abc_40319_new_n2488_));
OR2X2 OR2X2_663 ( .A(_abc_40319_new_n2477_), .B(_abc_40319_new_n2488_), .Y(n1206));
OR2X2 OR2X2_664 ( .A(_abc_40319_new_n985_), .B(_abc_40319_new_n2491_), .Y(_abc_40319_new_n2492_));
OR2X2 OR2X2_665 ( .A(_abc_40319_new_n984_), .B(_abc_40319_new_n2490_), .Y(_abc_40319_new_n2493_));
OR2X2 OR2X2_666 ( .A(_abc_40319_new_n2496_), .B(_abc_40319_new_n2497_), .Y(_abc_40319_new_n2498_));
OR2X2 OR2X2_667 ( .A(_abc_40319_new_n2502_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n2503_));
OR2X2 OR2X2_668 ( .A(_abc_40319_new_n2501_), .B(_abc_40319_new_n2503_), .Y(_abc_40319_new_n2504_));
OR2X2 OR2X2_669 ( .A(_abc_40319_new_n2500_), .B(_abc_40319_new_n2504_), .Y(_abc_40319_new_n2505_));
OR2X2 OR2X2_67 ( .A(_abc_40319_new_n811_), .B(_abc_40319_new_n812_), .Y(_abc_40319_new_n813_));
OR2X2 OR2X2_670 ( .A(_abc_40319_new_n2505_), .B(_abc_40319_new_n2499_), .Y(_abc_40319_new_n2506_));
OR2X2 OR2X2_671 ( .A(_abc_40319_new_n2495_), .B(_abc_40319_new_n2506_), .Y(n1201));
OR2X2 OR2X2_672 ( .A(_abc_40319_new_n2509_), .B(_abc_40319_new_n1299_), .Y(_abc_40319_new_n2510_));
OR2X2 OR2X2_673 ( .A(_abc_40319_new_n2508_), .B(_abc_40319_new_n2510_), .Y(_abc_40319_new_n2511_));
OR2X2 OR2X2_674 ( .A(_abc_40319_new_n2514_), .B(_abc_40319_new_n2513_), .Y(_abc_40319_new_n2515_));
OR2X2 OR2X2_675 ( .A(_abc_40319_new_n2512_), .B(_abc_40319_new_n2515_), .Y(_abc_40319_new_n2516_));
OR2X2 OR2X2_676 ( .A(_abc_40319_new_n2520_), .B(_abc_40319_new_n2519_), .Y(_abc_40319_new_n2521_));
OR2X2 OR2X2_677 ( .A(_abc_40319_new_n2525_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n2526_));
OR2X2 OR2X2_678 ( .A(_abc_40319_new_n2524_), .B(_abc_40319_new_n2526_), .Y(_abc_40319_new_n2527_));
OR2X2 OR2X2_679 ( .A(_abc_40319_new_n2523_), .B(_abc_40319_new_n2527_), .Y(_abc_40319_new_n2528_));
OR2X2 OR2X2_68 ( .A(_abc_40319_new_n628_), .B(_abc_40319_new_n638_), .Y(_abc_40319_new_n817_));
OR2X2 OR2X2_680 ( .A(_abc_40319_new_n2522_), .B(_abc_40319_new_n2528_), .Y(_abc_40319_new_n2529_));
OR2X2 OR2X2_681 ( .A(_abc_40319_new_n2518_), .B(_abc_40319_new_n2529_), .Y(n1196));
OR2X2 OR2X2_682 ( .A(_abc_40319_new_n1934_), .B(_abc_40319_new_n2532_), .Y(_abc_40319_new_n2533_));
OR2X2 OR2X2_683 ( .A(_abc_40319_new_n1800_), .B(_abc_40319_new_n2531_), .Y(_abc_40319_new_n2534_));
OR2X2 OR2X2_684 ( .A(_abc_40319_new_n2537_), .B(_abc_40319_new_n2538_), .Y(_abc_40319_new_n2539_));
OR2X2 OR2X2_685 ( .A(_abc_40319_new_n2542_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n2543_));
OR2X2 OR2X2_686 ( .A(_abc_40319_new_n2541_), .B(_abc_40319_new_n2543_), .Y(_abc_40319_new_n2544_));
OR2X2 OR2X2_687 ( .A(_abc_40319_new_n2545_), .B(_abc_40319_new_n2544_), .Y(_abc_40319_new_n2546_));
OR2X2 OR2X2_688 ( .A(_abc_40319_new_n2546_), .B(_abc_40319_new_n2540_), .Y(_abc_40319_new_n2547_));
OR2X2 OR2X2_689 ( .A(_abc_40319_new_n2536_), .B(_abc_40319_new_n2547_), .Y(n1191));
OR2X2 OR2X2_69 ( .A(_abc_40319_new_n815_), .B(_abc_40319_new_n818_), .Y(_abc_40319_new_n819_));
OR2X2 OR2X2_690 ( .A(_abc_40319_new_n2558_), .B(_abc_40319_new_n2557_), .Y(_abc_40319_new_n2559_));
OR2X2 OR2X2_691 ( .A(_abc_40319_new_n2559_), .B(_abc_40319_new_n2556_), .Y(_abc_40319_new_n2560_));
OR2X2 OR2X2_692 ( .A(_abc_40319_new_n2561_), .B(_abc_40319_new_n2554_), .Y(_abc_40319_new_n2562_));
OR2X2 OR2X2_693 ( .A(_abc_40319_new_n2564_), .B(_abc_40319_new_n2563_), .Y(_abc_40319_new_n2565_));
OR2X2 OR2X2_694 ( .A(_abc_40319_new_n2570_), .B(_abc_40319_new_n2571_), .Y(_abc_40319_new_n2572_));
OR2X2 OR2X2_695 ( .A(_abc_40319_new_n2572_), .B(_abc_40319_new_n2569_), .Y(_abc_40319_new_n2573_));
OR2X2 OR2X2_696 ( .A(_abc_40319_new_n2579_), .B(_abc_40319_new_n2577_), .Y(_abc_40319_new_n2580_));
OR2X2 OR2X2_697 ( .A(_abc_40319_new_n2586_), .B(_abc_40319_new_n2584_), .Y(_abc_40319_new_n2587_));
OR2X2 OR2X2_698 ( .A(_abc_40319_new_n2590_), .B(_abc_40319_new_n2591_), .Y(_abc_40319_new_n2592_));
OR2X2 OR2X2_699 ( .A(_abc_40319_new_n2592_), .B(_abc_40319_new_n2589_), .Y(_abc_40319_new_n2593_));
OR2X2 OR2X2_7 ( .A(_abc_40319_new_n572_), .B(_abc_40319_new_n573_), .Y(_abc_40319_new_n593_));
OR2X2 OR2X2_70 ( .A(_abc_40319_new_n822_), .B(_abc_40319_new_n823_), .Y(_abc_40319_new_n824_));
OR2X2 OR2X2_700 ( .A(_abc_40319_new_n2582_), .B(_abc_40319_new_n2595_), .Y(_abc_40319_new_n2596_));
OR2X2 OR2X2_701 ( .A(_abc_40319_new_n2599_), .B(_abc_40319_new_n2600_), .Y(_abc_40319_new_n2601_));
OR2X2 OR2X2_702 ( .A(_abc_40319_new_n2601_), .B(_abc_40319_new_n2598_), .Y(_abc_40319_new_n2602_));
OR2X2 OR2X2_703 ( .A(_abc_40319_new_n2606_), .B(_abc_40319_new_n2604_), .Y(_abc_40319_new_n2607_));
OR2X2 OR2X2_704 ( .A(_abc_40319_new_n2602_), .B(_abc_40319_new_n2607_), .Y(_abc_40319_new_n2608_));
OR2X2 OR2X2_705 ( .A(_abc_40319_new_n864_), .B(_abc_40319_new_n2611_), .Y(_abc_40319_new_n2612_));
OR2X2 OR2X2_706 ( .A(_abc_40319_new_n903_), .B(_abc_40319_new_n2549_), .Y(_abc_40319_new_n2615_));
OR2X2 OR2X2_707 ( .A(_abc_40319_new_n2620_), .B(_abc_40319_new_n2619_), .Y(_abc_40319_new_n2621_));
OR2X2 OR2X2_708 ( .A(_abc_40319_new_n2624_), .B(_abc_40319_new_n613_), .Y(_abc_40319_new_n2625_));
OR2X2 OR2X2_709 ( .A(_abc_40319_new_n2625_), .B(_abc_40319_new_n2626_), .Y(_abc_40319_new_n2627_));
OR2X2 OR2X2_71 ( .A(_abc_40319_new_n825_), .B(_abc_40319_new_n827_), .Y(_abc_40319_new_n828_));
OR2X2 OR2X2_710 ( .A(_abc_40319_new_n2627_), .B(_abc_40319_new_n2628_), .Y(_abc_40319_new_n2629_));
OR2X2 OR2X2_711 ( .A(_abc_40319_new_n2630_), .B(_abc_40319_new_n2631_), .Y(_abc_40319_new_n2632_));
OR2X2 OR2X2_712 ( .A(_abc_40319_new_n2632_), .B(_abc_40319_new_n2633_), .Y(_abc_40319_new_n2634_));
OR2X2 OR2X2_713 ( .A(_abc_40319_new_n2636_), .B(_abc_40319_new_n2637_), .Y(_abc_40319_new_n2638_));
OR2X2 OR2X2_714 ( .A(_abc_40319_new_n2640_), .B(_abc_40319_new_n613_), .Y(_abc_40319_new_n2641_));
OR2X2 OR2X2_715 ( .A(_abc_40319_new_n2641_), .B(_abc_40319_new_n2642_), .Y(_abc_40319_new_n2643_));
OR2X2 OR2X2_716 ( .A(_abc_40319_new_n2643_), .B(_abc_40319_new_n2644_), .Y(_abc_40319_new_n2645_));
OR2X2 OR2X2_717 ( .A(_abc_40319_new_n2645_), .B(_abc_40319_new_n2639_), .Y(_abc_40319_new_n2646_));
OR2X2 OR2X2_718 ( .A(_abc_40319_new_n2647_), .B(_abc_40319_new_n2629_), .Y(_abc_40319_new_n2648_));
OR2X2 OR2X2_719 ( .A(_abc_40319_new_n2650_), .B(_abc_40319_new_n2611_), .Y(_abc_40319_new_n2651_));
OR2X2 OR2X2_72 ( .A(_abc_40319_new_n824_), .B(_abc_40319_new_n828_), .Y(_abc_40319_new_n829_));
OR2X2 OR2X2_720 ( .A(_abc_40319_new_n819_), .B(_abc_40319_new_n2551_), .Y(_abc_40319_new_n2652_));
OR2X2 OR2X2_721 ( .A(_abc_40319_new_n864_), .B(_abc_40319_new_n2549_), .Y(_abc_40319_new_n2653_));
OR2X2 OR2X2_722 ( .A(_abc_40319_new_n829_), .B(_abc_40319_new_n2656_), .Y(_abc_40319_new_n2657_));
OR2X2 OR2X2_723 ( .A(_abc_40319_new_n820_), .B(_abc_40319_new_n2611_), .Y(_abc_40319_new_n2658_));
OR2X2 OR2X2_724 ( .A(_abc_40319_new_n2655_), .B(_abc_40319_new_n2659_), .Y(_abc_40319_new_n2660_));
OR2X2 OR2X2_725 ( .A(_abc_40319_new_n2662_), .B(_abc_40319_new_n613_), .Y(_abc_40319_new_n2663_));
OR2X2 OR2X2_726 ( .A(_abc_40319_new_n2663_), .B(_abc_40319_new_n2661_), .Y(_abc_40319_new_n2664_));
OR2X2 OR2X2_727 ( .A(_abc_40319_new_n2650_), .B(_abc_40319_new_n2549_), .Y(_abc_40319_new_n2669_));
OR2X2 OR2X2_728 ( .A(_abc_40319_new_n2671_), .B(_abc_40319_new_n2664_), .Y(_abc_40319_new_n2672_));
OR2X2 OR2X2_729 ( .A(_abc_40319_new_n954_), .B(_abc_40319_new_n646_), .Y(_abc_40319_new_n2673_));
OR2X2 OR2X2_73 ( .A(_abc_40319_new_n821_), .B(_abc_40319_new_n830_), .Y(_abc_40319_new_n831_));
OR2X2 OR2X2_730 ( .A(_abc_40319_new_n2691_), .B(_abc_40319_new_n2687_), .Y(_abc_40319_new_n2692_));
OR2X2 OR2X2_731 ( .A(_abc_40319_new_n2692_), .B(_abc_40319_new_n2686_), .Y(_abc_40319_new_n2693_));
OR2X2 OR2X2_732 ( .A(_abc_40319_new_n2684_), .B(_abc_40319_new_n2693_), .Y(_abc_40319_new_n2694_));
OR2X2 OR2X2_733 ( .A(_abc_40319_new_n2694_), .B(_abc_40319_new_n2610_), .Y(_abc_40319_new_n2695_));
OR2X2 OR2X2_734 ( .A(_abc_40319_new_n2697_), .B(_abc_40319_new_n2698_), .Y(_abc_40319_new_n2699_));
OR2X2 OR2X2_735 ( .A(_abc_40319_new_n2699_), .B(_abc_40319_new_n2696_), .Y(_abc_40319_new_n2700_));
OR2X2 OR2X2_736 ( .A(_abc_40319_new_n2704_), .B(_abc_40319_new_n2702_), .Y(_abc_40319_new_n2705_));
OR2X2 OR2X2_737 ( .A(_abc_40319_new_n2708_), .B(_abc_40319_new_n2709_), .Y(_abc_40319_new_n2710_));
OR2X2 OR2X2_738 ( .A(_abc_40319_new_n2710_), .B(_abc_40319_new_n2707_), .Y(_abc_40319_new_n2711_));
OR2X2 OR2X2_739 ( .A(_abc_40319_new_n2715_), .B(_abc_40319_new_n2713_), .Y(_abc_40319_new_n2716_));
OR2X2 OR2X2_74 ( .A(_abc_40319_new_n833_), .B(_abc_40319_new_n834_), .Y(_abc_40319_new_n835_));
OR2X2 OR2X2_740 ( .A(_abc_40319_new_n2706_), .B(_abc_40319_new_n2717_), .Y(_abc_40319_new_n2718_));
OR2X2 OR2X2_741 ( .A(_abc_40319_new_n2594_), .B(_abc_40319_new_n2588_), .Y(_abc_40319_new_n2720_));
OR2X2 OR2X2_742 ( .A(_abc_40319_new_n2720_), .B(_abc_40319_new_n2582_), .Y(_abc_40319_new_n2721_));
OR2X2 OR2X2_743 ( .A(_abc_40319_new_n2724_), .B(_abc_40319_new_n2725_), .Y(_abc_40319_new_n2726_));
OR2X2 OR2X2_744 ( .A(_abc_40319_new_n2726_), .B(_abc_40319_new_n2723_), .Y(_abc_40319_new_n2727_));
OR2X2 OR2X2_745 ( .A(_abc_40319_new_n2731_), .B(_abc_40319_new_n2729_), .Y(_abc_40319_new_n2732_));
OR2X2 OR2X2_746 ( .A(_abc_40319_new_n2722_), .B(_abc_40319_new_n2733_), .Y(_abc_40319_new_n2734_));
OR2X2 OR2X2_747 ( .A(_abc_40319_new_n2727_), .B(_abc_40319_new_n2732_), .Y(_abc_40319_new_n2743_));
OR2X2 OR2X2_748 ( .A(_abc_40319_new_n2718_), .B(_abc_40319_new_n2743_), .Y(_abc_40319_new_n2744_));
OR2X2 OR2X2_749 ( .A(_abc_40319_new_n2711_), .B(_abc_40319_new_n2716_), .Y(_abc_40319_new_n2745_));
OR2X2 OR2X2_75 ( .A(_abc_40319_new_n837_), .B(_abc_40319_new_n836_), .Y(_abc_40319_new_n838_));
OR2X2 OR2X2_750 ( .A(_abc_40319_new_n2745_), .B(_abc_40319_new_n2706_), .Y(_abc_40319_new_n2746_));
OR2X2 OR2X2_751 ( .A(_abc_40319_new_n2748_), .B(_abc_40319_new_n2749_), .Y(_abc_40319_new_n2750_));
OR2X2 OR2X2_752 ( .A(_abc_40319_new_n2750_), .B(_abc_40319_new_n2747_), .Y(_abc_40319_new_n2751_));
OR2X2 OR2X2_753 ( .A(_abc_40319_new_n2756_), .B(_abc_40319_new_n2754_), .Y(_abc_40319_new_n2757_));
OR2X2 OR2X2_754 ( .A(_abc_40319_new_n2763_), .B(_abc_40319_new_n2761_), .Y(_abc_40319_new_n2764_));
OR2X2 OR2X2_755 ( .A(_abc_40319_new_n2767_), .B(_abc_40319_new_n2768_), .Y(_abc_40319_new_n2769_));
OR2X2 OR2X2_756 ( .A(_abc_40319_new_n2769_), .B(_abc_40319_new_n2766_), .Y(_abc_40319_new_n2770_));
OR2X2 OR2X2_757 ( .A(_abc_40319_new_n2759_), .B(_abc_40319_new_n2772_), .Y(_abc_40319_new_n2773_));
OR2X2 OR2X2_758 ( .A(_abc_40319_new_n2700_), .B(_abc_40319_new_n2705_), .Y(_abc_40319_new_n2775_));
OR2X2 OR2X2_759 ( .A(_abc_40319_new_n2777_), .B(_abc_40319_new_n2778_), .Y(_abc_40319_new_n2779_));
OR2X2 OR2X2_76 ( .A(_abc_40319_new_n839_), .B(_abc_40319_new_n528_), .Y(_abc_40319_new_n840_));
OR2X2 OR2X2_760 ( .A(_abc_40319_new_n2779_), .B(_abc_40319_new_n2776_), .Y(_abc_40319_new_n2780_));
OR2X2 OR2X2_761 ( .A(_abc_40319_new_n2785_), .B(_abc_40319_new_n2783_), .Y(_abc_40319_new_n2786_));
OR2X2 OR2X2_762 ( .A(_abc_40319_new_n2742_), .B(_abc_40319_new_n2794_), .Y(_abc_40319_new_n2795_));
OR2X2 OR2X2_763 ( .A(_abc_40319_new_n2803_), .B(_abc_40319_new_n2804_), .Y(_abc_40319_new_n2805_));
OR2X2 OR2X2_764 ( .A(_abc_40319_new_n2805_), .B(_abc_40319_new_n2802_), .Y(_abc_40319_new_n2806_));
OR2X2 OR2X2_765 ( .A(_abc_40319_new_n2810_), .B(_abc_40319_new_n2808_), .Y(_abc_40319_new_n2811_));
OR2X2 OR2X2_766 ( .A(_abc_40319_new_n2801_), .B(_abc_40319_new_n2812_), .Y(_abc_40319_new_n2813_));
OR2X2 OR2X2_767 ( .A(_abc_40319_new_n2800_), .B(_abc_40319_new_n2813_), .Y(_abc_40319_new_n2814_));
OR2X2 OR2X2_768 ( .A(_abc_40319_new_n2797_), .B(_abc_40319_new_n2814_), .Y(_abc_40319_new_n2815_));
OR2X2 OR2X2_769 ( .A(_abc_40319_new_n2806_), .B(_abc_40319_new_n2811_), .Y(_abc_40319_new_n2818_));
OR2X2 OR2X2_77 ( .A(_abc_40319_new_n844_), .B(_abc_40319_new_n846_), .Y(_abc_40319_new_n847_));
OR2X2 OR2X2_770 ( .A(_abc_40319_new_n2820_), .B(_abc_40319_new_n2821_), .Y(_abc_40319_new_n2822_));
OR2X2 OR2X2_771 ( .A(_abc_40319_new_n2822_), .B(_abc_40319_new_n2819_), .Y(_abc_40319_new_n2823_));
OR2X2 OR2X2_772 ( .A(_abc_40319_new_n2828_), .B(_abc_40319_new_n2826_), .Y(_abc_40319_new_n2829_));
OR2X2 OR2X2_773 ( .A(_abc_40319_new_n2817_), .B(_abc_40319_new_n2834_), .Y(_abc_40319_new_n2835_));
OR2X2 OR2X2_774 ( .A(_abc_40319_new_n2838_), .B(_abc_40319_new_n2839_), .Y(_abc_40319_new_n2840_));
OR2X2 OR2X2_775 ( .A(_abc_40319_new_n2840_), .B(_abc_40319_new_n2837_), .Y(_abc_40319_new_n2841_));
OR2X2 OR2X2_776 ( .A(_abc_40319_new_n2845_), .B(_abc_40319_new_n2843_), .Y(_abc_40319_new_n2846_));
OR2X2 OR2X2_777 ( .A(_abc_40319_new_n2836_), .B(_abc_40319_new_n2847_), .Y(_abc_40319_new_n2848_));
OR2X2 OR2X2_778 ( .A(_abc_40319_new_n2841_), .B(_abc_40319_new_n2846_), .Y(_abc_40319_new_n2851_));
OR2X2 OR2X2_779 ( .A(_abc_40319_new_n2853_), .B(_abc_40319_new_n2854_), .Y(_abc_40319_new_n2855_));
OR2X2 OR2X2_78 ( .A(_abc_40319_new_n716_), .B(_abc_40319_new_n732_), .Y(_abc_40319_new_n851_));
OR2X2 OR2X2_780 ( .A(_abc_40319_new_n2855_), .B(_abc_40319_new_n2852_), .Y(_abc_40319_new_n2856_));
OR2X2 OR2X2_781 ( .A(_abc_40319_new_n2861_), .B(_abc_40319_new_n2859_), .Y(_abc_40319_new_n2862_));
OR2X2 OR2X2_782 ( .A(_abc_40319_new_n2850_), .B(_abc_40319_new_n2867_), .Y(_abc_40319_new_n2868_));
OR2X2 OR2X2_783 ( .A(_abc_40319_new_n2871_), .B(_abc_40319_new_n2872_), .Y(_abc_40319_new_n2873_));
OR2X2 OR2X2_784 ( .A(_abc_40319_new_n2873_), .B(_abc_40319_new_n2870_), .Y(_abc_40319_new_n2874_));
OR2X2 OR2X2_785 ( .A(_abc_40319_new_n2876_), .B(_abc_40319_new_n2878_), .Y(_abc_40319_new_n2879_));
OR2X2 OR2X2_786 ( .A(_abc_40319_new_n2880_), .B(_abc_40319_new_n2869_), .Y(_abc_40319_new_n2881_));
OR2X2 OR2X2_787 ( .A(_abc_40319_new_n2879_), .B(_abc_40319_new_n2874_), .Y(_abc_40319_new_n2884_));
OR2X2 OR2X2_788 ( .A(_abc_40319_new_n2887_), .B(_abc_40319_new_n2886_), .Y(_abc_40319_new_n2888_));
OR2X2 OR2X2_789 ( .A(_abc_40319_new_n2888_), .B(_abc_40319_new_n2885_), .Y(_abc_40319_new_n2889_));
OR2X2 OR2X2_79 ( .A(_abc_40319_new_n851_), .B(_abc_40319_new_n850_), .Y(_abc_40319_new_n852_));
OR2X2 OR2X2_790 ( .A(_abc_40319_new_n2892_), .B(_abc_40319_new_n2894_), .Y(_abc_40319_new_n2895_));
OR2X2 OR2X2_791 ( .A(_abc_40319_new_n2883_), .B(_abc_40319_new_n2900_), .Y(_abc_40319_new_n2901_));
OR2X2 OR2X2_792 ( .A(_abc_40319_new_n2905_), .B(_abc_40319_new_n2904_), .Y(_abc_40319_new_n2906_));
OR2X2 OR2X2_793 ( .A(_abc_40319_new_n2906_), .B(_abc_40319_new_n2903_), .Y(_abc_40319_new_n2907_));
OR2X2 OR2X2_794 ( .A(_abc_40319_new_n2909_), .B(_abc_40319_new_n2911_), .Y(_abc_40319_new_n2912_));
OR2X2 OR2X2_795 ( .A(_abc_40319_new_n2902_), .B(_abc_40319_new_n2913_), .Y(_abc_40319_new_n2914_));
OR2X2 OR2X2_796 ( .A(_abc_40319_new_n2907_), .B(_abc_40319_new_n2912_), .Y(_abc_40319_new_n2917_));
OR2X2 OR2X2_797 ( .A(_abc_40319_new_n2920_), .B(_abc_40319_new_n2919_), .Y(_abc_40319_new_n2921_));
OR2X2 OR2X2_798 ( .A(_abc_40319_new_n2921_), .B(_abc_40319_new_n2918_), .Y(_abc_40319_new_n2922_));
OR2X2 OR2X2_799 ( .A(_abc_40319_new_n2925_), .B(_abc_40319_new_n2927_), .Y(_abc_40319_new_n2928_));
OR2X2 OR2X2_8 ( .A(_abc_40319_new_n594_), .B(_abc_40319_new_n524_), .Y(_abc_40319_new_n595_));
OR2X2 OR2X2_80 ( .A(_abc_40319_new_n729_), .B(_abc_40319_new_n732_), .Y(_abc_40319_new_n854_));
OR2X2 OR2X2_800 ( .A(_abc_40319_new_n2916_), .B(_abc_40319_new_n2933_), .Y(_abc_40319_new_n2934_));
OR2X2 OR2X2_801 ( .A(_abc_40319_new_n2938_), .B(_abc_40319_new_n2937_), .Y(_abc_40319_new_n2939_));
OR2X2 OR2X2_802 ( .A(_abc_40319_new_n2939_), .B(_abc_40319_new_n2936_), .Y(_abc_40319_new_n2940_));
OR2X2 OR2X2_803 ( .A(_abc_40319_new_n2942_), .B(_abc_40319_new_n2944_), .Y(_abc_40319_new_n2945_));
OR2X2 OR2X2_804 ( .A(_abc_40319_new_n2946_), .B(_abc_40319_new_n2935_), .Y(_abc_40319_new_n2947_));
OR2X2 OR2X2_805 ( .A(_abc_40319_new_n2945_), .B(_abc_40319_new_n2940_), .Y(_abc_40319_new_n2950_));
OR2X2 OR2X2_806 ( .A(_abc_40319_new_n2953_), .B(_abc_40319_new_n2952_), .Y(_abc_40319_new_n2954_));
OR2X2 OR2X2_807 ( .A(_abc_40319_new_n2954_), .B(_abc_40319_new_n2951_), .Y(_abc_40319_new_n2955_));
OR2X2 OR2X2_808 ( .A(_abc_40319_new_n2958_), .B(_abc_40319_new_n2960_), .Y(_abc_40319_new_n2961_));
OR2X2 OR2X2_809 ( .A(_abc_40319_new_n2949_), .B(_abc_40319_new_n2966_), .Y(_abc_40319_new_n2967_));
OR2X2 OR2X2_81 ( .A(_abc_40319_new_n854_), .B(_abc_40319_new_n853_), .Y(_abc_40319_new_n855_));
OR2X2 OR2X2_810 ( .A(_abc_40319_new_n2971_), .B(_abc_40319_new_n2970_), .Y(_abc_40319_new_n2972_));
OR2X2 OR2X2_811 ( .A(_abc_40319_new_n2972_), .B(_abc_40319_new_n2969_), .Y(_abc_40319_new_n2973_));
OR2X2 OR2X2_812 ( .A(_abc_40319_new_n2975_), .B(_abc_40319_new_n2977_), .Y(_abc_40319_new_n2978_));
OR2X2 OR2X2_813 ( .A(_abc_40319_new_n2979_), .B(_abc_40319_new_n2968_), .Y(_abc_40319_new_n2980_));
OR2X2 OR2X2_814 ( .A(_abc_40319_new_n2978_), .B(_abc_40319_new_n2973_), .Y(_abc_40319_new_n2983_));
OR2X2 OR2X2_815 ( .A(_abc_40319_new_n2986_), .B(_abc_40319_new_n2985_), .Y(_abc_40319_new_n2987_));
OR2X2 OR2X2_816 ( .A(_abc_40319_new_n2987_), .B(_abc_40319_new_n2984_), .Y(_abc_40319_new_n2988_));
OR2X2 OR2X2_817 ( .A(_abc_40319_new_n2991_), .B(_abc_40319_new_n2993_), .Y(_abc_40319_new_n2994_));
OR2X2 OR2X2_818 ( .A(_abc_40319_new_n2982_), .B(_abc_40319_new_n2999_), .Y(_abc_40319_new_n3000_));
OR2X2 OR2X2_819 ( .A(_abc_40319_new_n3004_), .B(_abc_40319_new_n3003_), .Y(_abc_40319_new_n3005_));
OR2X2 OR2X2_82 ( .A(_abc_40319_new_n729_), .B(_abc_40319_new_n721_), .Y(_abc_40319_new_n858_));
OR2X2 OR2X2_820 ( .A(_abc_40319_new_n3005_), .B(_abc_40319_new_n3002_), .Y(_abc_40319_new_n3006_));
OR2X2 OR2X2_821 ( .A(_abc_40319_new_n3008_), .B(_abc_40319_new_n3010_), .Y(_abc_40319_new_n3011_));
OR2X2 OR2X2_822 ( .A(_abc_40319_new_n3012_), .B(_abc_40319_new_n3001_), .Y(_abc_40319_new_n3013_));
OR2X2 OR2X2_823 ( .A(_abc_40319_new_n3011_), .B(_abc_40319_new_n3006_), .Y(_abc_40319_new_n3016_));
OR2X2 OR2X2_824 ( .A(_abc_40319_new_n3019_), .B(_abc_40319_new_n3018_), .Y(_abc_40319_new_n3020_));
OR2X2 OR2X2_825 ( .A(_abc_40319_new_n3020_), .B(_abc_40319_new_n3017_), .Y(_abc_40319_new_n3021_));
OR2X2 OR2X2_826 ( .A(_abc_40319_new_n3024_), .B(_abc_40319_new_n3026_), .Y(_abc_40319_new_n3027_));
OR2X2 OR2X2_827 ( .A(_abc_40319_new_n3015_), .B(_abc_40319_new_n3032_), .Y(_abc_40319_new_n3033_));
OR2X2 OR2X2_828 ( .A(_abc_40319_new_n3037_), .B(_abc_40319_new_n3036_), .Y(_abc_40319_new_n3038_));
OR2X2 OR2X2_829 ( .A(_abc_40319_new_n3035_), .B(_abc_40319_new_n3038_), .Y(_abc_40319_new_n3039_));
OR2X2 OR2X2_83 ( .A(_abc_40319_new_n858_), .B(_abc_40319_new_n857_), .Y(_abc_40319_new_n859_));
OR2X2 OR2X2_830 ( .A(_abc_40319_new_n3041_), .B(_abc_40319_new_n3043_), .Y(_abc_40319_new_n3044_));
OR2X2 OR2X2_831 ( .A(_abc_40319_new_n3045_), .B(_abc_40319_new_n3034_), .Y(_abc_40319_new_n3046_));
OR2X2 OR2X2_832 ( .A(_abc_40319_new_n3044_), .B(_abc_40319_new_n3039_), .Y(_abc_40319_new_n3049_));
OR2X2 OR2X2_833 ( .A(_abc_40319_new_n3053_), .B(_abc_40319_new_n3052_), .Y(_abc_40319_new_n3054_));
OR2X2 OR2X2_834 ( .A(_abc_40319_new_n3050_), .B(_abc_40319_new_n3054_), .Y(_abc_40319_new_n3055_));
OR2X2 OR2X2_835 ( .A(_abc_40319_new_n3058_), .B(_abc_40319_new_n3060_), .Y(_abc_40319_new_n3061_));
OR2X2 OR2X2_836 ( .A(_abc_40319_new_n3048_), .B(_abc_40319_new_n3066_), .Y(_abc_40319_new_n3067_));
OR2X2 OR2X2_837 ( .A(_abc_40319_new_n3073_), .B(_abc_40319_new_n3072_), .Y(_abc_40319_new_n3074_));
OR2X2 OR2X2_838 ( .A(_abc_40319_new_n3074_), .B(_abc_40319_new_n3071_), .Y(_abc_40319_new_n3075_));
OR2X2 OR2X2_839 ( .A(_abc_40319_new_n3076_), .B(_abc_40319_new_n3070_), .Y(_abc_40319_new_n3077_));
OR2X2 OR2X2_84 ( .A(_abc_40319_new_n716_), .B(_abc_40319_new_n721_), .Y(_abc_40319_new_n861_));
OR2X2 OR2X2_840 ( .A(_abc_40319_new_n3080_), .B(_abc_40319_new_n3081_), .Y(_abc_40319_new_n3082_));
OR2X2 OR2X2_841 ( .A(_abc_40319_new_n3082_), .B(_abc_40319_new_n3079_), .Y(_abc_40319_new_n3083_));
OR2X2 OR2X2_842 ( .A(_abc_40319_new_n3068_), .B(_abc_40319_new_n3085_), .Y(_abc_40319_new_n3086_));
OR2X2 OR2X2_843 ( .A(_abc_40319_new_n3084_), .B(_abc_40319_new_n3077_), .Y(_abc_40319_new_n3089_));
OR2X2 OR2X2_844 ( .A(_abc_40319_new_n2566_), .B(_abc_40319_new_n2562_), .Y(_abc_40319_new_n3090_));
OR2X2 OR2X2_845 ( .A(_abc_40319_new_n3088_), .B(_abc_40319_new_n3092_), .Y(_abc_40319_new_n3093_));
OR2X2 OR2X2_846 ( .A(_abc_40319_new_n3094_), .B(_abc_40319_new_n1115_), .Y(_abc_40319_new_n3095_));
OR2X2 OR2X2_847 ( .A(_abc_40319_new_n3105_), .B(_abc_40319_new_n3104_), .Y(_abc_40319_new_n3106_));
OR2X2 OR2X2_848 ( .A(_abc_40319_new_n3108_), .B(_abc_40319_new_n3109_), .Y(_abc_40319_new_n3110_));
OR2X2 OR2X2_849 ( .A(_abc_40319_new_n3111_), .B(_abc_40319_new_n3112_), .Y(_abc_40319_new_n3113_));
OR2X2 OR2X2_85 ( .A(_abc_40319_new_n861_), .B(_abc_40319_new_n860_), .Y(_abc_40319_new_n862_));
OR2X2 OR2X2_850 ( .A(_abc_40319_new_n903_), .B(_abc_40319_new_n891_), .Y(_abc_40319_new_n3115_));
OR2X2 OR2X2_851 ( .A(_abc_40319_new_n3116_), .B(_abc_40319_new_n3117_), .Y(_abc_40319_new_n3118_));
OR2X2 OR2X2_852 ( .A(_abc_40319_new_n3121_), .B(_abc_40319_new_n3122_), .Y(_abc_40319_new_n3123_));
OR2X2 OR2X2_853 ( .A(_abc_40319_new_n3125_), .B(_abc_40319_new_n3126_), .Y(_abc_40319_new_n3127_));
OR2X2 OR2X2_854 ( .A(_abc_40319_new_n3132_), .B(_abc_40319_new_n3131_), .Y(_abc_40319_new_n3133_));
OR2X2 OR2X2_855 ( .A(_abc_40319_new_n3135_), .B(_abc_40319_new_n3136_), .Y(_abc_40319_new_n3137_));
OR2X2 OR2X2_856 ( .A(_abc_40319_new_n3140_), .B(_abc_40319_new_n3141_), .Y(_abc_40319_new_n3142_));
OR2X2 OR2X2_857 ( .A(_abc_40319_new_n3144_), .B(_abc_40319_new_n3145_), .Y(_abc_40319_new_n3146_));
OR2X2 OR2X2_858 ( .A(_abc_40319_new_n3152_), .B(_abc_40319_new_n3151_), .Y(_abc_40319_new_n3153_));
OR2X2 OR2X2_859 ( .A(_abc_40319_new_n3155_), .B(_abc_40319_new_n3156_), .Y(_abc_40319_new_n3157_));
OR2X2 OR2X2_86 ( .A(_abc_40319_new_n866_), .B(_abc_40319_new_n849_), .Y(_abc_40319_new_n867_));
OR2X2 OR2X2_860 ( .A(_abc_40319_new_n3174_), .B(_abc_40319_new_n3175_), .Y(_abc_40319_new_n3176_));
OR2X2 OR2X2_861 ( .A(_abc_40319_new_n3183_), .B(_abc_40319_new_n3184_), .Y(_abc_40319_new_n3185_));
OR2X2 OR2X2_862 ( .A(_abc_40319_new_n3188_), .B(_abc_40319_new_n3187_), .Y(_abc_40319_new_n3189_));
OR2X2 OR2X2_863 ( .A(_abc_40319_new_n3193_), .B(_abc_40319_new_n3194_), .Y(_abc_40319_new_n3195_));
OR2X2 OR2X2_864 ( .A(_abc_40319_new_n3198_), .B(_abc_40319_new_n3197_), .Y(_abc_40319_new_n3199_));
OR2X2 OR2X2_865 ( .A(_abc_40319_new_n3202_), .B(_abc_40319_new_n3201_), .Y(_abc_40319_new_n3203_));
OR2X2 OR2X2_866 ( .A(_abc_40319_new_n3205_), .B(_abc_40319_new_n3206_), .Y(_abc_40319_new_n3207_));
OR2X2 OR2X2_867 ( .A(_abc_40319_new_n3209_), .B(_abc_40319_new_n3210_), .Y(_abc_40319_new_n3211_));
OR2X2 OR2X2_868 ( .A(_abc_40319_new_n3213_), .B(_abc_40319_new_n3214_), .Y(_abc_40319_new_n3215_));
OR2X2 OR2X2_869 ( .A(_abc_40319_new_n3219_), .B(_abc_40319_new_n3221_), .Y(_abc_40319_new_n3222_));
OR2X2 OR2X2_87 ( .A(_abc_40319_new_n868_), .B(_abc_40319_new_n869_), .Y(_abc_40319_new_n870_));
OR2X2 OR2X2_870 ( .A(_abc_40319_new_n3224_), .B(_abc_40319_new_n3225_), .Y(_abc_40319_new_n3226_));
OR2X2 OR2X2_871 ( .A(_abc_40319_new_n3229_), .B(_abc_40319_new_n3230_), .Y(_abc_40319_new_n3231_));
OR2X2 OR2X2_872 ( .A(_abc_40319_new_n3233_), .B(_abc_40319_new_n3234_), .Y(_abc_40319_new_n3235_));
OR2X2 OR2X2_873 ( .A(_abc_40319_new_n3248_), .B(_abc_40319_new_n3247_), .Y(_abc_40319_new_n3249_));
OR2X2 OR2X2_874 ( .A(_abc_40319_new_n3252_), .B(_abc_40319_new_n3251_), .Y(_abc_40319_new_n3253_));
OR2X2 OR2X2_875 ( .A(_abc_40319_new_n3256_), .B(_abc_40319_new_n3255_), .Y(_abc_40319_new_n3257_));
OR2X2 OR2X2_876 ( .A(_abc_40319_new_n3259_), .B(_abc_40319_new_n3260_), .Y(_abc_40319_new_n3261_));
OR2X2 OR2X2_877 ( .A(_abc_40319_new_n3255_), .B(_abc_40319_new_n3194_), .Y(_abc_40319_new_n3281_));
OR2X2 OR2X2_878 ( .A(_abc_40319_new_n3281_), .B(_abc_40319_new_n3104_), .Y(_abc_40319_new_n3282_));
OR2X2 OR2X2_879 ( .A(_abc_40319_new_n3282_), .B(_abc_40319_new_n3280_), .Y(_abc_40319_new_n3283_));
OR2X2 OR2X2_88 ( .A(_abc_40319_new_n870_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n871_));
OR2X2 OR2X2_880 ( .A(_abc_40319_new_n3294_), .B(_abc_40319_new_n3296_), .Y(_abc_40319_new_n3297_));
OR2X2 OR2X2_881 ( .A(_abc_40319_new_n3300_), .B(_abc_40319_new_n3188_), .Y(_abc_40319_new_n3301_));
OR2X2 OR2X2_882 ( .A(_abc_40319_new_n3313_), .B(_abc_40319_new_n3234_), .Y(_abc_40319_new_n3314_));
OR2X2 OR2X2_883 ( .A(_abc_40319_new_n3323_), .B(_abc_40319_new_n3302_), .Y(_abc_40319_new_n3324_));
OR2X2 OR2X2_884 ( .A(_abc_40319_new_n3332_), .B(_abc_40319_new_n3214_), .Y(_abc_40319_new_n3333_));
OR2X2 OR2X2_885 ( .A(_abc_40319_new_n1166_), .B(_abc_40319_new_n655_), .Y(_abc_40319_new_n3342_));
OR2X2 OR2X2_886 ( .A(_abc_40319_new_n3136_), .B(_abc_40319_new_n3342_), .Y(_abc_40319_new_n3343_));
OR2X2 OR2X2_887 ( .A(_abc_40319_new_n3116_), .B(_abc_40319_new_n3135_), .Y(_abc_40319_new_n3344_));
OR2X2 OR2X2_888 ( .A(_abc_40319_new_n3341_), .B(_abc_40319_new_n3352_), .Y(_abc_40319_new_n3353_));
OR2X2 OR2X2_889 ( .A(_abc_40319_new_n3360_), .B(_abc_40319_new_n3362_), .Y(_abc_40319_new_n3363_));
OR2X2 OR2X2_89 ( .A(_abc_40319_new_n874_), .B(_abc_40319_new_n768_), .Y(_abc_40319_new_n875_));
OR2X2 OR2X2_890 ( .A(_abc_40319_new_n3363_), .B(_abc_40319_new_n3357_), .Y(_abc_40319_new_n3364_));
OR2X2 OR2X2_891 ( .A(_abc_40319_new_n3367_), .B(_abc_40319_new_n3366_), .Y(_abc_40319_new_n3368_));
OR2X2 OR2X2_892 ( .A(_abc_40319_new_n3369_), .B(_abc_40319_new_n3371_), .Y(_abc_40319_new_n3372_));
OR2X2 OR2X2_893 ( .A(_abc_40319_new_n3380_), .B(_abc_40319_new_n3104_), .Y(_abc_40319_new_n3381_));
OR2X2 OR2X2_894 ( .A(_abc_40319_new_n3395_), .B(_abc_40319_new_n3274_), .Y(_abc_40319_new_n3396_));
OR2X2 OR2X2_895 ( .A(_abc_40319_new_n3248_), .B(_abc_40319_new_n3252_), .Y(_abc_40319_new_n3397_));
OR2X2 OR2X2_896 ( .A(_abc_40319_new_n3294_), .B(_abc_40319_new_n3403_), .Y(_abc_40319_new_n3404_));
OR2X2 OR2X2_897 ( .A(_abc_40319_new_n3404_), .B(_abc_40319_new_n3401_), .Y(_abc_40319_new_n3405_));
OR2X2 OR2X2_898 ( .A(_abc_40319_new_n3397_), .B(_abc_40319_new_n3410_), .Y(_abc_40319_new_n3411_));
OR2X2 OR2X2_899 ( .A(_abc_40319_new_n3412_), .B(_abc_40319_new_n3101_), .Y(_abc_40319_new_n3413_));
OR2X2 OR2X2_9 ( .A(IR_REG_19_), .B(IR_REG_18_), .Y(_abc_40319_new_n604_));
OR2X2 OR2X2_90 ( .A(_abc_40319_new_n877_), .B(_abc_40319_new_n838_), .Y(_abc_40319_new_n878_));
OR2X2 OR2X2_900 ( .A(_abc_40319_new_n3414_), .B(_abc_40319_new_n3167_), .Y(_abc_40319_new_n3415_));
OR2X2 OR2X2_901 ( .A(_abc_40319_new_n3421_), .B(_abc_40319_new_n3417_), .Y(_abc_40319_new_n3422_));
OR2X2 OR2X2_902 ( .A(_abc_40319_new_n3426_), .B(_abc_40319_new_n3163_), .Y(_abc_40319_new_n3427_));
OR2X2 OR2X2_903 ( .A(_abc_40319_new_n3431_), .B(_abc_40319_new_n3435_), .Y(_abc_40319_new_n3436_));
OR2X2 OR2X2_904 ( .A(_abc_40319_new_n3436_), .B(_abc_40319_new_n3427_), .Y(_abc_40319_new_n3437_));
OR2X2 OR2X2_905 ( .A(_abc_40319_new_n3437_), .B(_abc_40319_new_n3423_), .Y(_abc_40319_new_n3438_));
OR2X2 OR2X2_906 ( .A(_abc_40319_new_n3416_), .B(_abc_40319_new_n3438_), .Y(_abc_40319_new_n3439_));
OR2X2 OR2X2_907 ( .A(_abc_40319_new_n3442_), .B(_abc_40319_new_n656_), .Y(_abc_40319_new_n3443_));
OR2X2 OR2X2_908 ( .A(_abc_40319_new_n3445_), .B(_abc_40319_new_n3267_), .Y(_abc_40319_new_n3446_));
OR2X2 OR2X2_909 ( .A(_abc_40319_new_n3446_), .B(_abc_40319_new_n3097_), .Y(_abc_40319_new_n3447_));
OR2X2 OR2X2_91 ( .A(_abc_40319_new_n879_), .B(_abc_40319_new_n880_), .Y(_abc_40319_new_n881_));
OR2X2 OR2X2_910 ( .A(_abc_40319_new_n3451_), .B(_abc_40319_new_n3453_), .Y(_abc_40319_new_n3454_));
OR2X2 OR2X2_911 ( .A(_abc_40319_new_n3078_), .B(_abc_40319_new_n3169_), .Y(_abc_40319_new_n3458_));
OR2X2 OR2X2_912 ( .A(_abc_40319_new_n3461_), .B(_abc_40319_new_n3160_), .Y(_abc_40319_new_n3462_));
OR2X2 OR2X2_913 ( .A(_abc_40319_new_n3460_), .B(_abc_40319_new_n3462_), .Y(_abc_40319_new_n3463_));
OR2X2 OR2X2_914 ( .A(_abc_40319_new_n3260_), .B(_abc_40319_new_n3197_), .Y(_abc_40319_new_n3469_));
OR2X2 OR2X2_915 ( .A(_abc_40319_new_n3488_), .B(_abc_40319_new_n3225_), .Y(_abc_40319_new_n3489_));
OR2X2 OR2X2_916 ( .A(_abc_40319_new_n3117_), .B(_abc_40319_new_n3136_), .Y(_abc_40319_new_n3490_));
OR2X2 OR2X2_917 ( .A(_abc_40319_new_n3491_), .B(_abc_40319_new_n3126_), .Y(_abc_40319_new_n3492_));
OR2X2 OR2X2_918 ( .A(_abc_40319_new_n3494_), .B(_abc_40319_new_n3131_), .Y(_abc_40319_new_n3495_));
OR2X2 OR2X2_919 ( .A(_abc_40319_new_n3214_), .B(_abc_40319_new_n3122_), .Y(_abc_40319_new_n3497_));
OR2X2 OR2X2_92 ( .A(_abc_40319_new_n884_), .B(_abc_40319_new_n885_), .Y(_abc_40319_new_n886_));
OR2X2 OR2X2_920 ( .A(_abc_40319_new_n3495_), .B(_abc_40319_new_n3500_), .Y(_abc_40319_new_n3501_));
OR2X2 OR2X2_921 ( .A(_abc_40319_new_n3502_), .B(_abc_40319_new_n3497_), .Y(_abc_40319_new_n3503_));
OR2X2 OR2X2_922 ( .A(_abc_40319_new_n3505_), .B(_abc_40319_new_n3210_), .Y(_abc_40319_new_n3506_));
OR2X2 OR2X2_923 ( .A(_abc_40319_new_n3508_), .B(_abc_40319_new_n3175_), .Y(_abc_40319_new_n3509_));
OR2X2 OR2X2_924 ( .A(_abc_40319_new_n3509_), .B(_abc_40319_new_n3512_), .Y(_abc_40319_new_n3513_));
OR2X2 OR2X2_925 ( .A(_abc_40319_new_n3514_), .B(_abc_40319_new_n3234_), .Y(_abc_40319_new_n3515_));
OR2X2 OR2X2_926 ( .A(_abc_40319_new_n3516_), .B(_abc_40319_new_n3141_), .Y(_abc_40319_new_n3517_));
OR2X2 OR2X2_927 ( .A(_abc_40319_new_n3518_), .B(_abc_40319_new_n3481_), .Y(_abc_40319_new_n3519_));
OR2X2 OR2X2_928 ( .A(_abc_40319_new_n3307_), .B(_abc_40319_new_n3230_), .Y(_abc_40319_new_n3522_));
OR2X2 OR2X2_929 ( .A(_abc_40319_new_n3525_), .B(_abc_40319_new_n3183_), .Y(_abc_40319_new_n3526_));
OR2X2 OR2X2_93 ( .A(_abc_40319_new_n817_), .B(_abc_40319_new_n886_), .Y(_abc_40319_new_n887_));
OR2X2 OR2X2_930 ( .A(_abc_40319_new_n3529_), .B(_abc_40319_new_n3475_), .Y(_abc_40319_new_n3530_));
OR2X2 OR2X2_931 ( .A(_abc_40319_new_n3531_), .B(_abc_40319_new_n3408_), .Y(_abc_40319_new_n3532_));
OR2X2 OR2X2_932 ( .A(_abc_40319_new_n3534_), .B(_abc_40319_new_n3281_), .Y(_abc_40319_new_n3535_));
OR2X2 OR2X2_933 ( .A(_abc_40319_new_n3536_), .B(_abc_40319_new_n3468_), .Y(_abc_40319_new_n3537_));
OR2X2 OR2X2_934 ( .A(_abc_40319_new_n3538_), .B(_abc_40319_new_n3247_), .Y(_abc_40319_new_n3539_));
OR2X2 OR2X2_935 ( .A(_abc_40319_new_n3540_), .B(_abc_40319_new_n3463_), .Y(_abc_40319_new_n3541_));
OR2X2 OR2X2_936 ( .A(_abc_40319_new_n3548_), .B(_abc_40319_new_n3546_), .Y(_abc_40319_new_n3549_));
OR2X2 OR2X2_937 ( .A(_abc_40319_new_n3549_), .B(_abc_40319_new_n3543_), .Y(_abc_40319_new_n3550_));
OR2X2 OR2X2_938 ( .A(_abc_40319_new_n3550_), .B(_abc_40319_new_n3455_), .Y(_abc_40319_new_n3551_));
OR2X2 OR2X2_939 ( .A(_abc_40319_new_n3551_), .B(_abc_40319_new_n3449_), .Y(_abc_40319_new_n3552_));
OR2X2 OR2X2_94 ( .A(_abc_40319_new_n905_), .B(_abc_40319_new_n892_), .Y(_abc_40319_new_n906_));
OR2X2 OR2X2_940 ( .A(_abc_40319_new_n3448_), .B(_abc_40319_new_n3552_), .Y(_abc_40319_new_n3553_));
OR2X2 OR2X2_941 ( .A(_abc_40319_new_n3559_), .B(_abc_40319_new_n617_), .Y(_abc_40319_new_n3560_));
OR2X2 OR2X2_942 ( .A(_abc_40319_new_n3560_), .B(_abc_40319_new_n614_), .Y(_abc_40319_new_n3561_));
OR2X2 OR2X2_943 ( .A(_abc_40319_new_n3558_), .B(_abc_40319_new_n3561_), .Y(_abc_40319_new_n3562_));
OR2X2 OR2X2_944 ( .A(_abc_40319_new_n3563_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n3564_));
OR2X2 OR2X2_945 ( .A(_abc_40319_new_n3554_), .B(_abc_40319_new_n3564_), .Y(n1186));
OR2X2 OR2X2_946 ( .A(IR_REG_0_), .B(REG1_REG_0_), .Y(_abc_40319_new_n3566_));
OR2X2 OR2X2_947 ( .A(IR_REG_0_), .B(REG2_REG_0_), .Y(_abc_40319_new_n3572_));
OR2X2 OR2X2_948 ( .A(_abc_40319_new_n3576_), .B(_abc_40319_new_n3571_), .Y(_abc_40319_new_n3577_));
OR2X2 OR2X2_949 ( .A(_abc_40319_new_n3577_), .B(_abc_40319_new_n3570_), .Y(_abc_40319_new_n3578_));
OR2X2 OR2X2_95 ( .A(_abc_40319_new_n903_), .B(_abc_40319_new_n909_), .Y(_abc_40319_new_n910_));
OR2X2 OR2X2_950 ( .A(_abc_40319_new_n3579_), .B(_abc_40319_new_n3580_), .Y(_abc_40319_new_n3581_));
OR2X2 OR2X2_951 ( .A(_abc_40319_new_n2363_), .B(_abc_40319_new_n1173_), .Y(_abc_40319_new_n3583_));
OR2X2 OR2X2_952 ( .A(n1341), .B(_abc_40319_new_n614_), .Y(_abc_40319_new_n3584_));
OR2X2 OR2X2_953 ( .A(_abc_40319_new_n3586_), .B(_abc_40319_new_n3583_), .Y(_abc_40319_new_n3587_));
OR2X2 OR2X2_954 ( .A(_abc_40319_new_n3587_), .B(_abc_40319_new_n3582_), .Y(n1054));
OR2X2 OR2X2_955 ( .A(_abc_40319_new_n886_), .B(_abc_40319_new_n3594_), .Y(_abc_40319_new_n3595_));
OR2X2 OR2X2_956 ( .A(_abc_40319_new_n3596_), .B(_abc_40319_new_n3597_), .Y(_abc_40319_new_n3598_));
OR2X2 OR2X2_957 ( .A(_abc_40319_new_n886_), .B(_abc_40319_new_n3606_), .Y(_abc_40319_new_n3607_));
OR2X2 OR2X2_958 ( .A(_abc_40319_new_n3596_), .B(_abc_40319_new_n3608_), .Y(_abc_40319_new_n3609_));
OR2X2 OR2X2_959 ( .A(_abc_40319_new_n3611_), .B(_abc_40319_new_n3612_), .Y(_abc_40319_new_n3613_));
OR2X2 OR2X2_96 ( .A(_abc_40319_new_n912_), .B(_abc_40319_new_n757_), .Y(_abc_40319_new_n913_));
OR2X2 OR2X2_960 ( .A(_abc_40319_new_n3613_), .B(_abc_40319_new_n3600_), .Y(_abc_40319_new_n3614_));
OR2X2 OR2X2_961 ( .A(_abc_40319_new_n3616_), .B(_abc_40319_new_n2168_), .Y(_abc_40319_new_n3617_));
OR2X2 OR2X2_962 ( .A(_abc_40319_new_n3617_), .B(_abc_40319_new_n3615_), .Y(n1050));
OR2X2 OR2X2_963 ( .A(_abc_40319_new_n3620_), .B(_abc_40319_new_n3577_), .Y(_abc_40319_new_n3621_));
OR2X2 OR2X2_964 ( .A(_abc_40319_new_n3623_), .B(_abc_40319_new_n2467_), .Y(_abc_40319_new_n3624_));
OR2X2 OR2X2_965 ( .A(_abc_40319_new_n3632_), .B(_abc_40319_new_n3590_), .Y(_abc_40319_new_n3633_));
OR2X2 OR2X2_966 ( .A(_abc_40319_new_n3631_), .B(_abc_40319_new_n3633_), .Y(_abc_40319_new_n3634_));
OR2X2 OR2X2_967 ( .A(_abc_40319_new_n3630_), .B(_abc_40319_new_n3635_), .Y(_abc_40319_new_n3636_));
OR2X2 OR2X2_968 ( .A(_abc_40319_new_n3645_), .B(_abc_40319_new_n3601_), .Y(_abc_40319_new_n3646_));
OR2X2 OR2X2_969 ( .A(_abc_40319_new_n3644_), .B(_abc_40319_new_n3647_), .Y(_abc_40319_new_n3648_));
OR2X2 OR2X2_97 ( .A(_abc_40319_new_n911_), .B(_abc_40319_new_n768_), .Y(_abc_40319_new_n914_));
OR2X2 OR2X2_970 ( .A(_abc_40319_new_n3643_), .B(_abc_40319_new_n3646_), .Y(_abc_40319_new_n3649_));
OR2X2 OR2X2_971 ( .A(_abc_40319_new_n3651_), .B(_abc_40319_new_n3652_), .Y(_abc_40319_new_n3653_));
OR2X2 OR2X2_972 ( .A(_abc_40319_new_n3653_), .B(_abc_40319_new_n3638_), .Y(_abc_40319_new_n3654_));
OR2X2 OR2X2_973 ( .A(_abc_40319_new_n3655_), .B(_abc_40319_new_n3656_), .Y(_abc_40319_new_n3657_));
OR2X2 OR2X2_974 ( .A(_abc_40319_new_n3624_), .B(_abc_40319_new_n3657_), .Y(_abc_40319_new_n3658_));
OR2X2 OR2X2_975 ( .A(_abc_40319_new_n3622_), .B(_abc_40319_new_n3658_), .Y(n1046));
OR2X2 OR2X2_976 ( .A(_abc_40319_new_n3661_), .B(_abc_40319_new_n3626_), .Y(_abc_40319_new_n3662_));
OR2X2 OR2X2_977 ( .A(_abc_40319_new_n3667_), .B(_abc_40319_new_n3660_), .Y(_abc_40319_new_n3668_));
OR2X2 OR2X2_978 ( .A(_abc_40319_new_n3670_), .B(_abc_40319_new_n3662_), .Y(_abc_40319_new_n3671_));
OR2X2 OR2X2_979 ( .A(_abc_40319_new_n3675_), .B(_abc_40319_new_n3641_), .Y(_abc_40319_new_n3676_));
OR2X2 OR2X2_98 ( .A(_abc_40319_new_n915_), .B(_abc_40319_new_n906_), .Y(_abc_40319_new_n916_));
OR2X2 OR2X2_980 ( .A(_abc_40319_new_n3684_), .B(_abc_40319_new_n3685_), .Y(_abc_40319_new_n3686_));
OR2X2 OR2X2_981 ( .A(_abc_40319_new_n3687_), .B(_abc_40319_new_n3688_), .Y(_abc_40319_new_n3689_));
OR2X2 OR2X2_982 ( .A(_abc_40319_new_n3689_), .B(_abc_40319_new_n3673_), .Y(_abc_40319_new_n3690_));
OR2X2 OR2X2_983 ( .A(_abc_40319_new_n3692_), .B(_abc_40319_new_n2064_), .Y(_abc_40319_new_n3693_));
OR2X2 OR2X2_984 ( .A(_abc_40319_new_n3693_), .B(_abc_40319_new_n3691_), .Y(n1042));
OR2X2 OR2X2_985 ( .A(_abc_40319_new_n3703_), .B(_abc_40319_new_n3701_), .Y(_abc_40319_new_n3704_));
OR2X2 OR2X2_986 ( .A(_abc_40319_new_n3706_), .B(_abc_40319_new_n3696_), .Y(_abc_40319_new_n3707_));
OR2X2 OR2X2_987 ( .A(_abc_40319_new_n3678_), .B(_abc_40319_new_n814_), .Y(_abc_40319_new_n3711_));
OR2X2 OR2X2_988 ( .A(_abc_40319_new_n3712_), .B(_abc_40319_new_n3714_), .Y(_abc_40319_new_n3715_));
OR2X2 OR2X2_989 ( .A(_abc_40319_new_n3715_), .B(_abc_40319_new_n3710_), .Y(_abc_40319_new_n3716_));
OR2X2 OR2X2_99 ( .A(_abc_40319_new_n919_), .B(_abc_40319_new_n918_), .Y(_abc_40319_new_n920_));
OR2X2 OR2X2_990 ( .A(_abc_40319_new_n3720_), .B(_abc_40319_new_n3717_), .Y(_abc_40319_new_n3721_));
OR2X2 OR2X2_991 ( .A(_abc_40319_new_n3723_), .B(_abc_40319_new_n3724_), .Y(_abc_40319_new_n3725_));
OR2X2 OR2X2_992 ( .A(_abc_40319_new_n3709_), .B(_abc_40319_new_n3725_), .Y(_abc_40319_new_n3726_));
OR2X2 OR2X2_993 ( .A(_abc_40319_new_n3695_), .B(_abc_40319_new_n3727_), .Y(_abc_40319_new_n3728_));
OR2X2 OR2X2_994 ( .A(_abc_40319_new_n3729_), .B(_abc_40319_new_n2334_), .Y(_abc_40319_new_n3730_));
OR2X2 OR2X2_995 ( .A(_abc_40319_new_n3728_), .B(_abc_40319_new_n3730_), .Y(_abc_40319_new_n3731_));
OR2X2 OR2X2_996 ( .A(_abc_40319_new_n3622_), .B(_abc_40319_new_n3731_), .Y(n1038));
OR2X2 OR2X2_997 ( .A(_abc_40319_new_n3741_), .B(_abc_40319_new_n685_), .Y(_abc_40319_new_n3742_));
OR2X2 OR2X2_998 ( .A(_abc_40319_new_n3740_), .B(_abc_40319_new_n684_), .Y(_abc_40319_new_n3743_));
OR2X2 OR2X2_999 ( .A(_abc_40319_new_n3756_), .B(_abc_40319_new_n3753_), .Y(_abc_40319_new_n3757_));


endmodule