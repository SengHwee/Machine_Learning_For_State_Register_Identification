module FSM(clk, reset, \codif[0] , \codif[1] , \codif[2] , \codif[3] , \codif[4] , \codif[5] , \codif[6] , \codif[7] , \codif[8] , \codif[9] , \codif[10] , \codif[11] , busy_mem, done_mem, aligned_mem, done_exec, is_exec, \W_R_mem[0] , \W_R_mem[1] , \wordsize_mem[0] , \wordsize_mem[1] , sign_mem, en_mem, enable_exec, enable_exec_mem, trap, enable_pc);
  output \W_R_mem[0] ;
  output \W_R_mem[1] ;
  wire W_R_mem_0__FF_INPUT;
  wire W_R_mem_1__FF_INPUT;
  wire _abc_818_n100;
  wire _abc_818_n103;
  wire _abc_818_n118;
  wire _abc_818_n66;
  wire _abc_818_n72;
  wire _abc_818_n89;
  wire _abc_818_n92;
  wire _abc_953_n100;
  wire _abc_953_n101;
  wire _abc_953_n102;
  wire _abc_953_n104;
  wire _abc_953_n105;
  wire _abc_953_n106;
  wire _abc_953_n107;
  wire _abc_953_n109;
  wire _abc_953_n110;
  wire _abc_953_n111;
  wire _abc_953_n112;
  wire _abc_953_n113;
  wire _abc_953_n114_1;
  wire _abc_953_n116;
  wire _abc_953_n117;
  wire _abc_953_n118;
  wire _abc_953_n119;
  wire _abc_953_n121;
  wire _abc_953_n123;
  wire _abc_953_n124_1;
  wire _abc_953_n125_1;
  wire _abc_953_n126;
  wire _abc_953_n127;
  wire _abc_953_n128;
  wire _abc_953_n129;
  wire _abc_953_n130;
  wire _abc_953_n131;
  wire _abc_953_n132;
  wire _abc_953_n133;
  wire _abc_953_n134_1;
  wire _abc_953_n135_1;
  wire _abc_953_n136;
  wire _abc_953_n137_1;
  wire _abc_953_n138;
  wire _abc_953_n139_1;
  wire _abc_953_n140;
  wire _abc_953_n142;
  wire _abc_953_n143;
  wire _abc_953_n144;
  wire _abc_953_n145;
  wire _abc_953_n146;
  wire _abc_953_n147_1;
  wire _abc_953_n148_1;
  wire _abc_953_n149;
  wire _abc_953_n150;
  wire _abc_953_n153;
  wire _abc_953_n154;
  wire _abc_953_n155;
  wire _abc_953_n156;
  wire _abc_953_n157_1;
  wire _abc_953_n158;
  wire _abc_953_n160;
  wire _abc_953_n161;
  wire _abc_953_n162;
  wire _abc_953_n163_1;
  wire _abc_953_n165;
  wire _abc_953_n167;
  wire _abc_953_n168;
  wire _abc_953_n169;
  wire _abc_953_n170;
  wire _abc_953_n171;
  wire _abc_953_n172;
  wire _abc_953_n173;
  wire _abc_953_n174;
  wire _abc_953_n175;
  wire _abc_953_n176;
  wire _abc_953_n177;
  wire _abc_953_n179;
  wire _abc_953_n180;
  wire _abc_953_n181;
  wire _abc_953_n183;
  wire _abc_953_n184;
  wire _abc_953_n185;
  wire _abc_953_n186;
  wire _abc_953_n187;
  wire _abc_953_n188;
  wire _abc_953_n49;
  wire _abc_953_n50;
  wire _abc_953_n51;
  wire _abc_953_n52_1;
  wire _abc_953_n53;
  wire _abc_953_n54;
  wire _abc_953_n55;
  wire _abc_953_n56;
  wire _abc_953_n57;
  wire _abc_953_n58;
  wire _abc_953_n59;
  wire _abc_953_n60_1;
  wire _abc_953_n61_1;
  wire _abc_953_n62;
  wire _abc_953_n63;
  wire _abc_953_n64;
  wire _abc_953_n65;
  wire _abc_953_n66;
  wire _abc_953_n67_1;
  wire _abc_953_n68;
  wire _abc_953_n69;
  wire _abc_953_n70;
  wire _abc_953_n71;
  wire _abc_953_n72;
  wire _abc_953_n73;
  wire _abc_953_n74;
  wire _abc_953_n75;
  wire _abc_953_n77_1;
  wire _abc_953_n78_1;
  wire _abc_953_n79;
  wire _abc_953_n80;
  wire _abc_953_n82_1;
  wire _abc_953_n83;
  wire _abc_953_n84;
  wire _abc_953_n85;
  wire _abc_953_n86_1;
  wire _abc_953_n87;
  wire _abc_953_n88;
  wire _abc_953_n89;
  wire _abc_953_n90;
  wire _abc_953_n91;
  wire _abc_953_n92_1;
  wire _abc_953_n93_1;
  wire _abc_953_n94_1;
  wire _abc_953_n95;
  wire _abc_953_n96_1;
  wire _abc_953_n97_1;
  wire _abc_953_n98_1;
  input aligned_mem;
  input busy_mem;
  input clk;
  input \codif[0] ;
  input \codif[10] ;
  input \codif[11] ;
  input \codif[1] ;
  input \codif[2] ;
  input \codif[3] ;
  input \codif[4] ;
  input \codif[5] ;
  input \codif[6] ;
  input \codif[7] ;
  input \codif[8] ;
  input \codif[9] ;
  input done_exec;
  input done_mem;
  output en_mem;
  wire en_mem_FF_INPUT;
  output enable_exec;
  wire enable_exec_FF_INPUT;
  output enable_exec_mem;
  wire enable_exec_mem_FF_INPUT;
  output enable_pc;
  wire enable_pc_aux;
  wire enable_pc_aux_FF_INPUT;
  wire enable_pc_fsm;
  wire enable_pc_fsm_FF_INPUT;
  input is_exec;
  input reset;
  output sign_mem;
  wire state_0_;
  wire state_1_;
  wire state_2_;
  wire state_3_;
  wire state_4_;
  wire state_5_;
  wire state_6_;
  output trap;
  wire trap_FF_INPUT;
  output \wordsize_mem[0] ;
  output \wordsize_mem[1] ;
  AND2X2 AND2X2_1 ( .A(_abc_953_n94_1), .B(state_3_), .Y(_abc_953_n95) );
  AND2X2 AND2X2_10 ( .A(_abc_953_n83), .B(_abc_953_n112), .Y(_abc_953_n113) );
  AND2X2 AND2X2_11 ( .A(_abc_953_n113), .B(_abc_953_n73), .Y(_abc_953_n114_1) );
  AND2X2 AND2X2_12 ( .A(_abc_953_n77_1), .B(en_mem), .Y(_abc_953_n116) );
  AND2X2 AND2X2_13 ( .A(_abc_953_n116), .B(state_0_), .Y(_abc_953_n117) );
  AND2X2 AND2X2_14 ( .A(_abc_953_n77_1), .B(state_5_), .Y(_abc_953_n118) );
  AND2X2 AND2X2_15 ( .A(_abc_953_n119), .B(_abc_953_n73), .Y(_abc_818_n118) );
  AND2X2 AND2X2_16 ( .A(_abc_953_n121), .B(enable_pc_fsm), .Y(enable_pc) );
  AND2X2 AND2X2_17 ( .A(_abc_953_n77_1), .B(\W_R_mem[0] ), .Y(_abc_953_n124_1) );
  AND2X2 AND2X2_18 ( .A(_abc_953_n124_1), .B(_abc_953_n123), .Y(_abc_953_n125_1) );
  AND2X2 AND2X2_19 ( .A(_abc_953_n128), .B(state_6_), .Y(_abc_953_n129) );
  AND2X2 AND2X2_2 ( .A(_abc_953_n88), .B(state_0_), .Y(_abc_953_n100) );
  AND2X2 AND2X2_20 ( .A(_abc_953_n130), .B(_abc_953_n126), .Y(_abc_953_n131) );
  AND2X2 AND2X2_21 ( .A(_abc_953_n132), .B(_abc_953_n73), .Y(_abc_953_n133) );
  AND2X2 AND2X2_22 ( .A(_abc_953_n134_1), .B(_abc_953_n136), .Y(_abc_953_n137_1) );
  AND2X2 AND2X2_23 ( .A(_abc_953_n138), .B(reset), .Y(_abc_953_n139_1) );
  AND2X2 AND2X2_24 ( .A(_abc_953_n139_1), .B(\W_R_mem[0] ), .Y(_abc_953_n140) );
  AND2X2 AND2X2_25 ( .A(_abc_953_n139_1), .B(\W_R_mem[1] ), .Y(_abc_953_n142) );
  AND2X2 AND2X2_26 ( .A(_abc_953_n143), .B(\W_R_mem[1] ), .Y(_abc_953_n144) );
  AND2X2 AND2X2_27 ( .A(_abc_953_n123), .B(_abc_953_n77_1), .Y(_abc_953_n145) );
  AND2X2 AND2X2_28 ( .A(_abc_953_n147_1), .B(_abc_953_n144), .Y(_abc_953_n148_1) );
  AND2X2 AND2X2_29 ( .A(_abc_953_n149), .B(_abc_953_n73), .Y(_abc_953_n150) );
  AND2X2 AND2X2_3 ( .A(done_mem), .B(state_5_), .Y(_abc_953_n101) );
  AND2X2 AND2X2_30 ( .A(_abc_953_n109), .B(state_4_), .Y(_abc_953_n153) );
  AND2X2 AND2X2_31 ( .A(_abc_953_n155), .B(_abc_953_n156), .Y(_abc_953_n157_1) );
  AND2X2 AND2X2_32 ( .A(reset), .B(enable_pc_fsm), .Y(enable_pc_aux_FF_INPUT) );
  AND2X2 AND2X2_33 ( .A(_abc_953_n158), .B(enable_pc_aux_FF_INPUT), .Y(_abc_953_n160) );
  AND2X2 AND2X2_34 ( .A(_abc_953_n161), .B(_abc_953_n73), .Y(_abc_953_n162) );
  AND2X2 AND2X2_35 ( .A(_abc_953_n154), .B(_abc_953_n163_1), .Y(enable_pc_fsm_FF_INPUT) );
  AND2X2 AND2X2_36 ( .A(_abc_953_n165), .B(reset), .Y(trap_FF_INPUT) );
  AND2X2 AND2X2_37 ( .A(reset), .B(enable_exec_mem), .Y(_abc_953_n172) );
  AND2X2 AND2X2_38 ( .A(_abc_953_n171), .B(_abc_953_n172), .Y(_abc_953_n173) );
  AND2X2 AND2X2_39 ( .A(_abc_953_n173), .B(_abc_953_n170), .Y(_abc_953_n174) );
  AND2X2 AND2X2_4 ( .A(_abc_953_n73), .B(_abc_953_n101), .Y(_abc_953_n102) );
  AND2X2 AND2X2_40 ( .A(_abc_953_n143), .B(_abc_953_n73), .Y(_abc_953_n175) );
  AND2X2 AND2X2_41 ( .A(_abc_953_n129), .B(_abc_953_n175), .Y(_abc_953_n176) );
  AND2X2 AND2X2_42 ( .A(_abc_953_n177), .B(_abc_953_n167), .Y(enable_exec_mem_FF_INPUT) );
  AND2X2 AND2X2_43 ( .A(_abc_953_n158), .B(reset), .Y(_abc_953_n179) );
  AND2X2 AND2X2_44 ( .A(_abc_953_n180), .B(enable_exec), .Y(_abc_953_n181) );
  AND2X2 AND2X2_45 ( .A(reset), .B(en_mem), .Y(_abc_953_n183) );
  AND2X2 AND2X2_46 ( .A(_abc_953_n138), .B(_abc_953_n183), .Y(_abc_953_n184) );
  AND2X2 AND2X2_47 ( .A(_abc_953_n135_1), .B(_abc_953_n90), .Y(_abc_953_n185) );
  AND2X2 AND2X2_48 ( .A(_abc_953_n116), .B(_abc_953_n123), .Y(_abc_953_n186) );
  AND2X2 AND2X2_49 ( .A(_abc_953_n187), .B(_abc_953_n73), .Y(_abc_953_n188) );
  AND2X2 AND2X2_5 ( .A(_abc_953_n104), .B(_abc_953_n84), .Y(_abc_953_n105) );
  AND2X2 AND2X2_50 ( .A(_abc_953_n50), .B(reset), .Y(_abc_953_n51) );
  AND2X2 AND2X2_51 ( .A(\codif[6] ), .B(\codif[4] ), .Y(_abc_953_n52_1) );
  AND2X2 AND2X2_52 ( .A(\codif[7] ), .B(\codif[5] ), .Y(_abc_953_n53) );
  AND2X2 AND2X2_53 ( .A(_abc_953_n52_1), .B(_abc_953_n53), .Y(_abc_953_n54) );
  AND2X2 AND2X2_54 ( .A(\codif[10] ), .B(\codif[11] ), .Y(_abc_953_n55) );
  AND2X2 AND2X2_55 ( .A(\codif[2] ), .B(\codif[3] ), .Y(_abc_953_n56) );
  AND2X2 AND2X2_56 ( .A(_abc_953_n55), .B(_abc_953_n56), .Y(_abc_953_n57) );
  AND2X2 AND2X2_57 ( .A(\codif[0] ), .B(\codif[1] ), .Y(_abc_953_n58) );
  AND2X2 AND2X2_58 ( .A(\codif[8] ), .B(\codif[9] ), .Y(_abc_953_n59) );
  AND2X2 AND2X2_59 ( .A(_abc_953_n58), .B(_abc_953_n59), .Y(_abc_953_n60_1) );
  AND2X2 AND2X2_6 ( .A(_abc_953_n90), .B(state_6_), .Y(_abc_953_n106) );
  AND2X2 AND2X2_60 ( .A(_abc_953_n57), .B(_abc_953_n60_1), .Y(_abc_953_n61_1) );
  AND2X2 AND2X2_61 ( .A(_abc_953_n65), .B(_abc_953_n69), .Y(_abc_953_n70) );
  AND2X2 AND2X2_62 ( .A(_abc_953_n71), .B(_abc_953_n54), .Y(_abc_953_n72) );
  AND2X2 AND2X2_63 ( .A(reset), .B(aligned_mem), .Y(_abc_953_n73) );
  AND2X2 AND2X2_64 ( .A(_abc_953_n73), .B(state_4_), .Y(_abc_953_n74) );
  AND2X2 AND2X2_65 ( .A(_abc_953_n72), .B(_abc_953_n74), .Y(_abc_953_n75) );
  AND2X2 AND2X2_66 ( .A(_abc_953_n73), .B(_abc_953_n77_1), .Y(_abc_953_n78_1) );
  AND2X2 AND2X2_67 ( .A(state_6_), .B(en_mem), .Y(_abc_953_n79) );
  AND2X2 AND2X2_68 ( .A(_abc_953_n80), .B(_abc_953_n78_1), .Y(_abc_818_n72) );
  AND2X2 AND2X2_69 ( .A(_abc_953_n73), .B(state_2_), .Y(_abc_953_n84) );
  AND2X2 AND2X2_7 ( .A(_abc_953_n106), .B(_abc_953_n73), .Y(_abc_953_n107) );
  AND2X2 AND2X2_70 ( .A(_abc_953_n84), .B(done_exec), .Y(_abc_953_n85) );
  AND2X2 AND2X2_71 ( .A(_abc_953_n83), .B(_abc_953_n85), .Y(_abc_953_n86_1) );
  AND2X2 AND2X2_72 ( .A(en_mem), .B(done_mem), .Y(_abc_953_n87) );
  AND2X2 AND2X2_73 ( .A(_abc_953_n73), .B(_abc_953_n87), .Y(_abc_953_n88) );
  AND2X2 AND2X2_74 ( .A(_abc_953_n88), .B(state_6_), .Y(_abc_953_n89) );
  AND2X2 AND2X2_75 ( .A(_abc_953_n90), .B(state_0_), .Y(_abc_953_n91) );
  AND2X2 AND2X2_76 ( .A(_abc_953_n91), .B(_abc_953_n73), .Y(_abc_953_n92_1) );
  AND2X2 AND2X2_77 ( .A(aligned_mem), .B(done_mem), .Y(_abc_953_n94_1) );
  AND2X2 AND2X2_8 ( .A(_abc_953_n109), .B(_abc_953_n74), .Y(_abc_953_n110) );
  AND2X2 AND2X2_9 ( .A(_abc_953_n111), .B(state_2_), .Y(_abc_953_n112) );
  DFFPOSX1 DFFPOSX1_1 ( .CLK(clk), .D(_abc_818_n89), .Q(state_0_) );
  DFFPOSX1 DFFPOSX1_10 ( .CLK(clk), .D(en_mem_FF_INPUT), .Q(en_mem) );
  DFFPOSX1 DFFPOSX1_11 ( .CLK(clk), .D(enable_exec_FF_INPUT), .Q(enable_exec) );
  DFFPOSX1 DFFPOSX1_12 ( .CLK(clk), .D(enable_exec_mem_FF_INPUT), .Q(enable_exec_mem) );
  DFFPOSX1 DFFPOSX1_13 ( .CLK(clk), .D(trap_FF_INPUT), .Q(trap) );
  DFFPOSX1 DFFPOSX1_14 ( .CLK(clk), .D(enable_pc_fsm_FF_INPUT), .Q(enable_pc_fsm) );
  DFFPOSX1 DFFPOSX1_15 ( .CLK(clk), .D(enable_pc_aux_FF_INPUT), .Q(enable_pc_aux) );
  DFFPOSX1 DFFPOSX1_2 ( .CLK(clk), .D(_abc_818_n66), .Q(state_1_) );
  DFFPOSX1 DFFPOSX1_3 ( .CLK(clk), .D(_abc_818_n103), .Q(state_2_) );
  DFFPOSX1 DFFPOSX1_4 ( .CLK(clk), .D(_abc_818_n72), .Q(state_3_) );
  DFFPOSX1 DFFPOSX1_5 ( .CLK(clk), .D(_abc_818_n92), .Q(state_4_) );
  DFFPOSX1 DFFPOSX1_6 ( .CLK(clk), .D(_abc_818_n118), .Q(state_5_) );
  DFFPOSX1 DFFPOSX1_7 ( .CLK(clk), .D(_abc_818_n100), .Q(state_6_) );
  DFFPOSX1 DFFPOSX1_8 ( .CLK(clk), .D(W_R_mem_0__FF_INPUT), .Q(\W_R_mem[0] ) );
  DFFPOSX1 DFFPOSX1_9 ( .CLK(clk), .D(W_R_mem_1__FF_INPUT), .Q(\W_R_mem[1] ) );
  INVX1 INVX1_1 ( .A(_abc_953_n83), .Y(_abc_953_n104) );
  INVX1 INVX1_10 ( .A(state_4_), .Y(_abc_953_n155) );
  INVX1 INVX1_11 ( .A(state_2_), .Y(_abc_953_n156) );
  INVX1 INVX1_12 ( .A(state_6_), .Y(_abc_953_n168) );
  INVX1 INVX1_13 ( .A(_abc_953_n95), .Y(_abc_953_n171) );
  INVX1 INVX1_14 ( .A(_abc_953_n58), .Y(_abc_953_n62) );
  INVX1 INVX1_15 ( .A(_abc_953_n64), .Y(_abc_953_n65) );
  INVX1 INVX1_16 ( .A(_abc_953_n68), .Y(_abc_953_n69) );
  INVX1 INVX1_17 ( .A(reset), .Y(_abc_953_n93_1) );
  INVX1 INVX1_2 ( .A(_abc_953_n72), .Y(_abc_953_n109) );
  INVX1 INVX1_3 ( .A(done_exec), .Y(_abc_953_n111) );
  INVX1 INVX1_4 ( .A(enable_pc_aux), .Y(_abc_953_n121) );
  INVX1 INVX1_5 ( .A(\codif[5] ), .Y(_abc_953_n127) );
  INVX1 INVX1_6 ( .A(_abc_953_n123), .Y(_abc_953_n134_1) );
  INVX1 INVX1_7 ( .A(_abc_953_n135_1), .Y(_abc_953_n136) );
  INVX1 INVX1_8 ( .A(_abc_953_n87), .Y(_abc_953_n143) );
  INVX1 INVX1_9 ( .A(\codif[9] ), .Y(sign_mem) );
  INVX2 INVX2_1 ( .A(aligned_mem), .Y(_abc_953_n49) );
  INVX2 INVX2_2 ( .A(done_mem), .Y(_abc_953_n77_1) );
  INVX2 INVX2_3 ( .A(en_mem), .Y(_abc_953_n90) );
  OR2X2 OR2X2_1 ( .A(_abc_953_n95), .B(_abc_953_n93_1), .Y(_abc_953_n96_1) );
  OR2X2 OR2X2_10 ( .A(_abc_953_n124_1), .B(_abc_953_n90), .Y(_abc_953_n126) );
  OR2X2 OR2X2_11 ( .A(_abc_953_n127), .B(en_mem), .Y(_abc_953_n128) );
  OR2X2 OR2X2_12 ( .A(_abc_953_n129), .B(state_0_), .Y(_abc_953_n130) );
  OR2X2 OR2X2_13 ( .A(_abc_953_n131), .B(_abc_953_n125_1), .Y(_abc_953_n132) );
  OR2X2 OR2X2_14 ( .A(state_6_), .B(state_0_), .Y(_abc_953_n135_1) );
  OR2X2 OR2X2_15 ( .A(_abc_953_n137_1), .B(_abc_953_n49), .Y(_abc_953_n138) );
  OR2X2 OR2X2_16 ( .A(_abc_953_n133), .B(_abc_953_n140), .Y(W_R_mem_0__FF_INPUT) );
  OR2X2 OR2X2_17 ( .A(_abc_953_n79), .B(state_0_), .Y(_abc_953_n146) );
  OR2X2 OR2X2_18 ( .A(_abc_953_n145), .B(_abc_953_n146), .Y(_abc_953_n147_1) );
  OR2X2 OR2X2_19 ( .A(_abc_953_n148_1), .B(_abc_953_n91), .Y(_abc_953_n149) );
  OR2X2 OR2X2_2 ( .A(_abc_953_n96_1), .B(_abc_953_n92_1), .Y(_abc_953_n97_1) );
  OR2X2 OR2X2_20 ( .A(_abc_953_n150), .B(_abc_953_n142), .Y(W_R_mem_1__FF_INPUT) );
  OR2X2 OR2X2_21 ( .A(_abc_953_n153), .B(enable_pc_fsm), .Y(_abc_953_n154) );
  OR2X2 OR2X2_22 ( .A(_abc_953_n157_1), .B(_abc_953_n49), .Y(_abc_953_n158) );
  OR2X2 OR2X2_23 ( .A(_abc_953_n113), .B(state_4_), .Y(_abc_953_n161) );
  OR2X2 OR2X2_24 ( .A(_abc_953_n162), .B(_abc_953_n160), .Y(_abc_953_n163_1) );
  OR2X2 OR2X2_25 ( .A(_abc_953_n50), .B(trap), .Y(_abc_953_n165) );
  OR2X2 OR2X2_26 ( .A(_abc_953_n90), .B(enable_exec_mem), .Y(_abc_953_n167) );
  OR2X2 OR2X2_27 ( .A(_abc_953_n49), .B(state_3_), .Y(_abc_953_n169) );
  OR2X2 OR2X2_28 ( .A(_abc_953_n169), .B(_abc_953_n168), .Y(_abc_953_n170) );
  OR2X2 OR2X2_29 ( .A(_abc_953_n174), .B(_abc_953_n176), .Y(_abc_953_n177) );
  OR2X2 OR2X2_3 ( .A(_abc_953_n97_1), .B(_abc_953_n89), .Y(_abc_953_n98_1) );
  OR2X2 OR2X2_30 ( .A(_abc_953_n162), .B(_abc_953_n179), .Y(_abc_953_n180) );
  OR2X2 OR2X2_31 ( .A(_abc_953_n181), .B(_abc_953_n110), .Y(enable_exec_FF_INPUT) );
  OR2X2 OR2X2_32 ( .A(_abc_953_n186), .B(_abc_953_n185), .Y(_abc_953_n187) );
  OR2X2 OR2X2_33 ( .A(_abc_953_n184), .B(_abc_953_n188), .Y(en_mem_FF_INPUT) );
  OR2X2 OR2X2_34 ( .A(_abc_953_n49), .B(state_1_), .Y(_abc_953_n50) );
  OR2X2 OR2X2_35 ( .A(\codif[2] ), .B(\codif[3] ), .Y(_abc_953_n63) );
  OR2X2 OR2X2_36 ( .A(_abc_953_n62), .B(_abc_953_n63), .Y(_abc_953_n64) );
  OR2X2 OR2X2_37 ( .A(\codif[8] ), .B(\codif[9] ), .Y(_abc_953_n66) );
  OR2X2 OR2X2_38 ( .A(\codif[10] ), .B(\codif[11] ), .Y(_abc_953_n67_1) );
  OR2X2 OR2X2_39 ( .A(_abc_953_n66), .B(_abc_953_n67_1), .Y(_abc_953_n68) );
  OR2X2 OR2X2_4 ( .A(_abc_953_n98_1), .B(_abc_953_n86_1), .Y(_abc_818_n89) );
  OR2X2 OR2X2_40 ( .A(_abc_953_n70), .B(_abc_953_n61_1), .Y(_abc_953_n71) );
  OR2X2 OR2X2_41 ( .A(_abc_953_n75), .B(_abc_953_n51), .Y(_abc_818_n66) );
  OR2X2 OR2X2_42 ( .A(_abc_953_n79), .B(state_3_), .Y(_abc_953_n80) );
  OR2X2 OR2X2_43 ( .A(\codif[6] ), .B(\codif[4] ), .Y(_abc_953_n82_1) );
  OR2X2 OR2X2_44 ( .A(_abc_953_n64), .B(_abc_953_n82_1), .Y(_abc_953_n83) );
  OR2X2 OR2X2_5 ( .A(_abc_953_n100), .B(_abc_953_n102), .Y(_abc_818_n92) );
  OR2X2 OR2X2_6 ( .A(_abc_953_n105), .B(_abc_953_n107), .Y(_abc_818_n100) );
  OR2X2 OR2X2_7 ( .A(_abc_953_n110), .B(_abc_953_n114_1), .Y(_abc_818_n103) );
  OR2X2 OR2X2_8 ( .A(_abc_953_n117), .B(_abc_953_n118), .Y(_abc_953_n119) );
  OR2X2 OR2X2_9 ( .A(state_3_), .B(state_5_), .Y(_abc_953_n123) );
  assign \wordsize_mem[0]  = \codif[7] ;
  assign \wordsize_mem[1]  = \codif[8] ;
endmodule