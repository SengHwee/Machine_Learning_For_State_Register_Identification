module sha1_core(clk, reset_n, init, next, \block[0] , \block[1] , \block[2] , \block[3] , \block[4] , \block[5] , \block[6] , \block[7] , \block[8] , \block[9] , \block[10] , \block[11] , \block[12] , \block[13] , \block[14] , \block[15] , \block[16] , \block[17] , \block[18] , \block[19] , \block[20] , \block[21] , \block[22] , \block[23] , \block[24] , \block[25] , \block[26] , \block[27] , \block[28] , \block[29] , \block[30] , \block[31] , \block[32] , \block[33] , \block[34] , \block[35] , \block[36] , \block[37] , \block[38] , \block[39] , \block[40] , \block[41] , \block[42] , \block[43] , \block[44] , \block[45] , \block[46] , \block[47] , \block[48] , \block[49] , \block[50] , \block[51] , \block[52] , \block[53] , \block[54] , \block[55] , \block[56] , \block[57] , \block[58] , \block[59] , \block[60] , \block[61] , \block[62] , \block[63] , \block[64] , \block[65] , \block[66] , \block[67] , \block[68] , \block[69] , \block[70] , \block[71] , \block[72] , \block[73] , \block[74] , \block[75] , \block[76] , \block[77] , \block[78] , \block[79] , \block[80] , \block[81] , \block[82] , \block[83] , \block[84] , \block[85] , \block[86] , \block[87] , \block[88] , \block[89] , \block[90] , \block[91] , \block[92] , \block[93] , \block[94] , \block[95] , \block[96] , \block[97] , \block[98] , \block[99] , \block[100] , \block[101] , \block[102] , \block[103] , \block[104] , \block[105] , \block[106] , \block[107] , \block[108] , \block[109] , \block[110] , \block[111] , \block[112] , \block[113] , \block[114] , \block[115] , \block[116] , \block[117] , \block[118] , \block[119] , \block[120] , \block[121] , \block[122] , \block[123] , \block[124] , \block[125] , \block[126] , \block[127] , \block[128] , \block[129] , \block[130] , \block[131] , \block[132] , \block[133] , \block[134] , \block[135] , \block[136] , \block[137] , \block[138] , \block[139] , \block[140] , \block[141] , \block[142] , \block[143] , \block[144] , \block[145] , \block[146] , \block[147] , \block[148] , \block[149] , \block[150] , \block[151] , \block[152] , \block[153] , \block[154] , \block[155] , \block[156] , \block[157] , \block[158] , \block[159] , \block[160] , \block[161] , \block[162] , \block[163] , \block[164] , \block[165] , \block[166] , \block[167] , \block[168] , \block[169] , \block[170] , \block[171] , \block[172] , \block[173] , \block[174] , \block[175] , \block[176] , \block[177] , \block[178] , \block[179] , \block[180] , \block[181] , \block[182] , \block[183] , \block[184] , \block[185] , \block[186] , \block[187] , \block[188] , \block[189] , \block[190] , \block[191] , \block[192] , \block[193] , \block[194] , \block[195] , \block[196] , \block[197] , \block[198] , \block[199] , \block[200] , \block[201] , \block[202] , \block[203] , \block[204] , \block[205] , \block[206] , \block[207] , \block[208] , \block[209] , \block[210] , \block[211] , \block[212] , \block[213] , \block[214] , \block[215] , \block[216] , \block[217] , \block[218] , \block[219] , \block[220] , \block[221] , \block[222] , \block[223] , \block[224] , \block[225] , \block[226] , \block[227] , \block[228] , \block[229] , \block[230] , \block[231] , \block[232] , \block[233] , \block[234] , \block[235] , \block[236] , \block[237] , \block[238] , \block[239] , \block[240] , \block[241] , \block[242] , \block[243] , \block[244] , \block[245] , \block[246] , \block[247] , \block[248] , \block[249] , \block[250] , \block[251] , \block[252] , \block[253] , \block[254] , \block[255] , \block[256] , \block[257] , \block[258] , \block[259] , \block[260] , \block[261] , \block[262] , \block[263] , \block[264] , \block[265] , \block[266] , \block[267] , \block[268] , \block[269] , \block[270] , \block[271] , \block[272] , \block[273] , \block[274] , \block[275] , \block[276] , \block[277] , \block[278] , \block[279] , \block[280] , \block[281] , \block[282] , \block[283] , \block[284] , \block[285] , \block[286] , \block[287] , \block[288] , \block[289] , \block[290] , \block[291] , \block[292] , \block[293] , \block[294] , \block[295] , \block[296] , \block[297] , \block[298] , \block[299] , \block[300] , \block[301] , \block[302] , \block[303] , \block[304] , \block[305] , \block[306] , \block[307] , \block[308] , \block[309] , \block[310] , \block[311] , \block[312] , \block[313] , \block[314] , \block[315] , \block[316] , \block[317] , \block[318] , \block[319] , \block[320] , \block[321] , \block[322] , \block[323] , \block[324] , \block[325] , \block[326] , \block[327] , \block[328] , \block[329] , \block[330] , \block[331] , \block[332] , \block[333] , \block[334] , \block[335] , \block[336] , \block[337] , \block[338] , \block[339] , \block[340] , \block[341] , \block[342] , \block[343] , \block[344] , \block[345] , \block[346] , \block[347] , \block[348] , \block[349] , \block[350] , \block[351] , \block[352] , \block[353] , \block[354] , \block[355] , \block[356] , \block[357] , \block[358] , \block[359] , \block[360] , \block[361] , \block[362] , \block[363] , \block[364] , \block[365] , \block[366] , \block[367] , \block[368] , \block[369] , \block[370] , \block[371] , \block[372] , \block[373] , \block[374] , \block[375] , \block[376] , \block[377] , \block[378] , \block[379] , \block[380] , \block[381] , \block[382] , \block[383] , \block[384] , \block[385] , \block[386] , \block[387] , \block[388] , \block[389] , \block[390] , \block[391] , \block[392] , \block[393] , \block[394] , \block[395] , \block[396] , \block[397] , \block[398] , \block[399] , \block[400] , \block[401] , \block[402] , \block[403] , \block[404] , \block[405] , \block[406] , \block[407] , \block[408] , \block[409] , \block[410] , \block[411] , \block[412] , \block[413] , \block[414] , \block[415] , \block[416] , \block[417] , \block[418] , \block[419] , \block[420] , \block[421] , \block[422] , \block[423] , \block[424] , \block[425] , \block[426] , \block[427] , \block[428] , \block[429] , \block[430] , \block[431] , \block[432] , \block[433] , \block[434] , \block[435] , \block[436] , \block[437] , \block[438] , \block[439] , \block[440] , \block[441] , \block[442] , \block[443] , \block[444] , \block[445] , \block[446] , \block[447] , \block[448] , \block[449] , \block[450] , \block[451] , \block[452] , \block[453] , \block[454] , \block[455] , \block[456] , \block[457] , \block[458] , \block[459] , \block[460] , \block[461] , \block[462] , \block[463] , \block[464] , \block[465] , \block[466] , \block[467] , \block[468] , \block[469] , \block[470] , \block[471] , \block[472] , \block[473] , \block[474] , \block[475] , \block[476] , \block[477] , \block[478] , \block[479] , \block[480] , \block[481] , \block[482] , \block[483] , \block[484] , \block[485] , \block[486] , \block[487] , \block[488] , \block[489] , \block[490] , \block[491] , \block[492] , \block[493] , \block[494] , \block[495] , \block[496] , \block[497] , \block[498] , \block[499] , \block[500] , \block[501] , \block[502] , \block[503] , \block[504] , \block[505] , \block[506] , \block[507] , \block[508] , \block[509] , \block[510] , \block[511] , ready, \digest[0] , \digest[1] , \digest[2] , \digest[3] , \digest[4] , \digest[5] , \digest[6] , \digest[7] , \digest[8] , \digest[9] , \digest[10] , \digest[11] , \digest[12] , \digest[13] , \digest[14] , \digest[15] , \digest[16] , \digest[17] , \digest[18] , \digest[19] , \digest[20] , \digest[21] , \digest[22] , \digest[23] , \digest[24] , \digest[25] , \digest[26] , \digest[27] , \digest[28] , \digest[29] , \digest[30] , \digest[31] , \digest[32] , \digest[33] , \digest[34] , \digest[35] , \digest[36] , \digest[37] , \digest[38] , \digest[39] , \digest[40] , \digest[41] , \digest[42] , \digest[43] , \digest[44] , \digest[45] , \digest[46] , \digest[47] , \digest[48] , \digest[49] , \digest[50] , \digest[51] , \digest[52] , \digest[53] , \digest[54] , \digest[55] , \digest[56] , \digest[57] , \digest[58] , \digest[59] , \digest[60] , \digest[61] , \digest[62] , \digest[63] , \digest[64] , \digest[65] , \digest[66] , \digest[67] , \digest[68] , \digest[69] , \digest[70] , \digest[71] , \digest[72] , \digest[73] , \digest[74] , \digest[75] , \digest[76] , \digest[77] , \digest[78] , \digest[79] , \digest[80] , \digest[81] , \digest[82] , \digest[83] , \digest[84] , \digest[85] , \digest[86] , \digest[87] , \digest[88] , \digest[89] , \digest[90] , \digest[91] , \digest[92] , \digest[93] , \digest[94] , \digest[95] , \digest[96] , \digest[97] , \digest[98] , \digest[99] , \digest[100] , \digest[101] , \digest[102] , \digest[103] , \digest[104] , \digest[105] , \digest[106] , \digest[107] , \digest[108] , \digest[109] , \digest[110] , \digest[111] , \digest[112] , \digest[113] , \digest[114] , \digest[115] , \digest[116] , \digest[117] , \digest[118] , \digest[119] , \digest[120] , \digest[121] , \digest[122] , \digest[123] , \digest[124] , \digest[125] , \digest[126] , \digest[127] , \digest[128] , \digest[129] , \digest[130] , \digest[131] , \digest[132] , \digest[133] , \digest[134] , \digest[135] , \digest[136] , \digest[137] , \digest[138] , \digest[139] , \digest[140] , \digest[141] , \digest[142] , \digest[143] , \digest[144] , \digest[145] , \digest[146] , \digest[147] , \digest[148] , \digest[149] , \digest[150] , \digest[151] , \digest[152] , \digest[153] , \digest[154] , \digest[155] , \digest[156] , \digest[157] , \digest[158] , \digest[159] , digest_valid);

wire _0H0_reg_31_0__0_; 
wire _0H0_reg_31_0__10_; 
wire _0H0_reg_31_0__11_; 
wire _0H0_reg_31_0__12_; 
wire _0H0_reg_31_0__13_; 
wire _0H0_reg_31_0__14_; 
wire _0H0_reg_31_0__15_; 
wire _0H0_reg_31_0__16_; 
wire _0H0_reg_31_0__17_; 
wire _0H0_reg_31_0__18_; 
wire _0H0_reg_31_0__19_; 
wire _0H0_reg_31_0__1_; 
wire _0H0_reg_31_0__20_; 
wire _0H0_reg_31_0__21_; 
wire _0H0_reg_31_0__22_; 
wire _0H0_reg_31_0__23_; 
wire _0H0_reg_31_0__24_; 
wire _0H0_reg_31_0__25_; 
wire _0H0_reg_31_0__26_; 
wire _0H0_reg_31_0__27_; 
wire _0H0_reg_31_0__28_; 
wire _0H0_reg_31_0__29_; 
wire _0H0_reg_31_0__2_; 
wire _0H0_reg_31_0__30_; 
wire _0H0_reg_31_0__31_; 
wire _0H0_reg_31_0__3_; 
wire _0H0_reg_31_0__4_; 
wire _0H0_reg_31_0__5_; 
wire _0H0_reg_31_0__6_; 
wire _0H0_reg_31_0__7_; 
wire _0H0_reg_31_0__8_; 
wire _0H0_reg_31_0__9_; 
wire _0H1_reg_31_0__0_; 
wire _0H1_reg_31_0__10_; 
wire _0H1_reg_31_0__11_; 
wire _0H1_reg_31_0__12_; 
wire _0H1_reg_31_0__13_; 
wire _0H1_reg_31_0__14_; 
wire _0H1_reg_31_0__15_; 
wire _0H1_reg_31_0__16_; 
wire _0H1_reg_31_0__17_; 
wire _0H1_reg_31_0__18_; 
wire _0H1_reg_31_0__19_; 
wire _0H1_reg_31_0__1_; 
wire _0H1_reg_31_0__20_; 
wire _0H1_reg_31_0__21_; 
wire _0H1_reg_31_0__22_; 
wire _0H1_reg_31_0__23_; 
wire _0H1_reg_31_0__24_; 
wire _0H1_reg_31_0__25_; 
wire _0H1_reg_31_0__26_; 
wire _0H1_reg_31_0__27_; 
wire _0H1_reg_31_0__28_; 
wire _0H1_reg_31_0__29_; 
wire _0H1_reg_31_0__2_; 
wire _0H1_reg_31_0__30_; 
wire _0H1_reg_31_0__31_; 
wire _0H1_reg_31_0__3_; 
wire _0H1_reg_31_0__4_; 
wire _0H1_reg_31_0__5_; 
wire _0H1_reg_31_0__6_; 
wire _0H1_reg_31_0__7_; 
wire _0H1_reg_31_0__8_; 
wire _0H1_reg_31_0__9_; 
wire _0H2_reg_31_0__0_; 
wire _0H2_reg_31_0__10_; 
wire _0H2_reg_31_0__11_; 
wire _0H2_reg_31_0__12_; 
wire _0H2_reg_31_0__13_; 
wire _0H2_reg_31_0__14_; 
wire _0H2_reg_31_0__15_; 
wire _0H2_reg_31_0__16_; 
wire _0H2_reg_31_0__17_; 
wire _0H2_reg_31_0__18_; 
wire _0H2_reg_31_0__19_; 
wire _0H2_reg_31_0__1_; 
wire _0H2_reg_31_0__20_; 
wire _0H2_reg_31_0__21_; 
wire _0H2_reg_31_0__22_; 
wire _0H2_reg_31_0__23_; 
wire _0H2_reg_31_0__24_; 
wire _0H2_reg_31_0__25_; 
wire _0H2_reg_31_0__26_; 
wire _0H2_reg_31_0__27_; 
wire _0H2_reg_31_0__28_; 
wire _0H2_reg_31_0__29_; 
wire _0H2_reg_31_0__2_; 
wire _0H2_reg_31_0__30_; 
wire _0H2_reg_31_0__31_; 
wire _0H2_reg_31_0__3_; 
wire _0H2_reg_31_0__4_; 
wire _0H2_reg_31_0__5_; 
wire _0H2_reg_31_0__6_; 
wire _0H2_reg_31_0__7_; 
wire _0H2_reg_31_0__8_; 
wire _0H2_reg_31_0__9_; 
wire _0H3_reg_31_0__0_; 
wire _0H3_reg_31_0__10_; 
wire _0H3_reg_31_0__11_; 
wire _0H3_reg_31_0__12_; 
wire _0H3_reg_31_0__13_; 
wire _0H3_reg_31_0__14_; 
wire _0H3_reg_31_0__15_; 
wire _0H3_reg_31_0__16_; 
wire _0H3_reg_31_0__17_; 
wire _0H3_reg_31_0__18_; 
wire _0H3_reg_31_0__19_; 
wire _0H3_reg_31_0__1_; 
wire _0H3_reg_31_0__20_; 
wire _0H3_reg_31_0__21_; 
wire _0H3_reg_31_0__22_; 
wire _0H3_reg_31_0__23_; 
wire _0H3_reg_31_0__24_; 
wire _0H3_reg_31_0__25_; 
wire _0H3_reg_31_0__26_; 
wire _0H3_reg_31_0__27_; 
wire _0H3_reg_31_0__28_; 
wire _0H3_reg_31_0__29_; 
wire _0H3_reg_31_0__2_; 
wire _0H3_reg_31_0__30_; 
wire _0H3_reg_31_0__31_; 
wire _0H3_reg_31_0__3_; 
wire _0H3_reg_31_0__4_; 
wire _0H3_reg_31_0__5_; 
wire _0H3_reg_31_0__6_; 
wire _0H3_reg_31_0__7_; 
wire _0H3_reg_31_0__8_; 
wire _0H3_reg_31_0__9_; 
wire _0H4_reg_31_0__0_; 
wire _0H4_reg_31_0__10_; 
wire _0H4_reg_31_0__11_; 
wire _0H4_reg_31_0__12_; 
wire _0H4_reg_31_0__13_; 
wire _0H4_reg_31_0__14_; 
wire _0H4_reg_31_0__15_; 
wire _0H4_reg_31_0__16_; 
wire _0H4_reg_31_0__17_; 
wire _0H4_reg_31_0__18_; 
wire _0H4_reg_31_0__19_; 
wire _0H4_reg_31_0__1_; 
wire _0H4_reg_31_0__20_; 
wire _0H4_reg_31_0__21_; 
wire _0H4_reg_31_0__22_; 
wire _0H4_reg_31_0__23_; 
wire _0H4_reg_31_0__24_; 
wire _0H4_reg_31_0__25_; 
wire _0H4_reg_31_0__26_; 
wire _0H4_reg_31_0__27_; 
wire _0H4_reg_31_0__28_; 
wire _0H4_reg_31_0__29_; 
wire _0H4_reg_31_0__2_; 
wire _0H4_reg_31_0__30_; 
wire _0H4_reg_31_0__31_; 
wire _0H4_reg_31_0__3_; 
wire _0H4_reg_31_0__4_; 
wire _0H4_reg_31_0__5_; 
wire _0H4_reg_31_0__6_; 
wire _0H4_reg_31_0__7_; 
wire _0H4_reg_31_0__8_; 
wire _0H4_reg_31_0__9_; 
wire _0a_reg_31_0__0_; 
wire _0a_reg_31_0__10_; 
wire _0a_reg_31_0__11_; 
wire _0a_reg_31_0__12_; 
wire _0a_reg_31_0__13_; 
wire _0a_reg_31_0__14_; 
wire _0a_reg_31_0__15_; 
wire _0a_reg_31_0__16_; 
wire _0a_reg_31_0__17_; 
wire _0a_reg_31_0__18_; 
wire _0a_reg_31_0__19_; 
wire _0a_reg_31_0__1_; 
wire _0a_reg_31_0__20_; 
wire _0a_reg_31_0__21_; 
wire _0a_reg_31_0__22_; 
wire _0a_reg_31_0__23_; 
wire _0a_reg_31_0__24_; 
wire _0a_reg_31_0__25_; 
wire _0a_reg_31_0__26_; 
wire _0a_reg_31_0__27_; 
wire _0a_reg_31_0__28_; 
wire _0a_reg_31_0__29_; 
wire _0a_reg_31_0__2_; 
wire _0a_reg_31_0__30_; 
wire _0a_reg_31_0__31_; 
wire _0a_reg_31_0__3_; 
wire _0a_reg_31_0__4_; 
wire _0a_reg_31_0__5_; 
wire _0a_reg_31_0__6_; 
wire _0a_reg_31_0__7_; 
wire _0a_reg_31_0__8_; 
wire _0a_reg_31_0__9_; 
wire _0b_reg_31_0__0_; 
wire _0b_reg_31_0__10_; 
wire _0b_reg_31_0__11_; 
wire _0b_reg_31_0__12_; 
wire _0b_reg_31_0__13_; 
wire _0b_reg_31_0__14_; 
wire _0b_reg_31_0__15_; 
wire _0b_reg_31_0__16_; 
wire _0b_reg_31_0__17_; 
wire _0b_reg_31_0__18_; 
wire _0b_reg_31_0__19_; 
wire _0b_reg_31_0__1_; 
wire _0b_reg_31_0__20_; 
wire _0b_reg_31_0__21_; 
wire _0b_reg_31_0__22_; 
wire _0b_reg_31_0__23_; 
wire _0b_reg_31_0__24_; 
wire _0b_reg_31_0__25_; 
wire _0b_reg_31_0__26_; 
wire _0b_reg_31_0__27_; 
wire _0b_reg_31_0__28_; 
wire _0b_reg_31_0__29_; 
wire _0b_reg_31_0__2_; 
wire _0b_reg_31_0__30_; 
wire _0b_reg_31_0__31_; 
wire _0b_reg_31_0__3_; 
wire _0b_reg_31_0__4_; 
wire _0b_reg_31_0__5_; 
wire _0b_reg_31_0__6_; 
wire _0b_reg_31_0__7_; 
wire _0b_reg_31_0__8_; 
wire _0b_reg_31_0__9_; 
wire _0c_reg_31_0__0_; 
wire _0c_reg_31_0__10_; 
wire _0c_reg_31_0__11_; 
wire _0c_reg_31_0__12_; 
wire _0c_reg_31_0__13_; 
wire _0c_reg_31_0__14_; 
wire _0c_reg_31_0__15_; 
wire _0c_reg_31_0__16_; 
wire _0c_reg_31_0__17_; 
wire _0c_reg_31_0__18_; 
wire _0c_reg_31_0__19_; 
wire _0c_reg_31_0__1_; 
wire _0c_reg_31_0__20_; 
wire _0c_reg_31_0__21_; 
wire _0c_reg_31_0__22_; 
wire _0c_reg_31_0__23_; 
wire _0c_reg_31_0__24_; 
wire _0c_reg_31_0__25_; 
wire _0c_reg_31_0__26_; 
wire _0c_reg_31_0__27_; 
wire _0c_reg_31_0__28_; 
wire _0c_reg_31_0__29_; 
wire _0c_reg_31_0__2_; 
wire _0c_reg_31_0__30_; 
wire _0c_reg_31_0__31_; 
wire _0c_reg_31_0__3_; 
wire _0c_reg_31_0__4_; 
wire _0c_reg_31_0__5_; 
wire _0c_reg_31_0__6_; 
wire _0c_reg_31_0__7_; 
wire _0c_reg_31_0__8_; 
wire _0c_reg_31_0__9_; 
wire _0d_reg_31_0__0_; 
wire _0d_reg_31_0__10_; 
wire _0d_reg_31_0__11_; 
wire _0d_reg_31_0__12_; 
wire _0d_reg_31_0__13_; 
wire _0d_reg_31_0__14_; 
wire _0d_reg_31_0__15_; 
wire _0d_reg_31_0__16_; 
wire _0d_reg_31_0__17_; 
wire _0d_reg_31_0__18_; 
wire _0d_reg_31_0__19_; 
wire _0d_reg_31_0__1_; 
wire _0d_reg_31_0__20_; 
wire _0d_reg_31_0__21_; 
wire _0d_reg_31_0__22_; 
wire _0d_reg_31_0__23_; 
wire _0d_reg_31_0__24_; 
wire _0d_reg_31_0__25_; 
wire _0d_reg_31_0__26_; 
wire _0d_reg_31_0__27_; 
wire _0d_reg_31_0__28_; 
wire _0d_reg_31_0__29_; 
wire _0d_reg_31_0__2_; 
wire _0d_reg_31_0__30_; 
wire _0d_reg_31_0__31_; 
wire _0d_reg_31_0__3_; 
wire _0d_reg_31_0__4_; 
wire _0d_reg_31_0__5_; 
wire _0d_reg_31_0__6_; 
wire _0d_reg_31_0__7_; 
wire _0d_reg_31_0__8_; 
wire _0d_reg_31_0__9_; 
wire _0digest_valid_reg_0_0_; 
wire _0e_reg_31_0__0_; 
wire _0e_reg_31_0__10_; 
wire _0e_reg_31_0__11_; 
wire _0e_reg_31_0__12_; 
wire _0e_reg_31_0__13_; 
wire _0e_reg_31_0__14_; 
wire _0e_reg_31_0__15_; 
wire _0e_reg_31_0__16_; 
wire _0e_reg_31_0__17_; 
wire _0e_reg_31_0__18_; 
wire _0e_reg_31_0__19_; 
wire _0e_reg_31_0__1_; 
wire _0e_reg_31_0__20_; 
wire _0e_reg_31_0__21_; 
wire _0e_reg_31_0__22_; 
wire _0e_reg_31_0__23_; 
wire _0e_reg_31_0__24_; 
wire _0e_reg_31_0__25_; 
wire _0e_reg_31_0__26_; 
wire _0e_reg_31_0__27_; 
wire _0e_reg_31_0__28_; 
wire _0e_reg_31_0__29_; 
wire _0e_reg_31_0__2_; 
wire _0e_reg_31_0__30_; 
wire _0e_reg_31_0__31_; 
wire _0e_reg_31_0__3_; 
wire _0e_reg_31_0__4_; 
wire _0e_reg_31_0__5_; 
wire _0e_reg_31_0__6_; 
wire _0e_reg_31_0__7_; 
wire _0e_reg_31_0__8_; 
wire _0e_reg_31_0__9_; 
wire _0round_ctr_reg_6_0__0_; 
wire _0round_ctr_reg_6_0__1_; 
wire _0round_ctr_reg_6_0__2_; 
wire _0round_ctr_reg_6_0__3_; 
wire _0round_ctr_reg_6_0__4_; 
wire _0round_ctr_reg_6_0__5_; 
wire _0round_ctr_reg_6_0__6_; 
wire _abc_15497_abc_9717_auto_fsm_map_cc_118_implement_pattern_cache_863; 
wire _abc_15497_abc_9717_auto_fsm_map_cc_170_map_fsm_844_0_; 
wire _abc_15497_abc_9717_auto_fsm_map_cc_170_map_fsm_844_2_; 
wire _abc_15497_new_n1000_; 
wire _abc_15497_new_n1001_; 
wire _abc_15497_new_n1002_; 
wire _abc_15497_new_n1003_; 
wire _abc_15497_new_n1005_; 
wire _abc_15497_new_n1006_; 
wire _abc_15497_new_n1007_; 
wire _abc_15497_new_n1008_; 
wire _abc_15497_new_n1009_; 
wire _abc_15497_new_n1010_; 
wire _abc_15497_new_n1011_; 
wire _abc_15497_new_n1012_; 
wire _abc_15497_new_n1013_; 
wire _abc_15497_new_n1014_; 
wire _abc_15497_new_n1015_; 
wire _abc_15497_new_n1016_; 
wire _abc_15497_new_n1017_; 
wire _abc_15497_new_n1018_; 
wire _abc_15497_new_n1019_; 
wire _abc_15497_new_n1020_; 
wire _abc_15497_new_n1021_; 
wire _abc_15497_new_n1022_; 
wire _abc_15497_new_n1024_; 
wire _abc_15497_new_n1025_; 
wire _abc_15497_new_n1026_; 
wire _abc_15497_new_n1027_; 
wire _abc_15497_new_n1028_; 
wire _abc_15497_new_n1029_; 
wire _abc_15497_new_n1030_; 
wire _abc_15497_new_n1031_; 
wire _abc_15497_new_n1033_; 
wire _abc_15497_new_n1034_; 
wire _abc_15497_new_n1035_; 
wire _abc_15497_new_n1036_; 
wire _abc_15497_new_n1037_; 
wire _abc_15497_new_n1038_; 
wire _abc_15497_new_n1039_; 
wire _abc_15497_new_n1040_; 
wire _abc_15497_new_n1041_; 
wire _abc_15497_new_n1042_; 
wire _abc_15497_new_n1043_; 
wire _abc_15497_new_n1044_; 
wire _abc_15497_new_n1045_; 
wire _abc_15497_new_n1046_; 
wire _abc_15497_new_n1048_; 
wire _abc_15497_new_n1049_; 
wire _abc_15497_new_n1050_; 
wire _abc_15497_new_n1051_; 
wire _abc_15497_new_n1052_; 
wire _abc_15497_new_n1053_; 
wire _abc_15497_new_n1054_; 
wire _abc_15497_new_n1055_; 
wire _abc_15497_new_n1057_; 
wire _abc_15497_new_n1058_; 
wire _abc_15497_new_n1059_; 
wire _abc_15497_new_n1060_; 
wire _abc_15497_new_n1061_; 
wire _abc_15497_new_n1062_; 
wire _abc_15497_new_n1063_; 
wire _abc_15497_new_n1064_; 
wire _abc_15497_new_n1065_; 
wire _abc_15497_new_n1066_; 
wire _abc_15497_new_n1067_; 
wire _abc_15497_new_n1068_; 
wire _abc_15497_new_n1069_; 
wire _abc_15497_new_n1071_; 
wire _abc_15497_new_n1072_; 
wire _abc_15497_new_n1073_; 
wire _abc_15497_new_n1074_; 
wire _abc_15497_new_n1075_; 
wire _abc_15497_new_n1076_; 
wire _abc_15497_new_n1077_; 
wire _abc_15497_new_n1079_; 
wire _abc_15497_new_n1080_; 
wire _abc_15497_new_n1081_; 
wire _abc_15497_new_n1082_; 
wire _abc_15497_new_n1083_; 
wire _abc_15497_new_n1084_; 
wire _abc_15497_new_n1085_; 
wire _abc_15497_new_n1086_; 
wire _abc_15497_new_n1087_; 
wire _abc_15497_new_n1088_; 
wire _abc_15497_new_n1089_; 
wire _abc_15497_new_n1090_; 
wire _abc_15497_new_n1091_; 
wire _abc_15497_new_n1093_; 
wire _abc_15497_new_n1094_; 
wire _abc_15497_new_n1095_; 
wire _abc_15497_new_n1096_; 
wire _abc_15497_new_n1097_; 
wire _abc_15497_new_n1098_; 
wire _abc_15497_new_n1099_; 
wire _abc_15497_new_n1101_; 
wire _abc_15497_new_n1102_; 
wire _abc_15497_new_n1103_; 
wire _abc_15497_new_n1104_; 
wire _abc_15497_new_n1105_; 
wire _abc_15497_new_n1106_; 
wire _abc_15497_new_n1107_; 
wire _abc_15497_new_n1108_; 
wire _abc_15497_new_n1109_; 
wire _abc_15497_new_n1110_; 
wire _abc_15497_new_n1111_; 
wire _abc_15497_new_n1112_; 
wire _abc_15497_new_n1113_; 
wire _abc_15497_new_n1114_; 
wire _abc_15497_new_n1115_; 
wire _abc_15497_new_n1116_; 
wire _abc_15497_new_n1117_; 
wire _abc_15497_new_n1119_; 
wire _abc_15497_new_n1120_; 
wire _abc_15497_new_n1121_; 
wire _abc_15497_new_n1122_; 
wire _abc_15497_new_n1123_; 
wire _abc_15497_new_n1124_; 
wire _abc_15497_new_n1125_; 
wire _abc_15497_new_n1126_; 
wire _abc_15497_new_n1128_; 
wire _abc_15497_new_n1129_; 
wire _abc_15497_new_n1130_; 
wire _abc_15497_new_n1131_; 
wire _abc_15497_new_n1132_; 
wire _abc_15497_new_n1133_; 
wire _abc_15497_new_n1134_; 
wire _abc_15497_new_n1135_; 
wire _abc_15497_new_n1136_; 
wire _abc_15497_new_n1137_; 
wire _abc_15497_new_n1138_; 
wire _abc_15497_new_n1139_; 
wire _abc_15497_new_n1140_; 
wire _abc_15497_new_n1142_; 
wire _abc_15497_new_n1143_; 
wire _abc_15497_new_n1144_; 
wire _abc_15497_new_n1145_; 
wire _abc_15497_new_n1146_; 
wire _abc_15497_new_n1147_; 
wire _abc_15497_new_n1148_; 
wire _abc_15497_new_n1149_; 
wire _abc_15497_new_n1151_; 
wire _abc_15497_new_n1152_; 
wire _abc_15497_new_n1153_; 
wire _abc_15497_new_n1154_; 
wire _abc_15497_new_n1155_; 
wire _abc_15497_new_n1156_; 
wire _abc_15497_new_n1157_; 
wire _abc_15497_new_n1158_; 
wire _abc_15497_new_n1159_; 
wire _abc_15497_new_n1160_; 
wire _abc_15497_new_n1161_; 
wire _abc_15497_new_n1162_; 
wire _abc_15497_new_n1163_; 
wire _abc_15497_new_n1164_; 
wire _abc_15497_new_n1165_; 
wire _abc_15497_new_n1166_; 
wire _abc_15497_new_n1167_; 
wire _abc_15497_new_n1168_; 
wire _abc_15497_new_n1169_; 
wire _abc_15497_new_n1171_; 
wire _abc_15497_new_n1172_; 
wire _abc_15497_new_n1173_; 
wire _abc_15497_new_n1174_; 
wire _abc_15497_new_n1175_; 
wire _abc_15497_new_n1176_; 
wire _abc_15497_new_n1177_; 
wire _abc_15497_new_n1179_; 
wire _abc_15497_new_n1180_; 
wire _abc_15497_new_n1181_; 
wire _abc_15497_new_n1182_; 
wire _abc_15497_new_n1183_; 
wire _abc_15497_new_n1184_; 
wire _abc_15497_new_n1185_; 
wire _abc_15497_new_n1186_; 
wire _abc_15497_new_n1187_; 
wire _abc_15497_new_n1188_; 
wire _abc_15497_new_n1189_; 
wire _abc_15497_new_n1190_; 
wire _abc_15497_new_n1191_; 
wire _abc_15497_new_n1193_; 
wire _abc_15497_new_n1194_; 
wire _abc_15497_new_n1195_; 
wire _abc_15497_new_n1196_; 
wire _abc_15497_new_n1197_; 
wire _abc_15497_new_n1198_; 
wire _abc_15497_new_n1199_; 
wire _abc_15497_new_n1201_; 
wire _abc_15497_new_n1202_; 
wire _abc_15497_new_n1203_; 
wire _abc_15497_new_n1204_; 
wire _abc_15497_new_n1205_; 
wire _abc_15497_new_n1206_; 
wire _abc_15497_new_n1207_; 
wire _abc_15497_new_n1208_; 
wire _abc_15497_new_n1209_; 
wire _abc_15497_new_n1210_; 
wire _abc_15497_new_n1211_; 
wire _abc_15497_new_n1212_; 
wire _abc_15497_new_n1213_; 
wire _abc_15497_new_n1214_; 
wire _abc_15497_new_n1215_; 
wire _abc_15497_new_n1216_; 
wire _abc_15497_new_n1217_; 
wire _abc_15497_new_n1218_; 
wire _abc_15497_new_n1219_; 
wire _abc_15497_new_n1220_; 
wire _abc_15497_new_n1222_; 
wire _abc_15497_new_n1223_; 
wire _abc_15497_new_n1224_; 
wire _abc_15497_new_n1225_; 
wire _abc_15497_new_n1226_; 
wire _abc_15497_new_n1227_; 
wire _abc_15497_new_n1228_; 
wire _abc_15497_new_n1229_; 
wire _abc_15497_new_n1231_; 
wire _abc_15497_new_n1232_; 
wire _abc_15497_new_n1233_; 
wire _abc_15497_new_n1234_; 
wire _abc_15497_new_n1235_; 
wire _abc_15497_new_n1236_; 
wire _abc_15497_new_n1237_; 
wire _abc_15497_new_n1238_; 
wire _abc_15497_new_n1239_; 
wire _abc_15497_new_n1240_; 
wire _abc_15497_new_n1241_; 
wire _abc_15497_new_n1242_; 
wire _abc_15497_new_n1243_; 
wire _abc_15497_new_n1244_; 
wire _abc_15497_new_n1245_; 
wire _abc_15497_new_n1247_; 
wire _abc_15497_new_n1248_; 
wire _abc_15497_new_n1249_; 
wire _abc_15497_new_n1250_; 
wire _abc_15497_new_n1251_; 
wire _abc_15497_new_n1252_; 
wire _abc_15497_new_n1253_; 
wire _abc_15497_new_n1254_; 
wire _abc_15497_new_n1255_; 
wire _abc_15497_new_n1256_; 
wire _abc_15497_new_n1258_; 
wire _abc_15497_new_n1259_; 
wire _abc_15497_new_n1260_; 
wire _abc_15497_new_n1261_; 
wire _abc_15497_new_n1262_; 
wire _abc_15497_new_n1263_; 
wire _abc_15497_new_n1264_; 
wire _abc_15497_new_n1265_; 
wire _abc_15497_new_n1266_; 
wire _abc_15497_new_n1267_; 
wire _abc_15497_new_n1269_; 
wire _abc_15497_new_n1270_; 
wire _abc_15497_new_n1271_; 
wire _abc_15497_new_n1272_; 
wire _abc_15497_new_n1273_; 
wire _abc_15497_new_n1274_; 
wire _abc_15497_new_n1275_; 
wire _abc_15497_new_n1276_; 
wire _abc_15497_new_n1277_; 
wire _abc_15497_new_n1278_; 
wire _abc_15497_new_n1280_; 
wire _abc_15497_new_n1281_; 
wire _abc_15497_new_n1282_; 
wire _abc_15497_new_n1283_; 
wire _abc_15497_new_n1284_; 
wire _abc_15497_new_n1285_; 
wire _abc_15497_new_n1286_; 
wire _abc_15497_new_n1287_; 
wire _abc_15497_new_n1288_; 
wire _abc_15497_new_n1290_; 
wire _abc_15497_new_n1291_; 
wire _abc_15497_new_n1292_; 
wire _abc_15497_new_n1293_; 
wire _abc_15497_new_n1294_; 
wire _abc_15497_new_n1295_; 
wire _abc_15497_new_n1296_; 
wire _abc_15497_new_n1298_; 
wire _abc_15497_new_n1299_; 
wire _abc_15497_new_n1300_; 
wire _abc_15497_new_n1301_; 
wire _abc_15497_new_n1303_; 
wire _abc_15497_new_n1304_; 
wire _abc_15497_new_n1305_; 
wire _abc_15497_new_n1307_; 
wire _abc_15497_new_n1308_; 
wire _abc_15497_new_n1309_; 
wire _abc_15497_new_n1310_; 
wire _abc_15497_new_n1311_; 
wire _abc_15497_new_n1312_; 
wire _abc_15497_new_n1313_; 
wire _abc_15497_new_n1314_; 
wire _abc_15497_new_n1315_; 
wire _abc_15497_new_n1317_; 
wire _abc_15497_new_n1318_; 
wire _abc_15497_new_n1319_; 
wire _abc_15497_new_n1320_; 
wire _abc_15497_new_n1321_; 
wire _abc_15497_new_n1322_; 
wire _abc_15497_new_n1323_; 
wire _abc_15497_new_n1324_; 
wire _abc_15497_new_n1326_; 
wire _abc_15497_new_n1327_; 
wire _abc_15497_new_n1328_; 
wire _abc_15497_new_n1329_; 
wire _abc_15497_new_n1330_; 
wire _abc_15497_new_n1332_; 
wire _abc_15497_new_n1333_; 
wire _abc_15497_new_n1334_; 
wire _abc_15497_new_n1335_; 
wire _abc_15497_new_n1336_; 
wire _abc_15497_new_n1337_; 
wire _abc_15497_new_n1338_; 
wire _abc_15497_new_n1339_; 
wire _abc_15497_new_n1340_; 
wire _abc_15497_new_n1342_; 
wire _abc_15497_new_n1343_; 
wire _abc_15497_new_n1344_; 
wire _abc_15497_new_n1345_; 
wire _abc_15497_new_n1346_; 
wire _abc_15497_new_n1347_; 
wire _abc_15497_new_n1348_; 
wire _abc_15497_new_n1349_; 
wire _abc_15497_new_n1351_; 
wire _abc_15497_new_n1352_; 
wire _abc_15497_new_n1353_; 
wire _abc_15497_new_n1354_; 
wire _abc_15497_new_n1355_; 
wire _abc_15497_new_n1356_; 
wire _abc_15497_new_n1357_; 
wire _abc_15497_new_n1358_; 
wire _abc_15497_new_n1359_; 
wire _abc_15497_new_n1361_; 
wire _abc_15497_new_n1362_; 
wire _abc_15497_new_n1363_; 
wire _abc_15497_new_n1364_; 
wire _abc_15497_new_n1365_; 
wire _abc_15497_new_n1366_; 
wire _abc_15497_new_n1367_; 
wire _abc_15497_new_n1368_; 
wire _abc_15497_new_n1369_; 
wire _abc_15497_new_n1371_; 
wire _abc_15497_new_n1372_; 
wire _abc_15497_new_n1373_; 
wire _abc_15497_new_n1374_; 
wire _abc_15497_new_n1375_; 
wire _abc_15497_new_n1376_; 
wire _abc_15497_new_n1377_; 
wire _abc_15497_new_n1378_; 
wire _abc_15497_new_n1379_; 
wire _abc_15497_new_n1380_; 
wire _abc_15497_new_n1382_; 
wire _abc_15497_new_n1383_; 
wire _abc_15497_new_n1384_; 
wire _abc_15497_new_n1385_; 
wire _abc_15497_new_n1386_; 
wire _abc_15497_new_n1387_; 
wire _abc_15497_new_n1388_; 
wire _abc_15497_new_n1389_; 
wire _abc_15497_new_n1390_; 
wire _abc_15497_new_n1391_; 
wire _abc_15497_new_n1392_; 
wire _abc_15497_new_n1393_; 
wire _abc_15497_new_n1395_; 
wire _abc_15497_new_n1396_; 
wire _abc_15497_new_n1397_; 
wire _abc_15497_new_n1398_; 
wire _abc_15497_new_n1399_; 
wire _abc_15497_new_n1400_; 
wire _abc_15497_new_n1401_; 
wire _abc_15497_new_n1402_; 
wire _abc_15497_new_n1403_; 
wire _abc_15497_new_n1405_; 
wire _abc_15497_new_n1406_; 
wire _abc_15497_new_n1407_; 
wire _abc_15497_new_n1408_; 
wire _abc_15497_new_n1409_; 
wire _abc_15497_new_n1410_; 
wire _abc_15497_new_n1411_; 
wire _abc_15497_new_n1412_; 
wire _abc_15497_new_n1413_; 
wire _abc_15497_new_n1414_; 
wire _abc_15497_new_n1415_; 
wire _abc_15497_new_n1416_; 
wire _abc_15497_new_n1417_; 
wire _abc_15497_new_n1418_; 
wire _abc_15497_new_n1419_; 
wire _abc_15497_new_n1420_; 
wire _abc_15497_new_n1422_; 
wire _abc_15497_new_n1423_; 
wire _abc_15497_new_n1424_; 
wire _abc_15497_new_n1425_; 
wire _abc_15497_new_n1426_; 
wire _abc_15497_new_n1427_; 
wire _abc_15497_new_n1428_; 
wire _abc_15497_new_n1429_; 
wire _abc_15497_new_n1430_; 
wire _abc_15497_new_n1432_; 
wire _abc_15497_new_n1433_; 
wire _abc_15497_new_n1434_; 
wire _abc_15497_new_n1435_; 
wire _abc_15497_new_n1436_; 
wire _abc_15497_new_n1437_; 
wire _abc_15497_new_n1438_; 
wire _abc_15497_new_n1439_; 
wire _abc_15497_new_n1440_; 
wire _abc_15497_new_n1441_; 
wire _abc_15497_new_n1442_; 
wire _abc_15497_new_n1444_; 
wire _abc_15497_new_n1445_; 
wire _abc_15497_new_n1446_; 
wire _abc_15497_new_n1447_; 
wire _abc_15497_new_n1448_; 
wire _abc_15497_new_n1449_; 
wire _abc_15497_new_n1450_; 
wire _abc_15497_new_n1452_; 
wire _abc_15497_new_n1453_; 
wire _abc_15497_new_n1454_; 
wire _abc_15497_new_n1455_; 
wire _abc_15497_new_n1456_; 
wire _abc_15497_new_n1457_; 
wire _abc_15497_new_n1458_; 
wire _abc_15497_new_n1459_; 
wire _abc_15497_new_n1460_; 
wire _abc_15497_new_n1461_; 
wire _abc_15497_new_n1462_; 
wire _abc_15497_new_n1463_; 
wire _abc_15497_new_n1464_; 
wire _abc_15497_new_n1465_; 
wire _abc_15497_new_n1467_; 
wire _abc_15497_new_n1468_; 
wire _abc_15497_new_n1469_; 
wire _abc_15497_new_n1470_; 
wire _abc_15497_new_n1471_; 
wire _abc_15497_new_n1472_; 
wire _abc_15497_new_n1473_; 
wire _abc_15497_new_n1474_; 
wire _abc_15497_new_n1475_; 
wire _abc_15497_new_n1477_; 
wire _abc_15497_new_n1478_; 
wire _abc_15497_new_n1479_; 
wire _abc_15497_new_n1480_; 
wire _abc_15497_new_n1481_; 
wire _abc_15497_new_n1482_; 
wire _abc_15497_new_n1483_; 
wire _abc_15497_new_n1484_; 
wire _abc_15497_new_n1485_; 
wire _abc_15497_new_n1486_; 
wire _abc_15497_new_n1487_; 
wire _abc_15497_new_n1488_; 
wire _abc_15497_new_n1489_; 
wire _abc_15497_new_n1490_; 
wire _abc_15497_new_n1492_; 
wire _abc_15497_new_n1493_; 
wire _abc_15497_new_n1494_; 
wire _abc_15497_new_n1495_; 
wire _abc_15497_new_n1496_; 
wire _abc_15497_new_n1497_; 
wire _abc_15497_new_n1498_; 
wire _abc_15497_new_n1499_; 
wire _abc_15497_new_n1500_; 
wire _abc_15497_new_n1502_; 
wire _abc_15497_new_n1503_; 
wire _abc_15497_new_n1504_; 
wire _abc_15497_new_n1505_; 
wire _abc_15497_new_n1506_; 
wire _abc_15497_new_n1507_; 
wire _abc_15497_new_n1508_; 
wire _abc_15497_new_n1509_; 
wire _abc_15497_new_n1510_; 
wire _abc_15497_new_n1511_; 
wire _abc_15497_new_n1512_; 
wire _abc_15497_new_n1513_; 
wire _abc_15497_new_n1514_; 
wire _abc_15497_new_n1515_; 
wire _abc_15497_new_n1516_; 
wire _abc_15497_new_n1517_; 
wire _abc_15497_new_n1519_; 
wire _abc_15497_new_n1520_; 
wire _abc_15497_new_n1521_; 
wire _abc_15497_new_n1522_; 
wire _abc_15497_new_n1523_; 
wire _abc_15497_new_n1524_; 
wire _abc_15497_new_n1525_; 
wire _abc_15497_new_n1526_; 
wire _abc_15497_new_n1528_; 
wire _abc_15497_new_n1529_; 
wire _abc_15497_new_n1530_; 
wire _abc_15497_new_n1531_; 
wire _abc_15497_new_n1532_; 
wire _abc_15497_new_n1533_; 
wire _abc_15497_new_n1534_; 
wire _abc_15497_new_n1535_; 
wire _abc_15497_new_n1536_; 
wire _abc_15497_new_n1537_; 
wire _abc_15497_new_n1538_; 
wire _abc_15497_new_n1540_; 
wire _abc_15497_new_n1541_; 
wire _abc_15497_new_n1542_; 
wire _abc_15497_new_n1543_; 
wire _abc_15497_new_n1544_; 
wire _abc_15497_new_n1545_; 
wire _abc_15497_new_n1546_; 
wire _abc_15497_new_n1547_; 
wire _abc_15497_new_n1548_; 
wire _abc_15497_new_n1550_; 
wire _abc_15497_new_n1551_; 
wire _abc_15497_new_n1552_; 
wire _abc_15497_new_n1553_; 
wire _abc_15497_new_n1554_; 
wire _abc_15497_new_n1555_; 
wire _abc_15497_new_n1556_; 
wire _abc_15497_new_n1557_; 
wire _abc_15497_new_n1558_; 
wire _abc_15497_new_n1559_; 
wire _abc_15497_new_n1560_; 
wire _abc_15497_new_n1561_; 
wire _abc_15497_new_n1562_; 
wire _abc_15497_new_n1563_; 
wire _abc_15497_new_n1564_; 
wire _abc_15497_new_n1565_; 
wire _abc_15497_new_n1566_; 
wire _abc_15497_new_n1567_; 
wire _abc_15497_new_n1569_; 
wire _abc_15497_new_n1570_; 
wire _abc_15497_new_n1571_; 
wire _abc_15497_new_n1572_; 
wire _abc_15497_new_n1573_; 
wire _abc_15497_new_n1574_; 
wire _abc_15497_new_n1575_; 
wire _abc_15497_new_n1576_; 
wire _abc_15497_new_n1577_; 
wire _abc_15497_new_n1578_; 
wire _abc_15497_new_n1580_; 
wire _abc_15497_new_n1581_; 
wire _abc_15497_new_n1582_; 
wire _abc_15497_new_n1583_; 
wire _abc_15497_new_n1584_; 
wire _abc_15497_new_n1585_; 
wire _abc_15497_new_n1586_; 
wire _abc_15497_new_n1587_; 
wire _abc_15497_new_n1588_; 
wire _abc_15497_new_n1589_; 
wire _abc_15497_new_n1590_; 
wire _abc_15497_new_n1591_; 
wire _abc_15497_new_n1593_; 
wire _abc_15497_new_n1594_; 
wire _abc_15497_new_n1595_; 
wire _abc_15497_new_n1596_; 
wire _abc_15497_new_n1597_; 
wire _abc_15497_new_n1598_; 
wire _abc_15497_new_n1599_; 
wire _abc_15497_new_n1600_; 
wire _abc_15497_new_n1601_; 
wire _abc_15497_new_n1602_; 
wire _abc_15497_new_n1604_; 
wire _abc_15497_new_n1605_; 
wire _abc_15497_new_n1606_; 
wire _abc_15497_new_n1607_; 
wire _abc_15497_new_n1608_; 
wire _abc_15497_new_n1609_; 
wire _abc_15497_new_n1610_; 
wire _abc_15497_new_n1611_; 
wire _abc_15497_new_n1612_; 
wire _abc_15497_new_n1613_; 
wire _abc_15497_new_n1614_; 
wire _abc_15497_new_n1615_; 
wire _abc_15497_new_n1617_; 
wire _abc_15497_new_n1618_; 
wire _abc_15497_new_n1619_; 
wire _abc_15497_new_n1620_; 
wire _abc_15497_new_n1621_; 
wire _abc_15497_new_n1622_; 
wire _abc_15497_new_n1623_; 
wire _abc_15497_new_n1624_; 
wire _abc_15497_new_n1625_; 
wire _abc_15497_new_n1626_; 
wire _abc_15497_new_n1628_; 
wire _abc_15497_new_n1629_; 
wire _abc_15497_new_n1630_; 
wire _abc_15497_new_n1631_; 
wire _abc_15497_new_n1632_; 
wire _abc_15497_new_n1633_; 
wire _abc_15497_new_n1634_; 
wire _abc_15497_new_n1635_; 
wire _abc_15497_new_n1637_; 
wire _abc_15497_new_n1638_; 
wire _abc_15497_new_n1639_; 
wire _abc_15497_new_n1640_; 
wire _abc_15497_new_n1641_; 
wire _abc_15497_new_n1642_; 
wire _abc_15497_new_n1644_; 
wire _abc_15497_new_n1646_; 
wire _abc_15497_new_n1647_; 
wire _abc_15497_new_n1648_; 
wire _abc_15497_new_n1648__bF_buf0; 
wire _abc_15497_new_n1648__bF_buf1; 
wire _abc_15497_new_n1648__bF_buf2; 
wire _abc_15497_new_n1648__bF_buf3; 
wire _abc_15497_new_n1648__bF_buf4; 
wire _abc_15497_new_n1648__bF_buf5; 
wire _abc_15497_new_n1648__bF_buf6; 
wire _abc_15497_new_n1648__bF_buf7; 
wire _abc_15497_new_n1648__bF_buf8; 
wire _abc_15497_new_n1649_; 
wire _abc_15497_new_n1650_; 
wire _abc_15497_new_n1650__bF_buf0; 
wire _abc_15497_new_n1650__bF_buf1; 
wire _abc_15497_new_n1650__bF_buf2; 
wire _abc_15497_new_n1650__bF_buf3; 
wire _abc_15497_new_n1650__bF_buf4; 
wire _abc_15497_new_n1650__bF_buf5; 
wire _abc_15497_new_n1650__bF_buf6; 
wire _abc_15497_new_n1650__bF_buf7; 
wire _abc_15497_new_n1650__bF_buf8; 
wire _abc_15497_new_n1650__bF_buf9; 
wire _abc_15497_new_n1651_; 
wire _abc_15497_new_n1653_; 
wire _abc_15497_new_n1654_; 
wire _abc_15497_new_n1656_; 
wire _abc_15497_new_n1657_; 
wire _abc_15497_new_n1659_; 
wire _abc_15497_new_n1660_; 
wire _abc_15497_new_n1662_; 
wire _abc_15497_new_n1663_; 
wire _abc_15497_new_n1663__bF_buf0; 
wire _abc_15497_new_n1663__bF_buf1; 
wire _abc_15497_new_n1663__bF_buf2; 
wire _abc_15497_new_n1663__bF_buf3; 
wire _abc_15497_new_n1663__bF_buf4; 
wire _abc_15497_new_n1663__bF_buf5; 
wire _abc_15497_new_n1663__bF_buf6; 
wire _abc_15497_new_n1663__bF_buf7; 
wire _abc_15497_new_n1664_; 
wire _abc_15497_new_n1666_; 
wire _abc_15497_new_n1667_; 
wire _abc_15497_new_n1669_; 
wire _abc_15497_new_n1670_; 
wire _abc_15497_new_n1672_; 
wire _abc_15497_new_n1673_; 
wire _abc_15497_new_n1675_; 
wire _abc_15497_new_n1676_; 
wire _abc_15497_new_n1678_; 
wire _abc_15497_new_n1679_; 
wire _abc_15497_new_n1681_; 
wire _abc_15497_new_n1682_; 
wire _abc_15497_new_n1684_; 
wire _abc_15497_new_n1685_; 
wire _abc_15497_new_n1686_; 
wire _abc_15497_new_n1688_; 
wire _abc_15497_new_n1689_; 
wire _abc_15497_new_n1691_; 
wire _abc_15497_new_n1692_; 
wire _abc_15497_new_n1694_; 
wire _abc_15497_new_n1695_; 
wire _abc_15497_new_n1697_; 
wire _abc_15497_new_n1698_; 
wire _abc_15497_new_n1700_; 
wire _abc_15497_new_n1701_; 
wire _abc_15497_new_n1703_; 
wire _abc_15497_new_n1704_; 
wire _abc_15497_new_n1706_; 
wire _abc_15497_new_n1707_; 
wire _abc_15497_new_n1709_; 
wire _abc_15497_new_n1710_; 
wire _abc_15497_new_n1712_; 
wire _abc_15497_new_n1713_; 
wire _abc_15497_new_n1715_; 
wire _abc_15497_new_n1716_; 
wire _abc_15497_new_n1718_; 
wire _abc_15497_new_n1719_; 
wire _abc_15497_new_n1721_; 
wire _abc_15497_new_n1722_; 
wire _abc_15497_new_n1724_; 
wire _abc_15497_new_n1725_; 
wire _abc_15497_new_n1727_; 
wire _abc_15497_new_n1728_; 
wire _abc_15497_new_n1730_; 
wire _abc_15497_new_n1731_; 
wire _abc_15497_new_n1733_; 
wire _abc_15497_new_n1734_; 
wire _abc_15497_new_n1736_; 
wire _abc_15497_new_n1737_; 
wire _abc_15497_new_n1738_; 
wire _abc_15497_new_n1740_; 
wire _abc_15497_new_n1741_; 
wire _abc_15497_new_n1743_; 
wire _abc_15497_new_n1744_; 
wire _abc_15497_new_n1746_; 
wire _abc_15497_new_n1747_; 
wire _abc_15497_new_n1748_; 
wire _abc_15497_new_n1750_; 
wire _abc_15497_new_n1751_; 
wire _abc_15497_new_n1752_; 
wire _abc_15497_new_n1753_; 
wire _abc_15497_new_n1754_; 
wire _abc_15497_new_n1756_; 
wire _abc_15497_new_n1757_; 
wire _abc_15497_new_n1758_; 
wire _abc_15497_new_n1759_; 
wire _abc_15497_new_n1760_; 
wire _abc_15497_new_n1762_; 
wire _abc_15497_new_n1763_; 
wire _abc_15497_new_n1764_; 
wire _abc_15497_new_n1765_; 
wire _abc_15497_new_n1766_; 
wire _abc_15497_new_n1767_; 
wire _abc_15497_new_n1768_; 
wire _abc_15497_new_n1769_; 
wire _abc_15497_new_n1771_; 
wire _abc_15497_new_n1772_; 
wire _abc_15497_new_n1773_; 
wire _abc_15497_new_n1774_; 
wire _abc_15497_new_n1775_; 
wire _abc_15497_new_n1776_; 
wire _abc_15497_new_n1777_; 
wire _abc_15497_new_n1779_; 
wire _abc_15497_new_n1780_; 
wire _abc_15497_new_n1781_; 
wire _abc_15497_new_n1782_; 
wire _abc_15497_new_n1783_; 
wire _abc_15497_new_n1784_; 
wire _abc_15497_new_n1785_; 
wire _abc_15497_new_n1787_; 
wire _abc_15497_new_n1788_; 
wire _abc_15497_new_n1789_; 
wire _abc_15497_new_n1790_; 
wire _abc_15497_new_n1791_; 
wire _abc_15497_new_n1792_; 
wire _abc_15497_new_n1793_; 
wire _abc_15497_new_n1794_; 
wire _abc_15497_new_n1795_; 
wire _abc_15497_new_n1796_; 
wire _abc_15497_new_n1797_; 
wire _abc_15497_new_n1799_; 
wire _abc_15497_new_n1800_; 
wire _abc_15497_new_n1801_; 
wire _abc_15497_new_n1802_; 
wire _abc_15497_new_n1803_; 
wire _abc_15497_new_n1804_; 
wire _abc_15497_new_n1805_; 
wire _abc_15497_new_n1807_; 
wire _abc_15497_new_n1808_; 
wire _abc_15497_new_n1809_; 
wire _abc_15497_new_n1810_; 
wire _abc_15497_new_n1811_; 
wire _abc_15497_new_n1812_; 
wire _abc_15497_new_n1813_; 
wire _abc_15497_new_n1814_; 
wire _abc_15497_new_n1815_; 
wire _abc_15497_new_n1816_; 
wire _abc_15497_new_n1818_; 
wire _abc_15497_new_n1819_; 
wire _abc_15497_new_n1820_; 
wire _abc_15497_new_n1821_; 
wire _abc_15497_new_n1822_; 
wire _abc_15497_new_n1823_; 
wire _abc_15497_new_n1824_; 
wire _abc_15497_new_n1825_; 
wire _abc_15497_new_n1826_; 
wire _abc_15497_new_n1827_; 
wire _abc_15497_new_n1829_; 
wire _abc_15497_new_n1830_; 
wire _abc_15497_new_n1831_; 
wire _abc_15497_new_n1832_; 
wire _abc_15497_new_n1833_; 
wire _abc_15497_new_n1834_; 
wire _abc_15497_new_n1836_; 
wire _abc_15497_new_n1837_; 
wire _abc_15497_new_n1838_; 
wire _abc_15497_new_n1839_; 
wire _abc_15497_new_n1840_; 
wire _abc_15497_new_n1841_; 
wire _abc_15497_new_n1842_; 
wire _abc_15497_new_n1843_; 
wire _abc_15497_new_n1844_; 
wire _abc_15497_new_n1845_; 
wire _abc_15497_new_n1846_; 
wire _abc_15497_new_n1848_; 
wire _abc_15497_new_n1849_; 
wire _abc_15497_new_n1850_; 
wire _abc_15497_new_n1851_; 
wire _abc_15497_new_n1852_; 
wire _abc_15497_new_n1853_; 
wire _abc_15497_new_n1854_; 
wire _abc_15497_new_n1856_; 
wire _abc_15497_new_n1857_; 
wire _abc_15497_new_n1858_; 
wire _abc_15497_new_n1859_; 
wire _abc_15497_new_n1860_; 
wire _abc_15497_new_n1861_; 
wire _abc_15497_new_n1862_; 
wire _abc_15497_new_n1863_; 
wire _abc_15497_new_n1864_; 
wire _abc_15497_new_n1865_; 
wire _abc_15497_new_n1866_; 
wire _abc_15497_new_n1868_; 
wire _abc_15497_new_n1869_; 
wire _abc_15497_new_n1870_; 
wire _abc_15497_new_n1871_; 
wire _abc_15497_new_n1872_; 
wire _abc_15497_new_n1874_; 
wire _abc_15497_new_n1875_; 
wire _abc_15497_new_n1876_; 
wire _abc_15497_new_n1877_; 
wire _abc_15497_new_n1878_; 
wire _abc_15497_new_n1879_; 
wire _abc_15497_new_n1880_; 
wire _abc_15497_new_n1881_; 
wire _abc_15497_new_n1882_; 
wire _abc_15497_new_n1883_; 
wire _abc_15497_new_n1884_; 
wire _abc_15497_new_n1885_; 
wire _abc_15497_new_n1886_; 
wire _abc_15497_new_n1887_; 
wire _abc_15497_new_n1888_; 
wire _abc_15497_new_n1890_; 
wire _abc_15497_new_n1891_; 
wire _abc_15497_new_n1892_; 
wire _abc_15497_new_n1893_; 
wire _abc_15497_new_n1894_; 
wire _abc_15497_new_n1895_; 
wire _abc_15497_new_n1896_; 
wire _abc_15497_new_n1897_; 
wire _abc_15497_new_n1899_; 
wire _abc_15497_new_n1900_; 
wire _abc_15497_new_n1901_; 
wire _abc_15497_new_n1902_; 
wire _abc_15497_new_n1903_; 
wire _abc_15497_new_n1904_; 
wire _abc_15497_new_n1905_; 
wire _abc_15497_new_n1906_; 
wire _abc_15497_new_n1907_; 
wire _abc_15497_new_n1908_; 
wire _abc_15497_new_n1909_; 
wire _abc_15497_new_n1910_; 
wire _abc_15497_new_n1911_; 
wire _abc_15497_new_n1912_; 
wire _abc_15497_new_n1913_; 
wire _abc_15497_new_n1914_; 
wire _abc_15497_new_n1916_; 
wire _abc_15497_new_n1917_; 
wire _abc_15497_new_n1918_; 
wire _abc_15497_new_n1919_; 
wire _abc_15497_new_n1920_; 
wire _abc_15497_new_n1921_; 
wire _abc_15497_new_n1922_; 
wire _abc_15497_new_n1924_; 
wire _abc_15497_new_n1925_; 
wire _abc_15497_new_n1926_; 
wire _abc_15497_new_n1927_; 
wire _abc_15497_new_n1928_; 
wire _abc_15497_new_n1929_; 
wire _abc_15497_new_n1930_; 
wire _abc_15497_new_n1931_; 
wire _abc_15497_new_n1932_; 
wire _abc_15497_new_n1933_; 
wire _abc_15497_new_n1934_; 
wire _abc_15497_new_n1935_; 
wire _abc_15497_new_n1936_; 
wire _abc_15497_new_n1938_; 
wire _abc_15497_new_n1939_; 
wire _abc_15497_new_n1940_; 
wire _abc_15497_new_n1941_; 
wire _abc_15497_new_n1942_; 
wire _abc_15497_new_n1943_; 
wire _abc_15497_new_n1944_; 
wire _abc_15497_new_n1945_; 
wire _abc_15497_new_n1946_; 
wire _abc_15497_new_n1947_; 
wire _abc_15497_new_n1949_; 
wire _abc_15497_new_n1950_; 
wire _abc_15497_new_n1951_; 
wire _abc_15497_new_n1952_; 
wire _abc_15497_new_n1953_; 
wire _abc_15497_new_n1954_; 
wire _abc_15497_new_n1955_; 
wire _abc_15497_new_n1956_; 
wire _abc_15497_new_n1957_; 
wire _abc_15497_new_n1958_; 
wire _abc_15497_new_n1959_; 
wire _abc_15497_new_n1960_; 
wire _abc_15497_new_n1961_; 
wire _abc_15497_new_n1962_; 
wire _abc_15497_new_n1963_; 
wire _abc_15497_new_n1965_; 
wire _abc_15497_new_n1966_; 
wire _abc_15497_new_n1967_; 
wire _abc_15497_new_n1968_; 
wire _abc_15497_new_n1969_; 
wire _abc_15497_new_n1970_; 
wire _abc_15497_new_n1971_; 
wire _abc_15497_new_n1972_; 
wire _abc_15497_new_n1974_; 
wire _abc_15497_new_n1975_; 
wire _abc_15497_new_n1976_; 
wire _abc_15497_new_n1977_; 
wire _abc_15497_new_n1978_; 
wire _abc_15497_new_n1979_; 
wire _abc_15497_new_n1980_; 
wire _abc_15497_new_n1981_; 
wire _abc_15497_new_n1982_; 
wire _abc_15497_new_n1983_; 
wire _abc_15497_new_n1984_; 
wire _abc_15497_new_n1986_; 
wire _abc_15497_new_n1987_; 
wire _abc_15497_new_n1988_; 
wire _abc_15497_new_n1989_; 
wire _abc_15497_new_n1990_; 
wire _abc_15497_new_n1991_; 
wire _abc_15497_new_n1992_; 
wire _abc_15497_new_n1994_; 
wire _abc_15497_new_n1995_; 
wire _abc_15497_new_n1996_; 
wire _abc_15497_new_n1997_; 
wire _abc_15497_new_n1998_; 
wire _abc_15497_new_n1999_; 
wire _abc_15497_new_n2000_; 
wire _abc_15497_new_n2001_; 
wire _abc_15497_new_n2002_; 
wire _abc_15497_new_n2003_; 
wire _abc_15497_new_n2004_; 
wire _abc_15497_new_n2005_; 
wire _abc_15497_new_n2006_; 
wire _abc_15497_new_n2007_; 
wire _abc_15497_new_n2008_; 
wire _abc_15497_new_n2009_; 
wire _abc_15497_new_n2010_; 
wire _abc_15497_new_n2011_; 
wire _abc_15497_new_n2012_; 
wire _abc_15497_new_n2014_; 
wire _abc_15497_new_n2015_; 
wire _abc_15497_new_n2016_; 
wire _abc_15497_new_n2017_; 
wire _abc_15497_new_n2018_; 
wire _abc_15497_new_n2019_; 
wire _abc_15497_new_n2020_; 
wire _abc_15497_new_n2021_; 
wire _abc_15497_new_n2023_; 
wire _abc_15497_new_n2024_; 
wire _abc_15497_new_n2025_; 
wire _abc_15497_new_n2026_; 
wire _abc_15497_new_n2027_; 
wire _abc_15497_new_n2028_; 
wire _abc_15497_new_n2029_; 
wire _abc_15497_new_n2030_; 
wire _abc_15497_new_n2031_; 
wire _abc_15497_new_n2032_; 
wire _abc_15497_new_n2033_; 
wire _abc_15497_new_n2034_; 
wire _abc_15497_new_n2035_; 
wire _abc_15497_new_n2036_; 
wire _abc_15497_new_n2037_; 
wire _abc_15497_new_n2039_; 
wire _abc_15497_new_n2040_; 
wire _abc_15497_new_n2041_; 
wire _abc_15497_new_n2042_; 
wire _abc_15497_new_n2043_; 
wire _abc_15497_new_n2044_; 
wire _abc_15497_new_n2045_; 
wire _abc_15497_new_n2047_; 
wire _abc_15497_new_n2048_; 
wire _abc_15497_new_n2049_; 
wire _abc_15497_new_n2050_; 
wire _abc_15497_new_n2051_; 
wire _abc_15497_new_n2052_; 
wire _abc_15497_new_n2053_; 
wire _abc_15497_new_n2054_; 
wire _abc_15497_new_n2055_; 
wire _abc_15497_new_n2056_; 
wire _abc_15497_new_n2057_; 
wire _abc_15497_new_n2058_; 
wire _abc_15497_new_n2059_; 
wire _abc_15497_new_n2060_; 
wire _abc_15497_new_n2062_; 
wire _abc_15497_new_n2063_; 
wire _abc_15497_new_n2064_; 
wire _abc_15497_new_n2065_; 
wire _abc_15497_new_n2066_; 
wire _abc_15497_new_n2067_; 
wire _abc_15497_new_n2068_; 
wire _abc_15497_new_n2069_; 
wire _abc_15497_new_n2070_; 
wire _abc_15497_new_n2072_; 
wire _abc_15497_new_n2073_; 
wire _abc_15497_new_n2074_; 
wire _abc_15497_new_n2075_; 
wire _abc_15497_new_n2076_; 
wire _abc_15497_new_n2077_; 
wire _abc_15497_new_n2078_; 
wire _abc_15497_new_n2079_; 
wire _abc_15497_new_n2080_; 
wire _abc_15497_new_n2082_; 
wire _abc_15497_new_n2083_; 
wire _abc_15497_new_n2084_; 
wire _abc_15497_new_n2085_; 
wire _abc_15497_new_n2086_; 
wire _abc_15497_new_n2087_; 
wire _abc_15497_new_n2088_; 
wire _abc_15497_new_n2089_; 
wire _abc_15497_new_n2091_; 
wire _abc_15497_new_n2092_; 
wire _abc_15497_new_n2093_; 
wire _abc_15497_new_n2094_; 
wire _abc_15497_new_n2095_; 
wire _abc_15497_new_n2097_; 
wire _abc_15497_new_n2098_; 
wire _abc_15497_new_n2099_; 
wire _abc_15497_new_n2100_; 
wire _abc_15497_new_n2101_; 
wire _abc_15497_new_n2103_; 
wire _abc_15497_new_n2104_; 
wire _abc_15497_new_n2105_; 
wire _abc_15497_new_n2106_; 
wire _abc_15497_new_n2107_; 
wire _abc_15497_new_n2108_; 
wire _abc_15497_new_n2109_; 
wire _abc_15497_new_n2110_; 
wire _abc_15497_new_n2112_; 
wire _abc_15497_new_n2113_; 
wire _abc_15497_new_n2114_; 
wire _abc_15497_new_n2115_; 
wire _abc_15497_new_n2116_; 
wire _abc_15497_new_n2117_; 
wire _abc_15497_new_n2118_; 
wire _abc_15497_new_n2119_; 
wire _abc_15497_new_n2120_; 
wire _abc_15497_new_n2122_; 
wire _abc_15497_new_n2123_; 
wire _abc_15497_new_n2124_; 
wire _abc_15497_new_n2125_; 
wire _abc_15497_new_n2126_; 
wire _abc_15497_new_n2127_; 
wire _abc_15497_new_n2129_; 
wire _abc_15497_new_n2130_; 
wire _abc_15497_new_n2131_; 
wire _abc_15497_new_n2132_; 
wire _abc_15497_new_n2133_; 
wire _abc_15497_new_n2134_; 
wire _abc_15497_new_n2135_; 
wire _abc_15497_new_n2136_; 
wire _abc_15497_new_n2137_; 
wire _abc_15497_new_n2138_; 
wire _abc_15497_new_n2139_; 
wire _abc_15497_new_n2141_; 
wire _abc_15497_new_n2142_; 
wire _abc_15497_new_n2143_; 
wire _abc_15497_new_n2144_; 
wire _abc_15497_new_n2145_; 
wire _abc_15497_new_n2146_; 
wire _abc_15497_new_n2147_; 
wire _abc_15497_new_n2148_; 
wire _abc_15497_new_n2149_; 
wire _abc_15497_new_n2151_; 
wire _abc_15497_new_n2152_; 
wire _abc_15497_new_n2153_; 
wire _abc_15497_new_n2154_; 
wire _abc_15497_new_n2155_; 
wire _abc_15497_new_n2156_; 
wire _abc_15497_new_n2157_; 
wire _abc_15497_new_n2159_; 
wire _abc_15497_new_n2160_; 
wire _abc_15497_new_n2161_; 
wire _abc_15497_new_n2162_; 
wire _abc_15497_new_n2163_; 
wire _abc_15497_new_n2164_; 
wire _abc_15497_new_n2165_; 
wire _abc_15497_new_n2166_; 
wire _abc_15497_new_n2167_; 
wire _abc_15497_new_n2168_; 
wire _abc_15497_new_n2169_; 
wire _abc_15497_new_n2170_; 
wire _abc_15497_new_n2171_; 
wire _abc_15497_new_n2172_; 
wire _abc_15497_new_n2174_; 
wire _abc_15497_new_n2175_; 
wire _abc_15497_new_n2176_; 
wire _abc_15497_new_n2177_; 
wire _abc_15497_new_n2178_; 
wire _abc_15497_new_n2180_; 
wire _abc_15497_new_n2181_; 
wire _abc_15497_new_n2182_; 
wire _abc_15497_new_n2183_; 
wire _abc_15497_new_n2184_; 
wire _abc_15497_new_n2185_; 
wire _abc_15497_new_n2186_; 
wire _abc_15497_new_n2187_; 
wire _abc_15497_new_n2188_; 
wire _abc_15497_new_n2189_; 
wire _abc_15497_new_n2190_; 
wire _abc_15497_new_n2191_; 
wire _abc_15497_new_n2192_; 
wire _abc_15497_new_n2193_; 
wire _abc_15497_new_n2194_; 
wire _abc_15497_new_n2195_; 
wire _abc_15497_new_n2197_; 
wire _abc_15497_new_n2198_; 
wire _abc_15497_new_n2199_; 
wire _abc_15497_new_n2200_; 
wire _abc_15497_new_n2201_; 
wire _abc_15497_new_n2203_; 
wire _abc_15497_new_n2204_; 
wire _abc_15497_new_n2205_; 
wire _abc_15497_new_n2206_; 
wire _abc_15497_new_n2207_; 
wire _abc_15497_new_n2208_; 
wire _abc_15497_new_n2209_; 
wire _abc_15497_new_n2210_; 
wire _abc_15497_new_n2211_; 
wire _abc_15497_new_n2212_; 
wire _abc_15497_new_n2213_; 
wire _abc_15497_new_n2214_; 
wire _abc_15497_new_n2215_; 
wire _abc_15497_new_n2216_; 
wire _abc_15497_new_n2217_; 
wire _abc_15497_new_n2218_; 
wire _abc_15497_new_n2219_; 
wire _abc_15497_new_n2221_; 
wire _abc_15497_new_n2222_; 
wire _abc_15497_new_n2223_; 
wire _abc_15497_new_n2224_; 
wire _abc_15497_new_n2225_; 
wire _abc_15497_new_n2226_; 
wire _abc_15497_new_n2228_; 
wire _abc_15497_new_n2229_; 
wire _abc_15497_new_n2230_; 
wire _abc_15497_new_n2231_; 
wire _abc_15497_new_n2232_; 
wire _abc_15497_new_n2233_; 
wire _abc_15497_new_n2234_; 
wire _abc_15497_new_n2235_; 
wire _abc_15497_new_n2236_; 
wire _abc_15497_new_n2237_; 
wire _abc_15497_new_n2238_; 
wire _abc_15497_new_n2239_; 
wire _abc_15497_new_n2241_; 
wire _abc_15497_new_n2242_; 
wire _abc_15497_new_n2243_; 
wire _abc_15497_new_n2244_; 
wire _abc_15497_new_n2245_; 
wire _abc_15497_new_n2246_; 
wire _abc_15497_new_n2247_; 
wire _abc_15497_new_n2249_; 
wire _abc_15497_new_n2250_; 
wire _abc_15497_new_n2251_; 
wire _abc_15497_new_n2252_; 
wire _abc_15497_new_n2253_; 
wire _abc_15497_new_n2254_; 
wire _abc_15497_new_n2255_; 
wire _abc_15497_new_n2256_; 
wire _abc_15497_new_n2257_; 
wire _abc_15497_new_n2258_; 
wire _abc_15497_new_n2259_; 
wire _abc_15497_new_n2260_; 
wire _abc_15497_new_n2261_; 
wire _abc_15497_new_n2262_; 
wire _abc_15497_new_n2263_; 
wire _abc_15497_new_n2264_; 
wire _abc_15497_new_n2265_; 
wire _abc_15497_new_n2267_; 
wire _abc_15497_new_n2268_; 
wire _abc_15497_new_n2269_; 
wire _abc_15497_new_n2270_; 
wire _abc_15497_new_n2271_; 
wire _abc_15497_new_n2272_; 
wire _abc_15497_new_n2273_; 
wire _abc_15497_new_n2274_; 
wire _abc_15497_new_n2275_; 
wire _abc_15497_new_n2276_; 
wire _abc_15497_new_n2278_; 
wire _abc_15497_new_n2279_; 
wire _abc_15497_new_n2280_; 
wire _abc_15497_new_n2281_; 
wire _abc_15497_new_n2282_; 
wire _abc_15497_new_n2283_; 
wire _abc_15497_new_n2284_; 
wire _abc_15497_new_n2285_; 
wire _abc_15497_new_n2286_; 
wire _abc_15497_new_n2287_; 
wire _abc_15497_new_n2288_; 
wire _abc_15497_new_n2289_; 
wire _abc_15497_new_n2290_; 
wire _abc_15497_new_n2291_; 
wire _abc_15497_new_n2293_; 
wire _abc_15497_new_n2294_; 
wire _abc_15497_new_n2295_; 
wire _abc_15497_new_n2296_; 
wire _abc_15497_new_n2297_; 
wire _abc_15497_new_n2298_; 
wire _abc_15497_new_n2299_; 
wire _abc_15497_new_n2300_; 
wire _abc_15497_new_n2301_; 
wire _abc_15497_new_n2303_; 
wire _abc_15497_new_n2304_; 
wire _abc_15497_new_n2305_; 
wire _abc_15497_new_n2306_; 
wire _abc_15497_new_n2307_; 
wire _abc_15497_new_n2308_; 
wire _abc_15497_new_n2309_; 
wire _abc_15497_new_n2310_; 
wire _abc_15497_new_n2311_; 
wire _abc_15497_new_n2312_; 
wire _abc_15497_new_n2313_; 
wire _abc_15497_new_n2314_; 
wire _abc_15497_new_n2315_; 
wire _abc_15497_new_n2317_; 
wire _abc_15497_new_n2318_; 
wire _abc_15497_new_n2319_; 
wire _abc_15497_new_n2320_; 
wire _abc_15497_new_n2321_; 
wire _abc_15497_new_n2322_; 
wire _abc_15497_new_n2323_; 
wire _abc_15497_new_n2324_; 
wire _abc_15497_new_n2325_; 
wire _abc_15497_new_n2326_; 
wire _abc_15497_new_n2328_; 
wire _abc_15497_new_n2329_; 
wire _abc_15497_new_n2330_; 
wire _abc_15497_new_n2331_; 
wire _abc_15497_new_n2332_; 
wire _abc_15497_new_n2333_; 
wire _abc_15497_new_n2334_; 
wire _abc_15497_new_n2335_; 
wire _abc_15497_new_n2336_; 
wire _abc_15497_new_n2338_; 
wire _abc_15497_new_n2339_; 
wire _abc_15497_new_n2340_; 
wire _abc_15497_new_n2341_; 
wire _abc_15497_new_n2342_; 
wire _abc_15497_new_n2343_; 
wire _abc_15497_new_n2345_; 
wire _abc_15497_new_n2346_; 
wire _abc_15497_new_n2347_; 
wire _abc_15497_new_n2348_; 
wire _abc_15497_new_n2349_; 
wire _abc_15497_new_n2350_; 
wire _abc_15497_new_n2351_; 
wire _abc_15497_new_n2352_; 
wire _abc_15497_new_n2353_; 
wire _abc_15497_new_n2354_; 
wire _abc_15497_new_n2355_; 
wire _abc_15497_new_n2356_; 
wire _abc_15497_new_n2357_; 
wire _abc_15497_new_n2358_; 
wire _abc_15497_new_n2359_; 
wire _abc_15497_new_n2360_; 
wire _abc_15497_new_n2361_; 
wire _abc_15497_new_n2362_; 
wire _abc_15497_new_n2363_; 
wire _abc_15497_new_n2364_; 
wire _abc_15497_new_n2365_; 
wire _abc_15497_new_n2366_; 
wire _abc_15497_new_n2368_; 
wire _abc_15497_new_n2369_; 
wire _abc_15497_new_n2370_; 
wire _abc_15497_new_n2371_; 
wire _abc_15497_new_n2372_; 
wire _abc_15497_new_n2373_; 
wire _abc_15497_new_n2374_; 
wire _abc_15497_new_n2375_; 
wire _abc_15497_new_n2376_; 
wire _abc_15497_new_n2378_; 
wire _abc_15497_new_n2379_; 
wire _abc_15497_new_n2380_; 
wire _abc_15497_new_n2381_; 
wire _abc_15497_new_n2382_; 
wire _abc_15497_new_n2383_; 
wire _abc_15497_new_n2384_; 
wire _abc_15497_new_n2385_; 
wire _abc_15497_new_n2386_; 
wire _abc_15497_new_n2387_; 
wire _abc_15497_new_n2388_; 
wire _abc_15497_new_n2389_; 
wire _abc_15497_new_n2390_; 
wire _abc_15497_new_n2391_; 
wire _abc_15497_new_n2393_; 
wire _abc_15497_new_n2394_; 
wire _abc_15497_new_n2395_; 
wire _abc_15497_new_n2396_; 
wire _abc_15497_new_n2397_; 
wire _abc_15497_new_n2398_; 
wire _abc_15497_new_n2399_; 
wire _abc_15497_new_n2401_; 
wire _abc_15497_new_n2402_; 
wire _abc_15497_new_n2403_; 
wire _abc_15497_new_n2404_; 
wire _abc_15497_new_n2405_; 
wire _abc_15497_new_n2406_; 
wire _abc_15497_new_n2407_; 
wire _abc_15497_new_n2408_; 
wire _abc_15497_new_n2409_; 
wire _abc_15497_new_n2410_; 
wire _abc_15497_new_n2411_; 
wire _abc_15497_new_n2412_; 
wire _abc_15497_new_n2414_; 
wire _abc_15497_new_n2415_; 
wire _abc_15497_new_n2416_; 
wire _abc_15497_new_n2417_; 
wire _abc_15497_new_n2418_; 
wire _abc_15497_new_n2419_; 
wire _abc_15497_new_n2420_; 
wire _abc_15497_new_n2421_; 
wire _abc_15497_new_n2422_; 
wire _abc_15497_new_n2423_; 
wire _abc_15497_new_n2425_; 
wire _abc_15497_new_n2426_; 
wire _abc_15497_new_n2427_; 
wire _abc_15497_new_n2428_; 
wire _abc_15497_new_n2429_; 
wire _abc_15497_new_n2430_; 
wire _abc_15497_new_n2431_; 
wire _abc_15497_new_n2432_; 
wire _abc_15497_new_n2433_; 
wire _abc_15497_new_n2434_; 
wire _abc_15497_new_n2435_; 
wire _abc_15497_new_n2436_; 
wire _abc_15497_new_n2438_; 
wire _abc_15497_new_n2439_; 
wire _abc_15497_new_n2440_; 
wire _abc_15497_new_n2441_; 
wire _abc_15497_new_n2442_; 
wire _abc_15497_new_n2444_; 
wire _abc_15497_new_n2445_; 
wire _abc_15497_new_n2447_; 
wire _abc_15497_new_n2448_; 
wire _abc_15497_new_n2450_; 
wire _abc_15497_new_n2451_; 
wire _abc_15497_new_n2453_; 
wire _abc_15497_new_n2454_; 
wire _abc_15497_new_n2456_; 
wire _abc_15497_new_n2457_; 
wire _abc_15497_new_n2459_; 
wire _abc_15497_new_n2460_; 
wire _abc_15497_new_n2462_; 
wire _abc_15497_new_n2463_; 
wire _abc_15497_new_n2465_; 
wire _abc_15497_new_n2466_; 
wire _abc_15497_new_n2468_; 
wire _abc_15497_new_n2469_; 
wire _abc_15497_new_n2471_; 
wire _abc_15497_new_n2472_; 
wire _abc_15497_new_n2474_; 
wire _abc_15497_new_n2475_; 
wire _abc_15497_new_n2477_; 
wire _abc_15497_new_n2478_; 
wire _abc_15497_new_n2480_; 
wire _abc_15497_new_n2481_; 
wire _abc_15497_new_n2483_; 
wire _abc_15497_new_n2484_; 
wire _abc_15497_new_n2486_; 
wire _abc_15497_new_n2487_; 
wire _abc_15497_new_n2489_; 
wire _abc_15497_new_n2490_; 
wire _abc_15497_new_n2492_; 
wire _abc_15497_new_n2493_; 
wire _abc_15497_new_n2495_; 
wire _abc_15497_new_n2496_; 
wire _abc_15497_new_n2498_; 
wire _abc_15497_new_n2499_; 
wire _abc_15497_new_n2501_; 
wire _abc_15497_new_n2502_; 
wire _abc_15497_new_n2504_; 
wire _abc_15497_new_n2505_; 
wire _abc_15497_new_n2507_; 
wire _abc_15497_new_n2508_; 
wire _abc_15497_new_n2510_; 
wire _abc_15497_new_n2511_; 
wire _abc_15497_new_n2513_; 
wire _abc_15497_new_n2514_; 
wire _abc_15497_new_n2516_; 
wire _abc_15497_new_n2517_; 
wire _abc_15497_new_n2519_; 
wire _abc_15497_new_n2520_; 
wire _abc_15497_new_n2522_; 
wire _abc_15497_new_n2523_; 
wire _abc_15497_new_n2525_; 
wire _abc_15497_new_n2526_; 
wire _abc_15497_new_n2528_; 
wire _abc_15497_new_n2529_; 
wire _abc_15497_new_n2531_; 
wire _abc_15497_new_n2532_; 
wire _abc_15497_new_n2534_; 
wire _abc_15497_new_n2535_; 
wire _abc_15497_new_n2537_; 
wire _abc_15497_new_n2538_; 
wire _abc_15497_new_n2540_; 
wire _abc_15497_new_n2541_; 
wire _abc_15497_new_n2543_; 
wire _abc_15497_new_n2544_; 
wire _abc_15497_new_n2546_; 
wire _abc_15497_new_n2547_; 
wire _abc_15497_new_n2549_; 
wire _abc_15497_new_n2550_; 
wire _abc_15497_new_n2552_; 
wire _abc_15497_new_n2553_; 
wire _abc_15497_new_n2555_; 
wire _abc_15497_new_n2556_; 
wire _abc_15497_new_n2558_; 
wire _abc_15497_new_n2559_; 
wire _abc_15497_new_n2561_; 
wire _abc_15497_new_n2562_; 
wire _abc_15497_new_n2564_; 
wire _abc_15497_new_n2565_; 
wire _abc_15497_new_n2567_; 
wire _abc_15497_new_n2568_; 
wire _abc_15497_new_n2570_; 
wire _abc_15497_new_n2571_; 
wire _abc_15497_new_n2573_; 
wire _abc_15497_new_n2574_; 
wire _abc_15497_new_n2576_; 
wire _abc_15497_new_n2577_; 
wire _abc_15497_new_n2579_; 
wire _abc_15497_new_n2580_; 
wire _abc_15497_new_n2582_; 
wire _abc_15497_new_n2583_; 
wire _abc_15497_new_n2585_; 
wire _abc_15497_new_n2586_; 
wire _abc_15497_new_n2588_; 
wire _abc_15497_new_n2589_; 
wire _abc_15497_new_n2591_; 
wire _abc_15497_new_n2592_; 
wire _abc_15497_new_n2594_; 
wire _abc_15497_new_n2595_; 
wire _abc_15497_new_n2597_; 
wire _abc_15497_new_n2598_; 
wire _abc_15497_new_n2600_; 
wire _abc_15497_new_n2601_; 
wire _abc_15497_new_n2603_; 
wire _abc_15497_new_n2604_; 
wire _abc_15497_new_n2606_; 
wire _abc_15497_new_n2607_; 
wire _abc_15497_new_n2609_; 
wire _abc_15497_new_n2610_; 
wire _abc_15497_new_n2612_; 
wire _abc_15497_new_n2613_; 
wire _abc_15497_new_n2615_; 
wire _abc_15497_new_n2616_; 
wire _abc_15497_new_n2618_; 
wire _abc_15497_new_n2619_; 
wire _abc_15497_new_n2621_; 
wire _abc_15497_new_n2622_; 
wire _abc_15497_new_n2624_; 
wire _abc_15497_new_n2625_; 
wire _abc_15497_new_n2627_; 
wire _abc_15497_new_n2628_; 
wire _abc_15497_new_n2630_; 
wire _abc_15497_new_n2631_; 
wire _abc_15497_new_n2632_; 
wire _abc_15497_new_n2634_; 
wire _abc_15497_new_n2635_; 
wire _abc_15497_new_n2636_; 
wire _abc_15497_new_n2637_; 
wire _abc_15497_new_n2639_; 
wire _abc_15497_new_n2640_; 
wire _abc_15497_new_n2642_; 
wire _abc_15497_new_n2643_; 
wire _abc_15497_new_n2645_; 
wire _abc_15497_new_n2646_; 
wire _abc_15497_new_n2648_; 
wire _abc_15497_new_n2649_; 
wire _abc_15497_new_n2651_; 
wire _abc_15497_new_n2652_; 
wire _abc_15497_new_n2654_; 
wire _abc_15497_new_n2655_; 
wire _abc_15497_new_n2657_; 
wire _abc_15497_new_n2658_; 
wire _abc_15497_new_n2660_; 
wire _abc_15497_new_n2661_; 
wire _abc_15497_new_n2663_; 
wire _abc_15497_new_n2664_; 
wire _abc_15497_new_n2666_; 
wire _abc_15497_new_n2667_; 
wire _abc_15497_new_n2669_; 
wire _abc_15497_new_n2670_; 
wire _abc_15497_new_n2672_; 
wire _abc_15497_new_n2673_; 
wire _abc_15497_new_n2675_; 
wire _abc_15497_new_n2676_; 
wire _abc_15497_new_n2678_; 
wire _abc_15497_new_n2679_; 
wire _abc_15497_new_n2681_; 
wire _abc_15497_new_n2682_; 
wire _abc_15497_new_n2684_; 
wire _abc_15497_new_n2685_; 
wire _abc_15497_new_n2687_; 
wire _abc_15497_new_n2688_; 
wire _abc_15497_new_n2690_; 
wire _abc_15497_new_n2691_; 
wire _abc_15497_new_n2693_; 
wire _abc_15497_new_n2694_; 
wire _abc_15497_new_n2696_; 
wire _abc_15497_new_n2697_; 
wire _abc_15497_new_n2699_; 
wire _abc_15497_new_n2700_; 
wire _abc_15497_new_n2702_; 
wire _abc_15497_new_n2703_; 
wire _abc_15497_new_n2705_; 
wire _abc_15497_new_n2706_; 
wire _abc_15497_new_n2708_; 
wire _abc_15497_new_n2709_; 
wire _abc_15497_new_n2711_; 
wire _abc_15497_new_n2712_; 
wire _abc_15497_new_n2714_; 
wire _abc_15497_new_n2715_; 
wire _abc_15497_new_n2717_; 
wire _abc_15497_new_n2718_; 
wire _abc_15497_new_n2720_; 
wire _abc_15497_new_n2721_; 
wire _abc_15497_new_n2723_; 
wire _abc_15497_new_n2724_; 
wire _abc_15497_new_n2726_; 
wire _abc_15497_new_n2727_; 
wire _abc_15497_new_n2729_; 
wire _abc_15497_new_n2730_; 
wire _abc_15497_new_n2732_; 
wire _abc_15497_new_n2733_; 
wire _abc_15497_new_n2735_; 
wire _abc_15497_new_n2736_; 
wire _abc_15497_new_n2737_; 
wire _abc_15497_new_n2738_; 
wire _abc_15497_new_n2739_; 
wire _abc_15497_new_n2740_; 
wire _abc_15497_new_n2741_; 
wire _abc_15497_new_n2742_; 
wire _abc_15497_new_n2742__bF_buf0; 
wire _abc_15497_new_n2742__bF_buf1; 
wire _abc_15497_new_n2742__bF_buf2; 
wire _abc_15497_new_n2742__bF_buf3; 
wire _abc_15497_new_n2743_; 
wire _abc_15497_new_n2743__bF_buf0; 
wire _abc_15497_new_n2743__bF_buf1; 
wire _abc_15497_new_n2743__bF_buf2; 
wire _abc_15497_new_n2743__bF_buf3; 
wire _abc_15497_new_n2743__bF_buf4; 
wire _abc_15497_new_n2743__bF_buf5; 
wire _abc_15497_new_n2744_; 
wire _abc_15497_new_n2745_; 
wire _abc_15497_new_n2746_; 
wire _abc_15497_new_n2747_; 
wire _abc_15497_new_n2748_; 
wire _abc_15497_new_n2749_; 
wire _abc_15497_new_n2750_; 
wire _abc_15497_new_n2751_; 
wire _abc_15497_new_n2752_; 
wire _abc_15497_new_n2753_; 
wire _abc_15497_new_n2754_; 
wire _abc_15497_new_n2755_; 
wire _abc_15497_new_n2756_; 
wire _abc_15497_new_n2756__bF_buf0; 
wire _abc_15497_new_n2756__bF_buf1; 
wire _abc_15497_new_n2756__bF_buf2; 
wire _abc_15497_new_n2756__bF_buf3; 
wire _abc_15497_new_n2756__bF_buf4; 
wire _abc_15497_new_n2757_; 
wire _abc_15497_new_n2758_; 
wire _abc_15497_new_n2759_; 
wire _abc_15497_new_n2759__bF_buf0; 
wire _abc_15497_new_n2759__bF_buf1; 
wire _abc_15497_new_n2759__bF_buf2; 
wire _abc_15497_new_n2759__bF_buf3; 
wire _abc_15497_new_n2759__bF_buf4; 
wire _abc_15497_new_n2759__bF_buf5; 
wire _abc_15497_new_n2760_; 
wire _abc_15497_new_n2761_; 
wire _abc_15497_new_n2762_; 
wire _abc_15497_new_n2763_; 
wire _abc_15497_new_n2764_; 
wire _abc_15497_new_n2765_; 
wire _abc_15497_new_n2766_; 
wire _abc_15497_new_n2767_; 
wire _abc_15497_new_n2768_; 
wire _abc_15497_new_n2769_; 
wire _abc_15497_new_n2770_; 
wire _abc_15497_new_n2771_; 
wire _abc_15497_new_n2772_; 
wire _abc_15497_new_n2773_; 
wire _abc_15497_new_n2774_; 
wire _abc_15497_new_n2775_; 
wire _abc_15497_new_n2776_; 
wire _abc_15497_new_n2777_; 
wire _abc_15497_new_n2778_; 
wire _abc_15497_new_n2780_; 
wire _abc_15497_new_n2780__bF_buf0; 
wire _abc_15497_new_n2780__bF_buf1; 
wire _abc_15497_new_n2780__bF_buf2; 
wire _abc_15497_new_n2780__bF_buf3; 
wire _abc_15497_new_n2781_; 
wire _abc_15497_new_n2781__bF_buf0; 
wire _abc_15497_new_n2781__bF_buf1; 
wire _abc_15497_new_n2781__bF_buf2; 
wire _abc_15497_new_n2781__bF_buf3; 
wire _abc_15497_new_n2782_; 
wire _abc_15497_new_n2783_; 
wire _abc_15497_new_n2784_; 
wire _abc_15497_new_n2785_; 
wire _abc_15497_new_n2786_; 
wire _abc_15497_new_n2787_; 
wire _abc_15497_new_n2788_; 
wire _abc_15497_new_n2789_; 
wire _abc_15497_new_n2790_; 
wire _abc_15497_new_n2791_; 
wire _abc_15497_new_n2792_; 
wire _abc_15497_new_n2793_; 
wire _abc_15497_new_n2794_; 
wire _abc_15497_new_n2795_; 
wire _abc_15497_new_n2796_; 
wire _abc_15497_new_n2797_; 
wire _abc_15497_new_n2798_; 
wire _abc_15497_new_n2799_; 
wire _abc_15497_new_n2800_; 
wire _abc_15497_new_n2801_; 
wire _abc_15497_new_n2802_; 
wire _abc_15497_new_n2803_; 
wire _abc_15497_new_n2804_; 
wire _abc_15497_new_n2805_; 
wire _abc_15497_new_n2806_; 
wire _abc_15497_new_n2807_; 
wire _abc_15497_new_n2808_; 
wire _abc_15497_new_n2809_; 
wire _abc_15497_new_n2810_; 
wire _abc_15497_new_n2811_; 
wire _abc_15497_new_n2812_; 
wire _abc_15497_new_n2813_; 
wire _abc_15497_new_n2814_; 
wire _abc_15497_new_n2815_; 
wire _abc_15497_new_n2816_; 
wire _abc_15497_new_n2817_; 
wire _abc_15497_new_n2818_; 
wire _abc_15497_new_n2819_; 
wire _abc_15497_new_n2820_; 
wire _abc_15497_new_n2821_; 
wire _abc_15497_new_n2822_; 
wire _abc_15497_new_n2823_; 
wire _abc_15497_new_n2824_; 
wire _abc_15497_new_n2826_; 
wire _abc_15497_new_n2827_; 
wire _abc_15497_new_n2828_; 
wire _abc_15497_new_n2829_; 
wire _abc_15497_new_n2830_; 
wire _abc_15497_new_n2831_; 
wire _abc_15497_new_n2832_; 
wire _abc_15497_new_n2833_; 
wire _abc_15497_new_n2834_; 
wire _abc_15497_new_n2835_; 
wire _abc_15497_new_n2836_; 
wire _abc_15497_new_n2837_; 
wire _abc_15497_new_n2838_; 
wire _abc_15497_new_n2839_; 
wire _abc_15497_new_n2840_; 
wire _abc_15497_new_n2841_; 
wire _abc_15497_new_n2842_; 
wire _abc_15497_new_n2843_; 
wire _abc_15497_new_n2844_; 
wire _abc_15497_new_n2845_; 
wire _abc_15497_new_n2846_; 
wire _abc_15497_new_n2847_; 
wire _abc_15497_new_n2848_; 
wire _abc_15497_new_n2849_; 
wire _abc_15497_new_n2850_; 
wire _abc_15497_new_n2851_; 
wire _abc_15497_new_n2852_; 
wire _abc_15497_new_n2853_; 
wire _abc_15497_new_n2854_; 
wire _abc_15497_new_n2855_; 
wire _abc_15497_new_n2856_; 
wire _abc_15497_new_n2857_; 
wire _abc_15497_new_n2858_; 
wire _abc_15497_new_n2859_; 
wire _abc_15497_new_n2860_; 
wire _abc_15497_new_n2861_; 
wire _abc_15497_new_n2862_; 
wire _abc_15497_new_n2863_; 
wire _abc_15497_new_n2864_; 
wire _abc_15497_new_n2865_; 
wire _abc_15497_new_n2866_; 
wire _abc_15497_new_n2867_; 
wire _abc_15497_new_n2868_; 
wire _abc_15497_new_n2869_; 
wire _abc_15497_new_n2870_; 
wire _abc_15497_new_n2871_; 
wire _abc_15497_new_n2872_; 
wire _abc_15497_new_n2873_; 
wire _abc_15497_new_n2874_; 
wire _abc_15497_new_n2875_; 
wire _abc_15497_new_n2876_; 
wire _abc_15497_new_n2877_; 
wire _abc_15497_new_n2878_; 
wire _abc_15497_new_n2879_; 
wire _abc_15497_new_n2880_; 
wire _abc_15497_new_n2881_; 
wire _abc_15497_new_n2883_; 
wire _abc_15497_new_n2884_; 
wire _abc_15497_new_n2885_; 
wire _abc_15497_new_n2886_; 
wire _abc_15497_new_n2887_; 
wire _abc_15497_new_n2888_; 
wire _abc_15497_new_n2889_; 
wire _abc_15497_new_n2890_; 
wire _abc_15497_new_n2891_; 
wire _abc_15497_new_n2892_; 
wire _abc_15497_new_n2893_; 
wire _abc_15497_new_n2894_; 
wire _abc_15497_new_n2895_; 
wire _abc_15497_new_n2896_; 
wire _abc_15497_new_n2897_; 
wire _abc_15497_new_n2898_; 
wire _abc_15497_new_n2899_; 
wire _abc_15497_new_n2900_; 
wire _abc_15497_new_n2901_; 
wire _abc_15497_new_n2902_; 
wire _abc_15497_new_n2903_; 
wire _abc_15497_new_n2904_; 
wire _abc_15497_new_n2905_; 
wire _abc_15497_new_n2906_; 
wire _abc_15497_new_n2907_; 
wire _abc_15497_new_n2908_; 
wire _abc_15497_new_n2909_; 
wire _abc_15497_new_n2910_; 
wire _abc_15497_new_n2911_; 
wire _abc_15497_new_n2912_; 
wire _abc_15497_new_n2913_; 
wire _abc_15497_new_n2914_; 
wire _abc_15497_new_n2915_; 
wire _abc_15497_new_n2916_; 
wire _abc_15497_new_n2917_; 
wire _abc_15497_new_n2918_; 
wire _abc_15497_new_n2919_; 
wire _abc_15497_new_n2920_; 
wire _abc_15497_new_n2921_; 
wire _abc_15497_new_n2922_; 
wire _abc_15497_new_n2923_; 
wire _abc_15497_new_n2924_; 
wire _abc_15497_new_n2924__bF_buf0; 
wire _abc_15497_new_n2924__bF_buf1; 
wire _abc_15497_new_n2924__bF_buf2; 
wire _abc_15497_new_n2924__bF_buf3; 
wire _abc_15497_new_n2924__bF_buf4; 
wire _abc_15497_new_n2925_; 
wire _abc_15497_new_n2925__bF_buf0; 
wire _abc_15497_new_n2925__bF_buf1; 
wire _abc_15497_new_n2925__bF_buf2; 
wire _abc_15497_new_n2925__bF_buf3; 
wire _abc_15497_new_n2926_; 
wire _abc_15497_new_n2927_; 
wire _abc_15497_new_n2928_; 
wire _abc_15497_new_n2929_; 
wire _abc_15497_new_n2930_; 
wire _abc_15497_new_n2931_; 
wire _abc_15497_new_n2932_; 
wire _abc_15497_new_n2933_; 
wire _abc_15497_new_n2934_; 
wire _abc_15497_new_n2935_; 
wire _abc_15497_new_n2936_; 
wire _abc_15497_new_n2937_; 
wire _abc_15497_new_n2938_; 
wire _abc_15497_new_n2940_; 
wire _abc_15497_new_n2941_; 
wire _abc_15497_new_n2942_; 
wire _abc_15497_new_n2943_; 
wire _abc_15497_new_n2944_; 
wire _abc_15497_new_n2945_; 
wire _abc_15497_new_n2946_; 
wire _abc_15497_new_n2947_; 
wire _abc_15497_new_n2948_; 
wire _abc_15497_new_n2949_; 
wire _abc_15497_new_n2950_; 
wire _abc_15497_new_n2951_; 
wire _abc_15497_new_n2952_; 
wire _abc_15497_new_n2953_; 
wire _abc_15497_new_n2954_; 
wire _abc_15497_new_n2955_; 
wire _abc_15497_new_n2956_; 
wire _abc_15497_new_n2957_; 
wire _abc_15497_new_n2958_; 
wire _abc_15497_new_n2959_; 
wire _abc_15497_new_n2960_; 
wire _abc_15497_new_n2961_; 
wire _abc_15497_new_n2962_; 
wire _abc_15497_new_n2963_; 
wire _abc_15497_new_n2964_; 
wire _abc_15497_new_n2965_; 
wire _abc_15497_new_n2966_; 
wire _abc_15497_new_n2967_; 
wire _abc_15497_new_n2968_; 
wire _abc_15497_new_n2969_; 
wire _abc_15497_new_n2970_; 
wire _abc_15497_new_n2971_; 
wire _abc_15497_new_n2972_; 
wire _abc_15497_new_n2973_; 
wire _abc_15497_new_n2974_; 
wire _abc_15497_new_n2975_; 
wire _abc_15497_new_n2976_; 
wire _abc_15497_new_n2977_; 
wire _abc_15497_new_n2978_; 
wire _abc_15497_new_n2979_; 
wire _abc_15497_new_n2980_; 
wire _abc_15497_new_n2981_; 
wire _abc_15497_new_n2982_; 
wire _abc_15497_new_n2983_; 
wire _abc_15497_new_n2984_; 
wire _abc_15497_new_n2985_; 
wire _abc_15497_new_n2986_; 
wire _abc_15497_new_n2987_; 
wire _abc_15497_new_n2988_; 
wire _abc_15497_new_n2989_; 
wire _abc_15497_new_n2990_; 
wire _abc_15497_new_n2991_; 
wire _abc_15497_new_n2992_; 
wire _abc_15497_new_n2993_; 
wire _abc_15497_new_n2994_; 
wire _abc_15497_new_n2995_; 
wire _abc_15497_new_n2996_; 
wire _abc_15497_new_n2997_; 
wire _abc_15497_new_n2998_; 
wire _abc_15497_new_n2999_; 
wire _abc_15497_new_n3000_; 
wire _abc_15497_new_n3002_; 
wire _abc_15497_new_n3003_; 
wire _abc_15497_new_n3004_; 
wire _abc_15497_new_n3005_; 
wire _abc_15497_new_n3006_; 
wire _abc_15497_new_n3007_; 
wire _abc_15497_new_n3008_; 
wire _abc_15497_new_n3009_; 
wire _abc_15497_new_n3010_; 
wire _abc_15497_new_n3011_; 
wire _abc_15497_new_n3012_; 
wire _abc_15497_new_n3013_; 
wire _abc_15497_new_n3014_; 
wire _abc_15497_new_n3015_; 
wire _abc_15497_new_n3016_; 
wire _abc_15497_new_n3017_; 
wire _abc_15497_new_n3018_; 
wire _abc_15497_new_n3019_; 
wire _abc_15497_new_n3020_; 
wire _abc_15497_new_n3021_; 
wire _abc_15497_new_n3022_; 
wire _abc_15497_new_n3023_; 
wire _abc_15497_new_n3024_; 
wire _abc_15497_new_n3025_; 
wire _abc_15497_new_n3026_; 
wire _abc_15497_new_n3027_; 
wire _abc_15497_new_n3028_; 
wire _abc_15497_new_n3029_; 
wire _abc_15497_new_n3030_; 
wire _abc_15497_new_n3031_; 
wire _abc_15497_new_n3032_; 
wire _abc_15497_new_n3033_; 
wire _abc_15497_new_n3034_; 
wire _abc_15497_new_n3035_; 
wire _abc_15497_new_n3036_; 
wire _abc_15497_new_n3037_; 
wire _abc_15497_new_n3038_; 
wire _abc_15497_new_n3039_; 
wire _abc_15497_new_n3040_; 
wire _abc_15497_new_n3041_; 
wire _abc_15497_new_n3042_; 
wire _abc_15497_new_n3043_; 
wire _abc_15497_new_n3044_; 
wire _abc_15497_new_n3045_; 
wire _abc_15497_new_n3046_; 
wire _abc_15497_new_n3047_; 
wire _abc_15497_new_n3048_; 
wire _abc_15497_new_n3049_; 
wire _abc_15497_new_n3050_; 
wire _abc_15497_new_n3051_; 
wire _abc_15497_new_n3052_; 
wire _abc_15497_new_n3053_; 
wire _abc_15497_new_n3054_; 
wire _abc_15497_new_n3055_; 
wire _abc_15497_new_n3056_; 
wire _abc_15497_new_n3058_; 
wire _abc_15497_new_n3059_; 
wire _abc_15497_new_n3060_; 
wire _abc_15497_new_n3061_; 
wire _abc_15497_new_n3062_; 
wire _abc_15497_new_n3063_; 
wire _abc_15497_new_n3064_; 
wire _abc_15497_new_n3065_; 
wire _abc_15497_new_n3066_; 
wire _abc_15497_new_n3067_; 
wire _abc_15497_new_n3068_; 
wire _abc_15497_new_n3069_; 
wire _abc_15497_new_n3070_; 
wire _abc_15497_new_n3071_; 
wire _abc_15497_new_n3072_; 
wire _abc_15497_new_n3073_; 
wire _abc_15497_new_n3074_; 
wire _abc_15497_new_n3075_; 
wire _abc_15497_new_n3076_; 
wire _abc_15497_new_n3077_; 
wire _abc_15497_new_n3078_; 
wire _abc_15497_new_n3079_; 
wire _abc_15497_new_n3080_; 
wire _abc_15497_new_n3081_; 
wire _abc_15497_new_n3082_; 
wire _abc_15497_new_n3083_; 
wire _abc_15497_new_n3084_; 
wire _abc_15497_new_n3085_; 
wire _abc_15497_new_n3086_; 
wire _abc_15497_new_n3087_; 
wire _abc_15497_new_n3088_; 
wire _abc_15497_new_n3089_; 
wire _abc_15497_new_n3090_; 
wire _abc_15497_new_n3091_; 
wire _abc_15497_new_n3092_; 
wire _abc_15497_new_n3093_; 
wire _abc_15497_new_n3094_; 
wire _abc_15497_new_n3095_; 
wire _abc_15497_new_n3096_; 
wire _abc_15497_new_n3097_; 
wire _abc_15497_new_n3098_; 
wire _abc_15497_new_n3099_; 
wire _abc_15497_new_n3100_; 
wire _abc_15497_new_n3101_; 
wire _abc_15497_new_n3102_; 
wire _abc_15497_new_n3103_; 
wire _abc_15497_new_n3104_; 
wire _abc_15497_new_n3105_; 
wire _abc_15497_new_n3106_; 
wire _abc_15497_new_n3107_; 
wire _abc_15497_new_n3108_; 
wire _abc_15497_new_n3109_; 
wire _abc_15497_new_n3110_; 
wire _abc_15497_new_n3111_; 
wire _abc_15497_new_n3112_; 
wire _abc_15497_new_n3113_; 
wire _abc_15497_new_n3114_; 
wire _abc_15497_new_n3116_; 
wire _abc_15497_new_n3117_; 
wire _abc_15497_new_n3118_; 
wire _abc_15497_new_n3119_; 
wire _abc_15497_new_n3120_; 
wire _abc_15497_new_n3121_; 
wire _abc_15497_new_n3122_; 
wire _abc_15497_new_n3123_; 
wire _abc_15497_new_n3124_; 
wire _abc_15497_new_n3125_; 
wire _abc_15497_new_n3126_; 
wire _abc_15497_new_n3127_; 
wire _abc_15497_new_n3128_; 
wire _abc_15497_new_n3129_; 
wire _abc_15497_new_n3130_; 
wire _abc_15497_new_n3131_; 
wire _abc_15497_new_n3132_; 
wire _abc_15497_new_n3133_; 
wire _abc_15497_new_n3134_; 
wire _abc_15497_new_n3135_; 
wire _abc_15497_new_n3136_; 
wire _abc_15497_new_n3137_; 
wire _abc_15497_new_n3138_; 
wire _abc_15497_new_n3139_; 
wire _abc_15497_new_n3140_; 
wire _abc_15497_new_n3141_; 
wire _abc_15497_new_n3142_; 
wire _abc_15497_new_n3143_; 
wire _abc_15497_new_n3144_; 
wire _abc_15497_new_n3145_; 
wire _abc_15497_new_n3146_; 
wire _abc_15497_new_n3147_; 
wire _abc_15497_new_n3148_; 
wire _abc_15497_new_n3149_; 
wire _abc_15497_new_n3150_; 
wire _abc_15497_new_n3151_; 
wire _abc_15497_new_n3152_; 
wire _abc_15497_new_n3153_; 
wire _abc_15497_new_n3154_; 
wire _abc_15497_new_n3155_; 
wire _abc_15497_new_n3156_; 
wire _abc_15497_new_n3157_; 
wire _abc_15497_new_n3158_; 
wire _abc_15497_new_n3159_; 
wire _abc_15497_new_n3160_; 
wire _abc_15497_new_n3161_; 
wire _abc_15497_new_n3162_; 
wire _abc_15497_new_n3163_; 
wire _abc_15497_new_n3164_; 
wire _abc_15497_new_n3165_; 
wire _abc_15497_new_n3167_; 
wire _abc_15497_new_n3168_; 
wire _abc_15497_new_n3169_; 
wire _abc_15497_new_n3170_; 
wire _abc_15497_new_n3171_; 
wire _abc_15497_new_n3172_; 
wire _abc_15497_new_n3173_; 
wire _abc_15497_new_n3174_; 
wire _abc_15497_new_n3175_; 
wire _abc_15497_new_n3176_; 
wire _abc_15497_new_n3177_; 
wire _abc_15497_new_n3178_; 
wire _abc_15497_new_n3179_; 
wire _abc_15497_new_n3180_; 
wire _abc_15497_new_n3181_; 
wire _abc_15497_new_n3182_; 
wire _abc_15497_new_n3183_; 
wire _abc_15497_new_n3184_; 
wire _abc_15497_new_n3185_; 
wire _abc_15497_new_n3186_; 
wire _abc_15497_new_n3187_; 
wire _abc_15497_new_n3188_; 
wire _abc_15497_new_n3189_; 
wire _abc_15497_new_n3190_; 
wire _abc_15497_new_n3191_; 
wire _abc_15497_new_n3192_; 
wire _abc_15497_new_n3193_; 
wire _abc_15497_new_n3194_; 
wire _abc_15497_new_n3195_; 
wire _abc_15497_new_n3196_; 
wire _abc_15497_new_n3197_; 
wire _abc_15497_new_n3198_; 
wire _abc_15497_new_n3199_; 
wire _abc_15497_new_n3200_; 
wire _abc_15497_new_n3201_; 
wire _abc_15497_new_n3202_; 
wire _abc_15497_new_n3203_; 
wire _abc_15497_new_n3204_; 
wire _abc_15497_new_n3205_; 
wire _abc_15497_new_n3206_; 
wire _abc_15497_new_n3207_; 
wire _abc_15497_new_n3208_; 
wire _abc_15497_new_n3209_; 
wire _abc_15497_new_n3210_; 
wire _abc_15497_new_n3211_; 
wire _abc_15497_new_n3212_; 
wire _abc_15497_new_n3213_; 
wire _abc_15497_new_n3214_; 
wire _abc_15497_new_n3215_; 
wire _abc_15497_new_n3216_; 
wire _abc_15497_new_n3217_; 
wire _abc_15497_new_n3218_; 
wire _abc_15497_new_n3219_; 
wire _abc_15497_new_n3220_; 
wire _abc_15497_new_n3221_; 
wire _abc_15497_new_n3222_; 
wire _abc_15497_new_n3224_; 
wire _abc_15497_new_n3225_; 
wire _abc_15497_new_n3226_; 
wire _abc_15497_new_n3227_; 
wire _abc_15497_new_n3228_; 
wire _abc_15497_new_n3229_; 
wire _abc_15497_new_n3230_; 
wire _abc_15497_new_n3231_; 
wire _abc_15497_new_n3232_; 
wire _abc_15497_new_n3233_; 
wire _abc_15497_new_n3234_; 
wire _abc_15497_new_n3235_; 
wire _abc_15497_new_n3236_; 
wire _abc_15497_new_n3237_; 
wire _abc_15497_new_n3238_; 
wire _abc_15497_new_n3239_; 
wire _abc_15497_new_n3240_; 
wire _abc_15497_new_n3241_; 
wire _abc_15497_new_n3242_; 
wire _abc_15497_new_n3243_; 
wire _abc_15497_new_n3244_; 
wire _abc_15497_new_n3245_; 
wire _abc_15497_new_n3246_; 
wire _abc_15497_new_n3247_; 
wire _abc_15497_new_n3248_; 
wire _abc_15497_new_n3249_; 
wire _abc_15497_new_n3250_; 
wire _abc_15497_new_n3251_; 
wire _abc_15497_new_n3252_; 
wire _abc_15497_new_n3253_; 
wire _abc_15497_new_n3254_; 
wire _abc_15497_new_n3255_; 
wire _abc_15497_new_n3256_; 
wire _abc_15497_new_n3257_; 
wire _abc_15497_new_n3258_; 
wire _abc_15497_new_n3259_; 
wire _abc_15497_new_n3260_; 
wire _abc_15497_new_n3261_; 
wire _abc_15497_new_n3262_; 
wire _abc_15497_new_n3263_; 
wire _abc_15497_new_n3264_; 
wire _abc_15497_new_n3265_; 
wire _abc_15497_new_n3266_; 
wire _abc_15497_new_n3267_; 
wire _abc_15497_new_n3268_; 
wire _abc_15497_new_n3269_; 
wire _abc_15497_new_n3270_; 
wire _abc_15497_new_n3271_; 
wire _abc_15497_new_n3272_; 
wire _abc_15497_new_n3273_; 
wire _abc_15497_new_n3274_; 
wire _abc_15497_new_n3275_; 
wire _abc_15497_new_n3276_; 
wire _abc_15497_new_n3277_; 
wire _abc_15497_new_n3278_; 
wire _abc_15497_new_n3279_; 
wire _abc_15497_new_n3280_; 
wire _abc_15497_new_n3281_; 
wire _abc_15497_new_n3283_; 
wire _abc_15497_new_n3284_; 
wire _abc_15497_new_n3285_; 
wire _abc_15497_new_n3286_; 
wire _abc_15497_new_n3287_; 
wire _abc_15497_new_n3288_; 
wire _abc_15497_new_n3289_; 
wire _abc_15497_new_n3290_; 
wire _abc_15497_new_n3291_; 
wire _abc_15497_new_n3292_; 
wire _abc_15497_new_n3293_; 
wire _abc_15497_new_n3294_; 
wire _abc_15497_new_n3295_; 
wire _abc_15497_new_n3296_; 
wire _abc_15497_new_n3297_; 
wire _abc_15497_new_n3298_; 
wire _abc_15497_new_n3299_; 
wire _abc_15497_new_n3300_; 
wire _abc_15497_new_n3301_; 
wire _abc_15497_new_n3302_; 
wire _abc_15497_new_n3303_; 
wire _abc_15497_new_n3304_; 
wire _abc_15497_new_n3305_; 
wire _abc_15497_new_n3306_; 
wire _abc_15497_new_n3307_; 
wire _abc_15497_new_n3308_; 
wire _abc_15497_new_n3309_; 
wire _abc_15497_new_n3310_; 
wire _abc_15497_new_n3311_; 
wire _abc_15497_new_n3312_; 
wire _abc_15497_new_n3313_; 
wire _abc_15497_new_n3314_; 
wire _abc_15497_new_n3315_; 
wire _abc_15497_new_n3316_; 
wire _abc_15497_new_n3317_; 
wire _abc_15497_new_n3318_; 
wire _abc_15497_new_n3319_; 
wire _abc_15497_new_n3320_; 
wire _abc_15497_new_n3321_; 
wire _abc_15497_new_n3322_; 
wire _abc_15497_new_n3323_; 
wire _abc_15497_new_n3324_; 
wire _abc_15497_new_n3325_; 
wire _abc_15497_new_n3326_; 
wire _abc_15497_new_n3327_; 
wire _abc_15497_new_n3328_; 
wire _abc_15497_new_n3329_; 
wire _abc_15497_new_n3330_; 
wire _abc_15497_new_n3331_; 
wire _abc_15497_new_n3332_; 
wire _abc_15497_new_n3333_; 
wire _abc_15497_new_n3334_; 
wire _abc_15497_new_n3335_; 
wire _abc_15497_new_n3336_; 
wire _abc_15497_new_n3337_; 
wire _abc_15497_new_n3338_; 
wire _abc_15497_new_n3339_; 
wire _abc_15497_new_n3340_; 
wire _abc_15497_new_n3341_; 
wire _abc_15497_new_n3342_; 
wire _abc_15497_new_n3343_; 
wire _abc_15497_new_n3344_; 
wire _abc_15497_new_n3345_; 
wire _abc_15497_new_n3346_; 
wire _abc_15497_new_n3348_; 
wire _abc_15497_new_n3349_; 
wire _abc_15497_new_n3350_; 
wire _abc_15497_new_n3351_; 
wire _abc_15497_new_n3352_; 
wire _abc_15497_new_n3353_; 
wire _abc_15497_new_n3354_; 
wire _abc_15497_new_n3355_; 
wire _abc_15497_new_n3356_; 
wire _abc_15497_new_n3357_; 
wire _abc_15497_new_n3358_; 
wire _abc_15497_new_n3359_; 
wire _abc_15497_new_n3360_; 
wire _abc_15497_new_n3361_; 
wire _abc_15497_new_n3362_; 
wire _abc_15497_new_n3363_; 
wire _abc_15497_new_n3364_; 
wire _abc_15497_new_n3365_; 
wire _abc_15497_new_n3366_; 
wire _abc_15497_new_n3367_; 
wire _abc_15497_new_n3368_; 
wire _abc_15497_new_n3369_; 
wire _abc_15497_new_n3370_; 
wire _abc_15497_new_n3371_; 
wire _abc_15497_new_n3372_; 
wire _abc_15497_new_n3373_; 
wire _abc_15497_new_n3374_; 
wire _abc_15497_new_n3375_; 
wire _abc_15497_new_n3376_; 
wire _abc_15497_new_n3377_; 
wire _abc_15497_new_n3378_; 
wire _abc_15497_new_n3379_; 
wire _abc_15497_new_n3380_; 
wire _abc_15497_new_n3381_; 
wire _abc_15497_new_n3382_; 
wire _abc_15497_new_n3383_; 
wire _abc_15497_new_n3384_; 
wire _abc_15497_new_n3385_; 
wire _abc_15497_new_n3386_; 
wire _abc_15497_new_n3387_; 
wire _abc_15497_new_n3388_; 
wire _abc_15497_new_n3389_; 
wire _abc_15497_new_n3390_; 
wire _abc_15497_new_n3391_; 
wire _abc_15497_new_n3392_; 
wire _abc_15497_new_n3393_; 
wire _abc_15497_new_n3394_; 
wire _abc_15497_new_n3395_; 
wire _abc_15497_new_n3396_; 
wire _abc_15497_new_n3397_; 
wire _abc_15497_new_n3398_; 
wire _abc_15497_new_n3399_; 
wire _abc_15497_new_n3400_; 
wire _abc_15497_new_n3401_; 
wire _abc_15497_new_n3403_; 
wire _abc_15497_new_n3404_; 
wire _abc_15497_new_n3405_; 
wire _abc_15497_new_n3406_; 
wire _abc_15497_new_n3407_; 
wire _abc_15497_new_n3408_; 
wire _abc_15497_new_n3409_; 
wire _abc_15497_new_n3410_; 
wire _abc_15497_new_n3411_; 
wire _abc_15497_new_n3412_; 
wire _abc_15497_new_n3413_; 
wire _abc_15497_new_n3414_; 
wire _abc_15497_new_n3415_; 
wire _abc_15497_new_n3416_; 
wire _abc_15497_new_n3417_; 
wire _abc_15497_new_n3418_; 
wire _abc_15497_new_n3419_; 
wire _abc_15497_new_n3420_; 
wire _abc_15497_new_n3421_; 
wire _abc_15497_new_n3422_; 
wire _abc_15497_new_n3423_; 
wire _abc_15497_new_n3424_; 
wire _abc_15497_new_n3425_; 
wire _abc_15497_new_n3426_; 
wire _abc_15497_new_n3427_; 
wire _abc_15497_new_n3428_; 
wire _abc_15497_new_n3429_; 
wire _abc_15497_new_n3430_; 
wire _abc_15497_new_n3431_; 
wire _abc_15497_new_n3432_; 
wire _abc_15497_new_n3433_; 
wire _abc_15497_new_n3434_; 
wire _abc_15497_new_n3435_; 
wire _abc_15497_new_n3436_; 
wire _abc_15497_new_n3437_; 
wire _abc_15497_new_n3438_; 
wire _abc_15497_new_n3439_; 
wire _abc_15497_new_n3440_; 
wire _abc_15497_new_n3441_; 
wire _abc_15497_new_n3442_; 
wire _abc_15497_new_n3443_; 
wire _abc_15497_new_n3444_; 
wire _abc_15497_new_n3445_; 
wire _abc_15497_new_n3446_; 
wire _abc_15497_new_n3447_; 
wire _abc_15497_new_n3448_; 
wire _abc_15497_new_n3449_; 
wire _abc_15497_new_n3450_; 
wire _abc_15497_new_n3451_; 
wire _abc_15497_new_n3452_; 
wire _abc_15497_new_n3453_; 
wire _abc_15497_new_n3454_; 
wire _abc_15497_new_n3455_; 
wire _abc_15497_new_n3456_; 
wire _abc_15497_new_n3457_; 
wire _abc_15497_new_n3458_; 
wire _abc_15497_new_n3459_; 
wire _abc_15497_new_n3460_; 
wire _abc_15497_new_n3461_; 
wire _abc_15497_new_n3462_; 
wire _abc_15497_new_n3463_; 
wire _abc_15497_new_n3464_; 
wire _abc_15497_new_n3465_; 
wire _abc_15497_new_n3466_; 
wire _abc_15497_new_n3467_; 
wire _abc_15497_new_n3468_; 
wire _abc_15497_new_n3469_; 
wire _abc_15497_new_n3470_; 
wire _abc_15497_new_n3471_; 
wire _abc_15497_new_n3472_; 
wire _abc_15497_new_n3473_; 
wire _abc_15497_new_n3474_; 
wire _abc_15497_new_n3475_; 
wire _abc_15497_new_n3476_; 
wire _abc_15497_new_n3478_; 
wire _abc_15497_new_n3479_; 
wire _abc_15497_new_n3480_; 
wire _abc_15497_new_n3481_; 
wire _abc_15497_new_n3482_; 
wire _abc_15497_new_n3483_; 
wire _abc_15497_new_n3484_; 
wire _abc_15497_new_n3485_; 
wire _abc_15497_new_n3486_; 
wire _abc_15497_new_n3487_; 
wire _abc_15497_new_n3488_; 
wire _abc_15497_new_n3489_; 
wire _abc_15497_new_n3490_; 
wire _abc_15497_new_n3491_; 
wire _abc_15497_new_n3492_; 
wire _abc_15497_new_n3493_; 
wire _abc_15497_new_n3494_; 
wire _abc_15497_new_n3495_; 
wire _abc_15497_new_n3496_; 
wire _abc_15497_new_n3497_; 
wire _abc_15497_new_n3498_; 
wire _abc_15497_new_n3499_; 
wire _abc_15497_new_n3500_; 
wire _abc_15497_new_n3501_; 
wire _abc_15497_new_n3502_; 
wire _abc_15497_new_n3503_; 
wire _abc_15497_new_n3504_; 
wire _abc_15497_new_n3505_; 
wire _abc_15497_new_n3506_; 
wire _abc_15497_new_n3507_; 
wire _abc_15497_new_n3508_; 
wire _abc_15497_new_n3509_; 
wire _abc_15497_new_n3510_; 
wire _abc_15497_new_n3511_; 
wire _abc_15497_new_n3512_; 
wire _abc_15497_new_n3513_; 
wire _abc_15497_new_n3514_; 
wire _abc_15497_new_n3515_; 
wire _abc_15497_new_n3516_; 
wire _abc_15497_new_n3517_; 
wire _abc_15497_new_n3518_; 
wire _abc_15497_new_n3519_; 
wire _abc_15497_new_n3520_; 
wire _abc_15497_new_n3521_; 
wire _abc_15497_new_n3522_; 
wire _abc_15497_new_n3523_; 
wire _abc_15497_new_n3524_; 
wire _abc_15497_new_n3525_; 
wire _abc_15497_new_n3526_; 
wire _abc_15497_new_n3527_; 
wire _abc_15497_new_n3528_; 
wire _abc_15497_new_n3529_; 
wire _abc_15497_new_n3530_; 
wire _abc_15497_new_n3531_; 
wire _abc_15497_new_n3532_; 
wire _abc_15497_new_n3533_; 
wire _abc_15497_new_n3535_; 
wire _abc_15497_new_n3536_; 
wire _abc_15497_new_n3537_; 
wire _abc_15497_new_n3538_; 
wire _abc_15497_new_n3539_; 
wire _abc_15497_new_n3540_; 
wire _abc_15497_new_n3541_; 
wire _abc_15497_new_n3542_; 
wire _abc_15497_new_n3543_; 
wire _abc_15497_new_n3544_; 
wire _abc_15497_new_n3545_; 
wire _abc_15497_new_n3546_; 
wire _abc_15497_new_n3547_; 
wire _abc_15497_new_n3548_; 
wire _abc_15497_new_n3549_; 
wire _abc_15497_new_n3550_; 
wire _abc_15497_new_n3551_; 
wire _abc_15497_new_n3552_; 
wire _abc_15497_new_n3553_; 
wire _abc_15497_new_n3554_; 
wire _abc_15497_new_n3555_; 
wire _abc_15497_new_n3556_; 
wire _abc_15497_new_n3557_; 
wire _abc_15497_new_n3558_; 
wire _abc_15497_new_n3559_; 
wire _abc_15497_new_n3560_; 
wire _abc_15497_new_n3561_; 
wire _abc_15497_new_n3562_; 
wire _abc_15497_new_n3563_; 
wire _abc_15497_new_n3564_; 
wire _abc_15497_new_n3565_; 
wire _abc_15497_new_n3566_; 
wire _abc_15497_new_n3567_; 
wire _abc_15497_new_n3568_; 
wire _abc_15497_new_n3569_; 
wire _abc_15497_new_n3570_; 
wire _abc_15497_new_n3571_; 
wire _abc_15497_new_n3572_; 
wire _abc_15497_new_n3573_; 
wire _abc_15497_new_n3574_; 
wire _abc_15497_new_n3575_; 
wire _abc_15497_new_n3576_; 
wire _abc_15497_new_n3577_; 
wire _abc_15497_new_n3578_; 
wire _abc_15497_new_n3579_; 
wire _abc_15497_new_n3580_; 
wire _abc_15497_new_n3581_; 
wire _abc_15497_new_n3582_; 
wire _abc_15497_new_n3583_; 
wire _abc_15497_new_n3584_; 
wire _abc_15497_new_n3585_; 
wire _abc_15497_new_n3586_; 
wire _abc_15497_new_n3587_; 
wire _abc_15497_new_n3588_; 
wire _abc_15497_new_n3589_; 
wire _abc_15497_new_n3590_; 
wire _abc_15497_new_n3591_; 
wire _abc_15497_new_n3592_; 
wire _abc_15497_new_n3593_; 
wire _abc_15497_new_n3594_; 
wire _abc_15497_new_n3595_; 
wire _abc_15497_new_n3596_; 
wire _abc_15497_new_n3597_; 
wire _abc_15497_new_n3598_; 
wire _abc_15497_new_n3599_; 
wire _abc_15497_new_n3600_; 
wire _abc_15497_new_n3601_; 
wire _abc_15497_new_n3603_; 
wire _abc_15497_new_n3604_; 
wire _abc_15497_new_n3605_; 
wire _abc_15497_new_n3606_; 
wire _abc_15497_new_n3607_; 
wire _abc_15497_new_n3608_; 
wire _abc_15497_new_n3609_; 
wire _abc_15497_new_n3610_; 
wire _abc_15497_new_n3611_; 
wire _abc_15497_new_n3612_; 
wire _abc_15497_new_n3613_; 
wire _abc_15497_new_n3614_; 
wire _abc_15497_new_n3615_; 
wire _abc_15497_new_n3616_; 
wire _abc_15497_new_n3617_; 
wire _abc_15497_new_n3618_; 
wire _abc_15497_new_n3619_; 
wire _abc_15497_new_n3620_; 
wire _abc_15497_new_n3621_; 
wire _abc_15497_new_n3622_; 
wire _abc_15497_new_n3623_; 
wire _abc_15497_new_n3624_; 
wire _abc_15497_new_n3625_; 
wire _abc_15497_new_n3626_; 
wire _abc_15497_new_n3627_; 
wire _abc_15497_new_n3628_; 
wire _abc_15497_new_n3629_; 
wire _abc_15497_new_n3630_; 
wire _abc_15497_new_n3631_; 
wire _abc_15497_new_n3632_; 
wire _abc_15497_new_n3633_; 
wire _abc_15497_new_n3634_; 
wire _abc_15497_new_n3635_; 
wire _abc_15497_new_n3636_; 
wire _abc_15497_new_n3637_; 
wire _abc_15497_new_n3638_; 
wire _abc_15497_new_n3639_; 
wire _abc_15497_new_n3640_; 
wire _abc_15497_new_n3641_; 
wire _abc_15497_new_n3642_; 
wire _abc_15497_new_n3643_; 
wire _abc_15497_new_n3644_; 
wire _abc_15497_new_n3645_; 
wire _abc_15497_new_n3646_; 
wire _abc_15497_new_n3647_; 
wire _abc_15497_new_n3648_; 
wire _abc_15497_new_n3649_; 
wire _abc_15497_new_n3650_; 
wire _abc_15497_new_n3651_; 
wire _abc_15497_new_n3652_; 
wire _abc_15497_new_n3653_; 
wire _abc_15497_new_n3654_; 
wire _abc_15497_new_n3655_; 
wire _abc_15497_new_n3656_; 
wire _abc_15497_new_n3657_; 
wire _abc_15497_new_n3658_; 
wire _abc_15497_new_n3659_; 
wire _abc_15497_new_n3660_; 
wire _abc_15497_new_n3661_; 
wire _abc_15497_new_n3662_; 
wire _abc_15497_new_n3663_; 
wire _abc_15497_new_n3664_; 
wire _abc_15497_new_n3665_; 
wire _abc_15497_new_n3666_; 
wire _abc_15497_new_n3668_; 
wire _abc_15497_new_n3669_; 
wire _abc_15497_new_n3670_; 
wire _abc_15497_new_n3671_; 
wire _abc_15497_new_n3672_; 
wire _abc_15497_new_n3673_; 
wire _abc_15497_new_n3674_; 
wire _abc_15497_new_n3675_; 
wire _abc_15497_new_n3676_; 
wire _abc_15497_new_n3677_; 
wire _abc_15497_new_n3678_; 
wire _abc_15497_new_n3679_; 
wire _abc_15497_new_n3680_; 
wire _abc_15497_new_n3681_; 
wire _abc_15497_new_n3682_; 
wire _abc_15497_new_n3683_; 
wire _abc_15497_new_n3684_; 
wire _abc_15497_new_n3685_; 
wire _abc_15497_new_n3686_; 
wire _abc_15497_new_n3687_; 
wire _abc_15497_new_n3688_; 
wire _abc_15497_new_n3689_; 
wire _abc_15497_new_n3690_; 
wire _abc_15497_new_n3691_; 
wire _abc_15497_new_n3692_; 
wire _abc_15497_new_n3693_; 
wire _abc_15497_new_n3694_; 
wire _abc_15497_new_n3695_; 
wire _abc_15497_new_n3696_; 
wire _abc_15497_new_n3697_; 
wire _abc_15497_new_n3698_; 
wire _abc_15497_new_n3699_; 
wire _abc_15497_new_n3700_; 
wire _abc_15497_new_n3701_; 
wire _abc_15497_new_n3702_; 
wire _abc_15497_new_n3703_; 
wire _abc_15497_new_n3704_; 
wire _abc_15497_new_n3705_; 
wire _abc_15497_new_n3706_; 
wire _abc_15497_new_n3707_; 
wire _abc_15497_new_n3708_; 
wire _abc_15497_new_n3709_; 
wire _abc_15497_new_n3710_; 
wire _abc_15497_new_n3711_; 
wire _abc_15497_new_n3712_; 
wire _abc_15497_new_n3713_; 
wire _abc_15497_new_n3714_; 
wire _abc_15497_new_n3715_; 
wire _abc_15497_new_n3716_; 
wire _abc_15497_new_n3717_; 
wire _abc_15497_new_n3718_; 
wire _abc_15497_new_n3719_; 
wire _abc_15497_new_n3721_; 
wire _abc_15497_new_n3722_; 
wire _abc_15497_new_n3723_; 
wire _abc_15497_new_n3724_; 
wire _abc_15497_new_n3725_; 
wire _abc_15497_new_n3726_; 
wire _abc_15497_new_n3727_; 
wire _abc_15497_new_n3728_; 
wire _abc_15497_new_n3729_; 
wire _abc_15497_new_n3730_; 
wire _abc_15497_new_n3731_; 
wire _abc_15497_new_n3732_; 
wire _abc_15497_new_n3733_; 
wire _abc_15497_new_n3734_; 
wire _abc_15497_new_n3735_; 
wire _abc_15497_new_n3736_; 
wire _abc_15497_new_n3737_; 
wire _abc_15497_new_n3738_; 
wire _abc_15497_new_n3739_; 
wire _abc_15497_new_n3740_; 
wire _abc_15497_new_n3741_; 
wire _abc_15497_new_n3742_; 
wire _abc_15497_new_n3743_; 
wire _abc_15497_new_n3744_; 
wire _abc_15497_new_n3745_; 
wire _abc_15497_new_n3746_; 
wire _abc_15497_new_n3747_; 
wire _abc_15497_new_n3748_; 
wire _abc_15497_new_n3749_; 
wire _abc_15497_new_n3750_; 
wire _abc_15497_new_n3751_; 
wire _abc_15497_new_n3752_; 
wire _abc_15497_new_n3753_; 
wire _abc_15497_new_n3754_; 
wire _abc_15497_new_n3755_; 
wire _abc_15497_new_n3756_; 
wire _abc_15497_new_n3757_; 
wire _abc_15497_new_n3758_; 
wire _abc_15497_new_n3759_; 
wire _abc_15497_new_n3760_; 
wire _abc_15497_new_n3761_; 
wire _abc_15497_new_n3762_; 
wire _abc_15497_new_n3763_; 
wire _abc_15497_new_n3764_; 
wire _abc_15497_new_n3765_; 
wire _abc_15497_new_n3766_; 
wire _abc_15497_new_n3767_; 
wire _abc_15497_new_n3768_; 
wire _abc_15497_new_n3769_; 
wire _abc_15497_new_n3770_; 
wire _abc_15497_new_n3771_; 
wire _abc_15497_new_n3772_; 
wire _abc_15497_new_n3773_; 
wire _abc_15497_new_n3774_; 
wire _abc_15497_new_n3776_; 
wire _abc_15497_new_n3777_; 
wire _abc_15497_new_n3778_; 
wire _abc_15497_new_n3779_; 
wire _abc_15497_new_n3780_; 
wire _abc_15497_new_n3781_; 
wire _abc_15497_new_n3782_; 
wire _abc_15497_new_n3783_; 
wire _abc_15497_new_n3784_; 
wire _abc_15497_new_n3785_; 
wire _abc_15497_new_n3786_; 
wire _abc_15497_new_n3787_; 
wire _abc_15497_new_n3788_; 
wire _abc_15497_new_n3789_; 
wire _abc_15497_new_n3790_; 
wire _abc_15497_new_n3791_; 
wire _abc_15497_new_n3792_; 
wire _abc_15497_new_n3793_; 
wire _abc_15497_new_n3794_; 
wire _abc_15497_new_n3795_; 
wire _abc_15497_new_n3796_; 
wire _abc_15497_new_n3797_; 
wire _abc_15497_new_n3798_; 
wire _abc_15497_new_n3799_; 
wire _abc_15497_new_n3800_; 
wire _abc_15497_new_n3801_; 
wire _abc_15497_new_n3802_; 
wire _abc_15497_new_n3803_; 
wire _abc_15497_new_n3804_; 
wire _abc_15497_new_n3805_; 
wire _abc_15497_new_n3806_; 
wire _abc_15497_new_n3807_; 
wire _abc_15497_new_n3808_; 
wire _abc_15497_new_n3809_; 
wire _abc_15497_new_n3810_; 
wire _abc_15497_new_n3811_; 
wire _abc_15497_new_n3812_; 
wire _abc_15497_new_n3813_; 
wire _abc_15497_new_n3814_; 
wire _abc_15497_new_n3815_; 
wire _abc_15497_new_n3816_; 
wire _abc_15497_new_n3817_; 
wire _abc_15497_new_n3818_; 
wire _abc_15497_new_n3819_; 
wire _abc_15497_new_n3820_; 
wire _abc_15497_new_n3821_; 
wire _abc_15497_new_n3822_; 
wire _abc_15497_new_n3824_; 
wire _abc_15497_new_n3825_; 
wire _abc_15497_new_n3826_; 
wire _abc_15497_new_n3827_; 
wire _abc_15497_new_n3828_; 
wire _abc_15497_new_n3829_; 
wire _abc_15497_new_n3830_; 
wire _abc_15497_new_n3831_; 
wire _abc_15497_new_n3832_; 
wire _abc_15497_new_n3833_; 
wire _abc_15497_new_n3834_; 
wire _abc_15497_new_n3835_; 
wire _abc_15497_new_n3836_; 
wire _abc_15497_new_n3837_; 
wire _abc_15497_new_n3838_; 
wire _abc_15497_new_n3839_; 
wire _abc_15497_new_n3840_; 
wire _abc_15497_new_n3841_; 
wire _abc_15497_new_n3842_; 
wire _abc_15497_new_n3843_; 
wire _abc_15497_new_n3844_; 
wire _abc_15497_new_n3845_; 
wire _abc_15497_new_n3846_; 
wire _abc_15497_new_n3847_; 
wire _abc_15497_new_n3848_; 
wire _abc_15497_new_n3849_; 
wire _abc_15497_new_n3850_; 
wire _abc_15497_new_n3851_; 
wire _abc_15497_new_n3852_; 
wire _abc_15497_new_n3853_; 
wire _abc_15497_new_n3854_; 
wire _abc_15497_new_n3855_; 
wire _abc_15497_new_n3856_; 
wire _abc_15497_new_n3857_; 
wire _abc_15497_new_n3858_; 
wire _abc_15497_new_n3859_; 
wire _abc_15497_new_n3860_; 
wire _abc_15497_new_n3861_; 
wire _abc_15497_new_n3862_; 
wire _abc_15497_new_n3863_; 
wire _abc_15497_new_n3864_; 
wire _abc_15497_new_n3865_; 
wire _abc_15497_new_n3866_; 
wire _abc_15497_new_n3867_; 
wire _abc_15497_new_n3868_; 
wire _abc_15497_new_n3870_; 
wire _abc_15497_new_n3871_; 
wire _abc_15497_new_n3872_; 
wire _abc_15497_new_n3873_; 
wire _abc_15497_new_n3874_; 
wire _abc_15497_new_n3875_; 
wire _abc_15497_new_n3876_; 
wire _abc_15497_new_n3877_; 
wire _abc_15497_new_n3878_; 
wire _abc_15497_new_n3879_; 
wire _abc_15497_new_n3880_; 
wire _abc_15497_new_n3881_; 
wire _abc_15497_new_n3882_; 
wire _abc_15497_new_n3883_; 
wire _abc_15497_new_n3884_; 
wire _abc_15497_new_n3885_; 
wire _abc_15497_new_n3886_; 
wire _abc_15497_new_n3887_; 
wire _abc_15497_new_n3888_; 
wire _abc_15497_new_n3889_; 
wire _abc_15497_new_n3890_; 
wire _abc_15497_new_n3891_; 
wire _abc_15497_new_n3892_; 
wire _abc_15497_new_n3893_; 
wire _abc_15497_new_n3894_; 
wire _abc_15497_new_n3895_; 
wire _abc_15497_new_n3896_; 
wire _abc_15497_new_n3897_; 
wire _abc_15497_new_n3898_; 
wire _abc_15497_new_n3899_; 
wire _abc_15497_new_n3900_; 
wire _abc_15497_new_n3901_; 
wire _abc_15497_new_n3902_; 
wire _abc_15497_new_n3903_; 
wire _abc_15497_new_n3904_; 
wire _abc_15497_new_n3905_; 
wire _abc_15497_new_n3906_; 
wire _abc_15497_new_n3907_; 
wire _abc_15497_new_n3908_; 
wire _abc_15497_new_n3909_; 
wire _abc_15497_new_n3910_; 
wire _abc_15497_new_n3911_; 
wire _abc_15497_new_n3912_; 
wire _abc_15497_new_n3913_; 
wire _abc_15497_new_n3914_; 
wire _abc_15497_new_n3915_; 
wire _abc_15497_new_n3916_; 
wire _abc_15497_new_n3917_; 
wire _abc_15497_new_n3918_; 
wire _abc_15497_new_n3919_; 
wire _abc_15497_new_n3920_; 
wire _abc_15497_new_n3921_; 
wire _abc_15497_new_n3922_; 
wire _abc_15497_new_n3923_; 
wire _abc_15497_new_n3924_; 
wire _abc_15497_new_n3925_; 
wire _abc_15497_new_n3926_; 
wire _abc_15497_new_n3927_; 
wire _abc_15497_new_n3928_; 
wire _abc_15497_new_n3929_; 
wire _abc_15497_new_n3930_; 
wire _abc_15497_new_n3931_; 
wire _abc_15497_new_n3932_; 
wire _abc_15497_new_n3933_; 
wire _abc_15497_new_n3935_; 
wire _abc_15497_new_n3936_; 
wire _abc_15497_new_n3937_; 
wire _abc_15497_new_n3938_; 
wire _abc_15497_new_n3939_; 
wire _abc_15497_new_n3940_; 
wire _abc_15497_new_n3941_; 
wire _abc_15497_new_n3942_; 
wire _abc_15497_new_n3943_; 
wire _abc_15497_new_n3944_; 
wire _abc_15497_new_n3945_; 
wire _abc_15497_new_n3946_; 
wire _abc_15497_new_n3947_; 
wire _abc_15497_new_n3948_; 
wire _abc_15497_new_n3949_; 
wire _abc_15497_new_n3950_; 
wire _abc_15497_new_n3951_; 
wire _abc_15497_new_n3952_; 
wire _abc_15497_new_n3953_; 
wire _abc_15497_new_n3954_; 
wire _abc_15497_new_n3955_; 
wire _abc_15497_new_n3956_; 
wire _abc_15497_new_n3957_; 
wire _abc_15497_new_n3958_; 
wire _abc_15497_new_n3959_; 
wire _abc_15497_new_n3960_; 
wire _abc_15497_new_n3961_; 
wire _abc_15497_new_n3962_; 
wire _abc_15497_new_n3963_; 
wire _abc_15497_new_n3964_; 
wire _abc_15497_new_n3965_; 
wire _abc_15497_new_n3966_; 
wire _abc_15497_new_n3967_; 
wire _abc_15497_new_n3968_; 
wire _abc_15497_new_n3969_; 
wire _abc_15497_new_n3970_; 
wire _abc_15497_new_n3971_; 
wire _abc_15497_new_n3972_; 
wire _abc_15497_new_n3973_; 
wire _abc_15497_new_n3974_; 
wire _abc_15497_new_n3975_; 
wire _abc_15497_new_n3976_; 
wire _abc_15497_new_n3977_; 
wire _abc_15497_new_n3978_; 
wire _abc_15497_new_n3979_; 
wire _abc_15497_new_n3980_; 
wire _abc_15497_new_n3981_; 
wire _abc_15497_new_n3982_; 
wire _abc_15497_new_n3983_; 
wire _abc_15497_new_n3984_; 
wire _abc_15497_new_n3986_; 
wire _abc_15497_new_n3987_; 
wire _abc_15497_new_n3988_; 
wire _abc_15497_new_n3989_; 
wire _abc_15497_new_n3990_; 
wire _abc_15497_new_n3991_; 
wire _abc_15497_new_n3992_; 
wire _abc_15497_new_n3993_; 
wire _abc_15497_new_n3994_; 
wire _abc_15497_new_n3995_; 
wire _abc_15497_new_n3996_; 
wire _abc_15497_new_n3997_; 
wire _abc_15497_new_n3998_; 
wire _abc_15497_new_n3999_; 
wire _abc_15497_new_n4000_; 
wire _abc_15497_new_n4001_; 
wire _abc_15497_new_n4002_; 
wire _abc_15497_new_n4003_; 
wire _abc_15497_new_n4004_; 
wire _abc_15497_new_n4005_; 
wire _abc_15497_new_n4006_; 
wire _abc_15497_new_n4007_; 
wire _abc_15497_new_n4008_; 
wire _abc_15497_new_n4009_; 
wire _abc_15497_new_n4010_; 
wire _abc_15497_new_n4011_; 
wire _abc_15497_new_n4012_; 
wire _abc_15497_new_n4013_; 
wire _abc_15497_new_n4014_; 
wire _abc_15497_new_n4015_; 
wire _abc_15497_new_n4016_; 
wire _abc_15497_new_n4017_; 
wire _abc_15497_new_n4018_; 
wire _abc_15497_new_n4019_; 
wire _abc_15497_new_n4020_; 
wire _abc_15497_new_n4021_; 
wire _abc_15497_new_n4022_; 
wire _abc_15497_new_n4023_; 
wire _abc_15497_new_n4024_; 
wire _abc_15497_new_n4025_; 
wire _abc_15497_new_n4026_; 
wire _abc_15497_new_n4027_; 
wire _abc_15497_new_n4028_; 
wire _abc_15497_new_n4029_; 
wire _abc_15497_new_n4030_; 
wire _abc_15497_new_n4031_; 
wire _abc_15497_new_n4032_; 
wire _abc_15497_new_n4033_; 
wire _abc_15497_new_n4034_; 
wire _abc_15497_new_n4035_; 
wire _abc_15497_new_n4036_; 
wire _abc_15497_new_n4037_; 
wire _abc_15497_new_n4038_; 
wire _abc_15497_new_n4039_; 
wire _abc_15497_new_n4041_; 
wire _abc_15497_new_n4042_; 
wire _abc_15497_new_n4043_; 
wire _abc_15497_new_n4044_; 
wire _abc_15497_new_n4045_; 
wire _abc_15497_new_n4046_; 
wire _abc_15497_new_n4047_; 
wire _abc_15497_new_n4048_; 
wire _abc_15497_new_n4049_; 
wire _abc_15497_new_n4050_; 
wire _abc_15497_new_n4051_; 
wire _abc_15497_new_n4052_; 
wire _abc_15497_new_n4053_; 
wire _abc_15497_new_n4054_; 
wire _abc_15497_new_n4055_; 
wire _abc_15497_new_n4056_; 
wire _abc_15497_new_n4057_; 
wire _abc_15497_new_n4058_; 
wire _abc_15497_new_n4059_; 
wire _abc_15497_new_n4060_; 
wire _abc_15497_new_n4061_; 
wire _abc_15497_new_n4062_; 
wire _abc_15497_new_n4063_; 
wire _abc_15497_new_n4064_; 
wire _abc_15497_new_n4065_; 
wire _abc_15497_new_n4066_; 
wire _abc_15497_new_n4067_; 
wire _abc_15497_new_n4068_; 
wire _abc_15497_new_n4069_; 
wire _abc_15497_new_n4070_; 
wire _abc_15497_new_n4071_; 
wire _abc_15497_new_n4072_; 
wire _abc_15497_new_n4073_; 
wire _abc_15497_new_n4074_; 
wire _abc_15497_new_n4075_; 
wire _abc_15497_new_n4076_; 
wire _abc_15497_new_n4077_; 
wire _abc_15497_new_n4078_; 
wire _abc_15497_new_n4079_; 
wire _abc_15497_new_n4080_; 
wire _abc_15497_new_n4081_; 
wire _abc_15497_new_n4082_; 
wire _abc_15497_new_n4083_; 
wire _abc_15497_new_n4084_; 
wire _abc_15497_new_n4085_; 
wire _abc_15497_new_n4086_; 
wire _abc_15497_new_n4087_; 
wire _abc_15497_new_n4088_; 
wire _abc_15497_new_n4089_; 
wire _abc_15497_new_n4090_; 
wire _abc_15497_new_n4091_; 
wire _abc_15497_new_n4092_; 
wire _abc_15497_new_n4093_; 
wire _abc_15497_new_n4094_; 
wire _abc_15497_new_n4095_; 
wire _abc_15497_new_n4097_; 
wire _abc_15497_new_n4098_; 
wire _abc_15497_new_n4099_; 
wire _abc_15497_new_n4100_; 
wire _abc_15497_new_n4101_; 
wire _abc_15497_new_n4102_; 
wire _abc_15497_new_n4103_; 
wire _abc_15497_new_n4104_; 
wire _abc_15497_new_n4105_; 
wire _abc_15497_new_n4106_; 
wire _abc_15497_new_n4107_; 
wire _abc_15497_new_n4108_; 
wire _abc_15497_new_n4109_; 
wire _abc_15497_new_n4110_; 
wire _abc_15497_new_n4111_; 
wire _abc_15497_new_n4112_; 
wire _abc_15497_new_n4113_; 
wire _abc_15497_new_n4114_; 
wire _abc_15497_new_n4115_; 
wire _abc_15497_new_n4116_; 
wire _abc_15497_new_n4117_; 
wire _abc_15497_new_n4118_; 
wire _abc_15497_new_n4119_; 
wire _abc_15497_new_n4120_; 
wire _abc_15497_new_n4121_; 
wire _abc_15497_new_n4122_; 
wire _abc_15497_new_n4123_; 
wire _abc_15497_new_n4124_; 
wire _abc_15497_new_n4125_; 
wire _abc_15497_new_n4126_; 
wire _abc_15497_new_n4127_; 
wire _abc_15497_new_n4128_; 
wire _abc_15497_new_n4129_; 
wire _abc_15497_new_n4130_; 
wire _abc_15497_new_n4131_; 
wire _abc_15497_new_n4132_; 
wire _abc_15497_new_n4133_; 
wire _abc_15497_new_n4134_; 
wire _abc_15497_new_n4135_; 
wire _abc_15497_new_n4136_; 
wire _abc_15497_new_n4137_; 
wire _abc_15497_new_n4138_; 
wire _abc_15497_new_n4139_; 
wire _abc_15497_new_n4140_; 
wire _abc_15497_new_n4141_; 
wire _abc_15497_new_n4142_; 
wire _abc_15497_new_n4143_; 
wire _abc_15497_new_n4144_; 
wire _abc_15497_new_n4145_; 
wire _abc_15497_new_n4146_; 
wire _abc_15497_new_n4147_; 
wire _abc_15497_new_n4149_; 
wire _abc_15497_new_n4150_; 
wire _abc_15497_new_n4151_; 
wire _abc_15497_new_n4152_; 
wire _abc_15497_new_n4153_; 
wire _abc_15497_new_n4154_; 
wire _abc_15497_new_n4155_; 
wire _abc_15497_new_n4156_; 
wire _abc_15497_new_n4157_; 
wire _abc_15497_new_n4158_; 
wire _abc_15497_new_n4159_; 
wire _abc_15497_new_n4160_; 
wire _abc_15497_new_n4161_; 
wire _abc_15497_new_n4162_; 
wire _abc_15497_new_n4163_; 
wire _abc_15497_new_n4164_; 
wire _abc_15497_new_n4165_; 
wire _abc_15497_new_n4166_; 
wire _abc_15497_new_n4167_; 
wire _abc_15497_new_n4168_; 
wire _abc_15497_new_n4169_; 
wire _abc_15497_new_n4170_; 
wire _abc_15497_new_n4171_; 
wire _abc_15497_new_n4172_; 
wire _abc_15497_new_n4173_; 
wire _abc_15497_new_n4174_; 
wire _abc_15497_new_n4175_; 
wire _abc_15497_new_n4176_; 
wire _abc_15497_new_n4177_; 
wire _abc_15497_new_n4178_; 
wire _abc_15497_new_n4179_; 
wire _abc_15497_new_n4180_; 
wire _abc_15497_new_n4181_; 
wire _abc_15497_new_n4182_; 
wire _abc_15497_new_n4183_; 
wire _abc_15497_new_n4184_; 
wire _abc_15497_new_n4185_; 
wire _abc_15497_new_n4187_; 
wire _abc_15497_new_n4188_; 
wire _abc_15497_new_n4189_; 
wire _abc_15497_new_n4190_; 
wire _abc_15497_new_n4191_; 
wire _abc_15497_new_n4192_; 
wire _abc_15497_new_n4193_; 
wire _abc_15497_new_n4194_; 
wire _abc_15497_new_n4195_; 
wire _abc_15497_new_n4196_; 
wire _abc_15497_new_n4197_; 
wire _abc_15497_new_n4198_; 
wire _abc_15497_new_n4199_; 
wire _abc_15497_new_n4200_; 
wire _abc_15497_new_n4201_; 
wire _abc_15497_new_n4202_; 
wire _abc_15497_new_n4203_; 
wire _abc_15497_new_n4204_; 
wire _abc_15497_new_n4205_; 
wire _abc_15497_new_n4206_; 
wire _abc_15497_new_n4207_; 
wire _abc_15497_new_n4208_; 
wire _abc_15497_new_n4209_; 
wire _abc_15497_new_n4210_; 
wire _abc_15497_new_n4211_; 
wire _abc_15497_new_n4212_; 
wire _abc_15497_new_n4213_; 
wire _abc_15497_new_n4214_; 
wire _abc_15497_new_n4215_; 
wire _abc_15497_new_n4216_; 
wire _abc_15497_new_n4217_; 
wire _abc_15497_new_n4218_; 
wire _abc_15497_new_n4219_; 
wire _abc_15497_new_n4220_; 
wire _abc_15497_new_n4221_; 
wire _abc_15497_new_n4222_; 
wire _abc_15497_new_n4223_; 
wire _abc_15497_new_n4224_; 
wire _abc_15497_new_n4225_; 
wire _abc_15497_new_n4226_; 
wire _abc_15497_new_n4227_; 
wire _abc_15497_new_n4228_; 
wire _abc_15497_new_n4229_; 
wire _abc_15497_new_n4231_; 
wire _abc_15497_new_n4232_; 
wire _abc_15497_new_n4233_; 
wire _abc_15497_new_n4234_; 
wire _abc_15497_new_n4235_; 
wire _abc_15497_new_n4236_; 
wire _abc_15497_new_n4237_; 
wire _abc_15497_new_n4238_; 
wire _abc_15497_new_n4239_; 
wire _abc_15497_new_n4240_; 
wire _abc_15497_new_n4241_; 
wire _abc_15497_new_n4242_; 
wire _abc_15497_new_n4243_; 
wire _abc_15497_new_n4244_; 
wire _abc_15497_new_n4245_; 
wire _abc_15497_new_n4246_; 
wire _abc_15497_new_n4247_; 
wire _abc_15497_new_n4248_; 
wire _abc_15497_new_n4249_; 
wire _abc_15497_new_n4250_; 
wire _abc_15497_new_n4251_; 
wire _abc_15497_new_n4252_; 
wire _abc_15497_new_n4253_; 
wire _abc_15497_new_n4254_; 
wire _abc_15497_new_n4255_; 
wire _abc_15497_new_n4256_; 
wire _abc_15497_new_n4257_; 
wire _abc_15497_new_n4258_; 
wire _abc_15497_new_n4259_; 
wire _abc_15497_new_n4260_; 
wire _abc_15497_new_n4261_; 
wire _abc_15497_new_n4262_; 
wire _abc_15497_new_n4263_; 
wire _abc_15497_new_n4264_; 
wire _abc_15497_new_n4265_; 
wire _abc_15497_new_n4266_; 
wire _abc_15497_new_n4267_; 
wire _abc_15497_new_n4269_; 
wire _abc_15497_new_n4270_; 
wire _abc_15497_new_n4271_; 
wire _abc_15497_new_n4272_; 
wire _abc_15497_new_n4273_; 
wire _abc_15497_new_n4274_; 
wire _abc_15497_new_n4275_; 
wire _abc_15497_new_n4276_; 
wire _abc_15497_new_n4277_; 
wire _abc_15497_new_n4278_; 
wire _abc_15497_new_n4279_; 
wire _abc_15497_new_n4280_; 
wire _abc_15497_new_n4281_; 
wire _abc_15497_new_n4282_; 
wire _abc_15497_new_n4283_; 
wire _abc_15497_new_n4284_; 
wire _abc_15497_new_n4285_; 
wire _abc_15497_new_n4286_; 
wire _abc_15497_new_n4287_; 
wire _abc_15497_new_n4288_; 
wire _abc_15497_new_n4289_; 
wire _abc_15497_new_n4290_; 
wire _abc_15497_new_n4291_; 
wire _abc_15497_new_n4292_; 
wire _abc_15497_new_n4293_; 
wire _abc_15497_new_n4294_; 
wire _abc_15497_new_n4295_; 
wire _abc_15497_new_n4296_; 
wire _abc_15497_new_n4297_; 
wire _abc_15497_new_n4298_; 
wire _abc_15497_new_n4299_; 
wire _abc_15497_new_n4300_; 
wire _abc_15497_new_n4301_; 
wire _abc_15497_new_n4302_; 
wire _abc_15497_new_n4303_; 
wire _abc_15497_new_n4304_; 
wire _abc_15497_new_n4305_; 
wire _abc_15497_new_n4306_; 
wire _abc_15497_new_n4307_; 
wire _abc_15497_new_n4308_; 
wire _abc_15497_new_n4309_; 
wire _abc_15497_new_n4310_; 
wire _abc_15497_new_n4311_; 
wire _abc_15497_new_n4312_; 
wire _abc_15497_new_n4313_; 
wire _abc_15497_new_n4314_; 
wire _abc_15497_new_n4315_; 
wire _abc_15497_new_n4316_; 
wire _abc_15497_new_n4317_; 
wire _abc_15497_new_n4318_; 
wire _abc_15497_new_n4319_; 
wire _abc_15497_new_n4320_; 
wire _abc_15497_new_n4321_; 
wire _abc_15497_new_n4322_; 
wire _abc_15497_new_n4324_; 
wire _abc_15497_new_n4325_; 
wire _abc_15497_new_n4326_; 
wire _abc_15497_new_n4327_; 
wire _abc_15497_new_n4328_; 
wire _abc_15497_new_n4329_; 
wire _abc_15497_new_n4330_; 
wire _abc_15497_new_n4331_; 
wire _abc_15497_new_n4332_; 
wire _abc_15497_new_n4333_; 
wire _abc_15497_new_n4334_; 
wire _abc_15497_new_n4335_; 
wire _abc_15497_new_n4336_; 
wire _abc_15497_new_n4337_; 
wire _abc_15497_new_n4338_; 
wire _abc_15497_new_n4339_; 
wire _abc_15497_new_n4340_; 
wire _abc_15497_new_n4341_; 
wire _abc_15497_new_n4342_; 
wire _abc_15497_new_n4343_; 
wire _abc_15497_new_n4344_; 
wire _abc_15497_new_n4345_; 
wire _abc_15497_new_n4346_; 
wire _abc_15497_new_n4347_; 
wire _abc_15497_new_n4348_; 
wire _abc_15497_new_n4349_; 
wire _abc_15497_new_n4350_; 
wire _abc_15497_new_n4351_; 
wire _abc_15497_new_n4352_; 
wire _abc_15497_new_n4353_; 
wire _abc_15497_new_n4354_; 
wire _abc_15497_new_n4355_; 
wire _abc_15497_new_n4356_; 
wire _abc_15497_new_n4357_; 
wire _abc_15497_new_n4358_; 
wire _abc_15497_new_n4359_; 
wire _abc_15497_new_n4360_; 
wire _abc_15497_new_n4361_; 
wire _abc_15497_new_n4362_; 
wire _abc_15497_new_n4363_; 
wire _abc_15497_new_n4365_; 
wire _abc_15497_new_n4366_; 
wire _abc_15497_new_n4367_; 
wire _abc_15497_new_n4368_; 
wire _abc_15497_new_n4369_; 
wire _abc_15497_new_n4370_; 
wire _abc_15497_new_n4371_; 
wire _abc_15497_new_n4372_; 
wire _abc_15497_new_n4373_; 
wire _abc_15497_new_n4374_; 
wire _abc_15497_new_n4375_; 
wire _abc_15497_new_n4376_; 
wire _abc_15497_new_n4377_; 
wire _abc_15497_new_n4378_; 
wire _abc_15497_new_n4379_; 
wire _abc_15497_new_n4380_; 
wire _abc_15497_new_n4381_; 
wire _abc_15497_new_n4382_; 
wire _abc_15497_new_n4383_; 
wire _abc_15497_new_n4384_; 
wire _abc_15497_new_n4385_; 
wire _abc_15497_new_n4386_; 
wire _abc_15497_new_n4387_; 
wire _abc_15497_new_n4388_; 
wire _abc_15497_new_n4389_; 
wire _abc_15497_new_n4390_; 
wire _abc_15497_new_n4391_; 
wire _abc_15497_new_n4392_; 
wire _abc_15497_new_n4393_; 
wire _abc_15497_new_n4394_; 
wire _abc_15497_new_n4395_; 
wire _abc_15497_new_n4396_; 
wire _abc_15497_new_n4397_; 
wire _abc_15497_new_n4398_; 
wire _abc_15497_new_n4399_; 
wire _abc_15497_new_n4400_; 
wire _abc_15497_new_n4401_; 
wire _abc_15497_new_n4402_; 
wire _abc_15497_new_n4403_; 
wire _abc_15497_new_n4404_; 
wire _abc_15497_new_n4406_; 
wire _abc_15497_new_n4407_; 
wire _abc_15497_new_n4408_; 
wire _abc_15497_new_n4409_; 
wire _abc_15497_new_n4410_; 
wire _abc_15497_new_n4411_; 
wire _abc_15497_new_n4412_; 
wire _abc_15497_new_n4413_; 
wire _abc_15497_new_n4414_; 
wire _abc_15497_new_n4415_; 
wire _abc_15497_new_n4416_; 
wire _abc_15497_new_n4417_; 
wire _abc_15497_new_n4418_; 
wire _abc_15497_new_n4419_; 
wire _abc_15497_new_n4420_; 
wire _abc_15497_new_n4421_; 
wire _abc_15497_new_n4422_; 
wire _abc_15497_new_n4423_; 
wire _abc_15497_new_n4424_; 
wire _abc_15497_new_n4425_; 
wire _abc_15497_new_n4426_; 
wire _abc_15497_new_n4427_; 
wire _abc_15497_new_n4428_; 
wire _abc_15497_new_n4429_; 
wire _abc_15497_new_n4430_; 
wire _abc_15497_new_n4431_; 
wire _abc_15497_new_n4432_; 
wire _abc_15497_new_n4433_; 
wire _abc_15497_new_n4434_; 
wire _abc_15497_new_n4435_; 
wire _abc_15497_new_n4436_; 
wire _abc_15497_new_n4437_; 
wire _abc_15497_new_n4438_; 
wire _abc_15497_new_n4439_; 
wire _abc_15497_new_n4441_; 
wire _abc_15497_new_n4442_; 
wire _abc_15497_new_n4443_; 
wire _abc_15497_new_n4444_; 
wire _abc_15497_new_n4445_; 
wire _abc_15497_new_n4446_; 
wire _abc_15497_new_n4447_; 
wire _abc_15497_new_n4449_; 
wire _abc_15497_new_n4451_; 
wire _abc_15497_new_n4453_; 
wire _abc_15497_new_n4455_; 
wire _abc_15497_new_n4456_; 
wire _abc_15497_new_n4458_; 
wire _abc_15497_new_n4459_; 
wire _abc_15497_new_n4460_; 
wire _abc_15497_new_n4462_; 
wire _abc_15497_new_n4463_; 
wire _abc_15497_new_n4464_; 
wire _abc_15497_new_n4466_; 
wire _abc_15497_new_n4468_; 
wire _abc_15497_new_n4469_; 
wire _abc_15497_new_n4470_; 
wire _abc_15497_new_n4472_; 
wire _abc_15497_new_n4474_; 
wire _abc_15497_new_n4476_; 
wire _abc_15497_new_n4477_; 
wire _abc_15497_new_n4479_; 
wire _abc_15497_new_n4480_; 
wire _abc_15497_new_n4482_; 
wire _abc_15497_new_n4483_; 
wire _abc_15497_new_n4485_; 
wire _abc_15497_new_n4486_; 
wire _abc_15497_new_n4487_; 
wire _abc_15497_new_n4488_; 
wire _abc_15497_new_n4490_; 
wire _abc_15497_new_n4491_; 
wire _abc_15497_new_n4493_; 
wire _abc_15497_new_n4494_; 
wire _abc_15497_new_n4495_; 
wire _abc_15497_new_n4496_; 
wire _abc_15497_new_n4497_; 
wire _abc_15497_new_n4499_; 
wire _abc_15497_new_n4500_; 
wire _abc_15497_new_n4501_; 
wire _abc_15497_new_n4502_; 
wire _abc_15497_new_n4503_; 
wire _abc_15497_new_n4504_; 
wire _abc_15497_new_n4505_; 
wire _abc_15497_new_n4507_; 
wire _abc_15497_new_n4508_; 
wire _abc_15497_new_n4509_; 
wire _abc_15497_new_n4511_; 
wire _abc_15497_new_n4512_; 
wire _abc_15497_new_n4513_; 
wire _abc_15497_new_n4515_; 
wire _abc_15497_new_n4516_; 
wire _abc_15497_new_n4517_; 
wire _abc_15497_new_n4519_; 
wire _abc_15497_new_n4520_; 
wire _abc_15497_new_n4521_; 
wire _abc_15497_new_n4522_; 
wire _abc_15497_new_n4523_; 
wire _abc_15497_new_n4524_; 
wire _abc_15497_new_n4526_; 
wire _abc_15497_new_n4527_; 
wire _abc_15497_new_n4528_; 
wire _abc_15497_new_n4530_; 
wire _abc_15497_new_n4531_; 
wire _abc_15497_new_n4532_; 
wire _abc_15497_new_n4533_; 
wire _abc_15497_new_n4535_; 
wire _abc_15497_new_n4536_; 
wire _abc_15497_new_n4537_; 
wire _abc_15497_new_n4539_; 
wire _abc_15497_new_n4540_; 
wire _abc_15497_new_n4541_; 
wire _abc_15497_new_n4542_; 
wire _abc_15497_new_n4543_; 
wire _abc_15497_new_n4545_; 
wire _abc_15497_new_n4546_; 
wire _abc_15497_new_n4547_; 
wire _abc_15497_new_n4549_; 
wire _abc_15497_new_n4550_; 
wire _abc_15497_new_n4551_; 
wire _abc_15497_new_n4553_; 
wire _abc_15497_new_n4554_; 
wire _abc_15497_new_n4555_; 
wire _abc_15497_new_n4557_; 
wire _abc_15497_new_n4558_; 
wire _abc_15497_new_n4560_; 
wire _abc_15497_new_n4561_; 
wire _abc_15497_new_n4562_; 
wire _abc_15497_new_n4564_; 
wire _abc_15497_new_n4565_; 
wire _abc_15497_new_n4566_; 
wire _abc_15497_new_n4567_; 
wire _abc_15497_new_n4568_; 
wire _abc_15497_new_n4569_; 
wire _abc_15497_new_n4571_; 
wire _abc_15497_new_n4572_; 
wire _abc_15497_new_n4573_; 
wire _abc_15497_new_n4574_; 
wire _abc_15497_new_n4575_; 
wire _abc_15497_new_n4577_; 
wire _abc_15497_new_n4578_; 
wire _abc_15497_new_n4579_; 
wire _abc_15497_new_n4580_; 
wire _abc_15497_new_n4582_; 
wire _abc_15497_new_n4583_; 
wire _abc_15497_new_n4584_; 
wire _abc_15497_new_n4585_; 
wire _abc_15497_new_n4586_; 
wire _abc_15497_new_n4588_; 
wire _abc_15497_new_n4589_; 
wire _abc_15497_new_n4591_; 
wire _abc_15497_new_n4592_; 
wire _abc_15497_new_n4593_; 
wire _abc_15497_new_n4594_; 
wire _abc_15497_new_n698_; 
wire _abc_15497_new_n699_; 
wire _abc_15497_new_n700_; 
wire _abc_15497_new_n701_; 
wire _abc_15497_new_n702_; 
wire _abc_15497_new_n703_; 
wire _abc_15497_new_n704_; 
wire _abc_15497_new_n705_; 
wire _abc_15497_new_n706_; 
wire _abc_15497_new_n707_; 
wire _abc_15497_new_n708_; 
wire _abc_15497_new_n709_; 
wire _abc_15497_new_n710_; 
wire _abc_15497_new_n711_; 
wire _abc_15497_new_n712_; 
wire _abc_15497_new_n713_; 
wire _abc_15497_new_n714_; 
wire _abc_15497_new_n715_; 
wire _abc_15497_new_n716_; 
wire _abc_15497_new_n717_; 
wire _abc_15497_new_n718_; 
wire _abc_15497_new_n719_; 
wire _abc_15497_new_n720_; 
wire _abc_15497_new_n721_; 
wire _abc_15497_new_n722_; 
wire _abc_15497_new_n723_; 
wire _abc_15497_new_n724_; 
wire _abc_15497_new_n725_; 
wire _abc_15497_new_n726_; 
wire _abc_15497_new_n727_; 
wire _abc_15497_new_n728_; 
wire _abc_15497_new_n729_; 
wire _abc_15497_new_n730_; 
wire _abc_15497_new_n731_; 
wire _abc_15497_new_n732_; 
wire _abc_15497_new_n733_; 
wire _abc_15497_new_n734_; 
wire _abc_15497_new_n735_; 
wire _abc_15497_new_n736_; 
wire _abc_15497_new_n737_; 
wire _abc_15497_new_n738_; 
wire _abc_15497_new_n739_; 
wire _abc_15497_new_n740_; 
wire _abc_15497_new_n741_; 
wire _abc_15497_new_n742_; 
wire _abc_15497_new_n743_; 
wire _abc_15497_new_n744_; 
wire _abc_15497_new_n745_; 
wire _abc_15497_new_n746_; 
wire _abc_15497_new_n747_; 
wire _abc_15497_new_n748_; 
wire _abc_15497_new_n749_; 
wire _abc_15497_new_n750_; 
wire _abc_15497_new_n751_; 
wire _abc_15497_new_n752_; 
wire _abc_15497_new_n753_; 
wire _abc_15497_new_n754_; 
wire _abc_15497_new_n755_; 
wire _abc_15497_new_n756_; 
wire _abc_15497_new_n757_; 
wire _abc_15497_new_n758_; 
wire _abc_15497_new_n759_; 
wire _abc_15497_new_n760_; 
wire _abc_15497_new_n761_; 
wire _abc_15497_new_n762_; 
wire _abc_15497_new_n763_; 
wire _abc_15497_new_n764_; 
wire _abc_15497_new_n765_; 
wire _abc_15497_new_n766_; 
wire _abc_15497_new_n767_; 
wire _abc_15497_new_n768_; 
wire _abc_15497_new_n769_; 
wire _abc_15497_new_n770_; 
wire _abc_15497_new_n771_; 
wire _abc_15497_new_n772_; 
wire _abc_15497_new_n773_; 
wire _abc_15497_new_n774_; 
wire _abc_15497_new_n775_; 
wire _abc_15497_new_n776_; 
wire _abc_15497_new_n777_; 
wire _abc_15497_new_n778_; 
wire _abc_15497_new_n779_; 
wire _abc_15497_new_n780_; 
wire _abc_15497_new_n781_; 
wire _abc_15497_new_n782_; 
wire _abc_15497_new_n783_; 
wire _abc_15497_new_n784_; 
wire _abc_15497_new_n785_; 
wire _abc_15497_new_n786_; 
wire _abc_15497_new_n787_; 
wire _abc_15497_new_n788_; 
wire _abc_15497_new_n789_; 
wire _abc_15497_new_n790_; 
wire _abc_15497_new_n791_; 
wire _abc_15497_new_n792_; 
wire _abc_15497_new_n793_; 
wire _abc_15497_new_n794_; 
wire _abc_15497_new_n795_; 
wire _abc_15497_new_n796_; 
wire _abc_15497_new_n797_; 
wire _abc_15497_new_n798_; 
wire _abc_15497_new_n799_; 
wire _abc_15497_new_n800_; 
wire _abc_15497_new_n801_; 
wire _abc_15497_new_n802_; 
wire _abc_15497_new_n803_; 
wire _abc_15497_new_n804_; 
wire _abc_15497_new_n805_; 
wire _abc_15497_new_n806_; 
wire _abc_15497_new_n807_; 
wire _abc_15497_new_n808_; 
wire _abc_15497_new_n809_; 
wire _abc_15497_new_n810_; 
wire _abc_15497_new_n811_; 
wire _abc_15497_new_n812_; 
wire _abc_15497_new_n813_; 
wire _abc_15497_new_n814_; 
wire _abc_15497_new_n815_; 
wire _abc_15497_new_n816_; 
wire _abc_15497_new_n817_; 
wire _abc_15497_new_n818_; 
wire _abc_15497_new_n819_; 
wire _abc_15497_new_n820_; 
wire _abc_15497_new_n821_; 
wire _abc_15497_new_n822_; 
wire _abc_15497_new_n823_; 
wire _abc_15497_new_n824_; 
wire _abc_15497_new_n825_; 
wire _abc_15497_new_n826_; 
wire _abc_15497_new_n827_; 
wire _abc_15497_new_n828_; 
wire _abc_15497_new_n829_; 
wire _abc_15497_new_n830_; 
wire _abc_15497_new_n831_; 
wire _abc_15497_new_n832_; 
wire _abc_15497_new_n833_; 
wire _abc_15497_new_n834_; 
wire _abc_15497_new_n835_; 
wire _abc_15497_new_n836_; 
wire _abc_15497_new_n837_; 
wire _abc_15497_new_n838_; 
wire _abc_15497_new_n839_; 
wire _abc_15497_new_n840_; 
wire _abc_15497_new_n841_; 
wire _abc_15497_new_n842_; 
wire _abc_15497_new_n843_; 
wire _abc_15497_new_n844_; 
wire _abc_15497_new_n845_; 
wire _abc_15497_new_n846_; 
wire _abc_15497_new_n847_; 
wire _abc_15497_new_n848_; 
wire _abc_15497_new_n849_; 
wire _abc_15497_new_n850_; 
wire _abc_15497_new_n851_; 
wire _abc_15497_new_n852_; 
wire _abc_15497_new_n853_; 
wire _abc_15497_new_n854_; 
wire _abc_15497_new_n855_; 
wire _abc_15497_new_n856_; 
wire _abc_15497_new_n857_; 
wire _abc_15497_new_n858_; 
wire _abc_15497_new_n859_; 
wire _abc_15497_new_n860_; 
wire _abc_15497_new_n861_; 
wire _abc_15497_new_n862_; 
wire _abc_15497_new_n863_; 
wire _abc_15497_new_n864_; 
wire _abc_15497_new_n865_; 
wire _abc_15497_new_n866_; 
wire _abc_15497_new_n867_; 
wire _abc_15497_new_n868_; 
wire _abc_15497_new_n869_; 
wire _abc_15497_new_n870_; 
wire _abc_15497_new_n870__bF_buf0; 
wire _abc_15497_new_n870__bF_buf1; 
wire _abc_15497_new_n870__bF_buf10; 
wire _abc_15497_new_n870__bF_buf11; 
wire _abc_15497_new_n870__bF_buf2; 
wire _abc_15497_new_n870__bF_buf3; 
wire _abc_15497_new_n870__bF_buf4; 
wire _abc_15497_new_n870__bF_buf5; 
wire _abc_15497_new_n870__bF_buf6; 
wire _abc_15497_new_n870__bF_buf7; 
wire _abc_15497_new_n870__bF_buf8; 
wire _abc_15497_new_n870__bF_buf9; 
wire _abc_15497_new_n871_; 
wire _abc_15497_new_n871__bF_buf0; 
wire _abc_15497_new_n871__bF_buf1; 
wire _abc_15497_new_n871__bF_buf2; 
wire _abc_15497_new_n871__bF_buf3; 
wire _abc_15497_new_n871__bF_buf4; 
wire _abc_15497_new_n872_; 
wire _abc_15497_new_n872__bF_buf0; 
wire _abc_15497_new_n872__bF_buf1; 
wire _abc_15497_new_n872__bF_buf2; 
wire _abc_15497_new_n872__bF_buf3; 
wire _abc_15497_new_n872__bF_buf4; 
wire _abc_15497_new_n873_; 
wire _abc_15497_new_n873__bF_buf0; 
wire _abc_15497_new_n873__bF_buf1; 
wire _abc_15497_new_n873__bF_buf2; 
wire _abc_15497_new_n873__bF_buf3; 
wire _abc_15497_new_n873__bF_buf4; 
wire _abc_15497_new_n873__bF_buf5; 
wire _abc_15497_new_n873__bF_buf6; 
wire _abc_15497_new_n873__bF_buf7; 
wire _abc_15497_new_n874_; 
wire _abc_15497_new_n875_; 
wire _abc_15497_new_n877_; 
wire _abc_15497_new_n878_; 
wire _abc_15497_new_n879_; 
wire _abc_15497_new_n880_; 
wire _abc_15497_new_n881_; 
wire _abc_15497_new_n882_; 
wire _abc_15497_new_n883_; 
wire _abc_15497_new_n883__bF_buf0; 
wire _abc_15497_new_n883__bF_buf1; 
wire _abc_15497_new_n883__bF_buf10; 
wire _abc_15497_new_n883__bF_buf11; 
wire _abc_15497_new_n883__bF_buf12; 
wire _abc_15497_new_n883__bF_buf13; 
wire _abc_15497_new_n883__bF_buf2; 
wire _abc_15497_new_n883__bF_buf3; 
wire _abc_15497_new_n883__bF_buf4; 
wire _abc_15497_new_n883__bF_buf5; 
wire _abc_15497_new_n883__bF_buf6; 
wire _abc_15497_new_n883__bF_buf7; 
wire _abc_15497_new_n883__bF_buf8; 
wire _abc_15497_new_n883__bF_buf9; 
wire _abc_15497_new_n884_; 
wire _abc_15497_new_n886_; 
wire _abc_15497_new_n887_; 
wire _abc_15497_new_n888_; 
wire _abc_15497_new_n889_; 
wire _abc_15497_new_n890_; 
wire _abc_15497_new_n891_; 
wire _abc_15497_new_n892_; 
wire _abc_15497_new_n893_; 
wire _abc_15497_new_n894_; 
wire _abc_15497_new_n895_; 
wire _abc_15497_new_n896_; 
wire _abc_15497_new_n897_; 
wire _abc_15497_new_n898_; 
wire _abc_15497_new_n899_; 
wire _abc_15497_new_n901_; 
wire _abc_15497_new_n902_; 
wire _abc_15497_new_n903_; 
wire _abc_15497_new_n904_; 
wire _abc_15497_new_n905_; 
wire _abc_15497_new_n906_; 
wire _abc_15497_new_n907_; 
wire _abc_15497_new_n908_; 
wire _abc_15497_new_n909_; 
wire _abc_15497_new_n911_; 
wire _abc_15497_new_n912_; 
wire _abc_15497_new_n913_; 
wire _abc_15497_new_n914_; 
wire _abc_15497_new_n915_; 
wire _abc_15497_new_n916_; 
wire _abc_15497_new_n917_; 
wire _abc_15497_new_n918_; 
wire _abc_15497_new_n919_; 
wire _abc_15497_new_n920_; 
wire _abc_15497_new_n921_; 
wire _abc_15497_new_n922_; 
wire _abc_15497_new_n923_; 
wire _abc_15497_new_n925_; 
wire _abc_15497_new_n926_; 
wire _abc_15497_new_n927_; 
wire _abc_15497_new_n928_; 
wire _abc_15497_new_n929_; 
wire _abc_15497_new_n930_; 
wire _abc_15497_new_n931_; 
wire _abc_15497_new_n932_; 
wire _abc_15497_new_n933_; 
wire _abc_15497_new_n934_; 
wire _abc_15497_new_n936_; 
wire _abc_15497_new_n937_; 
wire _abc_15497_new_n938_; 
wire _abc_15497_new_n939_; 
wire _abc_15497_new_n941_; 
wire _abc_15497_new_n942_; 
wire _abc_15497_new_n943_; 
wire _abc_15497_new_n944_; 
wire _abc_15497_new_n946_; 
wire _abc_15497_new_n947_; 
wire _abc_15497_new_n948_; 
wire _abc_15497_new_n949_; 
wire _abc_15497_new_n950_; 
wire _abc_15497_new_n951_; 
wire _abc_15497_new_n952_; 
wire _abc_15497_new_n953_; 
wire _abc_15497_new_n955_; 
wire _abc_15497_new_n956_; 
wire _abc_15497_new_n957_; 
wire _abc_15497_new_n958_; 
wire _abc_15497_new_n959_; 
wire _abc_15497_new_n960_; 
wire _abc_15497_new_n961_; 
wire _abc_15497_new_n962_; 
wire _abc_15497_new_n963_; 
wire _abc_15497_new_n964_; 
wire _abc_15497_new_n966_; 
wire _abc_15497_new_n967_; 
wire _abc_15497_new_n968_; 
wire _abc_15497_new_n969_; 
wire _abc_15497_new_n970_; 
wire _abc_15497_new_n971_; 
wire _abc_15497_new_n972_; 
wire _abc_15497_new_n973_; 
wire _abc_15497_new_n974_; 
wire _abc_15497_new_n976_; 
wire _abc_15497_new_n977_; 
wire _abc_15497_new_n978_; 
wire _abc_15497_new_n979_; 
wire _abc_15497_new_n980_; 
wire _abc_15497_new_n981_; 
wire _abc_15497_new_n982_; 
wire _abc_15497_new_n984_; 
wire _abc_15497_new_n985_; 
wire _abc_15497_new_n986_; 
wire _abc_15497_new_n987_; 
wire _abc_15497_new_n988_; 
wire _abc_15497_new_n989_; 
wire _abc_15497_new_n991_; 
wire _abc_15497_new_n992_; 
wire _abc_15497_new_n993_; 
wire _abc_15497_new_n994_; 
wire _abc_15497_new_n995_; 
wire _abc_15497_new_n996_; 
wire _abc_15497_new_n997_; 
wire _abc_15497_new_n998_; 
wire _abc_15497_new_n999_; 
wire _auto_iopadmap_cc_368_execute_22625_0_; 
wire _auto_iopadmap_cc_368_execute_22625_100_; 
wire _auto_iopadmap_cc_368_execute_22625_101_; 
wire _auto_iopadmap_cc_368_execute_22625_102_; 
wire _auto_iopadmap_cc_368_execute_22625_103_; 
wire _auto_iopadmap_cc_368_execute_22625_104_; 
wire _auto_iopadmap_cc_368_execute_22625_105_; 
wire _auto_iopadmap_cc_368_execute_22625_106_; 
wire _auto_iopadmap_cc_368_execute_22625_107_; 
wire _auto_iopadmap_cc_368_execute_22625_108_; 
wire _auto_iopadmap_cc_368_execute_22625_109_; 
wire _auto_iopadmap_cc_368_execute_22625_10_; 
wire _auto_iopadmap_cc_368_execute_22625_110_; 
wire _auto_iopadmap_cc_368_execute_22625_111_; 
wire _auto_iopadmap_cc_368_execute_22625_112_; 
wire _auto_iopadmap_cc_368_execute_22625_113_; 
wire _auto_iopadmap_cc_368_execute_22625_114_; 
wire _auto_iopadmap_cc_368_execute_22625_115_; 
wire _auto_iopadmap_cc_368_execute_22625_116_; 
wire _auto_iopadmap_cc_368_execute_22625_117_; 
wire _auto_iopadmap_cc_368_execute_22625_118_; 
wire _auto_iopadmap_cc_368_execute_22625_119_; 
wire _auto_iopadmap_cc_368_execute_22625_11_; 
wire _auto_iopadmap_cc_368_execute_22625_120_; 
wire _auto_iopadmap_cc_368_execute_22625_121_; 
wire _auto_iopadmap_cc_368_execute_22625_122_; 
wire _auto_iopadmap_cc_368_execute_22625_123_; 
wire _auto_iopadmap_cc_368_execute_22625_124_; 
wire _auto_iopadmap_cc_368_execute_22625_125_; 
wire _auto_iopadmap_cc_368_execute_22625_126_; 
wire _auto_iopadmap_cc_368_execute_22625_127_; 
wire _auto_iopadmap_cc_368_execute_22625_128_; 
wire _auto_iopadmap_cc_368_execute_22625_129_; 
wire _auto_iopadmap_cc_368_execute_22625_12_; 
wire _auto_iopadmap_cc_368_execute_22625_130_; 
wire _auto_iopadmap_cc_368_execute_22625_131_; 
wire _auto_iopadmap_cc_368_execute_22625_132_; 
wire _auto_iopadmap_cc_368_execute_22625_133_; 
wire _auto_iopadmap_cc_368_execute_22625_134_; 
wire _auto_iopadmap_cc_368_execute_22625_135_; 
wire _auto_iopadmap_cc_368_execute_22625_136_; 
wire _auto_iopadmap_cc_368_execute_22625_137_; 
wire _auto_iopadmap_cc_368_execute_22625_138_; 
wire _auto_iopadmap_cc_368_execute_22625_139_; 
wire _auto_iopadmap_cc_368_execute_22625_13_; 
wire _auto_iopadmap_cc_368_execute_22625_140_; 
wire _auto_iopadmap_cc_368_execute_22625_141_; 
wire _auto_iopadmap_cc_368_execute_22625_142_; 
wire _auto_iopadmap_cc_368_execute_22625_143_; 
wire _auto_iopadmap_cc_368_execute_22625_144_; 
wire _auto_iopadmap_cc_368_execute_22625_145_; 
wire _auto_iopadmap_cc_368_execute_22625_146_; 
wire _auto_iopadmap_cc_368_execute_22625_147_; 
wire _auto_iopadmap_cc_368_execute_22625_148_; 
wire _auto_iopadmap_cc_368_execute_22625_149_; 
wire _auto_iopadmap_cc_368_execute_22625_14_; 
wire _auto_iopadmap_cc_368_execute_22625_150_; 
wire _auto_iopadmap_cc_368_execute_22625_151_; 
wire _auto_iopadmap_cc_368_execute_22625_152_; 
wire _auto_iopadmap_cc_368_execute_22625_153_; 
wire _auto_iopadmap_cc_368_execute_22625_154_; 
wire _auto_iopadmap_cc_368_execute_22625_155_; 
wire _auto_iopadmap_cc_368_execute_22625_156_; 
wire _auto_iopadmap_cc_368_execute_22625_157_; 
wire _auto_iopadmap_cc_368_execute_22625_158_; 
wire _auto_iopadmap_cc_368_execute_22625_159_; 
wire _auto_iopadmap_cc_368_execute_22625_15_; 
wire _auto_iopadmap_cc_368_execute_22625_16_; 
wire _auto_iopadmap_cc_368_execute_22625_17_; 
wire _auto_iopadmap_cc_368_execute_22625_18_; 
wire _auto_iopadmap_cc_368_execute_22625_19_; 
wire _auto_iopadmap_cc_368_execute_22625_1_; 
wire _auto_iopadmap_cc_368_execute_22625_20_; 
wire _auto_iopadmap_cc_368_execute_22625_21_; 
wire _auto_iopadmap_cc_368_execute_22625_22_; 
wire _auto_iopadmap_cc_368_execute_22625_23_; 
wire _auto_iopadmap_cc_368_execute_22625_24_; 
wire _auto_iopadmap_cc_368_execute_22625_25_; 
wire _auto_iopadmap_cc_368_execute_22625_26_; 
wire _auto_iopadmap_cc_368_execute_22625_27_; 
wire _auto_iopadmap_cc_368_execute_22625_28_; 
wire _auto_iopadmap_cc_368_execute_22625_29_; 
wire _auto_iopadmap_cc_368_execute_22625_2_; 
wire _auto_iopadmap_cc_368_execute_22625_30_; 
wire _auto_iopadmap_cc_368_execute_22625_31_; 
wire _auto_iopadmap_cc_368_execute_22625_32_; 
wire _auto_iopadmap_cc_368_execute_22625_33_; 
wire _auto_iopadmap_cc_368_execute_22625_34_; 
wire _auto_iopadmap_cc_368_execute_22625_35_; 
wire _auto_iopadmap_cc_368_execute_22625_36_; 
wire _auto_iopadmap_cc_368_execute_22625_37_; 
wire _auto_iopadmap_cc_368_execute_22625_38_; 
wire _auto_iopadmap_cc_368_execute_22625_39_; 
wire _auto_iopadmap_cc_368_execute_22625_3_; 
wire _auto_iopadmap_cc_368_execute_22625_40_; 
wire _auto_iopadmap_cc_368_execute_22625_41_; 
wire _auto_iopadmap_cc_368_execute_22625_42_; 
wire _auto_iopadmap_cc_368_execute_22625_43_; 
wire _auto_iopadmap_cc_368_execute_22625_44_; 
wire _auto_iopadmap_cc_368_execute_22625_45_; 
wire _auto_iopadmap_cc_368_execute_22625_46_; 
wire _auto_iopadmap_cc_368_execute_22625_47_; 
wire _auto_iopadmap_cc_368_execute_22625_48_; 
wire _auto_iopadmap_cc_368_execute_22625_49_; 
wire _auto_iopadmap_cc_368_execute_22625_4_; 
wire _auto_iopadmap_cc_368_execute_22625_50_; 
wire _auto_iopadmap_cc_368_execute_22625_51_; 
wire _auto_iopadmap_cc_368_execute_22625_52_; 
wire _auto_iopadmap_cc_368_execute_22625_53_; 
wire _auto_iopadmap_cc_368_execute_22625_54_; 
wire _auto_iopadmap_cc_368_execute_22625_55_; 
wire _auto_iopadmap_cc_368_execute_22625_56_; 
wire _auto_iopadmap_cc_368_execute_22625_57_; 
wire _auto_iopadmap_cc_368_execute_22625_58_; 
wire _auto_iopadmap_cc_368_execute_22625_59_; 
wire _auto_iopadmap_cc_368_execute_22625_5_; 
wire _auto_iopadmap_cc_368_execute_22625_60_; 
wire _auto_iopadmap_cc_368_execute_22625_61_; 
wire _auto_iopadmap_cc_368_execute_22625_62_; 
wire _auto_iopadmap_cc_368_execute_22625_63_; 
wire _auto_iopadmap_cc_368_execute_22625_64_; 
wire _auto_iopadmap_cc_368_execute_22625_65_; 
wire _auto_iopadmap_cc_368_execute_22625_66_; 
wire _auto_iopadmap_cc_368_execute_22625_67_; 
wire _auto_iopadmap_cc_368_execute_22625_68_; 
wire _auto_iopadmap_cc_368_execute_22625_69_; 
wire _auto_iopadmap_cc_368_execute_22625_6_; 
wire _auto_iopadmap_cc_368_execute_22625_70_; 
wire _auto_iopadmap_cc_368_execute_22625_71_; 
wire _auto_iopadmap_cc_368_execute_22625_72_; 
wire _auto_iopadmap_cc_368_execute_22625_73_; 
wire _auto_iopadmap_cc_368_execute_22625_74_; 
wire _auto_iopadmap_cc_368_execute_22625_75_; 
wire _auto_iopadmap_cc_368_execute_22625_76_; 
wire _auto_iopadmap_cc_368_execute_22625_77_; 
wire _auto_iopadmap_cc_368_execute_22625_78_; 
wire _auto_iopadmap_cc_368_execute_22625_79_; 
wire _auto_iopadmap_cc_368_execute_22625_7_; 
wire _auto_iopadmap_cc_368_execute_22625_80_; 
wire _auto_iopadmap_cc_368_execute_22625_81_; 
wire _auto_iopadmap_cc_368_execute_22625_82_; 
wire _auto_iopadmap_cc_368_execute_22625_83_; 
wire _auto_iopadmap_cc_368_execute_22625_84_; 
wire _auto_iopadmap_cc_368_execute_22625_85_; 
wire _auto_iopadmap_cc_368_execute_22625_86_; 
wire _auto_iopadmap_cc_368_execute_22625_87_; 
wire _auto_iopadmap_cc_368_execute_22625_88_; 
wire _auto_iopadmap_cc_368_execute_22625_89_; 
wire _auto_iopadmap_cc_368_execute_22625_8_; 
wire _auto_iopadmap_cc_368_execute_22625_90_; 
wire _auto_iopadmap_cc_368_execute_22625_91_; 
wire _auto_iopadmap_cc_368_execute_22625_92_; 
wire _auto_iopadmap_cc_368_execute_22625_93_; 
wire _auto_iopadmap_cc_368_execute_22625_94_; 
wire _auto_iopadmap_cc_368_execute_22625_95_; 
wire _auto_iopadmap_cc_368_execute_22625_96_; 
wire _auto_iopadmap_cc_368_execute_22625_97_; 
wire _auto_iopadmap_cc_368_execute_22625_98_; 
wire _auto_iopadmap_cc_368_execute_22625_99_; 
wire _auto_iopadmap_cc_368_execute_22625_9_; 
wire _auto_iopadmap_cc_368_execute_22786; 
wire _auto_iopadmap_cc_368_execute_22788; 
wire a_reg_0_; 
wire a_reg_10_; 
wire a_reg_11_; 
wire a_reg_12_; 
wire a_reg_13_; 
wire a_reg_14_; 
wire a_reg_15_; 
wire a_reg_16_; 
wire a_reg_17_; 
wire a_reg_18_; 
wire a_reg_19_; 
wire a_reg_1_; 
wire a_reg_20_; 
wire a_reg_21_; 
wire a_reg_22_; 
wire a_reg_23_; 
wire a_reg_24_; 
wire a_reg_25_; 
wire a_reg_26_; 
wire a_reg_27_; 
wire a_reg_28_; 
wire a_reg_29_; 
wire a_reg_2_; 
wire a_reg_30_; 
wire a_reg_31_; 
wire a_reg_3_; 
wire a_reg_4_; 
wire a_reg_5_; 
wire a_reg_6_; 
wire a_reg_7_; 
wire a_reg_8_; 
wire a_reg_9_; 
wire b_reg_0_; 
wire b_reg_10_; 
wire b_reg_11_; 
wire b_reg_12_; 
wire b_reg_13_; 
wire b_reg_14_; 
wire b_reg_15_; 
wire b_reg_16_; 
wire b_reg_17_; 
wire b_reg_18_; 
wire b_reg_19_; 
wire b_reg_1_; 
wire b_reg_20_; 
wire b_reg_21_; 
wire b_reg_22_; 
wire b_reg_23_; 
wire b_reg_24_; 
wire b_reg_25_; 
wire b_reg_26_; 
wire b_reg_27_; 
wire b_reg_28_; 
wire b_reg_29_; 
wire b_reg_2_; 
wire b_reg_30_; 
wire b_reg_31_; 
wire b_reg_3_; 
wire b_reg_4_; 
wire b_reg_5_; 
wire b_reg_6_; 
wire b_reg_7_; 
wire b_reg_8_; 
wire b_reg_9_; 
input \block[0] ;
input \block[100] ;
input \block[101] ;
input \block[102] ;
input \block[103] ;
input \block[104] ;
input \block[105] ;
input \block[106] ;
input \block[107] ;
input \block[108] ;
input \block[109] ;
input \block[10] ;
input \block[110] ;
input \block[111] ;
input \block[112] ;
input \block[113] ;
input \block[114] ;
input \block[115] ;
input \block[116] ;
input \block[117] ;
input \block[118] ;
input \block[119] ;
input \block[11] ;
input \block[120] ;
input \block[121] ;
input \block[122] ;
input \block[123] ;
input \block[124] ;
input \block[125] ;
input \block[126] ;
input \block[127] ;
input \block[128] ;
input \block[129] ;
input \block[12] ;
input \block[130] ;
input \block[131] ;
input \block[132] ;
input \block[133] ;
input \block[134] ;
input \block[135] ;
input \block[136] ;
input \block[137] ;
input \block[138] ;
input \block[139] ;
input \block[13] ;
input \block[140] ;
input \block[141] ;
input \block[142] ;
input \block[143] ;
input \block[144] ;
input \block[145] ;
input \block[146] ;
input \block[147] ;
input \block[148] ;
input \block[149] ;
input \block[14] ;
input \block[150] ;
input \block[151] ;
input \block[152] ;
input \block[153] ;
input \block[154] ;
input \block[155] ;
input \block[156] ;
input \block[157] ;
input \block[158] ;
input \block[159] ;
input \block[15] ;
input \block[160] ;
input \block[161] ;
input \block[162] ;
input \block[163] ;
input \block[164] ;
input \block[165] ;
input \block[166] ;
input \block[167] ;
input \block[168] ;
input \block[169] ;
input \block[16] ;
input \block[170] ;
input \block[171] ;
input \block[172] ;
input \block[173] ;
input \block[174] ;
input \block[175] ;
input \block[176] ;
input \block[177] ;
input \block[178] ;
input \block[179] ;
input \block[17] ;
input \block[180] ;
input \block[181] ;
input \block[182] ;
input \block[183] ;
input \block[184] ;
input \block[185] ;
input \block[186] ;
input \block[187] ;
input \block[188] ;
input \block[189] ;
input \block[18] ;
input \block[190] ;
input \block[191] ;
input \block[192] ;
input \block[193] ;
input \block[194] ;
input \block[195] ;
input \block[196] ;
input \block[197] ;
input \block[198] ;
input \block[199] ;
input \block[19] ;
input \block[1] ;
input \block[200] ;
input \block[201] ;
input \block[202] ;
input \block[203] ;
input \block[204] ;
input \block[205] ;
input \block[206] ;
input \block[207] ;
input \block[208] ;
input \block[209] ;
input \block[20] ;
input \block[210] ;
input \block[211] ;
input \block[212] ;
input \block[213] ;
input \block[214] ;
input \block[215] ;
input \block[216] ;
input \block[217] ;
input \block[218] ;
input \block[219] ;
input \block[21] ;
input \block[220] ;
input \block[221] ;
input \block[222] ;
input \block[223] ;
input \block[224] ;
input \block[225] ;
input \block[226] ;
input \block[227] ;
input \block[228] ;
input \block[229] ;
input \block[22] ;
input \block[230] ;
input \block[231] ;
input \block[232] ;
input \block[233] ;
input \block[234] ;
input \block[235] ;
input \block[236] ;
input \block[237] ;
input \block[238] ;
input \block[239] ;
input \block[23] ;
input \block[240] ;
input \block[241] ;
input \block[242] ;
input \block[243] ;
input \block[244] ;
input \block[245] ;
input \block[246] ;
input \block[247] ;
input \block[248] ;
input \block[249] ;
input \block[24] ;
input \block[250] ;
input \block[251] ;
input \block[252] ;
input \block[253] ;
input \block[254] ;
input \block[255] ;
input \block[256] ;
input \block[257] ;
input \block[258] ;
input \block[259] ;
input \block[25] ;
input \block[260] ;
input \block[261] ;
input \block[262] ;
input \block[263] ;
input \block[264] ;
input \block[265] ;
input \block[266] ;
input \block[267] ;
input \block[268] ;
input \block[269] ;
input \block[26] ;
input \block[270] ;
input \block[271] ;
input \block[272] ;
input \block[273] ;
input \block[274] ;
input \block[275] ;
input \block[276] ;
input \block[277] ;
input \block[278] ;
input \block[279] ;
input \block[27] ;
input \block[280] ;
input \block[281] ;
input \block[282] ;
input \block[283] ;
input \block[284] ;
input \block[285] ;
input \block[286] ;
input \block[287] ;
input \block[288] ;
input \block[289] ;
input \block[28] ;
input \block[290] ;
input \block[291] ;
input \block[292] ;
input \block[293] ;
input \block[294] ;
input \block[295] ;
input \block[296] ;
input \block[297] ;
input \block[298] ;
input \block[299] ;
input \block[29] ;
input \block[2] ;
input \block[300] ;
input \block[301] ;
input \block[302] ;
input \block[303] ;
input \block[304] ;
input \block[305] ;
input \block[306] ;
input \block[307] ;
input \block[308] ;
input \block[309] ;
input \block[30] ;
input \block[310] ;
input \block[311] ;
input \block[312] ;
input \block[313] ;
input \block[314] ;
input \block[315] ;
input \block[316] ;
input \block[317] ;
input \block[318] ;
input \block[319] ;
input \block[31] ;
input \block[320] ;
input \block[321] ;
input \block[322] ;
input \block[323] ;
input \block[324] ;
input \block[325] ;
input \block[326] ;
input \block[327] ;
input \block[328] ;
input \block[329] ;
input \block[32] ;
input \block[330] ;
input \block[331] ;
input \block[332] ;
input \block[333] ;
input \block[334] ;
input \block[335] ;
input \block[336] ;
input \block[337] ;
input \block[338] ;
input \block[339] ;
input \block[33] ;
input \block[340] ;
input \block[341] ;
input \block[342] ;
input \block[343] ;
input \block[344] ;
input \block[345] ;
input \block[346] ;
input \block[347] ;
input \block[348] ;
input \block[349] ;
input \block[34] ;
input \block[350] ;
input \block[351] ;
input \block[352] ;
input \block[353] ;
input \block[354] ;
input \block[355] ;
input \block[356] ;
input \block[357] ;
input \block[358] ;
input \block[359] ;
input \block[35] ;
input \block[360] ;
input \block[361] ;
input \block[362] ;
input \block[363] ;
input \block[364] ;
input \block[365] ;
input \block[366] ;
input \block[367] ;
input \block[368] ;
input \block[369] ;
input \block[36] ;
input \block[370] ;
input \block[371] ;
input \block[372] ;
input \block[373] ;
input \block[374] ;
input \block[375] ;
input \block[376] ;
input \block[377] ;
input \block[378] ;
input \block[379] ;
input \block[37] ;
input \block[380] ;
input \block[381] ;
input \block[382] ;
input \block[383] ;
input \block[384] ;
input \block[385] ;
input \block[386] ;
input \block[387] ;
input \block[388] ;
input \block[389] ;
input \block[38] ;
input \block[390] ;
input \block[391] ;
input \block[392] ;
input \block[393] ;
input \block[394] ;
input \block[395] ;
input \block[396] ;
input \block[397] ;
input \block[398] ;
input \block[399] ;
input \block[39] ;
input \block[3] ;
input \block[400] ;
input \block[401] ;
input \block[402] ;
input \block[403] ;
input \block[404] ;
input \block[405] ;
input \block[406] ;
input \block[407] ;
input \block[408] ;
input \block[409] ;
input \block[40] ;
input \block[410] ;
input \block[411] ;
input \block[412] ;
input \block[413] ;
input \block[414] ;
input \block[415] ;
input \block[416] ;
input \block[417] ;
input \block[418] ;
input \block[419] ;
input \block[41] ;
input \block[420] ;
input \block[421] ;
input \block[422] ;
input \block[423] ;
input \block[424] ;
input \block[425] ;
input \block[426] ;
input \block[427] ;
input \block[428] ;
input \block[429] ;
input \block[42] ;
input \block[430] ;
input \block[431] ;
input \block[432] ;
input \block[433] ;
input \block[434] ;
input \block[435] ;
input \block[436] ;
input \block[437] ;
input \block[438] ;
input \block[439] ;
input \block[43] ;
input \block[440] ;
input \block[441] ;
input \block[442] ;
input \block[443] ;
input \block[444] ;
input \block[445] ;
input \block[446] ;
input \block[447] ;
input \block[448] ;
input \block[449] ;
input \block[44] ;
input \block[450] ;
input \block[451] ;
input \block[452] ;
input \block[453] ;
input \block[454] ;
input \block[455] ;
input \block[456] ;
input \block[457] ;
input \block[458] ;
input \block[459] ;
input \block[45] ;
input \block[460] ;
input \block[461] ;
input \block[462] ;
input \block[463] ;
input \block[464] ;
input \block[465] ;
input \block[466] ;
input \block[467] ;
input \block[468] ;
input \block[469] ;
input \block[46] ;
input \block[470] ;
input \block[471] ;
input \block[472] ;
input \block[473] ;
input \block[474] ;
input \block[475] ;
input \block[476] ;
input \block[477] ;
input \block[478] ;
input \block[479] ;
input \block[47] ;
input \block[480] ;
input \block[481] ;
input \block[482] ;
input \block[483] ;
input \block[484] ;
input \block[485] ;
input \block[486] ;
input \block[487] ;
input \block[488] ;
input \block[489] ;
input \block[48] ;
input \block[490] ;
input \block[491] ;
input \block[492] ;
input \block[493] ;
input \block[494] ;
input \block[495] ;
input \block[496] ;
input \block[497] ;
input \block[498] ;
input \block[499] ;
input \block[49] ;
input \block[4] ;
input \block[500] ;
input \block[501] ;
input \block[502] ;
input \block[503] ;
input \block[504] ;
input \block[505] ;
input \block[506] ;
input \block[507] ;
input \block[508] ;
input \block[509] ;
input \block[50] ;
input \block[510] ;
input \block[511] ;
input \block[51] ;
input \block[52] ;
input \block[53] ;
input \block[54] ;
input \block[55] ;
input \block[56] ;
input \block[57] ;
input \block[58] ;
input \block[59] ;
input \block[5] ;
input \block[60] ;
input \block[61] ;
input \block[62] ;
input \block[63] ;
input \block[64] ;
input \block[65] ;
input \block[66] ;
input \block[67] ;
input \block[68] ;
input \block[69] ;
input \block[6] ;
input \block[70] ;
input \block[71] ;
input \block[72] ;
input \block[73] ;
input \block[74] ;
input \block[75] ;
input \block[76] ;
input \block[77] ;
input \block[78] ;
input \block[79] ;
input \block[7] ;
input \block[80] ;
input \block[81] ;
input \block[82] ;
input \block[83] ;
input \block[84] ;
input \block[85] ;
input \block[86] ;
input \block[87] ;
input \block[88] ;
input \block[89] ;
input \block[8] ;
input \block[90] ;
input \block[91] ;
input \block[92] ;
input \block[93] ;
input \block[94] ;
input \block[95] ;
input \block[96] ;
input \block[97] ;
input \block[98] ;
input \block[99] ;
input \block[9] ;
wire c_reg_0_; 
wire c_reg_10_; 
wire c_reg_11_; 
wire c_reg_12_; 
wire c_reg_13_; 
wire c_reg_14_; 
wire c_reg_15_; 
wire c_reg_16_; 
wire c_reg_17_; 
wire c_reg_18_; 
wire c_reg_19_; 
wire c_reg_1_; 
wire c_reg_20_; 
wire c_reg_21_; 
wire c_reg_22_; 
wire c_reg_23_; 
wire c_reg_24_; 
wire c_reg_25_; 
wire c_reg_26_; 
wire c_reg_27_; 
wire c_reg_28_; 
wire c_reg_29_; 
wire c_reg_2_; 
wire c_reg_30_; 
wire c_reg_31_; 
wire c_reg_3_; 
wire c_reg_4_; 
wire c_reg_5_; 
wire c_reg_6_; 
wire c_reg_7_; 
wire c_reg_8_; 
wire c_reg_9_; 
input clk;
wire clk_bF_buf0; 
wire clk_bF_buf1; 
wire clk_bF_buf10; 
wire clk_bF_buf11; 
wire clk_bF_buf12; 
wire clk_bF_buf13; 
wire clk_bF_buf14; 
wire clk_bF_buf15; 
wire clk_bF_buf16; 
wire clk_bF_buf17; 
wire clk_bF_buf18; 
wire clk_bF_buf19; 
wire clk_bF_buf2; 
wire clk_bF_buf20; 
wire clk_bF_buf21; 
wire clk_bF_buf22; 
wire clk_bF_buf23; 
wire clk_bF_buf24; 
wire clk_bF_buf25; 
wire clk_bF_buf26; 
wire clk_bF_buf27; 
wire clk_bF_buf28; 
wire clk_bF_buf29; 
wire clk_bF_buf3; 
wire clk_bF_buf30; 
wire clk_bF_buf31; 
wire clk_bF_buf32; 
wire clk_bF_buf33; 
wire clk_bF_buf34; 
wire clk_bF_buf35; 
wire clk_bF_buf36; 
wire clk_bF_buf37; 
wire clk_bF_buf38; 
wire clk_bF_buf39; 
wire clk_bF_buf4; 
wire clk_bF_buf40; 
wire clk_bF_buf41; 
wire clk_bF_buf42; 
wire clk_bF_buf43; 
wire clk_bF_buf44; 
wire clk_bF_buf45; 
wire clk_bF_buf46; 
wire clk_bF_buf47; 
wire clk_bF_buf48; 
wire clk_bF_buf49; 
wire clk_bF_buf5; 
wire clk_bF_buf50; 
wire clk_bF_buf51; 
wire clk_bF_buf52; 
wire clk_bF_buf53; 
wire clk_bF_buf54; 
wire clk_bF_buf55; 
wire clk_bF_buf56; 
wire clk_bF_buf57; 
wire clk_bF_buf58; 
wire clk_bF_buf59; 
wire clk_bF_buf6; 
wire clk_bF_buf60; 
wire clk_bF_buf61; 
wire clk_bF_buf62; 
wire clk_bF_buf63; 
wire clk_bF_buf64; 
wire clk_bF_buf65; 
wire clk_bF_buf66; 
wire clk_bF_buf67; 
wire clk_bF_buf68; 
wire clk_bF_buf69; 
wire clk_bF_buf7; 
wire clk_bF_buf70; 
wire clk_bF_buf71; 
wire clk_bF_buf72; 
wire clk_bF_buf73; 
wire clk_bF_buf74; 
wire clk_bF_buf75; 
wire clk_bF_buf76; 
wire clk_bF_buf77; 
wire clk_bF_buf78; 
wire clk_bF_buf79; 
wire clk_bF_buf8; 
wire clk_bF_buf80; 
wire clk_bF_buf81; 
wire clk_bF_buf82; 
wire clk_bF_buf83; 
wire clk_bF_buf84; 
wire clk_bF_buf85; 
wire clk_bF_buf86; 
wire clk_bF_buf87; 
wire clk_bF_buf88; 
wire clk_bF_buf9; 
wire clk_hier0_bF_buf0; 
wire clk_hier0_bF_buf1; 
wire clk_hier0_bF_buf2; 
wire clk_hier0_bF_buf3; 
wire clk_hier0_bF_buf4; 
wire clk_hier0_bF_buf5; 
wire clk_hier0_bF_buf6; 
wire clk_hier0_bF_buf7; 
wire clk_hier0_bF_buf8; 
wire d_reg_0_; 
wire d_reg_10_; 
wire d_reg_11_; 
wire d_reg_12_; 
wire d_reg_13_; 
wire d_reg_14_; 
wire d_reg_15_; 
wire d_reg_16_; 
wire d_reg_17_; 
wire d_reg_18_; 
wire d_reg_19_; 
wire d_reg_1_; 
wire d_reg_20_; 
wire d_reg_21_; 
wire d_reg_22_; 
wire d_reg_23_; 
wire d_reg_24_; 
wire d_reg_25_; 
wire d_reg_26_; 
wire d_reg_27_; 
wire d_reg_28_; 
wire d_reg_29_; 
wire d_reg_2_; 
wire d_reg_30_; 
wire d_reg_31_; 
wire d_reg_3_; 
wire d_reg_4_; 
wire d_reg_5_; 
wire d_reg_6_; 
wire d_reg_7_; 
wire d_reg_8_; 
wire d_reg_9_; 
output \digest[0] ;
output \digest[100] ;
output \digest[101] ;
output \digest[102] ;
output \digest[103] ;
output \digest[104] ;
output \digest[105] ;
output \digest[106] ;
output \digest[107] ;
output \digest[108] ;
output \digest[109] ;
output \digest[10] ;
output \digest[110] ;
output \digest[111] ;
output \digest[112] ;
output \digest[113] ;
output \digest[114] ;
output \digest[115] ;
output \digest[116] ;
output \digest[117] ;
output \digest[118] ;
output \digest[119] ;
output \digest[11] ;
output \digest[120] ;
output \digest[121] ;
output \digest[122] ;
output \digest[123] ;
output \digest[124] ;
output \digest[125] ;
output \digest[126] ;
output \digest[127] ;
output \digest[128] ;
output \digest[129] ;
output \digest[12] ;
output \digest[130] ;
output \digest[131] ;
output \digest[132] ;
output \digest[133] ;
output \digest[134] ;
output \digest[135] ;
output \digest[136] ;
output \digest[137] ;
output \digest[138] ;
output \digest[139] ;
output \digest[13] ;
output \digest[140] ;
output \digest[141] ;
output \digest[142] ;
output \digest[143] ;
output \digest[144] ;
output \digest[145] ;
output \digest[146] ;
output \digest[147] ;
output \digest[148] ;
output \digest[149] ;
output \digest[14] ;
output \digest[150] ;
output \digest[151] ;
output \digest[152] ;
output \digest[153] ;
output \digest[154] ;
output \digest[155] ;
output \digest[156] ;
output \digest[157] ;
output \digest[158] ;
output \digest[159] ;
output \digest[15] ;
output \digest[16] ;
output \digest[17] ;
output \digest[18] ;
output \digest[19] ;
output \digest[1] ;
output \digest[20] ;
output \digest[21] ;
output \digest[22] ;
output \digest[23] ;
output \digest[24] ;
output \digest[25] ;
output \digest[26] ;
output \digest[27] ;
output \digest[28] ;
output \digest[29] ;
output \digest[2] ;
output \digest[30] ;
output \digest[31] ;
output \digest[32] ;
output \digest[33] ;
output \digest[34] ;
output \digest[35] ;
output \digest[36] ;
output \digest[37] ;
output \digest[38] ;
output \digest[39] ;
output \digest[3] ;
output \digest[40] ;
output \digest[41] ;
output \digest[42] ;
output \digest[43] ;
output \digest[44] ;
output \digest[45] ;
output \digest[46] ;
output \digest[47] ;
output \digest[48] ;
output \digest[49] ;
output \digest[4] ;
output \digest[50] ;
output \digest[51] ;
output \digest[52] ;
output \digest[53] ;
output \digest[54] ;
output \digest[55] ;
output \digest[56] ;
output \digest[57] ;
output \digest[58] ;
output \digest[59] ;
output \digest[5] ;
output \digest[60] ;
output \digest[61] ;
output \digest[62] ;
output \digest[63] ;
output \digest[64] ;
output \digest[65] ;
output \digest[66] ;
output \digest[67] ;
output \digest[68] ;
output \digest[69] ;
output \digest[6] ;
output \digest[70] ;
output \digest[71] ;
output \digest[72] ;
output \digest[73] ;
output \digest[74] ;
output \digest[75] ;
output \digest[76] ;
output \digest[77] ;
output \digest[78] ;
output \digest[79] ;
output \digest[7] ;
output \digest[80] ;
output \digest[81] ;
output \digest[82] ;
output \digest[83] ;
output \digest[84] ;
output \digest[85] ;
output \digest[86] ;
output \digest[87] ;
output \digest[88] ;
output \digest[89] ;
output \digest[8] ;
output \digest[90] ;
output \digest[91] ;
output \digest[92] ;
output \digest[93] ;
output \digest[94] ;
output \digest[95] ;
output \digest[96] ;
output \digest[97] ;
output \digest[98] ;
output \digest[99] ;
output \digest[9] ;
wire digest_update; 
wire digest_update_bF_buf0; 
wire digest_update_bF_buf1; 
wire digest_update_bF_buf2; 
wire digest_update_bF_buf3; 
wire digest_update_bF_buf4; 
wire digest_update_bF_buf5; 
wire digest_update_bF_buf6; 
wire digest_update_bF_buf7; 
wire digest_update_bF_buf8; 
output digest_valid;
wire e_reg_0_; 
wire e_reg_10_; 
wire e_reg_11_; 
wire e_reg_12_; 
wire e_reg_13_; 
wire e_reg_14_; 
wire e_reg_15_; 
wire e_reg_16_; 
wire e_reg_17_; 
wire e_reg_18_; 
wire e_reg_19_; 
wire e_reg_1_; 
wire e_reg_20_; 
wire e_reg_21_; 
wire e_reg_22_; 
wire e_reg_23_; 
wire e_reg_24_; 
wire e_reg_25_; 
wire e_reg_26_; 
wire e_reg_27_; 
wire e_reg_28_; 
wire e_reg_29_; 
wire e_reg_2_; 
wire e_reg_30_; 
wire e_reg_31_; 
wire e_reg_3_; 
wire e_reg_4_; 
wire e_reg_5_; 
wire e_reg_6_; 
wire e_reg_7_; 
wire e_reg_8_; 
wire e_reg_9_; 
input init;
input next;
output ready;
input reset_n;
wire reset_n_bF_buf0; 
wire reset_n_bF_buf1; 
wire reset_n_bF_buf10; 
wire reset_n_bF_buf11; 
wire reset_n_bF_buf12; 
wire reset_n_bF_buf13; 
wire reset_n_bF_buf14; 
wire reset_n_bF_buf15; 
wire reset_n_bF_buf16; 
wire reset_n_bF_buf17; 
wire reset_n_bF_buf18; 
wire reset_n_bF_buf19; 
wire reset_n_bF_buf2; 
wire reset_n_bF_buf20; 
wire reset_n_bF_buf21; 
wire reset_n_bF_buf22; 
wire reset_n_bF_buf23; 
wire reset_n_bF_buf24; 
wire reset_n_bF_buf25; 
wire reset_n_bF_buf26; 
wire reset_n_bF_buf27; 
wire reset_n_bF_buf28; 
wire reset_n_bF_buf29; 
wire reset_n_bF_buf3; 
wire reset_n_bF_buf30; 
wire reset_n_bF_buf31; 
wire reset_n_bF_buf32; 
wire reset_n_bF_buf33; 
wire reset_n_bF_buf34; 
wire reset_n_bF_buf35; 
wire reset_n_bF_buf36; 
wire reset_n_bF_buf37; 
wire reset_n_bF_buf38; 
wire reset_n_bF_buf39; 
wire reset_n_bF_buf4; 
wire reset_n_bF_buf40; 
wire reset_n_bF_buf41; 
wire reset_n_bF_buf42; 
wire reset_n_bF_buf43; 
wire reset_n_bF_buf44; 
wire reset_n_bF_buf45; 
wire reset_n_bF_buf46; 
wire reset_n_bF_buf47; 
wire reset_n_bF_buf48; 
wire reset_n_bF_buf49; 
wire reset_n_bF_buf5; 
wire reset_n_bF_buf50; 
wire reset_n_bF_buf51; 
wire reset_n_bF_buf52; 
wire reset_n_bF_buf53; 
wire reset_n_bF_buf54; 
wire reset_n_bF_buf55; 
wire reset_n_bF_buf56; 
wire reset_n_bF_buf57; 
wire reset_n_bF_buf58; 
wire reset_n_bF_buf59; 
wire reset_n_bF_buf6; 
wire reset_n_bF_buf60; 
wire reset_n_bF_buf61; 
wire reset_n_bF_buf62; 
wire reset_n_bF_buf63; 
wire reset_n_bF_buf64; 
wire reset_n_bF_buf65; 
wire reset_n_bF_buf66; 
wire reset_n_bF_buf67; 
wire reset_n_bF_buf68; 
wire reset_n_bF_buf69; 
wire reset_n_bF_buf7; 
wire reset_n_bF_buf70; 
wire reset_n_bF_buf71; 
wire reset_n_bF_buf72; 
wire reset_n_bF_buf73; 
wire reset_n_bF_buf74; 
wire reset_n_bF_buf75; 
wire reset_n_bF_buf76; 
wire reset_n_bF_buf77; 
wire reset_n_bF_buf78; 
wire reset_n_bF_buf79; 
wire reset_n_bF_buf8; 
wire reset_n_bF_buf80; 
wire reset_n_bF_buf81; 
wire reset_n_bF_buf82; 
wire reset_n_bF_buf83; 
wire reset_n_bF_buf84; 
wire reset_n_bF_buf85; 
wire reset_n_bF_buf86; 
wire reset_n_bF_buf87; 
wire reset_n_bF_buf88; 
wire reset_n_bF_buf9; 
wire reset_n_hier0_bF_buf0; 
wire reset_n_hier0_bF_buf1; 
wire reset_n_hier0_bF_buf2; 
wire reset_n_hier0_bF_buf3; 
wire reset_n_hier0_bF_buf4; 
wire reset_n_hier0_bF_buf5; 
wire reset_n_hier0_bF_buf6; 
wire reset_n_hier0_bF_buf7; 
wire reset_n_hier0_bF_buf8; 
wire round_ctr_inc; 
wire round_ctr_inc_bF_buf0; 
wire round_ctr_inc_bF_buf1; 
wire round_ctr_inc_bF_buf10; 
wire round_ctr_inc_bF_buf11; 
wire round_ctr_inc_bF_buf12; 
wire round_ctr_inc_bF_buf13; 
wire round_ctr_inc_bF_buf2; 
wire round_ctr_inc_bF_buf3; 
wire round_ctr_inc_bF_buf4; 
wire round_ctr_inc_bF_buf5; 
wire round_ctr_inc_bF_buf6; 
wire round_ctr_inc_bF_buf7; 
wire round_ctr_inc_bF_buf8; 
wire round_ctr_inc_bF_buf9; 
wire round_ctr_reg_0_; 
wire round_ctr_reg_1_; 
wire round_ctr_reg_2_; 
wire round_ctr_reg_3_; 
wire round_ctr_reg_4_; 
wire round_ctr_reg_5_; 
wire round_ctr_reg_6_; 
wire round_ctr_rst; 
wire round_ctr_rst_bF_buf0; 
wire round_ctr_rst_bF_buf1; 
wire round_ctr_rst_bF_buf2; 
wire round_ctr_rst_bF_buf3; 
wire round_ctr_rst_bF_buf4; 
wire round_ctr_rst_bF_buf5; 
wire round_ctr_rst_bF_buf6; 
wire round_ctr_rst_bF_buf7; 
wire round_ctr_rst_bF_buf8; 
wire w_0_; 
wire w_10_; 
wire w_11_; 
wire w_12_; 
wire w_13_; 
wire w_14_; 
wire w_15_; 
wire w_16_; 
wire w_17_; 
wire w_18_; 
wire w_19_; 
wire w_1_; 
wire w_20_; 
wire w_21_; 
wire w_22_; 
wire w_23_; 
wire w_24_; 
wire w_25_; 
wire w_26_; 
wire w_27_; 
wire w_28_; 
wire w_29_; 
wire w_2_; 
wire w_30_; 
wire w_31_; 
wire w_3_; 
wire w_4_; 
wire w_5_; 
wire w_6_; 
wire w_7_; 
wire w_8_; 
wire w_9_; 
wire w_mem_inst__0w_ctr_reg_6_0__0_; 
wire w_mem_inst__0w_ctr_reg_6_0__1_; 
wire w_mem_inst__0w_ctr_reg_6_0__2_; 
wire w_mem_inst__0w_ctr_reg_6_0__3_; 
wire w_mem_inst__0w_ctr_reg_6_0__4_; 
wire w_mem_inst__0w_ctr_reg_6_0__5_; 
wire w_mem_inst__0w_ctr_reg_6_0__6_; 
wire w_mem_inst__0w_mem_0__31_0__0_; 
wire w_mem_inst__0w_mem_0__31_0__10_; 
wire w_mem_inst__0w_mem_0__31_0__11_; 
wire w_mem_inst__0w_mem_0__31_0__12_; 
wire w_mem_inst__0w_mem_0__31_0__13_; 
wire w_mem_inst__0w_mem_0__31_0__14_; 
wire w_mem_inst__0w_mem_0__31_0__15_; 
wire w_mem_inst__0w_mem_0__31_0__16_; 
wire w_mem_inst__0w_mem_0__31_0__17_; 
wire w_mem_inst__0w_mem_0__31_0__18_; 
wire w_mem_inst__0w_mem_0__31_0__19_; 
wire w_mem_inst__0w_mem_0__31_0__1_; 
wire w_mem_inst__0w_mem_0__31_0__20_; 
wire w_mem_inst__0w_mem_0__31_0__21_; 
wire w_mem_inst__0w_mem_0__31_0__22_; 
wire w_mem_inst__0w_mem_0__31_0__23_; 
wire w_mem_inst__0w_mem_0__31_0__24_; 
wire w_mem_inst__0w_mem_0__31_0__25_; 
wire w_mem_inst__0w_mem_0__31_0__26_; 
wire w_mem_inst__0w_mem_0__31_0__27_; 
wire w_mem_inst__0w_mem_0__31_0__28_; 
wire w_mem_inst__0w_mem_0__31_0__29_; 
wire w_mem_inst__0w_mem_0__31_0__2_; 
wire w_mem_inst__0w_mem_0__31_0__30_; 
wire w_mem_inst__0w_mem_0__31_0__31_; 
wire w_mem_inst__0w_mem_0__31_0__3_; 
wire w_mem_inst__0w_mem_0__31_0__4_; 
wire w_mem_inst__0w_mem_0__31_0__5_; 
wire w_mem_inst__0w_mem_0__31_0__6_; 
wire w_mem_inst__0w_mem_0__31_0__7_; 
wire w_mem_inst__0w_mem_0__31_0__8_; 
wire w_mem_inst__0w_mem_0__31_0__9_; 
wire w_mem_inst__0w_mem_10__31_0__0_; 
wire w_mem_inst__0w_mem_10__31_0__10_; 
wire w_mem_inst__0w_mem_10__31_0__11_; 
wire w_mem_inst__0w_mem_10__31_0__12_; 
wire w_mem_inst__0w_mem_10__31_0__13_; 
wire w_mem_inst__0w_mem_10__31_0__14_; 
wire w_mem_inst__0w_mem_10__31_0__15_; 
wire w_mem_inst__0w_mem_10__31_0__16_; 
wire w_mem_inst__0w_mem_10__31_0__17_; 
wire w_mem_inst__0w_mem_10__31_0__18_; 
wire w_mem_inst__0w_mem_10__31_0__19_; 
wire w_mem_inst__0w_mem_10__31_0__1_; 
wire w_mem_inst__0w_mem_10__31_0__20_; 
wire w_mem_inst__0w_mem_10__31_0__21_; 
wire w_mem_inst__0w_mem_10__31_0__22_; 
wire w_mem_inst__0w_mem_10__31_0__23_; 
wire w_mem_inst__0w_mem_10__31_0__24_; 
wire w_mem_inst__0w_mem_10__31_0__25_; 
wire w_mem_inst__0w_mem_10__31_0__26_; 
wire w_mem_inst__0w_mem_10__31_0__27_; 
wire w_mem_inst__0w_mem_10__31_0__28_; 
wire w_mem_inst__0w_mem_10__31_0__29_; 
wire w_mem_inst__0w_mem_10__31_0__2_; 
wire w_mem_inst__0w_mem_10__31_0__30_; 
wire w_mem_inst__0w_mem_10__31_0__31_; 
wire w_mem_inst__0w_mem_10__31_0__3_; 
wire w_mem_inst__0w_mem_10__31_0__4_; 
wire w_mem_inst__0w_mem_10__31_0__5_; 
wire w_mem_inst__0w_mem_10__31_0__6_; 
wire w_mem_inst__0w_mem_10__31_0__7_; 
wire w_mem_inst__0w_mem_10__31_0__8_; 
wire w_mem_inst__0w_mem_10__31_0__9_; 
wire w_mem_inst__0w_mem_11__31_0__0_; 
wire w_mem_inst__0w_mem_11__31_0__10_; 
wire w_mem_inst__0w_mem_11__31_0__11_; 
wire w_mem_inst__0w_mem_11__31_0__12_; 
wire w_mem_inst__0w_mem_11__31_0__13_; 
wire w_mem_inst__0w_mem_11__31_0__14_; 
wire w_mem_inst__0w_mem_11__31_0__15_; 
wire w_mem_inst__0w_mem_11__31_0__16_; 
wire w_mem_inst__0w_mem_11__31_0__17_; 
wire w_mem_inst__0w_mem_11__31_0__18_; 
wire w_mem_inst__0w_mem_11__31_0__19_; 
wire w_mem_inst__0w_mem_11__31_0__1_; 
wire w_mem_inst__0w_mem_11__31_0__20_; 
wire w_mem_inst__0w_mem_11__31_0__21_; 
wire w_mem_inst__0w_mem_11__31_0__22_; 
wire w_mem_inst__0w_mem_11__31_0__23_; 
wire w_mem_inst__0w_mem_11__31_0__24_; 
wire w_mem_inst__0w_mem_11__31_0__25_; 
wire w_mem_inst__0w_mem_11__31_0__26_; 
wire w_mem_inst__0w_mem_11__31_0__27_; 
wire w_mem_inst__0w_mem_11__31_0__28_; 
wire w_mem_inst__0w_mem_11__31_0__29_; 
wire w_mem_inst__0w_mem_11__31_0__2_; 
wire w_mem_inst__0w_mem_11__31_0__30_; 
wire w_mem_inst__0w_mem_11__31_0__31_; 
wire w_mem_inst__0w_mem_11__31_0__3_; 
wire w_mem_inst__0w_mem_11__31_0__4_; 
wire w_mem_inst__0w_mem_11__31_0__5_; 
wire w_mem_inst__0w_mem_11__31_0__6_; 
wire w_mem_inst__0w_mem_11__31_0__7_; 
wire w_mem_inst__0w_mem_11__31_0__8_; 
wire w_mem_inst__0w_mem_11__31_0__9_; 
wire w_mem_inst__0w_mem_12__31_0__0_; 
wire w_mem_inst__0w_mem_12__31_0__10_; 
wire w_mem_inst__0w_mem_12__31_0__11_; 
wire w_mem_inst__0w_mem_12__31_0__12_; 
wire w_mem_inst__0w_mem_12__31_0__13_; 
wire w_mem_inst__0w_mem_12__31_0__14_; 
wire w_mem_inst__0w_mem_12__31_0__15_; 
wire w_mem_inst__0w_mem_12__31_0__16_; 
wire w_mem_inst__0w_mem_12__31_0__17_; 
wire w_mem_inst__0w_mem_12__31_0__18_; 
wire w_mem_inst__0w_mem_12__31_0__19_; 
wire w_mem_inst__0w_mem_12__31_0__1_; 
wire w_mem_inst__0w_mem_12__31_0__20_; 
wire w_mem_inst__0w_mem_12__31_0__21_; 
wire w_mem_inst__0w_mem_12__31_0__22_; 
wire w_mem_inst__0w_mem_12__31_0__23_; 
wire w_mem_inst__0w_mem_12__31_0__24_; 
wire w_mem_inst__0w_mem_12__31_0__25_; 
wire w_mem_inst__0w_mem_12__31_0__26_; 
wire w_mem_inst__0w_mem_12__31_0__27_; 
wire w_mem_inst__0w_mem_12__31_0__28_; 
wire w_mem_inst__0w_mem_12__31_0__29_; 
wire w_mem_inst__0w_mem_12__31_0__2_; 
wire w_mem_inst__0w_mem_12__31_0__30_; 
wire w_mem_inst__0w_mem_12__31_0__31_; 
wire w_mem_inst__0w_mem_12__31_0__3_; 
wire w_mem_inst__0w_mem_12__31_0__4_; 
wire w_mem_inst__0w_mem_12__31_0__5_; 
wire w_mem_inst__0w_mem_12__31_0__6_; 
wire w_mem_inst__0w_mem_12__31_0__7_; 
wire w_mem_inst__0w_mem_12__31_0__8_; 
wire w_mem_inst__0w_mem_12__31_0__9_; 
wire w_mem_inst__0w_mem_13__31_0__0_; 
wire w_mem_inst__0w_mem_13__31_0__10_; 
wire w_mem_inst__0w_mem_13__31_0__11_; 
wire w_mem_inst__0w_mem_13__31_0__12_; 
wire w_mem_inst__0w_mem_13__31_0__13_; 
wire w_mem_inst__0w_mem_13__31_0__14_; 
wire w_mem_inst__0w_mem_13__31_0__15_; 
wire w_mem_inst__0w_mem_13__31_0__16_; 
wire w_mem_inst__0w_mem_13__31_0__17_; 
wire w_mem_inst__0w_mem_13__31_0__18_; 
wire w_mem_inst__0w_mem_13__31_0__19_; 
wire w_mem_inst__0w_mem_13__31_0__1_; 
wire w_mem_inst__0w_mem_13__31_0__20_; 
wire w_mem_inst__0w_mem_13__31_0__21_; 
wire w_mem_inst__0w_mem_13__31_0__22_; 
wire w_mem_inst__0w_mem_13__31_0__23_; 
wire w_mem_inst__0w_mem_13__31_0__24_; 
wire w_mem_inst__0w_mem_13__31_0__25_; 
wire w_mem_inst__0w_mem_13__31_0__26_; 
wire w_mem_inst__0w_mem_13__31_0__27_; 
wire w_mem_inst__0w_mem_13__31_0__28_; 
wire w_mem_inst__0w_mem_13__31_0__29_; 
wire w_mem_inst__0w_mem_13__31_0__2_; 
wire w_mem_inst__0w_mem_13__31_0__30_; 
wire w_mem_inst__0w_mem_13__31_0__31_; 
wire w_mem_inst__0w_mem_13__31_0__3_; 
wire w_mem_inst__0w_mem_13__31_0__4_; 
wire w_mem_inst__0w_mem_13__31_0__5_; 
wire w_mem_inst__0w_mem_13__31_0__6_; 
wire w_mem_inst__0w_mem_13__31_0__7_; 
wire w_mem_inst__0w_mem_13__31_0__8_; 
wire w_mem_inst__0w_mem_13__31_0__9_; 
wire w_mem_inst__0w_mem_14__31_0__0_; 
wire w_mem_inst__0w_mem_14__31_0__10_; 
wire w_mem_inst__0w_mem_14__31_0__11_; 
wire w_mem_inst__0w_mem_14__31_0__12_; 
wire w_mem_inst__0w_mem_14__31_0__13_; 
wire w_mem_inst__0w_mem_14__31_0__14_; 
wire w_mem_inst__0w_mem_14__31_0__15_; 
wire w_mem_inst__0w_mem_14__31_0__16_; 
wire w_mem_inst__0w_mem_14__31_0__17_; 
wire w_mem_inst__0w_mem_14__31_0__18_; 
wire w_mem_inst__0w_mem_14__31_0__19_; 
wire w_mem_inst__0w_mem_14__31_0__1_; 
wire w_mem_inst__0w_mem_14__31_0__20_; 
wire w_mem_inst__0w_mem_14__31_0__21_; 
wire w_mem_inst__0w_mem_14__31_0__22_; 
wire w_mem_inst__0w_mem_14__31_0__23_; 
wire w_mem_inst__0w_mem_14__31_0__24_; 
wire w_mem_inst__0w_mem_14__31_0__25_; 
wire w_mem_inst__0w_mem_14__31_0__26_; 
wire w_mem_inst__0w_mem_14__31_0__27_; 
wire w_mem_inst__0w_mem_14__31_0__28_; 
wire w_mem_inst__0w_mem_14__31_0__29_; 
wire w_mem_inst__0w_mem_14__31_0__2_; 
wire w_mem_inst__0w_mem_14__31_0__30_; 
wire w_mem_inst__0w_mem_14__31_0__31_; 
wire w_mem_inst__0w_mem_14__31_0__3_; 
wire w_mem_inst__0w_mem_14__31_0__4_; 
wire w_mem_inst__0w_mem_14__31_0__5_; 
wire w_mem_inst__0w_mem_14__31_0__6_; 
wire w_mem_inst__0w_mem_14__31_0__7_; 
wire w_mem_inst__0w_mem_14__31_0__8_; 
wire w_mem_inst__0w_mem_14__31_0__9_; 
wire w_mem_inst__0w_mem_15__31_0__0_; 
wire w_mem_inst__0w_mem_15__31_0__10_; 
wire w_mem_inst__0w_mem_15__31_0__11_; 
wire w_mem_inst__0w_mem_15__31_0__12_; 
wire w_mem_inst__0w_mem_15__31_0__13_; 
wire w_mem_inst__0w_mem_15__31_0__14_; 
wire w_mem_inst__0w_mem_15__31_0__15_; 
wire w_mem_inst__0w_mem_15__31_0__16_; 
wire w_mem_inst__0w_mem_15__31_0__17_; 
wire w_mem_inst__0w_mem_15__31_0__18_; 
wire w_mem_inst__0w_mem_15__31_0__19_; 
wire w_mem_inst__0w_mem_15__31_0__1_; 
wire w_mem_inst__0w_mem_15__31_0__20_; 
wire w_mem_inst__0w_mem_15__31_0__21_; 
wire w_mem_inst__0w_mem_15__31_0__22_; 
wire w_mem_inst__0w_mem_15__31_0__23_; 
wire w_mem_inst__0w_mem_15__31_0__24_; 
wire w_mem_inst__0w_mem_15__31_0__25_; 
wire w_mem_inst__0w_mem_15__31_0__26_; 
wire w_mem_inst__0w_mem_15__31_0__27_; 
wire w_mem_inst__0w_mem_15__31_0__28_; 
wire w_mem_inst__0w_mem_15__31_0__29_; 
wire w_mem_inst__0w_mem_15__31_0__2_; 
wire w_mem_inst__0w_mem_15__31_0__30_; 
wire w_mem_inst__0w_mem_15__31_0__31_; 
wire w_mem_inst__0w_mem_15__31_0__3_; 
wire w_mem_inst__0w_mem_15__31_0__4_; 
wire w_mem_inst__0w_mem_15__31_0__5_; 
wire w_mem_inst__0w_mem_15__31_0__6_; 
wire w_mem_inst__0w_mem_15__31_0__7_; 
wire w_mem_inst__0w_mem_15__31_0__8_; 
wire w_mem_inst__0w_mem_15__31_0__9_; 
wire w_mem_inst__0w_mem_1__31_0__0_; 
wire w_mem_inst__0w_mem_1__31_0__10_; 
wire w_mem_inst__0w_mem_1__31_0__11_; 
wire w_mem_inst__0w_mem_1__31_0__12_; 
wire w_mem_inst__0w_mem_1__31_0__13_; 
wire w_mem_inst__0w_mem_1__31_0__14_; 
wire w_mem_inst__0w_mem_1__31_0__15_; 
wire w_mem_inst__0w_mem_1__31_0__16_; 
wire w_mem_inst__0w_mem_1__31_0__17_; 
wire w_mem_inst__0w_mem_1__31_0__18_; 
wire w_mem_inst__0w_mem_1__31_0__19_; 
wire w_mem_inst__0w_mem_1__31_0__1_; 
wire w_mem_inst__0w_mem_1__31_0__20_; 
wire w_mem_inst__0w_mem_1__31_0__21_; 
wire w_mem_inst__0w_mem_1__31_0__22_; 
wire w_mem_inst__0w_mem_1__31_0__23_; 
wire w_mem_inst__0w_mem_1__31_0__24_; 
wire w_mem_inst__0w_mem_1__31_0__25_; 
wire w_mem_inst__0w_mem_1__31_0__26_; 
wire w_mem_inst__0w_mem_1__31_0__27_; 
wire w_mem_inst__0w_mem_1__31_0__28_; 
wire w_mem_inst__0w_mem_1__31_0__29_; 
wire w_mem_inst__0w_mem_1__31_0__2_; 
wire w_mem_inst__0w_mem_1__31_0__30_; 
wire w_mem_inst__0w_mem_1__31_0__31_; 
wire w_mem_inst__0w_mem_1__31_0__3_; 
wire w_mem_inst__0w_mem_1__31_0__4_; 
wire w_mem_inst__0w_mem_1__31_0__5_; 
wire w_mem_inst__0w_mem_1__31_0__6_; 
wire w_mem_inst__0w_mem_1__31_0__7_; 
wire w_mem_inst__0w_mem_1__31_0__8_; 
wire w_mem_inst__0w_mem_1__31_0__9_; 
wire w_mem_inst__0w_mem_2__31_0__0_; 
wire w_mem_inst__0w_mem_2__31_0__10_; 
wire w_mem_inst__0w_mem_2__31_0__11_; 
wire w_mem_inst__0w_mem_2__31_0__12_; 
wire w_mem_inst__0w_mem_2__31_0__13_; 
wire w_mem_inst__0w_mem_2__31_0__14_; 
wire w_mem_inst__0w_mem_2__31_0__15_; 
wire w_mem_inst__0w_mem_2__31_0__16_; 
wire w_mem_inst__0w_mem_2__31_0__17_; 
wire w_mem_inst__0w_mem_2__31_0__18_; 
wire w_mem_inst__0w_mem_2__31_0__19_; 
wire w_mem_inst__0w_mem_2__31_0__1_; 
wire w_mem_inst__0w_mem_2__31_0__20_; 
wire w_mem_inst__0w_mem_2__31_0__21_; 
wire w_mem_inst__0w_mem_2__31_0__22_; 
wire w_mem_inst__0w_mem_2__31_0__23_; 
wire w_mem_inst__0w_mem_2__31_0__24_; 
wire w_mem_inst__0w_mem_2__31_0__25_; 
wire w_mem_inst__0w_mem_2__31_0__26_; 
wire w_mem_inst__0w_mem_2__31_0__27_; 
wire w_mem_inst__0w_mem_2__31_0__28_; 
wire w_mem_inst__0w_mem_2__31_0__29_; 
wire w_mem_inst__0w_mem_2__31_0__2_; 
wire w_mem_inst__0w_mem_2__31_0__30_; 
wire w_mem_inst__0w_mem_2__31_0__31_; 
wire w_mem_inst__0w_mem_2__31_0__3_; 
wire w_mem_inst__0w_mem_2__31_0__4_; 
wire w_mem_inst__0w_mem_2__31_0__5_; 
wire w_mem_inst__0w_mem_2__31_0__6_; 
wire w_mem_inst__0w_mem_2__31_0__7_; 
wire w_mem_inst__0w_mem_2__31_0__8_; 
wire w_mem_inst__0w_mem_2__31_0__9_; 
wire w_mem_inst__0w_mem_3__31_0__0_; 
wire w_mem_inst__0w_mem_3__31_0__10_; 
wire w_mem_inst__0w_mem_3__31_0__11_; 
wire w_mem_inst__0w_mem_3__31_0__12_; 
wire w_mem_inst__0w_mem_3__31_0__13_; 
wire w_mem_inst__0w_mem_3__31_0__14_; 
wire w_mem_inst__0w_mem_3__31_0__15_; 
wire w_mem_inst__0w_mem_3__31_0__16_; 
wire w_mem_inst__0w_mem_3__31_0__17_; 
wire w_mem_inst__0w_mem_3__31_0__18_; 
wire w_mem_inst__0w_mem_3__31_0__19_; 
wire w_mem_inst__0w_mem_3__31_0__1_; 
wire w_mem_inst__0w_mem_3__31_0__20_; 
wire w_mem_inst__0w_mem_3__31_0__21_; 
wire w_mem_inst__0w_mem_3__31_0__22_; 
wire w_mem_inst__0w_mem_3__31_0__23_; 
wire w_mem_inst__0w_mem_3__31_0__24_; 
wire w_mem_inst__0w_mem_3__31_0__25_; 
wire w_mem_inst__0w_mem_3__31_0__26_; 
wire w_mem_inst__0w_mem_3__31_0__27_; 
wire w_mem_inst__0w_mem_3__31_0__28_; 
wire w_mem_inst__0w_mem_3__31_0__29_; 
wire w_mem_inst__0w_mem_3__31_0__2_; 
wire w_mem_inst__0w_mem_3__31_0__30_; 
wire w_mem_inst__0w_mem_3__31_0__31_; 
wire w_mem_inst__0w_mem_3__31_0__3_; 
wire w_mem_inst__0w_mem_3__31_0__4_; 
wire w_mem_inst__0w_mem_3__31_0__5_; 
wire w_mem_inst__0w_mem_3__31_0__6_; 
wire w_mem_inst__0w_mem_3__31_0__7_; 
wire w_mem_inst__0w_mem_3__31_0__8_; 
wire w_mem_inst__0w_mem_3__31_0__9_; 
wire w_mem_inst__0w_mem_4__31_0__0_; 
wire w_mem_inst__0w_mem_4__31_0__10_; 
wire w_mem_inst__0w_mem_4__31_0__11_; 
wire w_mem_inst__0w_mem_4__31_0__12_; 
wire w_mem_inst__0w_mem_4__31_0__13_; 
wire w_mem_inst__0w_mem_4__31_0__14_; 
wire w_mem_inst__0w_mem_4__31_0__15_; 
wire w_mem_inst__0w_mem_4__31_0__16_; 
wire w_mem_inst__0w_mem_4__31_0__17_; 
wire w_mem_inst__0w_mem_4__31_0__18_; 
wire w_mem_inst__0w_mem_4__31_0__19_; 
wire w_mem_inst__0w_mem_4__31_0__1_; 
wire w_mem_inst__0w_mem_4__31_0__20_; 
wire w_mem_inst__0w_mem_4__31_0__21_; 
wire w_mem_inst__0w_mem_4__31_0__22_; 
wire w_mem_inst__0w_mem_4__31_0__23_; 
wire w_mem_inst__0w_mem_4__31_0__24_; 
wire w_mem_inst__0w_mem_4__31_0__25_; 
wire w_mem_inst__0w_mem_4__31_0__26_; 
wire w_mem_inst__0w_mem_4__31_0__27_; 
wire w_mem_inst__0w_mem_4__31_0__28_; 
wire w_mem_inst__0w_mem_4__31_0__29_; 
wire w_mem_inst__0w_mem_4__31_0__2_; 
wire w_mem_inst__0w_mem_4__31_0__30_; 
wire w_mem_inst__0w_mem_4__31_0__31_; 
wire w_mem_inst__0w_mem_4__31_0__3_; 
wire w_mem_inst__0w_mem_4__31_0__4_; 
wire w_mem_inst__0w_mem_4__31_0__5_; 
wire w_mem_inst__0w_mem_4__31_0__6_; 
wire w_mem_inst__0w_mem_4__31_0__7_; 
wire w_mem_inst__0w_mem_4__31_0__8_; 
wire w_mem_inst__0w_mem_4__31_0__9_; 
wire w_mem_inst__0w_mem_5__31_0__0_; 
wire w_mem_inst__0w_mem_5__31_0__10_; 
wire w_mem_inst__0w_mem_5__31_0__11_; 
wire w_mem_inst__0w_mem_5__31_0__12_; 
wire w_mem_inst__0w_mem_5__31_0__13_; 
wire w_mem_inst__0w_mem_5__31_0__14_; 
wire w_mem_inst__0w_mem_5__31_0__15_; 
wire w_mem_inst__0w_mem_5__31_0__16_; 
wire w_mem_inst__0w_mem_5__31_0__17_; 
wire w_mem_inst__0w_mem_5__31_0__18_; 
wire w_mem_inst__0w_mem_5__31_0__19_; 
wire w_mem_inst__0w_mem_5__31_0__1_; 
wire w_mem_inst__0w_mem_5__31_0__20_; 
wire w_mem_inst__0w_mem_5__31_0__21_; 
wire w_mem_inst__0w_mem_5__31_0__22_; 
wire w_mem_inst__0w_mem_5__31_0__23_; 
wire w_mem_inst__0w_mem_5__31_0__24_; 
wire w_mem_inst__0w_mem_5__31_0__25_; 
wire w_mem_inst__0w_mem_5__31_0__26_; 
wire w_mem_inst__0w_mem_5__31_0__27_; 
wire w_mem_inst__0w_mem_5__31_0__28_; 
wire w_mem_inst__0w_mem_5__31_0__29_; 
wire w_mem_inst__0w_mem_5__31_0__2_; 
wire w_mem_inst__0w_mem_5__31_0__30_; 
wire w_mem_inst__0w_mem_5__31_0__31_; 
wire w_mem_inst__0w_mem_5__31_0__3_; 
wire w_mem_inst__0w_mem_5__31_0__4_; 
wire w_mem_inst__0w_mem_5__31_0__5_; 
wire w_mem_inst__0w_mem_5__31_0__6_; 
wire w_mem_inst__0w_mem_5__31_0__7_; 
wire w_mem_inst__0w_mem_5__31_0__8_; 
wire w_mem_inst__0w_mem_5__31_0__9_; 
wire w_mem_inst__0w_mem_6__31_0__0_; 
wire w_mem_inst__0w_mem_6__31_0__10_; 
wire w_mem_inst__0w_mem_6__31_0__11_; 
wire w_mem_inst__0w_mem_6__31_0__12_; 
wire w_mem_inst__0w_mem_6__31_0__13_; 
wire w_mem_inst__0w_mem_6__31_0__14_; 
wire w_mem_inst__0w_mem_6__31_0__15_; 
wire w_mem_inst__0w_mem_6__31_0__16_; 
wire w_mem_inst__0w_mem_6__31_0__17_; 
wire w_mem_inst__0w_mem_6__31_0__18_; 
wire w_mem_inst__0w_mem_6__31_0__19_; 
wire w_mem_inst__0w_mem_6__31_0__1_; 
wire w_mem_inst__0w_mem_6__31_0__20_; 
wire w_mem_inst__0w_mem_6__31_0__21_; 
wire w_mem_inst__0w_mem_6__31_0__22_; 
wire w_mem_inst__0w_mem_6__31_0__23_; 
wire w_mem_inst__0w_mem_6__31_0__24_; 
wire w_mem_inst__0w_mem_6__31_0__25_; 
wire w_mem_inst__0w_mem_6__31_0__26_; 
wire w_mem_inst__0w_mem_6__31_0__27_; 
wire w_mem_inst__0w_mem_6__31_0__28_; 
wire w_mem_inst__0w_mem_6__31_0__29_; 
wire w_mem_inst__0w_mem_6__31_0__2_; 
wire w_mem_inst__0w_mem_6__31_0__30_; 
wire w_mem_inst__0w_mem_6__31_0__31_; 
wire w_mem_inst__0w_mem_6__31_0__3_; 
wire w_mem_inst__0w_mem_6__31_0__4_; 
wire w_mem_inst__0w_mem_6__31_0__5_; 
wire w_mem_inst__0w_mem_6__31_0__6_; 
wire w_mem_inst__0w_mem_6__31_0__7_; 
wire w_mem_inst__0w_mem_6__31_0__8_; 
wire w_mem_inst__0w_mem_6__31_0__9_; 
wire w_mem_inst__0w_mem_7__31_0__0_; 
wire w_mem_inst__0w_mem_7__31_0__10_; 
wire w_mem_inst__0w_mem_7__31_0__11_; 
wire w_mem_inst__0w_mem_7__31_0__12_; 
wire w_mem_inst__0w_mem_7__31_0__13_; 
wire w_mem_inst__0w_mem_7__31_0__14_; 
wire w_mem_inst__0w_mem_7__31_0__15_; 
wire w_mem_inst__0w_mem_7__31_0__16_; 
wire w_mem_inst__0w_mem_7__31_0__17_; 
wire w_mem_inst__0w_mem_7__31_0__18_; 
wire w_mem_inst__0w_mem_7__31_0__19_; 
wire w_mem_inst__0w_mem_7__31_0__1_; 
wire w_mem_inst__0w_mem_7__31_0__20_; 
wire w_mem_inst__0w_mem_7__31_0__21_; 
wire w_mem_inst__0w_mem_7__31_0__22_; 
wire w_mem_inst__0w_mem_7__31_0__23_; 
wire w_mem_inst__0w_mem_7__31_0__24_; 
wire w_mem_inst__0w_mem_7__31_0__25_; 
wire w_mem_inst__0w_mem_7__31_0__26_; 
wire w_mem_inst__0w_mem_7__31_0__27_; 
wire w_mem_inst__0w_mem_7__31_0__28_; 
wire w_mem_inst__0w_mem_7__31_0__29_; 
wire w_mem_inst__0w_mem_7__31_0__2_; 
wire w_mem_inst__0w_mem_7__31_0__30_; 
wire w_mem_inst__0w_mem_7__31_0__31_; 
wire w_mem_inst__0w_mem_7__31_0__3_; 
wire w_mem_inst__0w_mem_7__31_0__4_; 
wire w_mem_inst__0w_mem_7__31_0__5_; 
wire w_mem_inst__0w_mem_7__31_0__6_; 
wire w_mem_inst__0w_mem_7__31_0__7_; 
wire w_mem_inst__0w_mem_7__31_0__8_; 
wire w_mem_inst__0w_mem_7__31_0__9_; 
wire w_mem_inst__0w_mem_8__31_0__0_; 
wire w_mem_inst__0w_mem_8__31_0__10_; 
wire w_mem_inst__0w_mem_8__31_0__11_; 
wire w_mem_inst__0w_mem_8__31_0__12_; 
wire w_mem_inst__0w_mem_8__31_0__13_; 
wire w_mem_inst__0w_mem_8__31_0__14_; 
wire w_mem_inst__0w_mem_8__31_0__15_; 
wire w_mem_inst__0w_mem_8__31_0__16_; 
wire w_mem_inst__0w_mem_8__31_0__17_; 
wire w_mem_inst__0w_mem_8__31_0__18_; 
wire w_mem_inst__0w_mem_8__31_0__19_; 
wire w_mem_inst__0w_mem_8__31_0__1_; 
wire w_mem_inst__0w_mem_8__31_0__20_; 
wire w_mem_inst__0w_mem_8__31_0__21_; 
wire w_mem_inst__0w_mem_8__31_0__22_; 
wire w_mem_inst__0w_mem_8__31_0__23_; 
wire w_mem_inst__0w_mem_8__31_0__24_; 
wire w_mem_inst__0w_mem_8__31_0__25_; 
wire w_mem_inst__0w_mem_8__31_0__26_; 
wire w_mem_inst__0w_mem_8__31_0__27_; 
wire w_mem_inst__0w_mem_8__31_0__28_; 
wire w_mem_inst__0w_mem_8__31_0__29_; 
wire w_mem_inst__0w_mem_8__31_0__2_; 
wire w_mem_inst__0w_mem_8__31_0__30_; 
wire w_mem_inst__0w_mem_8__31_0__31_; 
wire w_mem_inst__0w_mem_8__31_0__3_; 
wire w_mem_inst__0w_mem_8__31_0__4_; 
wire w_mem_inst__0w_mem_8__31_0__5_; 
wire w_mem_inst__0w_mem_8__31_0__6_; 
wire w_mem_inst__0w_mem_8__31_0__7_; 
wire w_mem_inst__0w_mem_8__31_0__8_; 
wire w_mem_inst__0w_mem_8__31_0__9_; 
wire w_mem_inst__0w_mem_9__31_0__0_; 
wire w_mem_inst__0w_mem_9__31_0__10_; 
wire w_mem_inst__0w_mem_9__31_0__11_; 
wire w_mem_inst__0w_mem_9__31_0__12_; 
wire w_mem_inst__0w_mem_9__31_0__13_; 
wire w_mem_inst__0w_mem_9__31_0__14_; 
wire w_mem_inst__0w_mem_9__31_0__15_; 
wire w_mem_inst__0w_mem_9__31_0__16_; 
wire w_mem_inst__0w_mem_9__31_0__17_; 
wire w_mem_inst__0w_mem_9__31_0__18_; 
wire w_mem_inst__0w_mem_9__31_0__19_; 
wire w_mem_inst__0w_mem_9__31_0__1_; 
wire w_mem_inst__0w_mem_9__31_0__20_; 
wire w_mem_inst__0w_mem_9__31_0__21_; 
wire w_mem_inst__0w_mem_9__31_0__22_; 
wire w_mem_inst__0w_mem_9__31_0__23_; 
wire w_mem_inst__0w_mem_9__31_0__24_; 
wire w_mem_inst__0w_mem_9__31_0__25_; 
wire w_mem_inst__0w_mem_9__31_0__26_; 
wire w_mem_inst__0w_mem_9__31_0__27_; 
wire w_mem_inst__0w_mem_9__31_0__28_; 
wire w_mem_inst__0w_mem_9__31_0__29_; 
wire w_mem_inst__0w_mem_9__31_0__2_; 
wire w_mem_inst__0w_mem_9__31_0__30_; 
wire w_mem_inst__0w_mem_9__31_0__31_; 
wire w_mem_inst__0w_mem_9__31_0__3_; 
wire w_mem_inst__0w_mem_9__31_0__4_; 
wire w_mem_inst__0w_mem_9__31_0__5_; 
wire w_mem_inst__0w_mem_9__31_0__6_; 
wire w_mem_inst__0w_mem_9__31_0__7_; 
wire w_mem_inst__0w_mem_9__31_0__8_; 
wire w_mem_inst__0w_mem_9__31_0__9_; 
wire w_mem_inst__abc_19396_new_n1585_; 
wire w_mem_inst__abc_19396_new_n1586_; 
wire w_mem_inst__abc_19396_new_n1586__bF_buf0; 
wire w_mem_inst__abc_19396_new_n1586__bF_buf1; 
wire w_mem_inst__abc_19396_new_n1586__bF_buf2; 
wire w_mem_inst__abc_19396_new_n1586__bF_buf3; 
wire w_mem_inst__abc_19396_new_n1586__bF_buf4; 
wire w_mem_inst__abc_19396_new_n1587_; 
wire w_mem_inst__abc_19396_new_n1587__bF_buf0; 
wire w_mem_inst__abc_19396_new_n1587__bF_buf1; 
wire w_mem_inst__abc_19396_new_n1587__bF_buf2; 
wire w_mem_inst__abc_19396_new_n1587__bF_buf3; 
wire w_mem_inst__abc_19396_new_n1587__bF_buf4; 
wire w_mem_inst__abc_19396_new_n1588_; 
wire w_mem_inst__abc_19396_new_n1589_; 
wire w_mem_inst__abc_19396_new_n1590_; 
wire w_mem_inst__abc_19396_new_n1591_; 
wire w_mem_inst__abc_19396_new_n1592_; 
wire w_mem_inst__abc_19396_new_n1593_; 
wire w_mem_inst__abc_19396_new_n1594_; 
wire w_mem_inst__abc_19396_new_n1594__bF_buf0; 
wire w_mem_inst__abc_19396_new_n1594__bF_buf1; 
wire w_mem_inst__abc_19396_new_n1594__bF_buf2; 
wire w_mem_inst__abc_19396_new_n1594__bF_buf3; 
wire w_mem_inst__abc_19396_new_n1594__bF_buf4; 
wire w_mem_inst__abc_19396_new_n1594__bF_buf5; 
wire w_mem_inst__abc_19396_new_n1594__bF_buf6; 
wire w_mem_inst__abc_19396_new_n1594__bF_buf7; 
wire w_mem_inst__abc_19396_new_n1595_; 
wire w_mem_inst__abc_19396_new_n1596_; 
wire w_mem_inst__abc_19396_new_n1597_; 
wire w_mem_inst__abc_19396_new_n1598_; 
wire w_mem_inst__abc_19396_new_n1598__bF_buf0; 
wire w_mem_inst__abc_19396_new_n1598__bF_buf1; 
wire w_mem_inst__abc_19396_new_n1598__bF_buf2; 
wire w_mem_inst__abc_19396_new_n1598__bF_buf3; 
wire w_mem_inst__abc_19396_new_n1598__bF_buf4; 
wire w_mem_inst__abc_19396_new_n1599_; 
wire w_mem_inst__abc_19396_new_n1600_; 
wire w_mem_inst__abc_19396_new_n1601_; 
wire w_mem_inst__abc_19396_new_n1602_; 
wire w_mem_inst__abc_19396_new_n1603_; 
wire w_mem_inst__abc_19396_new_n1604_; 
wire w_mem_inst__abc_19396_new_n1604__bF_buf0; 
wire w_mem_inst__abc_19396_new_n1604__bF_buf1; 
wire w_mem_inst__abc_19396_new_n1604__bF_buf2; 
wire w_mem_inst__abc_19396_new_n1604__bF_buf3; 
wire w_mem_inst__abc_19396_new_n1604__bF_buf4; 
wire w_mem_inst__abc_19396_new_n1605_; 
wire w_mem_inst__abc_19396_new_n1606_; 
wire w_mem_inst__abc_19396_new_n1606__bF_buf0; 
wire w_mem_inst__abc_19396_new_n1606__bF_buf1; 
wire w_mem_inst__abc_19396_new_n1606__bF_buf2; 
wire w_mem_inst__abc_19396_new_n1606__bF_buf3; 
wire w_mem_inst__abc_19396_new_n1606__bF_buf4; 
wire w_mem_inst__abc_19396_new_n1607_; 
wire w_mem_inst__abc_19396_new_n1608_; 
wire w_mem_inst__abc_19396_new_n1609_; 
wire w_mem_inst__abc_19396_new_n1610_; 
wire w_mem_inst__abc_19396_new_n1611_; 
wire w_mem_inst__abc_19396_new_n1611__bF_buf0; 
wire w_mem_inst__abc_19396_new_n1611__bF_buf1; 
wire w_mem_inst__abc_19396_new_n1611__bF_buf2; 
wire w_mem_inst__abc_19396_new_n1611__bF_buf3; 
wire w_mem_inst__abc_19396_new_n1611__bF_buf4; 
wire w_mem_inst__abc_19396_new_n1612_; 
wire w_mem_inst__abc_19396_new_n1613_; 
wire w_mem_inst__abc_19396_new_n1613__bF_buf0; 
wire w_mem_inst__abc_19396_new_n1613__bF_buf1; 
wire w_mem_inst__abc_19396_new_n1613__bF_buf2; 
wire w_mem_inst__abc_19396_new_n1613__bF_buf3; 
wire w_mem_inst__abc_19396_new_n1613__bF_buf4; 
wire w_mem_inst__abc_19396_new_n1614_; 
wire w_mem_inst__abc_19396_new_n1615_; 
wire w_mem_inst__abc_19396_new_n1616_; 
wire w_mem_inst__abc_19396_new_n1617_; 
wire w_mem_inst__abc_19396_new_n1617__bF_buf0; 
wire w_mem_inst__abc_19396_new_n1617__bF_buf1; 
wire w_mem_inst__abc_19396_new_n1617__bF_buf2; 
wire w_mem_inst__abc_19396_new_n1617__bF_buf3; 
wire w_mem_inst__abc_19396_new_n1617__bF_buf4; 
wire w_mem_inst__abc_19396_new_n1617__bF_buf5; 
wire w_mem_inst__abc_19396_new_n1617__bF_buf6; 
wire w_mem_inst__abc_19396_new_n1617__bF_buf7; 
wire w_mem_inst__abc_19396_new_n1618_; 
wire w_mem_inst__abc_19396_new_n1619_; 
wire w_mem_inst__abc_19396_new_n1619__bF_buf0; 
wire w_mem_inst__abc_19396_new_n1619__bF_buf1; 
wire w_mem_inst__abc_19396_new_n1619__bF_buf2; 
wire w_mem_inst__abc_19396_new_n1619__bF_buf3; 
wire w_mem_inst__abc_19396_new_n1619__bF_buf4; 
wire w_mem_inst__abc_19396_new_n1620_; 
wire w_mem_inst__abc_19396_new_n1620__bF_buf0; 
wire w_mem_inst__abc_19396_new_n1620__bF_buf1; 
wire w_mem_inst__abc_19396_new_n1620__bF_buf2; 
wire w_mem_inst__abc_19396_new_n1620__bF_buf3; 
wire w_mem_inst__abc_19396_new_n1620__bF_buf4; 
wire w_mem_inst__abc_19396_new_n1620__bF_buf5; 
wire w_mem_inst__abc_19396_new_n1620__bF_buf6; 
wire w_mem_inst__abc_19396_new_n1620__bF_buf7; 
wire w_mem_inst__abc_19396_new_n1621_; 
wire w_mem_inst__abc_19396_new_n1621__bF_buf0; 
wire w_mem_inst__abc_19396_new_n1621__bF_buf1; 
wire w_mem_inst__abc_19396_new_n1621__bF_buf2; 
wire w_mem_inst__abc_19396_new_n1621__bF_buf3; 
wire w_mem_inst__abc_19396_new_n1621__bF_buf4; 
wire w_mem_inst__abc_19396_new_n1622_; 
wire w_mem_inst__abc_19396_new_n1623_; 
wire w_mem_inst__abc_19396_new_n1624_; 
wire w_mem_inst__abc_19396_new_n1625_; 
wire w_mem_inst__abc_19396_new_n1625__bF_buf0; 
wire w_mem_inst__abc_19396_new_n1625__bF_buf1; 
wire w_mem_inst__abc_19396_new_n1625__bF_buf2; 
wire w_mem_inst__abc_19396_new_n1625__bF_buf3; 
wire w_mem_inst__abc_19396_new_n1625__bF_buf4; 
wire w_mem_inst__abc_19396_new_n1626_; 
wire w_mem_inst__abc_19396_new_n1627_; 
wire w_mem_inst__abc_19396_new_n1628_; 
wire w_mem_inst__abc_19396_new_n1628__bF_buf0; 
wire w_mem_inst__abc_19396_new_n1628__bF_buf1; 
wire w_mem_inst__abc_19396_new_n1628__bF_buf2; 
wire w_mem_inst__abc_19396_new_n1628__bF_buf3; 
wire w_mem_inst__abc_19396_new_n1628__bF_buf4; 
wire w_mem_inst__abc_19396_new_n1629_; 
wire w_mem_inst__abc_19396_new_n1630_; 
wire w_mem_inst__abc_19396_new_n1630__bF_buf0; 
wire w_mem_inst__abc_19396_new_n1630__bF_buf1; 
wire w_mem_inst__abc_19396_new_n1630__bF_buf2; 
wire w_mem_inst__abc_19396_new_n1630__bF_buf3; 
wire w_mem_inst__abc_19396_new_n1630__bF_buf4; 
wire w_mem_inst__abc_19396_new_n1631_; 
wire w_mem_inst__abc_19396_new_n1631__bF_buf0; 
wire w_mem_inst__abc_19396_new_n1631__bF_buf1; 
wire w_mem_inst__abc_19396_new_n1631__bF_buf2; 
wire w_mem_inst__abc_19396_new_n1631__bF_buf3; 
wire w_mem_inst__abc_19396_new_n1631__bF_buf4; 
wire w_mem_inst__abc_19396_new_n1632_; 
wire w_mem_inst__abc_19396_new_n1633_; 
wire w_mem_inst__abc_19396_new_n1634_; 
wire w_mem_inst__abc_19396_new_n1635_; 
wire w_mem_inst__abc_19396_new_n1635__bF_buf0; 
wire w_mem_inst__abc_19396_new_n1635__bF_buf1; 
wire w_mem_inst__abc_19396_new_n1635__bF_buf2; 
wire w_mem_inst__abc_19396_new_n1635__bF_buf3; 
wire w_mem_inst__abc_19396_new_n1635__bF_buf4; 
wire w_mem_inst__abc_19396_new_n1636_; 
wire w_mem_inst__abc_19396_new_n1637_; 
wire w_mem_inst__abc_19396_new_n1637__bF_buf0; 
wire w_mem_inst__abc_19396_new_n1637__bF_buf1; 
wire w_mem_inst__abc_19396_new_n1637__bF_buf2; 
wire w_mem_inst__abc_19396_new_n1637__bF_buf3; 
wire w_mem_inst__abc_19396_new_n1637__bF_buf4; 
wire w_mem_inst__abc_19396_new_n1638_; 
wire w_mem_inst__abc_19396_new_n1638__bF_buf0; 
wire w_mem_inst__abc_19396_new_n1638__bF_buf1; 
wire w_mem_inst__abc_19396_new_n1638__bF_buf2; 
wire w_mem_inst__abc_19396_new_n1638__bF_buf3; 
wire w_mem_inst__abc_19396_new_n1638__bF_buf4; 
wire w_mem_inst__abc_19396_new_n1639_; 
wire w_mem_inst__abc_19396_new_n1640_; 
wire w_mem_inst__abc_19396_new_n1641_; 
wire w_mem_inst__abc_19396_new_n1643_; 
wire w_mem_inst__abc_19396_new_n1644_; 
wire w_mem_inst__abc_19396_new_n1645_; 
wire w_mem_inst__abc_19396_new_n1646_; 
wire w_mem_inst__abc_19396_new_n1647_; 
wire w_mem_inst__abc_19396_new_n1648_; 
wire w_mem_inst__abc_19396_new_n1649_; 
wire w_mem_inst__abc_19396_new_n1650_; 
wire w_mem_inst__abc_19396_new_n1651_; 
wire w_mem_inst__abc_19396_new_n1652_; 
wire w_mem_inst__abc_19396_new_n1653_; 
wire w_mem_inst__abc_19396_new_n1654_; 
wire w_mem_inst__abc_19396_new_n1655_; 
wire w_mem_inst__abc_19396_new_n1656_; 
wire w_mem_inst__abc_19396_new_n1657_; 
wire w_mem_inst__abc_19396_new_n1658_; 
wire w_mem_inst__abc_19396_new_n1659_; 
wire w_mem_inst__abc_19396_new_n1660_; 
wire w_mem_inst__abc_19396_new_n1661_; 
wire w_mem_inst__abc_19396_new_n1662_; 
wire w_mem_inst__abc_19396_new_n1663_; 
wire w_mem_inst__abc_19396_new_n1664_; 
wire w_mem_inst__abc_19396_new_n1665_; 
wire w_mem_inst__abc_19396_new_n1666_; 
wire w_mem_inst__abc_19396_new_n1668_; 
wire w_mem_inst__abc_19396_new_n1669_; 
wire w_mem_inst__abc_19396_new_n1670_; 
wire w_mem_inst__abc_19396_new_n1671_; 
wire w_mem_inst__abc_19396_new_n1672_; 
wire w_mem_inst__abc_19396_new_n1673_; 
wire w_mem_inst__abc_19396_new_n1674_; 
wire w_mem_inst__abc_19396_new_n1675_; 
wire w_mem_inst__abc_19396_new_n1676_; 
wire w_mem_inst__abc_19396_new_n1677_; 
wire w_mem_inst__abc_19396_new_n1678_; 
wire w_mem_inst__abc_19396_new_n1679_; 
wire w_mem_inst__abc_19396_new_n1680_; 
wire w_mem_inst__abc_19396_new_n1681_; 
wire w_mem_inst__abc_19396_new_n1682_; 
wire w_mem_inst__abc_19396_new_n1683_; 
wire w_mem_inst__abc_19396_new_n1684_; 
wire w_mem_inst__abc_19396_new_n1685_; 
wire w_mem_inst__abc_19396_new_n1686_; 
wire w_mem_inst__abc_19396_new_n1687_; 
wire w_mem_inst__abc_19396_new_n1688_; 
wire w_mem_inst__abc_19396_new_n1689_; 
wire w_mem_inst__abc_19396_new_n1690_; 
wire w_mem_inst__abc_19396_new_n1691_; 
wire w_mem_inst__abc_19396_new_n1693_; 
wire w_mem_inst__abc_19396_new_n1694_; 
wire w_mem_inst__abc_19396_new_n1695_; 
wire w_mem_inst__abc_19396_new_n1696_; 
wire w_mem_inst__abc_19396_new_n1697_; 
wire w_mem_inst__abc_19396_new_n1698_; 
wire w_mem_inst__abc_19396_new_n1699_; 
wire w_mem_inst__abc_19396_new_n1700_; 
wire w_mem_inst__abc_19396_new_n1701_; 
wire w_mem_inst__abc_19396_new_n1702_; 
wire w_mem_inst__abc_19396_new_n1703_; 
wire w_mem_inst__abc_19396_new_n1704_; 
wire w_mem_inst__abc_19396_new_n1705_; 
wire w_mem_inst__abc_19396_new_n1706_; 
wire w_mem_inst__abc_19396_new_n1707_; 
wire w_mem_inst__abc_19396_new_n1708_; 
wire w_mem_inst__abc_19396_new_n1709_; 
wire w_mem_inst__abc_19396_new_n1710_; 
wire w_mem_inst__abc_19396_new_n1711_; 
wire w_mem_inst__abc_19396_new_n1712_; 
wire w_mem_inst__abc_19396_new_n1713_; 
wire w_mem_inst__abc_19396_new_n1714_; 
wire w_mem_inst__abc_19396_new_n1715_; 
wire w_mem_inst__abc_19396_new_n1716_; 
wire w_mem_inst__abc_19396_new_n1718_; 
wire w_mem_inst__abc_19396_new_n1719_; 
wire w_mem_inst__abc_19396_new_n1720_; 
wire w_mem_inst__abc_19396_new_n1721_; 
wire w_mem_inst__abc_19396_new_n1722_; 
wire w_mem_inst__abc_19396_new_n1723_; 
wire w_mem_inst__abc_19396_new_n1724_; 
wire w_mem_inst__abc_19396_new_n1725_; 
wire w_mem_inst__abc_19396_new_n1726_; 
wire w_mem_inst__abc_19396_new_n1727_; 
wire w_mem_inst__abc_19396_new_n1728_; 
wire w_mem_inst__abc_19396_new_n1729_; 
wire w_mem_inst__abc_19396_new_n1730_; 
wire w_mem_inst__abc_19396_new_n1731_; 
wire w_mem_inst__abc_19396_new_n1732_; 
wire w_mem_inst__abc_19396_new_n1733_; 
wire w_mem_inst__abc_19396_new_n1734_; 
wire w_mem_inst__abc_19396_new_n1735_; 
wire w_mem_inst__abc_19396_new_n1736_; 
wire w_mem_inst__abc_19396_new_n1737_; 
wire w_mem_inst__abc_19396_new_n1738_; 
wire w_mem_inst__abc_19396_new_n1739_; 
wire w_mem_inst__abc_19396_new_n1740_; 
wire w_mem_inst__abc_19396_new_n1741_; 
wire w_mem_inst__abc_19396_new_n1743_; 
wire w_mem_inst__abc_19396_new_n1744_; 
wire w_mem_inst__abc_19396_new_n1745_; 
wire w_mem_inst__abc_19396_new_n1746_; 
wire w_mem_inst__abc_19396_new_n1747_; 
wire w_mem_inst__abc_19396_new_n1748_; 
wire w_mem_inst__abc_19396_new_n1749_; 
wire w_mem_inst__abc_19396_new_n1750_; 
wire w_mem_inst__abc_19396_new_n1751_; 
wire w_mem_inst__abc_19396_new_n1752_; 
wire w_mem_inst__abc_19396_new_n1753_; 
wire w_mem_inst__abc_19396_new_n1754_; 
wire w_mem_inst__abc_19396_new_n1755_; 
wire w_mem_inst__abc_19396_new_n1756_; 
wire w_mem_inst__abc_19396_new_n1757_; 
wire w_mem_inst__abc_19396_new_n1758_; 
wire w_mem_inst__abc_19396_new_n1759_; 
wire w_mem_inst__abc_19396_new_n1760_; 
wire w_mem_inst__abc_19396_new_n1761_; 
wire w_mem_inst__abc_19396_new_n1762_; 
wire w_mem_inst__abc_19396_new_n1763_; 
wire w_mem_inst__abc_19396_new_n1764_; 
wire w_mem_inst__abc_19396_new_n1765_; 
wire w_mem_inst__abc_19396_new_n1766_; 
wire w_mem_inst__abc_19396_new_n1768_; 
wire w_mem_inst__abc_19396_new_n1769_; 
wire w_mem_inst__abc_19396_new_n1770_; 
wire w_mem_inst__abc_19396_new_n1771_; 
wire w_mem_inst__abc_19396_new_n1772_; 
wire w_mem_inst__abc_19396_new_n1773_; 
wire w_mem_inst__abc_19396_new_n1774_; 
wire w_mem_inst__abc_19396_new_n1775_; 
wire w_mem_inst__abc_19396_new_n1776_; 
wire w_mem_inst__abc_19396_new_n1777_; 
wire w_mem_inst__abc_19396_new_n1778_; 
wire w_mem_inst__abc_19396_new_n1779_; 
wire w_mem_inst__abc_19396_new_n1780_; 
wire w_mem_inst__abc_19396_new_n1781_; 
wire w_mem_inst__abc_19396_new_n1782_; 
wire w_mem_inst__abc_19396_new_n1783_; 
wire w_mem_inst__abc_19396_new_n1784_; 
wire w_mem_inst__abc_19396_new_n1785_; 
wire w_mem_inst__abc_19396_new_n1786_; 
wire w_mem_inst__abc_19396_new_n1787_; 
wire w_mem_inst__abc_19396_new_n1788_; 
wire w_mem_inst__abc_19396_new_n1789_; 
wire w_mem_inst__abc_19396_new_n1790_; 
wire w_mem_inst__abc_19396_new_n1791_; 
wire w_mem_inst__abc_19396_new_n1793_; 
wire w_mem_inst__abc_19396_new_n1794_; 
wire w_mem_inst__abc_19396_new_n1795_; 
wire w_mem_inst__abc_19396_new_n1796_; 
wire w_mem_inst__abc_19396_new_n1797_; 
wire w_mem_inst__abc_19396_new_n1798_; 
wire w_mem_inst__abc_19396_new_n1799_; 
wire w_mem_inst__abc_19396_new_n1800_; 
wire w_mem_inst__abc_19396_new_n1801_; 
wire w_mem_inst__abc_19396_new_n1802_; 
wire w_mem_inst__abc_19396_new_n1803_; 
wire w_mem_inst__abc_19396_new_n1804_; 
wire w_mem_inst__abc_19396_new_n1805_; 
wire w_mem_inst__abc_19396_new_n1806_; 
wire w_mem_inst__abc_19396_new_n1807_; 
wire w_mem_inst__abc_19396_new_n1808_; 
wire w_mem_inst__abc_19396_new_n1809_; 
wire w_mem_inst__abc_19396_new_n1810_; 
wire w_mem_inst__abc_19396_new_n1811_; 
wire w_mem_inst__abc_19396_new_n1812_; 
wire w_mem_inst__abc_19396_new_n1813_; 
wire w_mem_inst__abc_19396_new_n1814_; 
wire w_mem_inst__abc_19396_new_n1815_; 
wire w_mem_inst__abc_19396_new_n1816_; 
wire w_mem_inst__abc_19396_new_n1818_; 
wire w_mem_inst__abc_19396_new_n1819_; 
wire w_mem_inst__abc_19396_new_n1820_; 
wire w_mem_inst__abc_19396_new_n1821_; 
wire w_mem_inst__abc_19396_new_n1822_; 
wire w_mem_inst__abc_19396_new_n1823_; 
wire w_mem_inst__abc_19396_new_n1824_; 
wire w_mem_inst__abc_19396_new_n1825_; 
wire w_mem_inst__abc_19396_new_n1826_; 
wire w_mem_inst__abc_19396_new_n1827_; 
wire w_mem_inst__abc_19396_new_n1828_; 
wire w_mem_inst__abc_19396_new_n1829_; 
wire w_mem_inst__abc_19396_new_n1830_; 
wire w_mem_inst__abc_19396_new_n1831_; 
wire w_mem_inst__abc_19396_new_n1832_; 
wire w_mem_inst__abc_19396_new_n1833_; 
wire w_mem_inst__abc_19396_new_n1834_; 
wire w_mem_inst__abc_19396_new_n1835_; 
wire w_mem_inst__abc_19396_new_n1836_; 
wire w_mem_inst__abc_19396_new_n1837_; 
wire w_mem_inst__abc_19396_new_n1838_; 
wire w_mem_inst__abc_19396_new_n1839_; 
wire w_mem_inst__abc_19396_new_n1840_; 
wire w_mem_inst__abc_19396_new_n1841_; 
wire w_mem_inst__abc_19396_new_n1843_; 
wire w_mem_inst__abc_19396_new_n1844_; 
wire w_mem_inst__abc_19396_new_n1845_; 
wire w_mem_inst__abc_19396_new_n1846_; 
wire w_mem_inst__abc_19396_new_n1847_; 
wire w_mem_inst__abc_19396_new_n1848_; 
wire w_mem_inst__abc_19396_new_n1849_; 
wire w_mem_inst__abc_19396_new_n1850_; 
wire w_mem_inst__abc_19396_new_n1851_; 
wire w_mem_inst__abc_19396_new_n1852_; 
wire w_mem_inst__abc_19396_new_n1853_; 
wire w_mem_inst__abc_19396_new_n1854_; 
wire w_mem_inst__abc_19396_new_n1855_; 
wire w_mem_inst__abc_19396_new_n1856_; 
wire w_mem_inst__abc_19396_new_n1857_; 
wire w_mem_inst__abc_19396_new_n1858_; 
wire w_mem_inst__abc_19396_new_n1859_; 
wire w_mem_inst__abc_19396_new_n1860_; 
wire w_mem_inst__abc_19396_new_n1861_; 
wire w_mem_inst__abc_19396_new_n1862_; 
wire w_mem_inst__abc_19396_new_n1863_; 
wire w_mem_inst__abc_19396_new_n1864_; 
wire w_mem_inst__abc_19396_new_n1865_; 
wire w_mem_inst__abc_19396_new_n1866_; 
wire w_mem_inst__abc_19396_new_n1868_; 
wire w_mem_inst__abc_19396_new_n1869_; 
wire w_mem_inst__abc_19396_new_n1870_; 
wire w_mem_inst__abc_19396_new_n1871_; 
wire w_mem_inst__abc_19396_new_n1872_; 
wire w_mem_inst__abc_19396_new_n1873_; 
wire w_mem_inst__abc_19396_new_n1874_; 
wire w_mem_inst__abc_19396_new_n1875_; 
wire w_mem_inst__abc_19396_new_n1876_; 
wire w_mem_inst__abc_19396_new_n1877_; 
wire w_mem_inst__abc_19396_new_n1878_; 
wire w_mem_inst__abc_19396_new_n1879_; 
wire w_mem_inst__abc_19396_new_n1880_; 
wire w_mem_inst__abc_19396_new_n1881_; 
wire w_mem_inst__abc_19396_new_n1882_; 
wire w_mem_inst__abc_19396_new_n1883_; 
wire w_mem_inst__abc_19396_new_n1884_; 
wire w_mem_inst__abc_19396_new_n1885_; 
wire w_mem_inst__abc_19396_new_n1886_; 
wire w_mem_inst__abc_19396_new_n1887_; 
wire w_mem_inst__abc_19396_new_n1888_; 
wire w_mem_inst__abc_19396_new_n1889_; 
wire w_mem_inst__abc_19396_new_n1890_; 
wire w_mem_inst__abc_19396_new_n1891_; 
wire w_mem_inst__abc_19396_new_n1893_; 
wire w_mem_inst__abc_19396_new_n1894_; 
wire w_mem_inst__abc_19396_new_n1895_; 
wire w_mem_inst__abc_19396_new_n1896_; 
wire w_mem_inst__abc_19396_new_n1897_; 
wire w_mem_inst__abc_19396_new_n1898_; 
wire w_mem_inst__abc_19396_new_n1899_; 
wire w_mem_inst__abc_19396_new_n1900_; 
wire w_mem_inst__abc_19396_new_n1901_; 
wire w_mem_inst__abc_19396_new_n1902_; 
wire w_mem_inst__abc_19396_new_n1903_; 
wire w_mem_inst__abc_19396_new_n1904_; 
wire w_mem_inst__abc_19396_new_n1905_; 
wire w_mem_inst__abc_19396_new_n1906_; 
wire w_mem_inst__abc_19396_new_n1907_; 
wire w_mem_inst__abc_19396_new_n1908_; 
wire w_mem_inst__abc_19396_new_n1909_; 
wire w_mem_inst__abc_19396_new_n1910_; 
wire w_mem_inst__abc_19396_new_n1911_; 
wire w_mem_inst__abc_19396_new_n1912_; 
wire w_mem_inst__abc_19396_new_n1913_; 
wire w_mem_inst__abc_19396_new_n1914_; 
wire w_mem_inst__abc_19396_new_n1915_; 
wire w_mem_inst__abc_19396_new_n1916_; 
wire w_mem_inst__abc_19396_new_n1918_; 
wire w_mem_inst__abc_19396_new_n1919_; 
wire w_mem_inst__abc_19396_new_n1920_; 
wire w_mem_inst__abc_19396_new_n1921_; 
wire w_mem_inst__abc_19396_new_n1922_; 
wire w_mem_inst__abc_19396_new_n1923_; 
wire w_mem_inst__abc_19396_new_n1924_; 
wire w_mem_inst__abc_19396_new_n1925_; 
wire w_mem_inst__abc_19396_new_n1926_; 
wire w_mem_inst__abc_19396_new_n1927_; 
wire w_mem_inst__abc_19396_new_n1928_; 
wire w_mem_inst__abc_19396_new_n1929_; 
wire w_mem_inst__abc_19396_new_n1930_; 
wire w_mem_inst__abc_19396_new_n1931_; 
wire w_mem_inst__abc_19396_new_n1932_; 
wire w_mem_inst__abc_19396_new_n1933_; 
wire w_mem_inst__abc_19396_new_n1934_; 
wire w_mem_inst__abc_19396_new_n1935_; 
wire w_mem_inst__abc_19396_new_n1936_; 
wire w_mem_inst__abc_19396_new_n1937_; 
wire w_mem_inst__abc_19396_new_n1938_; 
wire w_mem_inst__abc_19396_new_n1939_; 
wire w_mem_inst__abc_19396_new_n1940_; 
wire w_mem_inst__abc_19396_new_n1941_; 
wire w_mem_inst__abc_19396_new_n1943_; 
wire w_mem_inst__abc_19396_new_n1944_; 
wire w_mem_inst__abc_19396_new_n1945_; 
wire w_mem_inst__abc_19396_new_n1946_; 
wire w_mem_inst__abc_19396_new_n1947_; 
wire w_mem_inst__abc_19396_new_n1948_; 
wire w_mem_inst__abc_19396_new_n1949_; 
wire w_mem_inst__abc_19396_new_n1950_; 
wire w_mem_inst__abc_19396_new_n1951_; 
wire w_mem_inst__abc_19396_new_n1952_; 
wire w_mem_inst__abc_19396_new_n1953_; 
wire w_mem_inst__abc_19396_new_n1954_; 
wire w_mem_inst__abc_19396_new_n1955_; 
wire w_mem_inst__abc_19396_new_n1956_; 
wire w_mem_inst__abc_19396_new_n1957_; 
wire w_mem_inst__abc_19396_new_n1958_; 
wire w_mem_inst__abc_19396_new_n1959_; 
wire w_mem_inst__abc_19396_new_n1960_; 
wire w_mem_inst__abc_19396_new_n1961_; 
wire w_mem_inst__abc_19396_new_n1962_; 
wire w_mem_inst__abc_19396_new_n1963_; 
wire w_mem_inst__abc_19396_new_n1964_; 
wire w_mem_inst__abc_19396_new_n1965_; 
wire w_mem_inst__abc_19396_new_n1966_; 
wire w_mem_inst__abc_19396_new_n1968_; 
wire w_mem_inst__abc_19396_new_n1969_; 
wire w_mem_inst__abc_19396_new_n1970_; 
wire w_mem_inst__abc_19396_new_n1971_; 
wire w_mem_inst__abc_19396_new_n1972_; 
wire w_mem_inst__abc_19396_new_n1973_; 
wire w_mem_inst__abc_19396_new_n1974_; 
wire w_mem_inst__abc_19396_new_n1975_; 
wire w_mem_inst__abc_19396_new_n1976_; 
wire w_mem_inst__abc_19396_new_n1977_; 
wire w_mem_inst__abc_19396_new_n1978_; 
wire w_mem_inst__abc_19396_new_n1979_; 
wire w_mem_inst__abc_19396_new_n1980_; 
wire w_mem_inst__abc_19396_new_n1981_; 
wire w_mem_inst__abc_19396_new_n1982_; 
wire w_mem_inst__abc_19396_new_n1983_; 
wire w_mem_inst__abc_19396_new_n1984_; 
wire w_mem_inst__abc_19396_new_n1985_; 
wire w_mem_inst__abc_19396_new_n1986_; 
wire w_mem_inst__abc_19396_new_n1987_; 
wire w_mem_inst__abc_19396_new_n1988_; 
wire w_mem_inst__abc_19396_new_n1989_; 
wire w_mem_inst__abc_19396_new_n1990_; 
wire w_mem_inst__abc_19396_new_n1991_; 
wire w_mem_inst__abc_19396_new_n1993_; 
wire w_mem_inst__abc_19396_new_n1994_; 
wire w_mem_inst__abc_19396_new_n1995_; 
wire w_mem_inst__abc_19396_new_n1996_; 
wire w_mem_inst__abc_19396_new_n1997_; 
wire w_mem_inst__abc_19396_new_n1998_; 
wire w_mem_inst__abc_19396_new_n1999_; 
wire w_mem_inst__abc_19396_new_n2000_; 
wire w_mem_inst__abc_19396_new_n2001_; 
wire w_mem_inst__abc_19396_new_n2002_; 
wire w_mem_inst__abc_19396_new_n2003_; 
wire w_mem_inst__abc_19396_new_n2004_; 
wire w_mem_inst__abc_19396_new_n2005_; 
wire w_mem_inst__abc_19396_new_n2006_; 
wire w_mem_inst__abc_19396_new_n2007_; 
wire w_mem_inst__abc_19396_new_n2008_; 
wire w_mem_inst__abc_19396_new_n2009_; 
wire w_mem_inst__abc_19396_new_n2010_; 
wire w_mem_inst__abc_19396_new_n2011_; 
wire w_mem_inst__abc_19396_new_n2012_; 
wire w_mem_inst__abc_19396_new_n2013_; 
wire w_mem_inst__abc_19396_new_n2014_; 
wire w_mem_inst__abc_19396_new_n2015_; 
wire w_mem_inst__abc_19396_new_n2016_; 
wire w_mem_inst__abc_19396_new_n2018_; 
wire w_mem_inst__abc_19396_new_n2019_; 
wire w_mem_inst__abc_19396_new_n2020_; 
wire w_mem_inst__abc_19396_new_n2021_; 
wire w_mem_inst__abc_19396_new_n2022_; 
wire w_mem_inst__abc_19396_new_n2023_; 
wire w_mem_inst__abc_19396_new_n2024_; 
wire w_mem_inst__abc_19396_new_n2025_; 
wire w_mem_inst__abc_19396_new_n2026_; 
wire w_mem_inst__abc_19396_new_n2027_; 
wire w_mem_inst__abc_19396_new_n2028_; 
wire w_mem_inst__abc_19396_new_n2029_; 
wire w_mem_inst__abc_19396_new_n2030_; 
wire w_mem_inst__abc_19396_new_n2031_; 
wire w_mem_inst__abc_19396_new_n2032_; 
wire w_mem_inst__abc_19396_new_n2033_; 
wire w_mem_inst__abc_19396_new_n2034_; 
wire w_mem_inst__abc_19396_new_n2035_; 
wire w_mem_inst__abc_19396_new_n2036_; 
wire w_mem_inst__abc_19396_new_n2037_; 
wire w_mem_inst__abc_19396_new_n2038_; 
wire w_mem_inst__abc_19396_new_n2039_; 
wire w_mem_inst__abc_19396_new_n2040_; 
wire w_mem_inst__abc_19396_new_n2041_; 
wire w_mem_inst__abc_19396_new_n2043_; 
wire w_mem_inst__abc_19396_new_n2044_; 
wire w_mem_inst__abc_19396_new_n2045_; 
wire w_mem_inst__abc_19396_new_n2046_; 
wire w_mem_inst__abc_19396_new_n2047_; 
wire w_mem_inst__abc_19396_new_n2048_; 
wire w_mem_inst__abc_19396_new_n2049_; 
wire w_mem_inst__abc_19396_new_n2050_; 
wire w_mem_inst__abc_19396_new_n2051_; 
wire w_mem_inst__abc_19396_new_n2052_; 
wire w_mem_inst__abc_19396_new_n2053_; 
wire w_mem_inst__abc_19396_new_n2054_; 
wire w_mem_inst__abc_19396_new_n2055_; 
wire w_mem_inst__abc_19396_new_n2056_; 
wire w_mem_inst__abc_19396_new_n2057_; 
wire w_mem_inst__abc_19396_new_n2058_; 
wire w_mem_inst__abc_19396_new_n2059_; 
wire w_mem_inst__abc_19396_new_n2060_; 
wire w_mem_inst__abc_19396_new_n2061_; 
wire w_mem_inst__abc_19396_new_n2062_; 
wire w_mem_inst__abc_19396_new_n2063_; 
wire w_mem_inst__abc_19396_new_n2064_; 
wire w_mem_inst__abc_19396_new_n2065_; 
wire w_mem_inst__abc_19396_new_n2066_; 
wire w_mem_inst__abc_19396_new_n2068_; 
wire w_mem_inst__abc_19396_new_n2069_; 
wire w_mem_inst__abc_19396_new_n2070_; 
wire w_mem_inst__abc_19396_new_n2071_; 
wire w_mem_inst__abc_19396_new_n2072_; 
wire w_mem_inst__abc_19396_new_n2073_; 
wire w_mem_inst__abc_19396_new_n2074_; 
wire w_mem_inst__abc_19396_new_n2075_; 
wire w_mem_inst__abc_19396_new_n2076_; 
wire w_mem_inst__abc_19396_new_n2077_; 
wire w_mem_inst__abc_19396_new_n2078_; 
wire w_mem_inst__abc_19396_new_n2079_; 
wire w_mem_inst__abc_19396_new_n2080_; 
wire w_mem_inst__abc_19396_new_n2081_; 
wire w_mem_inst__abc_19396_new_n2082_; 
wire w_mem_inst__abc_19396_new_n2083_; 
wire w_mem_inst__abc_19396_new_n2084_; 
wire w_mem_inst__abc_19396_new_n2085_; 
wire w_mem_inst__abc_19396_new_n2086_; 
wire w_mem_inst__abc_19396_new_n2087_; 
wire w_mem_inst__abc_19396_new_n2088_; 
wire w_mem_inst__abc_19396_new_n2089_; 
wire w_mem_inst__abc_19396_new_n2090_; 
wire w_mem_inst__abc_19396_new_n2091_; 
wire w_mem_inst__abc_19396_new_n2093_; 
wire w_mem_inst__abc_19396_new_n2094_; 
wire w_mem_inst__abc_19396_new_n2095_; 
wire w_mem_inst__abc_19396_new_n2096_; 
wire w_mem_inst__abc_19396_new_n2097_; 
wire w_mem_inst__abc_19396_new_n2098_; 
wire w_mem_inst__abc_19396_new_n2099_; 
wire w_mem_inst__abc_19396_new_n2100_; 
wire w_mem_inst__abc_19396_new_n2101_; 
wire w_mem_inst__abc_19396_new_n2102_; 
wire w_mem_inst__abc_19396_new_n2103_; 
wire w_mem_inst__abc_19396_new_n2104_; 
wire w_mem_inst__abc_19396_new_n2105_; 
wire w_mem_inst__abc_19396_new_n2106_; 
wire w_mem_inst__abc_19396_new_n2107_; 
wire w_mem_inst__abc_19396_new_n2108_; 
wire w_mem_inst__abc_19396_new_n2109_; 
wire w_mem_inst__abc_19396_new_n2110_; 
wire w_mem_inst__abc_19396_new_n2111_; 
wire w_mem_inst__abc_19396_new_n2112_; 
wire w_mem_inst__abc_19396_new_n2113_; 
wire w_mem_inst__abc_19396_new_n2114_; 
wire w_mem_inst__abc_19396_new_n2115_; 
wire w_mem_inst__abc_19396_new_n2116_; 
wire w_mem_inst__abc_19396_new_n2118_; 
wire w_mem_inst__abc_19396_new_n2119_; 
wire w_mem_inst__abc_19396_new_n2120_; 
wire w_mem_inst__abc_19396_new_n2121_; 
wire w_mem_inst__abc_19396_new_n2122_; 
wire w_mem_inst__abc_19396_new_n2123_; 
wire w_mem_inst__abc_19396_new_n2124_; 
wire w_mem_inst__abc_19396_new_n2125_; 
wire w_mem_inst__abc_19396_new_n2126_; 
wire w_mem_inst__abc_19396_new_n2127_; 
wire w_mem_inst__abc_19396_new_n2128_; 
wire w_mem_inst__abc_19396_new_n2129_; 
wire w_mem_inst__abc_19396_new_n2130_; 
wire w_mem_inst__abc_19396_new_n2131_; 
wire w_mem_inst__abc_19396_new_n2132_; 
wire w_mem_inst__abc_19396_new_n2133_; 
wire w_mem_inst__abc_19396_new_n2134_; 
wire w_mem_inst__abc_19396_new_n2135_; 
wire w_mem_inst__abc_19396_new_n2136_; 
wire w_mem_inst__abc_19396_new_n2137_; 
wire w_mem_inst__abc_19396_new_n2138_; 
wire w_mem_inst__abc_19396_new_n2139_; 
wire w_mem_inst__abc_19396_new_n2140_; 
wire w_mem_inst__abc_19396_new_n2141_; 
wire w_mem_inst__abc_19396_new_n2143_; 
wire w_mem_inst__abc_19396_new_n2144_; 
wire w_mem_inst__abc_19396_new_n2145_; 
wire w_mem_inst__abc_19396_new_n2146_; 
wire w_mem_inst__abc_19396_new_n2147_; 
wire w_mem_inst__abc_19396_new_n2148_; 
wire w_mem_inst__abc_19396_new_n2149_; 
wire w_mem_inst__abc_19396_new_n2150_; 
wire w_mem_inst__abc_19396_new_n2151_; 
wire w_mem_inst__abc_19396_new_n2152_; 
wire w_mem_inst__abc_19396_new_n2153_; 
wire w_mem_inst__abc_19396_new_n2154_; 
wire w_mem_inst__abc_19396_new_n2155_; 
wire w_mem_inst__abc_19396_new_n2156_; 
wire w_mem_inst__abc_19396_new_n2157_; 
wire w_mem_inst__abc_19396_new_n2158_; 
wire w_mem_inst__abc_19396_new_n2159_; 
wire w_mem_inst__abc_19396_new_n2160_; 
wire w_mem_inst__abc_19396_new_n2161_; 
wire w_mem_inst__abc_19396_new_n2162_; 
wire w_mem_inst__abc_19396_new_n2163_; 
wire w_mem_inst__abc_19396_new_n2164_; 
wire w_mem_inst__abc_19396_new_n2165_; 
wire w_mem_inst__abc_19396_new_n2166_; 
wire w_mem_inst__abc_19396_new_n2168_; 
wire w_mem_inst__abc_19396_new_n2169_; 
wire w_mem_inst__abc_19396_new_n2170_; 
wire w_mem_inst__abc_19396_new_n2171_; 
wire w_mem_inst__abc_19396_new_n2172_; 
wire w_mem_inst__abc_19396_new_n2173_; 
wire w_mem_inst__abc_19396_new_n2174_; 
wire w_mem_inst__abc_19396_new_n2175_; 
wire w_mem_inst__abc_19396_new_n2176_; 
wire w_mem_inst__abc_19396_new_n2177_; 
wire w_mem_inst__abc_19396_new_n2178_; 
wire w_mem_inst__abc_19396_new_n2179_; 
wire w_mem_inst__abc_19396_new_n2180_; 
wire w_mem_inst__abc_19396_new_n2181_; 
wire w_mem_inst__abc_19396_new_n2182_; 
wire w_mem_inst__abc_19396_new_n2183_; 
wire w_mem_inst__abc_19396_new_n2184_; 
wire w_mem_inst__abc_19396_new_n2185_; 
wire w_mem_inst__abc_19396_new_n2186_; 
wire w_mem_inst__abc_19396_new_n2187_; 
wire w_mem_inst__abc_19396_new_n2188_; 
wire w_mem_inst__abc_19396_new_n2189_; 
wire w_mem_inst__abc_19396_new_n2190_; 
wire w_mem_inst__abc_19396_new_n2191_; 
wire w_mem_inst__abc_19396_new_n2193_; 
wire w_mem_inst__abc_19396_new_n2194_; 
wire w_mem_inst__abc_19396_new_n2195_; 
wire w_mem_inst__abc_19396_new_n2196_; 
wire w_mem_inst__abc_19396_new_n2197_; 
wire w_mem_inst__abc_19396_new_n2198_; 
wire w_mem_inst__abc_19396_new_n2199_; 
wire w_mem_inst__abc_19396_new_n2200_; 
wire w_mem_inst__abc_19396_new_n2201_; 
wire w_mem_inst__abc_19396_new_n2202_; 
wire w_mem_inst__abc_19396_new_n2203_; 
wire w_mem_inst__abc_19396_new_n2204_; 
wire w_mem_inst__abc_19396_new_n2205_; 
wire w_mem_inst__abc_19396_new_n2206_; 
wire w_mem_inst__abc_19396_new_n2207_; 
wire w_mem_inst__abc_19396_new_n2208_; 
wire w_mem_inst__abc_19396_new_n2209_; 
wire w_mem_inst__abc_19396_new_n2210_; 
wire w_mem_inst__abc_19396_new_n2211_; 
wire w_mem_inst__abc_19396_new_n2212_; 
wire w_mem_inst__abc_19396_new_n2213_; 
wire w_mem_inst__abc_19396_new_n2214_; 
wire w_mem_inst__abc_19396_new_n2215_; 
wire w_mem_inst__abc_19396_new_n2216_; 
wire w_mem_inst__abc_19396_new_n2218_; 
wire w_mem_inst__abc_19396_new_n2219_; 
wire w_mem_inst__abc_19396_new_n2220_; 
wire w_mem_inst__abc_19396_new_n2221_; 
wire w_mem_inst__abc_19396_new_n2222_; 
wire w_mem_inst__abc_19396_new_n2223_; 
wire w_mem_inst__abc_19396_new_n2224_; 
wire w_mem_inst__abc_19396_new_n2225_; 
wire w_mem_inst__abc_19396_new_n2226_; 
wire w_mem_inst__abc_19396_new_n2227_; 
wire w_mem_inst__abc_19396_new_n2228_; 
wire w_mem_inst__abc_19396_new_n2229_; 
wire w_mem_inst__abc_19396_new_n2230_; 
wire w_mem_inst__abc_19396_new_n2231_; 
wire w_mem_inst__abc_19396_new_n2232_; 
wire w_mem_inst__abc_19396_new_n2233_; 
wire w_mem_inst__abc_19396_new_n2234_; 
wire w_mem_inst__abc_19396_new_n2235_; 
wire w_mem_inst__abc_19396_new_n2236_; 
wire w_mem_inst__abc_19396_new_n2237_; 
wire w_mem_inst__abc_19396_new_n2238_; 
wire w_mem_inst__abc_19396_new_n2239_; 
wire w_mem_inst__abc_19396_new_n2240_; 
wire w_mem_inst__abc_19396_new_n2241_; 
wire w_mem_inst__abc_19396_new_n2243_; 
wire w_mem_inst__abc_19396_new_n2244_; 
wire w_mem_inst__abc_19396_new_n2245_; 
wire w_mem_inst__abc_19396_new_n2246_; 
wire w_mem_inst__abc_19396_new_n2247_; 
wire w_mem_inst__abc_19396_new_n2248_; 
wire w_mem_inst__abc_19396_new_n2249_; 
wire w_mem_inst__abc_19396_new_n2250_; 
wire w_mem_inst__abc_19396_new_n2251_; 
wire w_mem_inst__abc_19396_new_n2252_; 
wire w_mem_inst__abc_19396_new_n2253_; 
wire w_mem_inst__abc_19396_new_n2254_; 
wire w_mem_inst__abc_19396_new_n2255_; 
wire w_mem_inst__abc_19396_new_n2256_; 
wire w_mem_inst__abc_19396_new_n2257_; 
wire w_mem_inst__abc_19396_new_n2258_; 
wire w_mem_inst__abc_19396_new_n2259_; 
wire w_mem_inst__abc_19396_new_n2260_; 
wire w_mem_inst__abc_19396_new_n2261_; 
wire w_mem_inst__abc_19396_new_n2262_; 
wire w_mem_inst__abc_19396_new_n2263_; 
wire w_mem_inst__abc_19396_new_n2264_; 
wire w_mem_inst__abc_19396_new_n2265_; 
wire w_mem_inst__abc_19396_new_n2266_; 
wire w_mem_inst__abc_19396_new_n2268_; 
wire w_mem_inst__abc_19396_new_n2269_; 
wire w_mem_inst__abc_19396_new_n2270_; 
wire w_mem_inst__abc_19396_new_n2271_; 
wire w_mem_inst__abc_19396_new_n2272_; 
wire w_mem_inst__abc_19396_new_n2273_; 
wire w_mem_inst__abc_19396_new_n2274_; 
wire w_mem_inst__abc_19396_new_n2275_; 
wire w_mem_inst__abc_19396_new_n2276_; 
wire w_mem_inst__abc_19396_new_n2277_; 
wire w_mem_inst__abc_19396_new_n2278_; 
wire w_mem_inst__abc_19396_new_n2279_; 
wire w_mem_inst__abc_19396_new_n2280_; 
wire w_mem_inst__abc_19396_new_n2281_; 
wire w_mem_inst__abc_19396_new_n2282_; 
wire w_mem_inst__abc_19396_new_n2283_; 
wire w_mem_inst__abc_19396_new_n2284_; 
wire w_mem_inst__abc_19396_new_n2285_; 
wire w_mem_inst__abc_19396_new_n2286_; 
wire w_mem_inst__abc_19396_new_n2287_; 
wire w_mem_inst__abc_19396_new_n2288_; 
wire w_mem_inst__abc_19396_new_n2289_; 
wire w_mem_inst__abc_19396_new_n2290_; 
wire w_mem_inst__abc_19396_new_n2291_; 
wire w_mem_inst__abc_19396_new_n2293_; 
wire w_mem_inst__abc_19396_new_n2294_; 
wire w_mem_inst__abc_19396_new_n2295_; 
wire w_mem_inst__abc_19396_new_n2296_; 
wire w_mem_inst__abc_19396_new_n2297_; 
wire w_mem_inst__abc_19396_new_n2298_; 
wire w_mem_inst__abc_19396_new_n2299_; 
wire w_mem_inst__abc_19396_new_n2300_; 
wire w_mem_inst__abc_19396_new_n2301_; 
wire w_mem_inst__abc_19396_new_n2302_; 
wire w_mem_inst__abc_19396_new_n2303_; 
wire w_mem_inst__abc_19396_new_n2304_; 
wire w_mem_inst__abc_19396_new_n2305_; 
wire w_mem_inst__abc_19396_new_n2306_; 
wire w_mem_inst__abc_19396_new_n2307_; 
wire w_mem_inst__abc_19396_new_n2308_; 
wire w_mem_inst__abc_19396_new_n2309_; 
wire w_mem_inst__abc_19396_new_n2310_; 
wire w_mem_inst__abc_19396_new_n2311_; 
wire w_mem_inst__abc_19396_new_n2312_; 
wire w_mem_inst__abc_19396_new_n2313_; 
wire w_mem_inst__abc_19396_new_n2314_; 
wire w_mem_inst__abc_19396_new_n2315_; 
wire w_mem_inst__abc_19396_new_n2316_; 
wire w_mem_inst__abc_19396_new_n2318_; 
wire w_mem_inst__abc_19396_new_n2319_; 
wire w_mem_inst__abc_19396_new_n2320_; 
wire w_mem_inst__abc_19396_new_n2321_; 
wire w_mem_inst__abc_19396_new_n2322_; 
wire w_mem_inst__abc_19396_new_n2323_; 
wire w_mem_inst__abc_19396_new_n2324_; 
wire w_mem_inst__abc_19396_new_n2325_; 
wire w_mem_inst__abc_19396_new_n2326_; 
wire w_mem_inst__abc_19396_new_n2327_; 
wire w_mem_inst__abc_19396_new_n2328_; 
wire w_mem_inst__abc_19396_new_n2329_; 
wire w_mem_inst__abc_19396_new_n2330_; 
wire w_mem_inst__abc_19396_new_n2331_; 
wire w_mem_inst__abc_19396_new_n2332_; 
wire w_mem_inst__abc_19396_new_n2333_; 
wire w_mem_inst__abc_19396_new_n2334_; 
wire w_mem_inst__abc_19396_new_n2335_; 
wire w_mem_inst__abc_19396_new_n2336_; 
wire w_mem_inst__abc_19396_new_n2337_; 
wire w_mem_inst__abc_19396_new_n2338_; 
wire w_mem_inst__abc_19396_new_n2339_; 
wire w_mem_inst__abc_19396_new_n2340_; 
wire w_mem_inst__abc_19396_new_n2341_; 
wire w_mem_inst__abc_19396_new_n2343_; 
wire w_mem_inst__abc_19396_new_n2344_; 
wire w_mem_inst__abc_19396_new_n2345_; 
wire w_mem_inst__abc_19396_new_n2346_; 
wire w_mem_inst__abc_19396_new_n2347_; 
wire w_mem_inst__abc_19396_new_n2348_; 
wire w_mem_inst__abc_19396_new_n2349_; 
wire w_mem_inst__abc_19396_new_n2350_; 
wire w_mem_inst__abc_19396_new_n2351_; 
wire w_mem_inst__abc_19396_new_n2352_; 
wire w_mem_inst__abc_19396_new_n2353_; 
wire w_mem_inst__abc_19396_new_n2354_; 
wire w_mem_inst__abc_19396_new_n2355_; 
wire w_mem_inst__abc_19396_new_n2356_; 
wire w_mem_inst__abc_19396_new_n2357_; 
wire w_mem_inst__abc_19396_new_n2358_; 
wire w_mem_inst__abc_19396_new_n2359_; 
wire w_mem_inst__abc_19396_new_n2360_; 
wire w_mem_inst__abc_19396_new_n2361_; 
wire w_mem_inst__abc_19396_new_n2362_; 
wire w_mem_inst__abc_19396_new_n2363_; 
wire w_mem_inst__abc_19396_new_n2364_; 
wire w_mem_inst__abc_19396_new_n2365_; 
wire w_mem_inst__abc_19396_new_n2366_; 
wire w_mem_inst__abc_19396_new_n2368_; 
wire w_mem_inst__abc_19396_new_n2369_; 
wire w_mem_inst__abc_19396_new_n2370_; 
wire w_mem_inst__abc_19396_new_n2371_; 
wire w_mem_inst__abc_19396_new_n2372_; 
wire w_mem_inst__abc_19396_new_n2373_; 
wire w_mem_inst__abc_19396_new_n2374_; 
wire w_mem_inst__abc_19396_new_n2375_; 
wire w_mem_inst__abc_19396_new_n2376_; 
wire w_mem_inst__abc_19396_new_n2377_; 
wire w_mem_inst__abc_19396_new_n2378_; 
wire w_mem_inst__abc_19396_new_n2379_; 
wire w_mem_inst__abc_19396_new_n2380_; 
wire w_mem_inst__abc_19396_new_n2381_; 
wire w_mem_inst__abc_19396_new_n2382_; 
wire w_mem_inst__abc_19396_new_n2383_; 
wire w_mem_inst__abc_19396_new_n2384_; 
wire w_mem_inst__abc_19396_new_n2385_; 
wire w_mem_inst__abc_19396_new_n2386_; 
wire w_mem_inst__abc_19396_new_n2387_; 
wire w_mem_inst__abc_19396_new_n2388_; 
wire w_mem_inst__abc_19396_new_n2389_; 
wire w_mem_inst__abc_19396_new_n2390_; 
wire w_mem_inst__abc_19396_new_n2391_; 
wire w_mem_inst__abc_19396_new_n2393_; 
wire w_mem_inst__abc_19396_new_n2394_; 
wire w_mem_inst__abc_19396_new_n2395_; 
wire w_mem_inst__abc_19396_new_n2396_; 
wire w_mem_inst__abc_19396_new_n2397_; 
wire w_mem_inst__abc_19396_new_n2398_; 
wire w_mem_inst__abc_19396_new_n2399_; 
wire w_mem_inst__abc_19396_new_n2400_; 
wire w_mem_inst__abc_19396_new_n2401_; 
wire w_mem_inst__abc_19396_new_n2402_; 
wire w_mem_inst__abc_19396_new_n2403_; 
wire w_mem_inst__abc_19396_new_n2404_; 
wire w_mem_inst__abc_19396_new_n2405_; 
wire w_mem_inst__abc_19396_new_n2406_; 
wire w_mem_inst__abc_19396_new_n2407_; 
wire w_mem_inst__abc_19396_new_n2408_; 
wire w_mem_inst__abc_19396_new_n2409_; 
wire w_mem_inst__abc_19396_new_n2410_; 
wire w_mem_inst__abc_19396_new_n2411_; 
wire w_mem_inst__abc_19396_new_n2412_; 
wire w_mem_inst__abc_19396_new_n2413_; 
wire w_mem_inst__abc_19396_new_n2414_; 
wire w_mem_inst__abc_19396_new_n2415_; 
wire w_mem_inst__abc_19396_new_n2416_; 
wire w_mem_inst__abc_19396_new_n2418_; 
wire w_mem_inst__abc_19396_new_n2419_; 
wire w_mem_inst__abc_19396_new_n2420_; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf0; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf1; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf10; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf11; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf12; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf13; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf14; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf15; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf16; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf17; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf18; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf19; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf2; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf20; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf21; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf22; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf23; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf24; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf25; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf26; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf27; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf28; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf29; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf3; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf30; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf31; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf32; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf33; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf34; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf35; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf36; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf37; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf38; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf39; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf4; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf40; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf41; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf42; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf43; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf44; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf45; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf46; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf47; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf48; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf49; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf5; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf50; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf51; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf52; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf53; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf54; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf55; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf56; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf57; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf58; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf59; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf6; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf60; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf7; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf8; 
wire w_mem_inst__abc_19396_new_n2420__bF_buf9; 
wire w_mem_inst__abc_19396_new_n2420__hier0_bF_buf0; 
wire w_mem_inst__abc_19396_new_n2420__hier0_bF_buf1; 
wire w_mem_inst__abc_19396_new_n2420__hier0_bF_buf2; 
wire w_mem_inst__abc_19396_new_n2420__hier0_bF_buf3; 
wire w_mem_inst__abc_19396_new_n2420__hier0_bF_buf4; 
wire w_mem_inst__abc_19396_new_n2420__hier0_bF_buf5; 
wire w_mem_inst__abc_19396_new_n2420__hier0_bF_buf6; 
wire w_mem_inst__abc_19396_new_n2421_; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf0; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf1; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf10; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf11; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf12; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf13; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf14; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf15; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf16; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf17; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf18; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf19; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf2; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf20; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf21; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf22; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf23; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf24; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf25; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf26; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf27; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf28; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf29; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf3; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf30; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf31; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf32; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf33; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf34; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf35; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf36; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf37; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf38; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf39; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf4; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf40; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf41; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf42; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf43; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf44; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf45; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf46; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf47; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf48; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf49; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf5; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf50; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf51; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf52; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf53; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf54; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf55; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf56; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf57; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf58; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf59; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf6; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf60; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf7; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf8; 
wire w_mem_inst__abc_19396_new_n2421__bF_buf9; 
wire w_mem_inst__abc_19396_new_n2421__hier0_bF_buf0; 
wire w_mem_inst__abc_19396_new_n2421__hier0_bF_buf1; 
wire w_mem_inst__abc_19396_new_n2421__hier0_bF_buf2; 
wire w_mem_inst__abc_19396_new_n2421__hier0_bF_buf3; 
wire w_mem_inst__abc_19396_new_n2421__hier0_bF_buf4; 
wire w_mem_inst__abc_19396_new_n2421__hier0_bF_buf5; 
wire w_mem_inst__abc_19396_new_n2421__hier0_bF_buf6; 
wire w_mem_inst__abc_19396_new_n2422_; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf0; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf1; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf10; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf11; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf12; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf13; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf14; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf15; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf16; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf17; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf18; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf19; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf2; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf20; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf21; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf22; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf23; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf24; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf25; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf26; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf27; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf28; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf29; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf3; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf30; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf31; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf32; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf33; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf34; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf35; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf36; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf37; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf38; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf39; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf4; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf40; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf41; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf42; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf43; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf44; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf45; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf46; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf47; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf48; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf49; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf5; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf50; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf51; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf52; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf53; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf54; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf55; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf56; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf57; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf58; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf59; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf6; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf60; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf61; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf62; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf63; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf64; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf65; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf66; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf67; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf68; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf69; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf7; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf70; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf71; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf72; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf73; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf74; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf75; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf76; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf77; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf78; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf79; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf8; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf80; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf81; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf82; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf83; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf84; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf85; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf86; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf87; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf88; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf89; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf9; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf90; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf91; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf92; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf93; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf94; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf95; 
wire w_mem_inst__abc_19396_new_n2422__bF_buf96; 
wire w_mem_inst__abc_19396_new_n2422__hier0_bF_buf0; 
wire w_mem_inst__abc_19396_new_n2422__hier0_bF_buf1; 
wire w_mem_inst__abc_19396_new_n2422__hier0_bF_buf2; 
wire w_mem_inst__abc_19396_new_n2422__hier0_bF_buf3; 
wire w_mem_inst__abc_19396_new_n2422__hier0_bF_buf4; 
wire w_mem_inst__abc_19396_new_n2422__hier0_bF_buf5; 
wire w_mem_inst__abc_19396_new_n2422__hier0_bF_buf6; 
wire w_mem_inst__abc_19396_new_n2422__hier0_bF_buf7; 
wire w_mem_inst__abc_19396_new_n2422__hier0_bF_buf8; 
wire w_mem_inst__abc_19396_new_n2423_; 
wire w_mem_inst__abc_19396_new_n2424_; 
wire w_mem_inst__abc_19396_new_n2425_; 
wire w_mem_inst__abc_19396_new_n2427_; 
wire w_mem_inst__abc_19396_new_n2428_; 
wire w_mem_inst__abc_19396_new_n2429_; 
wire w_mem_inst__abc_19396_new_n2430_; 
wire w_mem_inst__abc_19396_new_n2432_; 
wire w_mem_inst__abc_19396_new_n2433_; 
wire w_mem_inst__abc_19396_new_n2434_; 
wire w_mem_inst__abc_19396_new_n2435_; 
wire w_mem_inst__abc_19396_new_n2437_; 
wire w_mem_inst__abc_19396_new_n2438_; 
wire w_mem_inst__abc_19396_new_n2439_; 
wire w_mem_inst__abc_19396_new_n2440_; 
wire w_mem_inst__abc_19396_new_n2442_; 
wire w_mem_inst__abc_19396_new_n2443_; 
wire w_mem_inst__abc_19396_new_n2444_; 
wire w_mem_inst__abc_19396_new_n2445_; 
wire w_mem_inst__abc_19396_new_n2447_; 
wire w_mem_inst__abc_19396_new_n2448_; 
wire w_mem_inst__abc_19396_new_n2449_; 
wire w_mem_inst__abc_19396_new_n2450_; 
wire w_mem_inst__abc_19396_new_n2452_; 
wire w_mem_inst__abc_19396_new_n2453_; 
wire w_mem_inst__abc_19396_new_n2454_; 
wire w_mem_inst__abc_19396_new_n2455_; 
wire w_mem_inst__abc_19396_new_n2457_; 
wire w_mem_inst__abc_19396_new_n2458_; 
wire w_mem_inst__abc_19396_new_n2459_; 
wire w_mem_inst__abc_19396_new_n2460_; 
wire w_mem_inst__abc_19396_new_n2462_; 
wire w_mem_inst__abc_19396_new_n2463_; 
wire w_mem_inst__abc_19396_new_n2464_; 
wire w_mem_inst__abc_19396_new_n2465_; 
wire w_mem_inst__abc_19396_new_n2467_; 
wire w_mem_inst__abc_19396_new_n2468_; 
wire w_mem_inst__abc_19396_new_n2469_; 
wire w_mem_inst__abc_19396_new_n2470_; 
wire w_mem_inst__abc_19396_new_n2472_; 
wire w_mem_inst__abc_19396_new_n2473_; 
wire w_mem_inst__abc_19396_new_n2474_; 
wire w_mem_inst__abc_19396_new_n2475_; 
wire w_mem_inst__abc_19396_new_n2477_; 
wire w_mem_inst__abc_19396_new_n2478_; 
wire w_mem_inst__abc_19396_new_n2479_; 
wire w_mem_inst__abc_19396_new_n2480_; 
wire w_mem_inst__abc_19396_new_n2482_; 
wire w_mem_inst__abc_19396_new_n2483_; 
wire w_mem_inst__abc_19396_new_n2484_; 
wire w_mem_inst__abc_19396_new_n2485_; 
wire w_mem_inst__abc_19396_new_n2487_; 
wire w_mem_inst__abc_19396_new_n2488_; 
wire w_mem_inst__abc_19396_new_n2489_; 
wire w_mem_inst__abc_19396_new_n2490_; 
wire w_mem_inst__abc_19396_new_n2492_; 
wire w_mem_inst__abc_19396_new_n2493_; 
wire w_mem_inst__abc_19396_new_n2494_; 
wire w_mem_inst__abc_19396_new_n2495_; 
wire w_mem_inst__abc_19396_new_n2497_; 
wire w_mem_inst__abc_19396_new_n2498_; 
wire w_mem_inst__abc_19396_new_n2499_; 
wire w_mem_inst__abc_19396_new_n2500_; 
wire w_mem_inst__abc_19396_new_n2502_; 
wire w_mem_inst__abc_19396_new_n2503_; 
wire w_mem_inst__abc_19396_new_n2504_; 
wire w_mem_inst__abc_19396_new_n2505_; 
wire w_mem_inst__abc_19396_new_n2507_; 
wire w_mem_inst__abc_19396_new_n2508_; 
wire w_mem_inst__abc_19396_new_n2509_; 
wire w_mem_inst__abc_19396_new_n2510_; 
wire w_mem_inst__abc_19396_new_n2512_; 
wire w_mem_inst__abc_19396_new_n2513_; 
wire w_mem_inst__abc_19396_new_n2514_; 
wire w_mem_inst__abc_19396_new_n2515_; 
wire w_mem_inst__abc_19396_new_n2517_; 
wire w_mem_inst__abc_19396_new_n2518_; 
wire w_mem_inst__abc_19396_new_n2519_; 
wire w_mem_inst__abc_19396_new_n2520_; 
wire w_mem_inst__abc_19396_new_n2522_; 
wire w_mem_inst__abc_19396_new_n2523_; 
wire w_mem_inst__abc_19396_new_n2524_; 
wire w_mem_inst__abc_19396_new_n2525_; 
wire w_mem_inst__abc_19396_new_n2527_; 
wire w_mem_inst__abc_19396_new_n2528_; 
wire w_mem_inst__abc_19396_new_n2529_; 
wire w_mem_inst__abc_19396_new_n2530_; 
wire w_mem_inst__abc_19396_new_n2532_; 
wire w_mem_inst__abc_19396_new_n2533_; 
wire w_mem_inst__abc_19396_new_n2534_; 
wire w_mem_inst__abc_19396_new_n2535_; 
wire w_mem_inst__abc_19396_new_n2537_; 
wire w_mem_inst__abc_19396_new_n2538_; 
wire w_mem_inst__abc_19396_new_n2539_; 
wire w_mem_inst__abc_19396_new_n2540_; 
wire w_mem_inst__abc_19396_new_n2542_; 
wire w_mem_inst__abc_19396_new_n2543_; 
wire w_mem_inst__abc_19396_new_n2544_; 
wire w_mem_inst__abc_19396_new_n2545_; 
wire w_mem_inst__abc_19396_new_n2547_; 
wire w_mem_inst__abc_19396_new_n2548_; 
wire w_mem_inst__abc_19396_new_n2549_; 
wire w_mem_inst__abc_19396_new_n2550_; 
wire w_mem_inst__abc_19396_new_n2552_; 
wire w_mem_inst__abc_19396_new_n2553_; 
wire w_mem_inst__abc_19396_new_n2554_; 
wire w_mem_inst__abc_19396_new_n2555_; 
wire w_mem_inst__abc_19396_new_n2557_; 
wire w_mem_inst__abc_19396_new_n2558_; 
wire w_mem_inst__abc_19396_new_n2559_; 
wire w_mem_inst__abc_19396_new_n2560_; 
wire w_mem_inst__abc_19396_new_n2562_; 
wire w_mem_inst__abc_19396_new_n2563_; 
wire w_mem_inst__abc_19396_new_n2564_; 
wire w_mem_inst__abc_19396_new_n2565_; 
wire w_mem_inst__abc_19396_new_n2567_; 
wire w_mem_inst__abc_19396_new_n2568_; 
wire w_mem_inst__abc_19396_new_n2569_; 
wire w_mem_inst__abc_19396_new_n2570_; 
wire w_mem_inst__abc_19396_new_n2572_; 
wire w_mem_inst__abc_19396_new_n2573_; 
wire w_mem_inst__abc_19396_new_n2574_; 
wire w_mem_inst__abc_19396_new_n2575_; 
wire w_mem_inst__abc_19396_new_n2577_; 
wire w_mem_inst__abc_19396_new_n2578_; 
wire w_mem_inst__abc_19396_new_n2579_; 
wire w_mem_inst__abc_19396_new_n2580_; 
wire w_mem_inst__abc_19396_new_n2582_; 
wire w_mem_inst__abc_19396_new_n2582__bF_buf0; 
wire w_mem_inst__abc_19396_new_n2582__bF_buf1; 
wire w_mem_inst__abc_19396_new_n2582__bF_buf2; 
wire w_mem_inst__abc_19396_new_n2582__bF_buf3; 
wire w_mem_inst__abc_19396_new_n2582__bF_buf4; 
wire w_mem_inst__abc_19396_new_n2583_; 
wire w_mem_inst__abc_19396_new_n2585_; 
wire w_mem_inst__abc_19396_new_n2587_; 
wire w_mem_inst__abc_19396_new_n2589_; 
wire w_mem_inst__abc_19396_new_n2591_; 
wire w_mem_inst__abc_19396_new_n2593_; 
wire w_mem_inst__abc_19396_new_n2595_; 
wire w_mem_inst__abc_19396_new_n2597_; 
wire w_mem_inst__abc_19396_new_n2599_; 
wire w_mem_inst__abc_19396_new_n2601_; 
wire w_mem_inst__abc_19396_new_n2603_; 
wire w_mem_inst__abc_19396_new_n2605_; 
wire w_mem_inst__abc_19396_new_n2607_; 
wire w_mem_inst__abc_19396_new_n2609_; 
wire w_mem_inst__abc_19396_new_n2611_; 
wire w_mem_inst__abc_19396_new_n2613_; 
wire w_mem_inst__abc_19396_new_n2615_; 
wire w_mem_inst__abc_19396_new_n2617_; 
wire w_mem_inst__abc_19396_new_n2619_; 
wire w_mem_inst__abc_19396_new_n2621_; 
wire w_mem_inst__abc_19396_new_n2623_; 
wire w_mem_inst__abc_19396_new_n2625_; 
wire w_mem_inst__abc_19396_new_n2627_; 
wire w_mem_inst__abc_19396_new_n2629_; 
wire w_mem_inst__abc_19396_new_n2631_; 
wire w_mem_inst__abc_19396_new_n2633_; 
wire w_mem_inst__abc_19396_new_n2635_; 
wire w_mem_inst__abc_19396_new_n2637_; 
wire w_mem_inst__abc_19396_new_n2639_; 
wire w_mem_inst__abc_19396_new_n2641_; 
wire w_mem_inst__abc_19396_new_n2643_; 
wire w_mem_inst__abc_19396_new_n2645_; 
wire w_mem_inst__abc_19396_new_n2647_; 
wire w_mem_inst__abc_19396_new_n2648_; 
wire w_mem_inst__abc_19396_new_n2649_; 
wire w_mem_inst__abc_19396_new_n2650_; 
wire w_mem_inst__abc_19396_new_n2652_; 
wire w_mem_inst__abc_19396_new_n2653_; 
wire w_mem_inst__abc_19396_new_n2654_; 
wire w_mem_inst__abc_19396_new_n2655_; 
wire w_mem_inst__abc_19396_new_n2657_; 
wire w_mem_inst__abc_19396_new_n2658_; 
wire w_mem_inst__abc_19396_new_n2659_; 
wire w_mem_inst__abc_19396_new_n2660_; 
wire w_mem_inst__abc_19396_new_n2662_; 
wire w_mem_inst__abc_19396_new_n2663_; 
wire w_mem_inst__abc_19396_new_n2664_; 
wire w_mem_inst__abc_19396_new_n2665_; 
wire w_mem_inst__abc_19396_new_n2667_; 
wire w_mem_inst__abc_19396_new_n2668_; 
wire w_mem_inst__abc_19396_new_n2669_; 
wire w_mem_inst__abc_19396_new_n2670_; 
wire w_mem_inst__abc_19396_new_n2672_; 
wire w_mem_inst__abc_19396_new_n2673_; 
wire w_mem_inst__abc_19396_new_n2674_; 
wire w_mem_inst__abc_19396_new_n2675_; 
wire w_mem_inst__abc_19396_new_n2677_; 
wire w_mem_inst__abc_19396_new_n2678_; 
wire w_mem_inst__abc_19396_new_n2679_; 
wire w_mem_inst__abc_19396_new_n2680_; 
wire w_mem_inst__abc_19396_new_n2682_; 
wire w_mem_inst__abc_19396_new_n2683_; 
wire w_mem_inst__abc_19396_new_n2684_; 
wire w_mem_inst__abc_19396_new_n2685_; 
wire w_mem_inst__abc_19396_new_n2687_; 
wire w_mem_inst__abc_19396_new_n2688_; 
wire w_mem_inst__abc_19396_new_n2689_; 
wire w_mem_inst__abc_19396_new_n2690_; 
wire w_mem_inst__abc_19396_new_n2692_; 
wire w_mem_inst__abc_19396_new_n2693_; 
wire w_mem_inst__abc_19396_new_n2694_; 
wire w_mem_inst__abc_19396_new_n2695_; 
wire w_mem_inst__abc_19396_new_n2697_; 
wire w_mem_inst__abc_19396_new_n2698_; 
wire w_mem_inst__abc_19396_new_n2699_; 
wire w_mem_inst__abc_19396_new_n2700_; 
wire w_mem_inst__abc_19396_new_n2702_; 
wire w_mem_inst__abc_19396_new_n2703_; 
wire w_mem_inst__abc_19396_new_n2704_; 
wire w_mem_inst__abc_19396_new_n2705_; 
wire w_mem_inst__abc_19396_new_n2707_; 
wire w_mem_inst__abc_19396_new_n2708_; 
wire w_mem_inst__abc_19396_new_n2709_; 
wire w_mem_inst__abc_19396_new_n2710_; 
wire w_mem_inst__abc_19396_new_n2712_; 
wire w_mem_inst__abc_19396_new_n2713_; 
wire w_mem_inst__abc_19396_new_n2714_; 
wire w_mem_inst__abc_19396_new_n2715_; 
wire w_mem_inst__abc_19396_new_n2717_; 
wire w_mem_inst__abc_19396_new_n2718_; 
wire w_mem_inst__abc_19396_new_n2719_; 
wire w_mem_inst__abc_19396_new_n2720_; 
wire w_mem_inst__abc_19396_new_n2722_; 
wire w_mem_inst__abc_19396_new_n2723_; 
wire w_mem_inst__abc_19396_new_n2724_; 
wire w_mem_inst__abc_19396_new_n2725_; 
wire w_mem_inst__abc_19396_new_n2727_; 
wire w_mem_inst__abc_19396_new_n2728_; 
wire w_mem_inst__abc_19396_new_n2729_; 
wire w_mem_inst__abc_19396_new_n2730_; 
wire w_mem_inst__abc_19396_new_n2732_; 
wire w_mem_inst__abc_19396_new_n2733_; 
wire w_mem_inst__abc_19396_new_n2734_; 
wire w_mem_inst__abc_19396_new_n2735_; 
wire w_mem_inst__abc_19396_new_n2737_; 
wire w_mem_inst__abc_19396_new_n2738_; 
wire w_mem_inst__abc_19396_new_n2739_; 
wire w_mem_inst__abc_19396_new_n2740_; 
wire w_mem_inst__abc_19396_new_n2742_; 
wire w_mem_inst__abc_19396_new_n2743_; 
wire w_mem_inst__abc_19396_new_n2744_; 
wire w_mem_inst__abc_19396_new_n2745_; 
wire w_mem_inst__abc_19396_new_n2747_; 
wire w_mem_inst__abc_19396_new_n2748_; 
wire w_mem_inst__abc_19396_new_n2749_; 
wire w_mem_inst__abc_19396_new_n2750_; 
wire w_mem_inst__abc_19396_new_n2752_; 
wire w_mem_inst__abc_19396_new_n2753_; 
wire w_mem_inst__abc_19396_new_n2754_; 
wire w_mem_inst__abc_19396_new_n2755_; 
wire w_mem_inst__abc_19396_new_n2757_; 
wire w_mem_inst__abc_19396_new_n2758_; 
wire w_mem_inst__abc_19396_new_n2759_; 
wire w_mem_inst__abc_19396_new_n2760_; 
wire w_mem_inst__abc_19396_new_n2762_; 
wire w_mem_inst__abc_19396_new_n2763_; 
wire w_mem_inst__abc_19396_new_n2764_; 
wire w_mem_inst__abc_19396_new_n2765_; 
wire w_mem_inst__abc_19396_new_n2767_; 
wire w_mem_inst__abc_19396_new_n2768_; 
wire w_mem_inst__abc_19396_new_n2769_; 
wire w_mem_inst__abc_19396_new_n2770_; 
wire w_mem_inst__abc_19396_new_n2772_; 
wire w_mem_inst__abc_19396_new_n2773_; 
wire w_mem_inst__abc_19396_new_n2774_; 
wire w_mem_inst__abc_19396_new_n2775_; 
wire w_mem_inst__abc_19396_new_n2777_; 
wire w_mem_inst__abc_19396_new_n2778_; 
wire w_mem_inst__abc_19396_new_n2779_; 
wire w_mem_inst__abc_19396_new_n2780_; 
wire w_mem_inst__abc_19396_new_n2782_; 
wire w_mem_inst__abc_19396_new_n2783_; 
wire w_mem_inst__abc_19396_new_n2784_; 
wire w_mem_inst__abc_19396_new_n2785_; 
wire w_mem_inst__abc_19396_new_n2787_; 
wire w_mem_inst__abc_19396_new_n2788_; 
wire w_mem_inst__abc_19396_new_n2789_; 
wire w_mem_inst__abc_19396_new_n2790_; 
wire w_mem_inst__abc_19396_new_n2792_; 
wire w_mem_inst__abc_19396_new_n2793_; 
wire w_mem_inst__abc_19396_new_n2794_; 
wire w_mem_inst__abc_19396_new_n2795_; 
wire w_mem_inst__abc_19396_new_n2797_; 
wire w_mem_inst__abc_19396_new_n2798_; 
wire w_mem_inst__abc_19396_new_n2799_; 
wire w_mem_inst__abc_19396_new_n2800_; 
wire w_mem_inst__abc_19396_new_n2802_; 
wire w_mem_inst__abc_19396_new_n2803_; 
wire w_mem_inst__abc_19396_new_n2804_; 
wire w_mem_inst__abc_19396_new_n2805_; 
wire w_mem_inst__abc_19396_new_n2807_; 
wire w_mem_inst__abc_19396_new_n2808_; 
wire w_mem_inst__abc_19396_new_n2809_; 
wire w_mem_inst__abc_19396_new_n2810_; 
wire w_mem_inst__abc_19396_new_n2812_; 
wire w_mem_inst__abc_19396_new_n2813_; 
wire w_mem_inst__abc_19396_new_n2814_; 
wire w_mem_inst__abc_19396_new_n2815_; 
wire w_mem_inst__abc_19396_new_n2817_; 
wire w_mem_inst__abc_19396_new_n2818_; 
wire w_mem_inst__abc_19396_new_n2819_; 
wire w_mem_inst__abc_19396_new_n2820_; 
wire w_mem_inst__abc_19396_new_n2822_; 
wire w_mem_inst__abc_19396_new_n2823_; 
wire w_mem_inst__abc_19396_new_n2824_; 
wire w_mem_inst__abc_19396_new_n2825_; 
wire w_mem_inst__abc_19396_new_n2827_; 
wire w_mem_inst__abc_19396_new_n2828_; 
wire w_mem_inst__abc_19396_new_n2829_; 
wire w_mem_inst__abc_19396_new_n2830_; 
wire w_mem_inst__abc_19396_new_n2832_; 
wire w_mem_inst__abc_19396_new_n2833_; 
wire w_mem_inst__abc_19396_new_n2834_; 
wire w_mem_inst__abc_19396_new_n2835_; 
wire w_mem_inst__abc_19396_new_n2837_; 
wire w_mem_inst__abc_19396_new_n2838_; 
wire w_mem_inst__abc_19396_new_n2839_; 
wire w_mem_inst__abc_19396_new_n2840_; 
wire w_mem_inst__abc_19396_new_n2842_; 
wire w_mem_inst__abc_19396_new_n2843_; 
wire w_mem_inst__abc_19396_new_n2844_; 
wire w_mem_inst__abc_19396_new_n2845_; 
wire w_mem_inst__abc_19396_new_n2847_; 
wire w_mem_inst__abc_19396_new_n2848_; 
wire w_mem_inst__abc_19396_new_n2849_; 
wire w_mem_inst__abc_19396_new_n2850_; 
wire w_mem_inst__abc_19396_new_n2852_; 
wire w_mem_inst__abc_19396_new_n2853_; 
wire w_mem_inst__abc_19396_new_n2854_; 
wire w_mem_inst__abc_19396_new_n2855_; 
wire w_mem_inst__abc_19396_new_n2857_; 
wire w_mem_inst__abc_19396_new_n2858_; 
wire w_mem_inst__abc_19396_new_n2859_; 
wire w_mem_inst__abc_19396_new_n2860_; 
wire w_mem_inst__abc_19396_new_n2862_; 
wire w_mem_inst__abc_19396_new_n2863_; 
wire w_mem_inst__abc_19396_new_n2864_; 
wire w_mem_inst__abc_19396_new_n2865_; 
wire w_mem_inst__abc_19396_new_n2867_; 
wire w_mem_inst__abc_19396_new_n2868_; 
wire w_mem_inst__abc_19396_new_n2869_; 
wire w_mem_inst__abc_19396_new_n2870_; 
wire w_mem_inst__abc_19396_new_n2872_; 
wire w_mem_inst__abc_19396_new_n2873_; 
wire w_mem_inst__abc_19396_new_n2874_; 
wire w_mem_inst__abc_19396_new_n2875_; 
wire w_mem_inst__abc_19396_new_n2877_; 
wire w_mem_inst__abc_19396_new_n2878_; 
wire w_mem_inst__abc_19396_new_n2879_; 
wire w_mem_inst__abc_19396_new_n2880_; 
wire w_mem_inst__abc_19396_new_n2882_; 
wire w_mem_inst__abc_19396_new_n2883_; 
wire w_mem_inst__abc_19396_new_n2884_; 
wire w_mem_inst__abc_19396_new_n2885_; 
wire w_mem_inst__abc_19396_new_n2887_; 
wire w_mem_inst__abc_19396_new_n2888_; 
wire w_mem_inst__abc_19396_new_n2889_; 
wire w_mem_inst__abc_19396_new_n2890_; 
wire w_mem_inst__abc_19396_new_n2892_; 
wire w_mem_inst__abc_19396_new_n2893_; 
wire w_mem_inst__abc_19396_new_n2894_; 
wire w_mem_inst__abc_19396_new_n2895_; 
wire w_mem_inst__abc_19396_new_n2897_; 
wire w_mem_inst__abc_19396_new_n2898_; 
wire w_mem_inst__abc_19396_new_n2899_; 
wire w_mem_inst__abc_19396_new_n2900_; 
wire w_mem_inst__abc_19396_new_n2902_; 
wire w_mem_inst__abc_19396_new_n2903_; 
wire w_mem_inst__abc_19396_new_n2904_; 
wire w_mem_inst__abc_19396_new_n2905_; 
wire w_mem_inst__abc_19396_new_n2907_; 
wire w_mem_inst__abc_19396_new_n2908_; 
wire w_mem_inst__abc_19396_new_n2909_; 
wire w_mem_inst__abc_19396_new_n2910_; 
wire w_mem_inst__abc_19396_new_n2912_; 
wire w_mem_inst__abc_19396_new_n2913_; 
wire w_mem_inst__abc_19396_new_n2914_; 
wire w_mem_inst__abc_19396_new_n2915_; 
wire w_mem_inst__abc_19396_new_n2917_; 
wire w_mem_inst__abc_19396_new_n2918_; 
wire w_mem_inst__abc_19396_new_n2919_; 
wire w_mem_inst__abc_19396_new_n2920_; 
wire w_mem_inst__abc_19396_new_n2922_; 
wire w_mem_inst__abc_19396_new_n2923_; 
wire w_mem_inst__abc_19396_new_n2924_; 
wire w_mem_inst__abc_19396_new_n2925_; 
wire w_mem_inst__abc_19396_new_n2927_; 
wire w_mem_inst__abc_19396_new_n2928_; 
wire w_mem_inst__abc_19396_new_n2929_; 
wire w_mem_inst__abc_19396_new_n2930_; 
wire w_mem_inst__abc_19396_new_n2932_; 
wire w_mem_inst__abc_19396_new_n2933_; 
wire w_mem_inst__abc_19396_new_n2934_; 
wire w_mem_inst__abc_19396_new_n2935_; 
wire w_mem_inst__abc_19396_new_n2937_; 
wire w_mem_inst__abc_19396_new_n2938_; 
wire w_mem_inst__abc_19396_new_n2939_; 
wire w_mem_inst__abc_19396_new_n2940_; 
wire w_mem_inst__abc_19396_new_n2942_; 
wire w_mem_inst__abc_19396_new_n2943_; 
wire w_mem_inst__abc_19396_new_n2944_; 
wire w_mem_inst__abc_19396_new_n2945_; 
wire w_mem_inst__abc_19396_new_n2947_; 
wire w_mem_inst__abc_19396_new_n2948_; 
wire w_mem_inst__abc_19396_new_n2949_; 
wire w_mem_inst__abc_19396_new_n2950_; 
wire w_mem_inst__abc_19396_new_n2952_; 
wire w_mem_inst__abc_19396_new_n2953_; 
wire w_mem_inst__abc_19396_new_n2954_; 
wire w_mem_inst__abc_19396_new_n2955_; 
wire w_mem_inst__abc_19396_new_n2957_; 
wire w_mem_inst__abc_19396_new_n2958_; 
wire w_mem_inst__abc_19396_new_n2959_; 
wire w_mem_inst__abc_19396_new_n2960_; 
wire w_mem_inst__abc_19396_new_n2962_; 
wire w_mem_inst__abc_19396_new_n2963_; 
wire w_mem_inst__abc_19396_new_n2964_; 
wire w_mem_inst__abc_19396_new_n2965_; 
wire w_mem_inst__abc_19396_new_n2967_; 
wire w_mem_inst__abc_19396_new_n2968_; 
wire w_mem_inst__abc_19396_new_n2969_; 
wire w_mem_inst__abc_19396_new_n2970_; 
wire w_mem_inst__abc_19396_new_n2972_; 
wire w_mem_inst__abc_19396_new_n2973_; 
wire w_mem_inst__abc_19396_new_n2974_; 
wire w_mem_inst__abc_19396_new_n2975_; 
wire w_mem_inst__abc_19396_new_n2977_; 
wire w_mem_inst__abc_19396_new_n2978_; 
wire w_mem_inst__abc_19396_new_n2979_; 
wire w_mem_inst__abc_19396_new_n2980_; 
wire w_mem_inst__abc_19396_new_n2982_; 
wire w_mem_inst__abc_19396_new_n2983_; 
wire w_mem_inst__abc_19396_new_n2984_; 
wire w_mem_inst__abc_19396_new_n2985_; 
wire w_mem_inst__abc_19396_new_n2987_; 
wire w_mem_inst__abc_19396_new_n2988_; 
wire w_mem_inst__abc_19396_new_n2989_; 
wire w_mem_inst__abc_19396_new_n2990_; 
wire w_mem_inst__abc_19396_new_n2992_; 
wire w_mem_inst__abc_19396_new_n2993_; 
wire w_mem_inst__abc_19396_new_n2994_; 
wire w_mem_inst__abc_19396_new_n2995_; 
wire w_mem_inst__abc_19396_new_n2997_; 
wire w_mem_inst__abc_19396_new_n2998_; 
wire w_mem_inst__abc_19396_new_n2999_; 
wire w_mem_inst__abc_19396_new_n3000_; 
wire w_mem_inst__abc_19396_new_n3002_; 
wire w_mem_inst__abc_19396_new_n3003_; 
wire w_mem_inst__abc_19396_new_n3004_; 
wire w_mem_inst__abc_19396_new_n3005_; 
wire w_mem_inst__abc_19396_new_n3007_; 
wire w_mem_inst__abc_19396_new_n3008_; 
wire w_mem_inst__abc_19396_new_n3009_; 
wire w_mem_inst__abc_19396_new_n3010_; 
wire w_mem_inst__abc_19396_new_n3012_; 
wire w_mem_inst__abc_19396_new_n3013_; 
wire w_mem_inst__abc_19396_new_n3014_; 
wire w_mem_inst__abc_19396_new_n3015_; 
wire w_mem_inst__abc_19396_new_n3017_; 
wire w_mem_inst__abc_19396_new_n3018_; 
wire w_mem_inst__abc_19396_new_n3019_; 
wire w_mem_inst__abc_19396_new_n3020_; 
wire w_mem_inst__abc_19396_new_n3022_; 
wire w_mem_inst__abc_19396_new_n3023_; 
wire w_mem_inst__abc_19396_new_n3024_; 
wire w_mem_inst__abc_19396_new_n3025_; 
wire w_mem_inst__abc_19396_new_n3027_; 
wire w_mem_inst__abc_19396_new_n3028_; 
wire w_mem_inst__abc_19396_new_n3029_; 
wire w_mem_inst__abc_19396_new_n3030_; 
wire w_mem_inst__abc_19396_new_n3032_; 
wire w_mem_inst__abc_19396_new_n3033_; 
wire w_mem_inst__abc_19396_new_n3034_; 
wire w_mem_inst__abc_19396_new_n3035_; 
wire w_mem_inst__abc_19396_new_n3037_; 
wire w_mem_inst__abc_19396_new_n3038_; 
wire w_mem_inst__abc_19396_new_n3039_; 
wire w_mem_inst__abc_19396_new_n3040_; 
wire w_mem_inst__abc_19396_new_n3042_; 
wire w_mem_inst__abc_19396_new_n3043_; 
wire w_mem_inst__abc_19396_new_n3044_; 
wire w_mem_inst__abc_19396_new_n3045_; 
wire w_mem_inst__abc_19396_new_n3047_; 
wire w_mem_inst__abc_19396_new_n3048_; 
wire w_mem_inst__abc_19396_new_n3049_; 
wire w_mem_inst__abc_19396_new_n3050_; 
wire w_mem_inst__abc_19396_new_n3052_; 
wire w_mem_inst__abc_19396_new_n3053_; 
wire w_mem_inst__abc_19396_new_n3054_; 
wire w_mem_inst__abc_19396_new_n3055_; 
wire w_mem_inst__abc_19396_new_n3057_; 
wire w_mem_inst__abc_19396_new_n3058_; 
wire w_mem_inst__abc_19396_new_n3059_; 
wire w_mem_inst__abc_19396_new_n3060_; 
wire w_mem_inst__abc_19396_new_n3062_; 
wire w_mem_inst__abc_19396_new_n3063_; 
wire w_mem_inst__abc_19396_new_n3064_; 
wire w_mem_inst__abc_19396_new_n3065_; 
wire w_mem_inst__abc_19396_new_n3067_; 
wire w_mem_inst__abc_19396_new_n3068_; 
wire w_mem_inst__abc_19396_new_n3069_; 
wire w_mem_inst__abc_19396_new_n3070_; 
wire w_mem_inst__abc_19396_new_n3072_; 
wire w_mem_inst__abc_19396_new_n3073_; 
wire w_mem_inst__abc_19396_new_n3074_; 
wire w_mem_inst__abc_19396_new_n3075_; 
wire w_mem_inst__abc_19396_new_n3077_; 
wire w_mem_inst__abc_19396_new_n3078_; 
wire w_mem_inst__abc_19396_new_n3079_; 
wire w_mem_inst__abc_19396_new_n3080_; 
wire w_mem_inst__abc_19396_new_n3082_; 
wire w_mem_inst__abc_19396_new_n3083_; 
wire w_mem_inst__abc_19396_new_n3084_; 
wire w_mem_inst__abc_19396_new_n3085_; 
wire w_mem_inst__abc_19396_new_n3087_; 
wire w_mem_inst__abc_19396_new_n3088_; 
wire w_mem_inst__abc_19396_new_n3089_; 
wire w_mem_inst__abc_19396_new_n3090_; 
wire w_mem_inst__abc_19396_new_n3092_; 
wire w_mem_inst__abc_19396_new_n3093_; 
wire w_mem_inst__abc_19396_new_n3094_; 
wire w_mem_inst__abc_19396_new_n3095_; 
wire w_mem_inst__abc_19396_new_n3097_; 
wire w_mem_inst__abc_19396_new_n3098_; 
wire w_mem_inst__abc_19396_new_n3099_; 
wire w_mem_inst__abc_19396_new_n3100_; 
wire w_mem_inst__abc_19396_new_n3102_; 
wire w_mem_inst__abc_19396_new_n3103_; 
wire w_mem_inst__abc_19396_new_n3104_; 
wire w_mem_inst__abc_19396_new_n3105_; 
wire w_mem_inst__abc_19396_new_n3107_; 
wire w_mem_inst__abc_19396_new_n3108_; 
wire w_mem_inst__abc_19396_new_n3109_; 
wire w_mem_inst__abc_19396_new_n3110_; 
wire w_mem_inst__abc_19396_new_n3112_; 
wire w_mem_inst__abc_19396_new_n3113_; 
wire w_mem_inst__abc_19396_new_n3114_; 
wire w_mem_inst__abc_19396_new_n3115_; 
wire w_mem_inst__abc_19396_new_n3117_; 
wire w_mem_inst__abc_19396_new_n3118_; 
wire w_mem_inst__abc_19396_new_n3119_; 
wire w_mem_inst__abc_19396_new_n3120_; 
wire w_mem_inst__abc_19396_new_n3122_; 
wire w_mem_inst__abc_19396_new_n3123_; 
wire w_mem_inst__abc_19396_new_n3124_; 
wire w_mem_inst__abc_19396_new_n3125_; 
wire w_mem_inst__abc_19396_new_n3127_; 
wire w_mem_inst__abc_19396_new_n3128_; 
wire w_mem_inst__abc_19396_new_n3129_; 
wire w_mem_inst__abc_19396_new_n3130_; 
wire w_mem_inst__abc_19396_new_n3132_; 
wire w_mem_inst__abc_19396_new_n3133_; 
wire w_mem_inst__abc_19396_new_n3134_; 
wire w_mem_inst__abc_19396_new_n3135_; 
wire w_mem_inst__abc_19396_new_n3137_; 
wire w_mem_inst__abc_19396_new_n3138_; 
wire w_mem_inst__abc_19396_new_n3139_; 
wire w_mem_inst__abc_19396_new_n3140_; 
wire w_mem_inst__abc_19396_new_n3142_; 
wire w_mem_inst__abc_19396_new_n3143_; 
wire w_mem_inst__abc_19396_new_n3144_; 
wire w_mem_inst__abc_19396_new_n3145_; 
wire w_mem_inst__abc_19396_new_n3147_; 
wire w_mem_inst__abc_19396_new_n3148_; 
wire w_mem_inst__abc_19396_new_n3149_; 
wire w_mem_inst__abc_19396_new_n3150_; 
wire w_mem_inst__abc_19396_new_n3152_; 
wire w_mem_inst__abc_19396_new_n3153_; 
wire w_mem_inst__abc_19396_new_n3154_; 
wire w_mem_inst__abc_19396_new_n3155_; 
wire w_mem_inst__abc_19396_new_n3157_; 
wire w_mem_inst__abc_19396_new_n3158_; 
wire w_mem_inst__abc_19396_new_n3159_; 
wire w_mem_inst__abc_19396_new_n3160_; 
wire w_mem_inst__abc_19396_new_n3162_; 
wire w_mem_inst__abc_19396_new_n3163_; 
wire w_mem_inst__abc_19396_new_n3164_; 
wire w_mem_inst__abc_19396_new_n3165_; 
wire w_mem_inst__abc_19396_new_n3167_; 
wire w_mem_inst__abc_19396_new_n3168_; 
wire w_mem_inst__abc_19396_new_n3169_; 
wire w_mem_inst__abc_19396_new_n3170_; 
wire w_mem_inst__abc_19396_new_n3172_; 
wire w_mem_inst__abc_19396_new_n3173_; 
wire w_mem_inst__abc_19396_new_n3174_; 
wire w_mem_inst__abc_19396_new_n3175_; 
wire w_mem_inst__abc_19396_new_n3177_; 
wire w_mem_inst__abc_19396_new_n3178_; 
wire w_mem_inst__abc_19396_new_n3179_; 
wire w_mem_inst__abc_19396_new_n3180_; 
wire w_mem_inst__abc_19396_new_n3182_; 
wire w_mem_inst__abc_19396_new_n3183_; 
wire w_mem_inst__abc_19396_new_n3184_; 
wire w_mem_inst__abc_19396_new_n3185_; 
wire w_mem_inst__abc_19396_new_n3187_; 
wire w_mem_inst__abc_19396_new_n3188_; 
wire w_mem_inst__abc_19396_new_n3189_; 
wire w_mem_inst__abc_19396_new_n3190_; 
wire w_mem_inst__abc_19396_new_n3192_; 
wire w_mem_inst__abc_19396_new_n3193_; 
wire w_mem_inst__abc_19396_new_n3194_; 
wire w_mem_inst__abc_19396_new_n3195_; 
wire w_mem_inst__abc_19396_new_n3197_; 
wire w_mem_inst__abc_19396_new_n3198_; 
wire w_mem_inst__abc_19396_new_n3199_; 
wire w_mem_inst__abc_19396_new_n3200_; 
wire w_mem_inst__abc_19396_new_n3202_; 
wire w_mem_inst__abc_19396_new_n3203_; 
wire w_mem_inst__abc_19396_new_n3204_; 
wire w_mem_inst__abc_19396_new_n3205_; 
wire w_mem_inst__abc_19396_new_n3207_; 
wire w_mem_inst__abc_19396_new_n3208_; 
wire w_mem_inst__abc_19396_new_n3209_; 
wire w_mem_inst__abc_19396_new_n3210_; 
wire w_mem_inst__abc_19396_new_n3212_; 
wire w_mem_inst__abc_19396_new_n3213_; 
wire w_mem_inst__abc_19396_new_n3214_; 
wire w_mem_inst__abc_19396_new_n3215_; 
wire w_mem_inst__abc_19396_new_n3217_; 
wire w_mem_inst__abc_19396_new_n3218_; 
wire w_mem_inst__abc_19396_new_n3219_; 
wire w_mem_inst__abc_19396_new_n3220_; 
wire w_mem_inst__abc_19396_new_n3222_; 
wire w_mem_inst__abc_19396_new_n3223_; 
wire w_mem_inst__abc_19396_new_n3224_; 
wire w_mem_inst__abc_19396_new_n3225_; 
wire w_mem_inst__abc_19396_new_n3227_; 
wire w_mem_inst__abc_19396_new_n3228_; 
wire w_mem_inst__abc_19396_new_n3229_; 
wire w_mem_inst__abc_19396_new_n3230_; 
wire w_mem_inst__abc_19396_new_n3232_; 
wire w_mem_inst__abc_19396_new_n3233_; 
wire w_mem_inst__abc_19396_new_n3234_; 
wire w_mem_inst__abc_19396_new_n3235_; 
wire w_mem_inst__abc_19396_new_n3237_; 
wire w_mem_inst__abc_19396_new_n3238_; 
wire w_mem_inst__abc_19396_new_n3239_; 
wire w_mem_inst__abc_19396_new_n3240_; 
wire w_mem_inst__abc_19396_new_n3242_; 
wire w_mem_inst__abc_19396_new_n3243_; 
wire w_mem_inst__abc_19396_new_n3244_; 
wire w_mem_inst__abc_19396_new_n3245_; 
wire w_mem_inst__abc_19396_new_n3247_; 
wire w_mem_inst__abc_19396_new_n3248_; 
wire w_mem_inst__abc_19396_new_n3249_; 
wire w_mem_inst__abc_19396_new_n3250_; 
wire w_mem_inst__abc_19396_new_n3252_; 
wire w_mem_inst__abc_19396_new_n3253_; 
wire w_mem_inst__abc_19396_new_n3254_; 
wire w_mem_inst__abc_19396_new_n3255_; 
wire w_mem_inst__abc_19396_new_n3257_; 
wire w_mem_inst__abc_19396_new_n3258_; 
wire w_mem_inst__abc_19396_new_n3259_; 
wire w_mem_inst__abc_19396_new_n3260_; 
wire w_mem_inst__abc_19396_new_n3262_; 
wire w_mem_inst__abc_19396_new_n3263_; 
wire w_mem_inst__abc_19396_new_n3264_; 
wire w_mem_inst__abc_19396_new_n3265_; 
wire w_mem_inst__abc_19396_new_n3267_; 
wire w_mem_inst__abc_19396_new_n3268_; 
wire w_mem_inst__abc_19396_new_n3269_; 
wire w_mem_inst__abc_19396_new_n3270_; 
wire w_mem_inst__abc_19396_new_n3272_; 
wire w_mem_inst__abc_19396_new_n3273_; 
wire w_mem_inst__abc_19396_new_n3274_; 
wire w_mem_inst__abc_19396_new_n3275_; 
wire w_mem_inst__abc_19396_new_n3277_; 
wire w_mem_inst__abc_19396_new_n3278_; 
wire w_mem_inst__abc_19396_new_n3279_; 
wire w_mem_inst__abc_19396_new_n3280_; 
wire w_mem_inst__abc_19396_new_n3282_; 
wire w_mem_inst__abc_19396_new_n3283_; 
wire w_mem_inst__abc_19396_new_n3284_; 
wire w_mem_inst__abc_19396_new_n3285_; 
wire w_mem_inst__abc_19396_new_n3287_; 
wire w_mem_inst__abc_19396_new_n3288_; 
wire w_mem_inst__abc_19396_new_n3289_; 
wire w_mem_inst__abc_19396_new_n3291_; 
wire w_mem_inst__abc_19396_new_n3292_; 
wire w_mem_inst__abc_19396_new_n3293_; 
wire w_mem_inst__abc_19396_new_n3295_; 
wire w_mem_inst__abc_19396_new_n3296_; 
wire w_mem_inst__abc_19396_new_n3297_; 
wire w_mem_inst__abc_19396_new_n3299_; 
wire w_mem_inst__abc_19396_new_n3300_; 
wire w_mem_inst__abc_19396_new_n3301_; 
wire w_mem_inst__abc_19396_new_n3303_; 
wire w_mem_inst__abc_19396_new_n3304_; 
wire w_mem_inst__abc_19396_new_n3305_; 
wire w_mem_inst__abc_19396_new_n3307_; 
wire w_mem_inst__abc_19396_new_n3308_; 
wire w_mem_inst__abc_19396_new_n3309_; 
wire w_mem_inst__abc_19396_new_n3311_; 
wire w_mem_inst__abc_19396_new_n3312_; 
wire w_mem_inst__abc_19396_new_n3313_; 
wire w_mem_inst__abc_19396_new_n3315_; 
wire w_mem_inst__abc_19396_new_n3316_; 
wire w_mem_inst__abc_19396_new_n3317_; 
wire w_mem_inst__abc_19396_new_n3319_; 
wire w_mem_inst__abc_19396_new_n3320_; 
wire w_mem_inst__abc_19396_new_n3321_; 
wire w_mem_inst__abc_19396_new_n3323_; 
wire w_mem_inst__abc_19396_new_n3324_; 
wire w_mem_inst__abc_19396_new_n3325_; 
wire w_mem_inst__abc_19396_new_n3327_; 
wire w_mem_inst__abc_19396_new_n3328_; 
wire w_mem_inst__abc_19396_new_n3329_; 
wire w_mem_inst__abc_19396_new_n3331_; 
wire w_mem_inst__abc_19396_new_n3332_; 
wire w_mem_inst__abc_19396_new_n3333_; 
wire w_mem_inst__abc_19396_new_n3335_; 
wire w_mem_inst__abc_19396_new_n3336_; 
wire w_mem_inst__abc_19396_new_n3337_; 
wire w_mem_inst__abc_19396_new_n3339_; 
wire w_mem_inst__abc_19396_new_n3340_; 
wire w_mem_inst__abc_19396_new_n3341_; 
wire w_mem_inst__abc_19396_new_n3343_; 
wire w_mem_inst__abc_19396_new_n3344_; 
wire w_mem_inst__abc_19396_new_n3345_; 
wire w_mem_inst__abc_19396_new_n3347_; 
wire w_mem_inst__abc_19396_new_n3348_; 
wire w_mem_inst__abc_19396_new_n3349_; 
wire w_mem_inst__abc_19396_new_n3351_; 
wire w_mem_inst__abc_19396_new_n3352_; 
wire w_mem_inst__abc_19396_new_n3353_; 
wire w_mem_inst__abc_19396_new_n3355_; 
wire w_mem_inst__abc_19396_new_n3356_; 
wire w_mem_inst__abc_19396_new_n3357_; 
wire w_mem_inst__abc_19396_new_n3359_; 
wire w_mem_inst__abc_19396_new_n3360_; 
wire w_mem_inst__abc_19396_new_n3361_; 
wire w_mem_inst__abc_19396_new_n3363_; 
wire w_mem_inst__abc_19396_new_n3364_; 
wire w_mem_inst__abc_19396_new_n3365_; 
wire w_mem_inst__abc_19396_new_n3367_; 
wire w_mem_inst__abc_19396_new_n3368_; 
wire w_mem_inst__abc_19396_new_n3369_; 
wire w_mem_inst__abc_19396_new_n3371_; 
wire w_mem_inst__abc_19396_new_n3372_; 
wire w_mem_inst__abc_19396_new_n3373_; 
wire w_mem_inst__abc_19396_new_n3375_; 
wire w_mem_inst__abc_19396_new_n3376_; 
wire w_mem_inst__abc_19396_new_n3377_; 
wire w_mem_inst__abc_19396_new_n3379_; 
wire w_mem_inst__abc_19396_new_n3380_; 
wire w_mem_inst__abc_19396_new_n3381_; 
wire w_mem_inst__abc_19396_new_n3383_; 
wire w_mem_inst__abc_19396_new_n3384_; 
wire w_mem_inst__abc_19396_new_n3385_; 
wire w_mem_inst__abc_19396_new_n3387_; 
wire w_mem_inst__abc_19396_new_n3388_; 
wire w_mem_inst__abc_19396_new_n3389_; 
wire w_mem_inst__abc_19396_new_n3391_; 
wire w_mem_inst__abc_19396_new_n3392_; 
wire w_mem_inst__abc_19396_new_n3393_; 
wire w_mem_inst__abc_19396_new_n3395_; 
wire w_mem_inst__abc_19396_new_n3396_; 
wire w_mem_inst__abc_19396_new_n3397_; 
wire w_mem_inst__abc_19396_new_n3399_; 
wire w_mem_inst__abc_19396_new_n3400_; 
wire w_mem_inst__abc_19396_new_n3401_; 
wire w_mem_inst__abc_19396_new_n3403_; 
wire w_mem_inst__abc_19396_new_n3404_; 
wire w_mem_inst__abc_19396_new_n3405_; 
wire w_mem_inst__abc_19396_new_n3407_; 
wire w_mem_inst__abc_19396_new_n3408_; 
wire w_mem_inst__abc_19396_new_n3409_; 
wire w_mem_inst__abc_19396_new_n3411_; 
wire w_mem_inst__abc_19396_new_n3412_; 
wire w_mem_inst__abc_19396_new_n3413_; 
wire w_mem_inst__abc_19396_new_n3415_; 
wire w_mem_inst__abc_19396_new_n3416_; 
wire w_mem_inst__abc_19396_new_n3417_; 
wire w_mem_inst__abc_19396_new_n3418_; 
wire w_mem_inst__abc_19396_new_n3420_; 
wire w_mem_inst__abc_19396_new_n3421_; 
wire w_mem_inst__abc_19396_new_n3422_; 
wire w_mem_inst__abc_19396_new_n3423_; 
wire w_mem_inst__abc_19396_new_n3425_; 
wire w_mem_inst__abc_19396_new_n3426_; 
wire w_mem_inst__abc_19396_new_n3427_; 
wire w_mem_inst__abc_19396_new_n3428_; 
wire w_mem_inst__abc_19396_new_n3430_; 
wire w_mem_inst__abc_19396_new_n3431_; 
wire w_mem_inst__abc_19396_new_n3432_; 
wire w_mem_inst__abc_19396_new_n3433_; 
wire w_mem_inst__abc_19396_new_n3435_; 
wire w_mem_inst__abc_19396_new_n3436_; 
wire w_mem_inst__abc_19396_new_n3437_; 
wire w_mem_inst__abc_19396_new_n3438_; 
wire w_mem_inst__abc_19396_new_n3440_; 
wire w_mem_inst__abc_19396_new_n3441_; 
wire w_mem_inst__abc_19396_new_n3442_; 
wire w_mem_inst__abc_19396_new_n3443_; 
wire w_mem_inst__abc_19396_new_n3445_; 
wire w_mem_inst__abc_19396_new_n3446_; 
wire w_mem_inst__abc_19396_new_n3447_; 
wire w_mem_inst__abc_19396_new_n3448_; 
wire w_mem_inst__abc_19396_new_n3450_; 
wire w_mem_inst__abc_19396_new_n3451_; 
wire w_mem_inst__abc_19396_new_n3452_; 
wire w_mem_inst__abc_19396_new_n3453_; 
wire w_mem_inst__abc_19396_new_n3455_; 
wire w_mem_inst__abc_19396_new_n3456_; 
wire w_mem_inst__abc_19396_new_n3457_; 
wire w_mem_inst__abc_19396_new_n3458_; 
wire w_mem_inst__abc_19396_new_n3460_; 
wire w_mem_inst__abc_19396_new_n3461_; 
wire w_mem_inst__abc_19396_new_n3462_; 
wire w_mem_inst__abc_19396_new_n3463_; 
wire w_mem_inst__abc_19396_new_n3465_; 
wire w_mem_inst__abc_19396_new_n3466_; 
wire w_mem_inst__abc_19396_new_n3467_; 
wire w_mem_inst__abc_19396_new_n3468_; 
wire w_mem_inst__abc_19396_new_n3470_; 
wire w_mem_inst__abc_19396_new_n3471_; 
wire w_mem_inst__abc_19396_new_n3472_; 
wire w_mem_inst__abc_19396_new_n3473_; 
wire w_mem_inst__abc_19396_new_n3475_; 
wire w_mem_inst__abc_19396_new_n3476_; 
wire w_mem_inst__abc_19396_new_n3477_; 
wire w_mem_inst__abc_19396_new_n3478_; 
wire w_mem_inst__abc_19396_new_n3480_; 
wire w_mem_inst__abc_19396_new_n3481_; 
wire w_mem_inst__abc_19396_new_n3482_; 
wire w_mem_inst__abc_19396_new_n3483_; 
wire w_mem_inst__abc_19396_new_n3485_; 
wire w_mem_inst__abc_19396_new_n3486_; 
wire w_mem_inst__abc_19396_new_n3487_; 
wire w_mem_inst__abc_19396_new_n3488_; 
wire w_mem_inst__abc_19396_new_n3490_; 
wire w_mem_inst__abc_19396_new_n3491_; 
wire w_mem_inst__abc_19396_new_n3492_; 
wire w_mem_inst__abc_19396_new_n3493_; 
wire w_mem_inst__abc_19396_new_n3495_; 
wire w_mem_inst__abc_19396_new_n3496_; 
wire w_mem_inst__abc_19396_new_n3497_; 
wire w_mem_inst__abc_19396_new_n3498_; 
wire w_mem_inst__abc_19396_new_n3500_; 
wire w_mem_inst__abc_19396_new_n3501_; 
wire w_mem_inst__abc_19396_new_n3502_; 
wire w_mem_inst__abc_19396_new_n3503_; 
wire w_mem_inst__abc_19396_new_n3505_; 
wire w_mem_inst__abc_19396_new_n3506_; 
wire w_mem_inst__abc_19396_new_n3507_; 
wire w_mem_inst__abc_19396_new_n3508_; 
wire w_mem_inst__abc_19396_new_n3510_; 
wire w_mem_inst__abc_19396_new_n3511_; 
wire w_mem_inst__abc_19396_new_n3512_; 
wire w_mem_inst__abc_19396_new_n3513_; 
wire w_mem_inst__abc_19396_new_n3515_; 
wire w_mem_inst__abc_19396_new_n3516_; 
wire w_mem_inst__abc_19396_new_n3517_; 
wire w_mem_inst__abc_19396_new_n3518_; 
wire w_mem_inst__abc_19396_new_n3520_; 
wire w_mem_inst__abc_19396_new_n3521_; 
wire w_mem_inst__abc_19396_new_n3522_; 
wire w_mem_inst__abc_19396_new_n3523_; 
wire w_mem_inst__abc_19396_new_n3525_; 
wire w_mem_inst__abc_19396_new_n3526_; 
wire w_mem_inst__abc_19396_new_n3527_; 
wire w_mem_inst__abc_19396_new_n3528_; 
wire w_mem_inst__abc_19396_new_n3530_; 
wire w_mem_inst__abc_19396_new_n3531_; 
wire w_mem_inst__abc_19396_new_n3532_; 
wire w_mem_inst__abc_19396_new_n3533_; 
wire w_mem_inst__abc_19396_new_n3535_; 
wire w_mem_inst__abc_19396_new_n3536_; 
wire w_mem_inst__abc_19396_new_n3537_; 
wire w_mem_inst__abc_19396_new_n3538_; 
wire w_mem_inst__abc_19396_new_n3540_; 
wire w_mem_inst__abc_19396_new_n3541_; 
wire w_mem_inst__abc_19396_new_n3542_; 
wire w_mem_inst__abc_19396_new_n3543_; 
wire w_mem_inst__abc_19396_new_n3545_; 
wire w_mem_inst__abc_19396_new_n3546_; 
wire w_mem_inst__abc_19396_new_n3547_; 
wire w_mem_inst__abc_19396_new_n3548_; 
wire w_mem_inst__abc_19396_new_n3550_; 
wire w_mem_inst__abc_19396_new_n3551_; 
wire w_mem_inst__abc_19396_new_n3552_; 
wire w_mem_inst__abc_19396_new_n3553_; 
wire w_mem_inst__abc_19396_new_n3555_; 
wire w_mem_inst__abc_19396_new_n3556_; 
wire w_mem_inst__abc_19396_new_n3557_; 
wire w_mem_inst__abc_19396_new_n3558_; 
wire w_mem_inst__abc_19396_new_n3560_; 
wire w_mem_inst__abc_19396_new_n3561_; 
wire w_mem_inst__abc_19396_new_n3562_; 
wire w_mem_inst__abc_19396_new_n3563_; 
wire w_mem_inst__abc_19396_new_n3565_; 
wire w_mem_inst__abc_19396_new_n3566_; 
wire w_mem_inst__abc_19396_new_n3567_; 
wire w_mem_inst__abc_19396_new_n3568_; 
wire w_mem_inst__abc_19396_new_n3570_; 
wire w_mem_inst__abc_19396_new_n3571_; 
wire w_mem_inst__abc_19396_new_n3572_; 
wire w_mem_inst__abc_19396_new_n3573_; 
wire w_mem_inst__abc_19396_new_n3575_; 
wire w_mem_inst__abc_19396_new_n3576_; 
wire w_mem_inst__abc_19396_new_n3577_; 
wire w_mem_inst__abc_19396_new_n3579_; 
wire w_mem_inst__abc_19396_new_n3580_; 
wire w_mem_inst__abc_19396_new_n3581_; 
wire w_mem_inst__abc_19396_new_n3583_; 
wire w_mem_inst__abc_19396_new_n3584_; 
wire w_mem_inst__abc_19396_new_n3585_; 
wire w_mem_inst__abc_19396_new_n3587_; 
wire w_mem_inst__abc_19396_new_n3588_; 
wire w_mem_inst__abc_19396_new_n3589_; 
wire w_mem_inst__abc_19396_new_n3591_; 
wire w_mem_inst__abc_19396_new_n3592_; 
wire w_mem_inst__abc_19396_new_n3593_; 
wire w_mem_inst__abc_19396_new_n3595_; 
wire w_mem_inst__abc_19396_new_n3596_; 
wire w_mem_inst__abc_19396_new_n3597_; 
wire w_mem_inst__abc_19396_new_n3599_; 
wire w_mem_inst__abc_19396_new_n3600_; 
wire w_mem_inst__abc_19396_new_n3601_; 
wire w_mem_inst__abc_19396_new_n3603_; 
wire w_mem_inst__abc_19396_new_n3604_; 
wire w_mem_inst__abc_19396_new_n3605_; 
wire w_mem_inst__abc_19396_new_n3607_; 
wire w_mem_inst__abc_19396_new_n3608_; 
wire w_mem_inst__abc_19396_new_n3609_; 
wire w_mem_inst__abc_19396_new_n3611_; 
wire w_mem_inst__abc_19396_new_n3612_; 
wire w_mem_inst__abc_19396_new_n3613_; 
wire w_mem_inst__abc_19396_new_n3615_; 
wire w_mem_inst__abc_19396_new_n3616_; 
wire w_mem_inst__abc_19396_new_n3617_; 
wire w_mem_inst__abc_19396_new_n3619_; 
wire w_mem_inst__abc_19396_new_n3620_; 
wire w_mem_inst__abc_19396_new_n3621_; 
wire w_mem_inst__abc_19396_new_n3623_; 
wire w_mem_inst__abc_19396_new_n3624_; 
wire w_mem_inst__abc_19396_new_n3625_; 
wire w_mem_inst__abc_19396_new_n3627_; 
wire w_mem_inst__abc_19396_new_n3628_; 
wire w_mem_inst__abc_19396_new_n3629_; 
wire w_mem_inst__abc_19396_new_n3631_; 
wire w_mem_inst__abc_19396_new_n3632_; 
wire w_mem_inst__abc_19396_new_n3633_; 
wire w_mem_inst__abc_19396_new_n3635_; 
wire w_mem_inst__abc_19396_new_n3636_; 
wire w_mem_inst__abc_19396_new_n3637_; 
wire w_mem_inst__abc_19396_new_n3639_; 
wire w_mem_inst__abc_19396_new_n3640_; 
wire w_mem_inst__abc_19396_new_n3641_; 
wire w_mem_inst__abc_19396_new_n3643_; 
wire w_mem_inst__abc_19396_new_n3644_; 
wire w_mem_inst__abc_19396_new_n3645_; 
wire w_mem_inst__abc_19396_new_n3647_; 
wire w_mem_inst__abc_19396_new_n3648_; 
wire w_mem_inst__abc_19396_new_n3649_; 
wire w_mem_inst__abc_19396_new_n3651_; 
wire w_mem_inst__abc_19396_new_n3652_; 
wire w_mem_inst__abc_19396_new_n3653_; 
wire w_mem_inst__abc_19396_new_n3655_; 
wire w_mem_inst__abc_19396_new_n3656_; 
wire w_mem_inst__abc_19396_new_n3657_; 
wire w_mem_inst__abc_19396_new_n3659_; 
wire w_mem_inst__abc_19396_new_n3660_; 
wire w_mem_inst__abc_19396_new_n3661_; 
wire w_mem_inst__abc_19396_new_n3663_; 
wire w_mem_inst__abc_19396_new_n3664_; 
wire w_mem_inst__abc_19396_new_n3665_; 
wire w_mem_inst__abc_19396_new_n3667_; 
wire w_mem_inst__abc_19396_new_n3668_; 
wire w_mem_inst__abc_19396_new_n3669_; 
wire w_mem_inst__abc_19396_new_n3671_; 
wire w_mem_inst__abc_19396_new_n3672_; 
wire w_mem_inst__abc_19396_new_n3673_; 
wire w_mem_inst__abc_19396_new_n3675_; 
wire w_mem_inst__abc_19396_new_n3676_; 
wire w_mem_inst__abc_19396_new_n3677_; 
wire w_mem_inst__abc_19396_new_n3679_; 
wire w_mem_inst__abc_19396_new_n3680_; 
wire w_mem_inst__abc_19396_new_n3681_; 
wire w_mem_inst__abc_19396_new_n3683_; 
wire w_mem_inst__abc_19396_new_n3684_; 
wire w_mem_inst__abc_19396_new_n3685_; 
wire w_mem_inst__abc_19396_new_n3687_; 
wire w_mem_inst__abc_19396_new_n3688_; 
wire w_mem_inst__abc_19396_new_n3689_; 
wire w_mem_inst__abc_19396_new_n3691_; 
wire w_mem_inst__abc_19396_new_n3692_; 
wire w_mem_inst__abc_19396_new_n3693_; 
wire w_mem_inst__abc_19396_new_n3695_; 
wire w_mem_inst__abc_19396_new_n3696_; 
wire w_mem_inst__abc_19396_new_n3697_; 
wire w_mem_inst__abc_19396_new_n3699_; 
wire w_mem_inst__abc_19396_new_n3700_; 
wire w_mem_inst__abc_19396_new_n3701_; 
wire w_mem_inst__abc_19396_new_n3703_; 
wire w_mem_inst__abc_19396_new_n3704_; 
wire w_mem_inst__abc_19396_new_n3705_; 
wire w_mem_inst__abc_19396_new_n3706_; 
wire w_mem_inst__abc_19396_new_n3708_; 
wire w_mem_inst__abc_19396_new_n3709_; 
wire w_mem_inst__abc_19396_new_n3710_; 
wire w_mem_inst__abc_19396_new_n3711_; 
wire w_mem_inst__abc_19396_new_n3713_; 
wire w_mem_inst__abc_19396_new_n3714_; 
wire w_mem_inst__abc_19396_new_n3715_; 
wire w_mem_inst__abc_19396_new_n3716_; 
wire w_mem_inst__abc_19396_new_n3718_; 
wire w_mem_inst__abc_19396_new_n3719_; 
wire w_mem_inst__abc_19396_new_n3720_; 
wire w_mem_inst__abc_19396_new_n3721_; 
wire w_mem_inst__abc_19396_new_n3723_; 
wire w_mem_inst__abc_19396_new_n3724_; 
wire w_mem_inst__abc_19396_new_n3725_; 
wire w_mem_inst__abc_19396_new_n3726_; 
wire w_mem_inst__abc_19396_new_n3728_; 
wire w_mem_inst__abc_19396_new_n3729_; 
wire w_mem_inst__abc_19396_new_n3730_; 
wire w_mem_inst__abc_19396_new_n3731_; 
wire w_mem_inst__abc_19396_new_n3733_; 
wire w_mem_inst__abc_19396_new_n3734_; 
wire w_mem_inst__abc_19396_new_n3735_; 
wire w_mem_inst__abc_19396_new_n3736_; 
wire w_mem_inst__abc_19396_new_n3738_; 
wire w_mem_inst__abc_19396_new_n3739_; 
wire w_mem_inst__abc_19396_new_n3740_; 
wire w_mem_inst__abc_19396_new_n3741_; 
wire w_mem_inst__abc_19396_new_n3743_; 
wire w_mem_inst__abc_19396_new_n3744_; 
wire w_mem_inst__abc_19396_new_n3745_; 
wire w_mem_inst__abc_19396_new_n3746_; 
wire w_mem_inst__abc_19396_new_n3748_; 
wire w_mem_inst__abc_19396_new_n3749_; 
wire w_mem_inst__abc_19396_new_n3750_; 
wire w_mem_inst__abc_19396_new_n3751_; 
wire w_mem_inst__abc_19396_new_n3753_; 
wire w_mem_inst__abc_19396_new_n3754_; 
wire w_mem_inst__abc_19396_new_n3755_; 
wire w_mem_inst__abc_19396_new_n3756_; 
wire w_mem_inst__abc_19396_new_n3758_; 
wire w_mem_inst__abc_19396_new_n3759_; 
wire w_mem_inst__abc_19396_new_n3760_; 
wire w_mem_inst__abc_19396_new_n3761_; 
wire w_mem_inst__abc_19396_new_n3763_; 
wire w_mem_inst__abc_19396_new_n3764_; 
wire w_mem_inst__abc_19396_new_n3765_; 
wire w_mem_inst__abc_19396_new_n3766_; 
wire w_mem_inst__abc_19396_new_n3768_; 
wire w_mem_inst__abc_19396_new_n3769_; 
wire w_mem_inst__abc_19396_new_n3770_; 
wire w_mem_inst__abc_19396_new_n3771_; 
wire w_mem_inst__abc_19396_new_n3773_; 
wire w_mem_inst__abc_19396_new_n3774_; 
wire w_mem_inst__abc_19396_new_n3775_; 
wire w_mem_inst__abc_19396_new_n3776_; 
wire w_mem_inst__abc_19396_new_n3778_; 
wire w_mem_inst__abc_19396_new_n3779_; 
wire w_mem_inst__abc_19396_new_n3780_; 
wire w_mem_inst__abc_19396_new_n3781_; 
wire w_mem_inst__abc_19396_new_n3783_; 
wire w_mem_inst__abc_19396_new_n3784_; 
wire w_mem_inst__abc_19396_new_n3785_; 
wire w_mem_inst__abc_19396_new_n3786_; 
wire w_mem_inst__abc_19396_new_n3788_; 
wire w_mem_inst__abc_19396_new_n3789_; 
wire w_mem_inst__abc_19396_new_n3790_; 
wire w_mem_inst__abc_19396_new_n3791_; 
wire w_mem_inst__abc_19396_new_n3793_; 
wire w_mem_inst__abc_19396_new_n3794_; 
wire w_mem_inst__abc_19396_new_n3795_; 
wire w_mem_inst__abc_19396_new_n3796_; 
wire w_mem_inst__abc_19396_new_n3798_; 
wire w_mem_inst__abc_19396_new_n3799_; 
wire w_mem_inst__abc_19396_new_n3800_; 
wire w_mem_inst__abc_19396_new_n3801_; 
wire w_mem_inst__abc_19396_new_n3803_; 
wire w_mem_inst__abc_19396_new_n3804_; 
wire w_mem_inst__abc_19396_new_n3805_; 
wire w_mem_inst__abc_19396_new_n3806_; 
wire w_mem_inst__abc_19396_new_n3808_; 
wire w_mem_inst__abc_19396_new_n3809_; 
wire w_mem_inst__abc_19396_new_n3810_; 
wire w_mem_inst__abc_19396_new_n3811_; 
wire w_mem_inst__abc_19396_new_n3813_; 
wire w_mem_inst__abc_19396_new_n3814_; 
wire w_mem_inst__abc_19396_new_n3815_; 
wire w_mem_inst__abc_19396_new_n3816_; 
wire w_mem_inst__abc_19396_new_n3818_; 
wire w_mem_inst__abc_19396_new_n3819_; 
wire w_mem_inst__abc_19396_new_n3820_; 
wire w_mem_inst__abc_19396_new_n3821_; 
wire w_mem_inst__abc_19396_new_n3823_; 
wire w_mem_inst__abc_19396_new_n3824_; 
wire w_mem_inst__abc_19396_new_n3825_; 
wire w_mem_inst__abc_19396_new_n3826_; 
wire w_mem_inst__abc_19396_new_n3828_; 
wire w_mem_inst__abc_19396_new_n3829_; 
wire w_mem_inst__abc_19396_new_n3830_; 
wire w_mem_inst__abc_19396_new_n3831_; 
wire w_mem_inst__abc_19396_new_n3833_; 
wire w_mem_inst__abc_19396_new_n3834_; 
wire w_mem_inst__abc_19396_new_n3835_; 
wire w_mem_inst__abc_19396_new_n3836_; 
wire w_mem_inst__abc_19396_new_n3838_; 
wire w_mem_inst__abc_19396_new_n3839_; 
wire w_mem_inst__abc_19396_new_n3840_; 
wire w_mem_inst__abc_19396_new_n3841_; 
wire w_mem_inst__abc_19396_new_n3843_; 
wire w_mem_inst__abc_19396_new_n3844_; 
wire w_mem_inst__abc_19396_new_n3845_; 
wire w_mem_inst__abc_19396_new_n3846_; 
wire w_mem_inst__abc_19396_new_n3848_; 
wire w_mem_inst__abc_19396_new_n3849_; 
wire w_mem_inst__abc_19396_new_n3850_; 
wire w_mem_inst__abc_19396_new_n3851_; 
wire w_mem_inst__abc_19396_new_n3853_; 
wire w_mem_inst__abc_19396_new_n3854_; 
wire w_mem_inst__abc_19396_new_n3855_; 
wire w_mem_inst__abc_19396_new_n3856_; 
wire w_mem_inst__abc_19396_new_n3858_; 
wire w_mem_inst__abc_19396_new_n3859_; 
wire w_mem_inst__abc_19396_new_n3860_; 
wire w_mem_inst__abc_19396_new_n3861_; 
wire w_mem_inst__abc_19396_new_n3863_; 
wire w_mem_inst__abc_19396_new_n3864_; 
wire w_mem_inst__abc_19396_new_n3865_; 
wire w_mem_inst__abc_19396_new_n3866_; 
wire w_mem_inst__abc_19396_new_n3868_; 
wire w_mem_inst__abc_19396_new_n3869_; 
wire w_mem_inst__abc_19396_new_n3870_; 
wire w_mem_inst__abc_19396_new_n3871_; 
wire w_mem_inst__abc_19396_new_n3873_; 
wire w_mem_inst__abc_19396_new_n3874_; 
wire w_mem_inst__abc_19396_new_n3875_; 
wire w_mem_inst__abc_19396_new_n3876_; 
wire w_mem_inst__abc_19396_new_n3878_; 
wire w_mem_inst__abc_19396_new_n3879_; 
wire w_mem_inst__abc_19396_new_n3880_; 
wire w_mem_inst__abc_19396_new_n3881_; 
wire w_mem_inst__abc_19396_new_n3883_; 
wire w_mem_inst__abc_19396_new_n3884_; 
wire w_mem_inst__abc_19396_new_n3885_; 
wire w_mem_inst__abc_19396_new_n3886_; 
wire w_mem_inst__abc_19396_new_n3888_; 
wire w_mem_inst__abc_19396_new_n3889_; 
wire w_mem_inst__abc_19396_new_n3890_; 
wire w_mem_inst__abc_19396_new_n3891_; 
wire w_mem_inst__abc_19396_new_n3893_; 
wire w_mem_inst__abc_19396_new_n3894_; 
wire w_mem_inst__abc_19396_new_n3895_; 
wire w_mem_inst__abc_19396_new_n3896_; 
wire w_mem_inst__abc_19396_new_n3898_; 
wire w_mem_inst__abc_19396_new_n3899_; 
wire w_mem_inst__abc_19396_new_n3900_; 
wire w_mem_inst__abc_19396_new_n3901_; 
wire w_mem_inst__abc_19396_new_n3903_; 
wire w_mem_inst__abc_19396_new_n3904_; 
wire w_mem_inst__abc_19396_new_n3905_; 
wire w_mem_inst__abc_19396_new_n3906_; 
wire w_mem_inst__abc_19396_new_n3908_; 
wire w_mem_inst__abc_19396_new_n3909_; 
wire w_mem_inst__abc_19396_new_n3910_; 
wire w_mem_inst__abc_19396_new_n3911_; 
wire w_mem_inst__abc_19396_new_n3913_; 
wire w_mem_inst__abc_19396_new_n3914_; 
wire w_mem_inst__abc_19396_new_n3915_; 
wire w_mem_inst__abc_19396_new_n3916_; 
wire w_mem_inst__abc_19396_new_n3918_; 
wire w_mem_inst__abc_19396_new_n3919_; 
wire w_mem_inst__abc_19396_new_n3920_; 
wire w_mem_inst__abc_19396_new_n3921_; 
wire w_mem_inst__abc_19396_new_n3923_; 
wire w_mem_inst__abc_19396_new_n3924_; 
wire w_mem_inst__abc_19396_new_n3925_; 
wire w_mem_inst__abc_19396_new_n3926_; 
wire w_mem_inst__abc_19396_new_n3928_; 
wire w_mem_inst__abc_19396_new_n3929_; 
wire w_mem_inst__abc_19396_new_n3930_; 
wire w_mem_inst__abc_19396_new_n3931_; 
wire w_mem_inst__abc_19396_new_n3933_; 
wire w_mem_inst__abc_19396_new_n3934_; 
wire w_mem_inst__abc_19396_new_n3935_; 
wire w_mem_inst__abc_19396_new_n3936_; 
wire w_mem_inst__abc_19396_new_n3938_; 
wire w_mem_inst__abc_19396_new_n3939_; 
wire w_mem_inst__abc_19396_new_n3940_; 
wire w_mem_inst__abc_19396_new_n3941_; 
wire w_mem_inst__abc_19396_new_n3943_; 
wire w_mem_inst__abc_19396_new_n3944_; 
wire w_mem_inst__abc_19396_new_n3945_; 
wire w_mem_inst__abc_19396_new_n3946_; 
wire w_mem_inst__abc_19396_new_n3948_; 
wire w_mem_inst__abc_19396_new_n3949_; 
wire w_mem_inst__abc_19396_new_n3950_; 
wire w_mem_inst__abc_19396_new_n3951_; 
wire w_mem_inst__abc_19396_new_n3953_; 
wire w_mem_inst__abc_19396_new_n3954_; 
wire w_mem_inst__abc_19396_new_n3955_; 
wire w_mem_inst__abc_19396_new_n3956_; 
wire w_mem_inst__abc_19396_new_n3958_; 
wire w_mem_inst__abc_19396_new_n3959_; 
wire w_mem_inst__abc_19396_new_n3960_; 
wire w_mem_inst__abc_19396_new_n3961_; 
wire w_mem_inst__abc_19396_new_n3963_; 
wire w_mem_inst__abc_19396_new_n3964_; 
wire w_mem_inst__abc_19396_new_n3965_; 
wire w_mem_inst__abc_19396_new_n3966_; 
wire w_mem_inst__abc_19396_new_n3968_; 
wire w_mem_inst__abc_19396_new_n3969_; 
wire w_mem_inst__abc_19396_new_n3970_; 
wire w_mem_inst__abc_19396_new_n3971_; 
wire w_mem_inst__abc_19396_new_n3973_; 
wire w_mem_inst__abc_19396_new_n3974_; 
wire w_mem_inst__abc_19396_new_n3975_; 
wire w_mem_inst__abc_19396_new_n3976_; 
wire w_mem_inst__abc_19396_new_n3978_; 
wire w_mem_inst__abc_19396_new_n3979_; 
wire w_mem_inst__abc_19396_new_n3980_; 
wire w_mem_inst__abc_19396_new_n3981_; 
wire w_mem_inst__abc_19396_new_n3983_; 
wire w_mem_inst__abc_19396_new_n3984_; 
wire w_mem_inst__abc_19396_new_n3985_; 
wire w_mem_inst__abc_19396_new_n3986_; 
wire w_mem_inst__abc_19396_new_n3988_; 
wire w_mem_inst__abc_19396_new_n3989_; 
wire w_mem_inst__abc_19396_new_n3990_; 
wire w_mem_inst__abc_19396_new_n3991_; 
wire w_mem_inst__abc_19396_new_n3993_; 
wire w_mem_inst__abc_19396_new_n3994_; 
wire w_mem_inst__abc_19396_new_n3995_; 
wire w_mem_inst__abc_19396_new_n3996_; 
wire w_mem_inst__abc_19396_new_n3998_; 
wire w_mem_inst__abc_19396_new_n3999_; 
wire w_mem_inst__abc_19396_new_n4000_; 
wire w_mem_inst__abc_19396_new_n4001_; 
wire w_mem_inst__abc_19396_new_n4003_; 
wire w_mem_inst__abc_19396_new_n4004_; 
wire w_mem_inst__abc_19396_new_n4005_; 
wire w_mem_inst__abc_19396_new_n4006_; 
wire w_mem_inst__abc_19396_new_n4008_; 
wire w_mem_inst__abc_19396_new_n4009_; 
wire w_mem_inst__abc_19396_new_n4010_; 
wire w_mem_inst__abc_19396_new_n4011_; 
wire w_mem_inst__abc_19396_new_n4013_; 
wire w_mem_inst__abc_19396_new_n4014_; 
wire w_mem_inst__abc_19396_new_n4015_; 
wire w_mem_inst__abc_19396_new_n4016_; 
wire w_mem_inst__abc_19396_new_n4018_; 
wire w_mem_inst__abc_19396_new_n4019_; 
wire w_mem_inst__abc_19396_new_n4020_; 
wire w_mem_inst__abc_19396_new_n4021_; 
wire w_mem_inst__abc_19396_new_n4023_; 
wire w_mem_inst__abc_19396_new_n4024_; 
wire w_mem_inst__abc_19396_new_n4025_; 
wire w_mem_inst__abc_19396_new_n4027_; 
wire w_mem_inst__abc_19396_new_n4028_; 
wire w_mem_inst__abc_19396_new_n4029_; 
wire w_mem_inst__abc_19396_new_n4031_; 
wire w_mem_inst__abc_19396_new_n4032_; 
wire w_mem_inst__abc_19396_new_n4033_; 
wire w_mem_inst__abc_19396_new_n4035_; 
wire w_mem_inst__abc_19396_new_n4036_; 
wire w_mem_inst__abc_19396_new_n4037_; 
wire w_mem_inst__abc_19396_new_n4039_; 
wire w_mem_inst__abc_19396_new_n4040_; 
wire w_mem_inst__abc_19396_new_n4041_; 
wire w_mem_inst__abc_19396_new_n4043_; 
wire w_mem_inst__abc_19396_new_n4044_; 
wire w_mem_inst__abc_19396_new_n4045_; 
wire w_mem_inst__abc_19396_new_n4047_; 
wire w_mem_inst__abc_19396_new_n4048_; 
wire w_mem_inst__abc_19396_new_n4049_; 
wire w_mem_inst__abc_19396_new_n4051_; 
wire w_mem_inst__abc_19396_new_n4052_; 
wire w_mem_inst__abc_19396_new_n4053_; 
wire w_mem_inst__abc_19396_new_n4055_; 
wire w_mem_inst__abc_19396_new_n4056_; 
wire w_mem_inst__abc_19396_new_n4057_; 
wire w_mem_inst__abc_19396_new_n4059_; 
wire w_mem_inst__abc_19396_new_n4060_; 
wire w_mem_inst__abc_19396_new_n4061_; 
wire w_mem_inst__abc_19396_new_n4063_; 
wire w_mem_inst__abc_19396_new_n4064_; 
wire w_mem_inst__abc_19396_new_n4065_; 
wire w_mem_inst__abc_19396_new_n4067_; 
wire w_mem_inst__abc_19396_new_n4068_; 
wire w_mem_inst__abc_19396_new_n4069_; 
wire w_mem_inst__abc_19396_new_n4071_; 
wire w_mem_inst__abc_19396_new_n4072_; 
wire w_mem_inst__abc_19396_new_n4073_; 
wire w_mem_inst__abc_19396_new_n4075_; 
wire w_mem_inst__abc_19396_new_n4076_; 
wire w_mem_inst__abc_19396_new_n4077_; 
wire w_mem_inst__abc_19396_new_n4079_; 
wire w_mem_inst__abc_19396_new_n4080_; 
wire w_mem_inst__abc_19396_new_n4081_; 
wire w_mem_inst__abc_19396_new_n4083_; 
wire w_mem_inst__abc_19396_new_n4084_; 
wire w_mem_inst__abc_19396_new_n4085_; 
wire w_mem_inst__abc_19396_new_n4087_; 
wire w_mem_inst__abc_19396_new_n4088_; 
wire w_mem_inst__abc_19396_new_n4089_; 
wire w_mem_inst__abc_19396_new_n4091_; 
wire w_mem_inst__abc_19396_new_n4092_; 
wire w_mem_inst__abc_19396_new_n4093_; 
wire w_mem_inst__abc_19396_new_n4095_; 
wire w_mem_inst__abc_19396_new_n4096_; 
wire w_mem_inst__abc_19396_new_n4097_; 
wire w_mem_inst__abc_19396_new_n4099_; 
wire w_mem_inst__abc_19396_new_n4100_; 
wire w_mem_inst__abc_19396_new_n4101_; 
wire w_mem_inst__abc_19396_new_n4103_; 
wire w_mem_inst__abc_19396_new_n4104_; 
wire w_mem_inst__abc_19396_new_n4105_; 
wire w_mem_inst__abc_19396_new_n4107_; 
wire w_mem_inst__abc_19396_new_n4108_; 
wire w_mem_inst__abc_19396_new_n4109_; 
wire w_mem_inst__abc_19396_new_n4111_; 
wire w_mem_inst__abc_19396_new_n4112_; 
wire w_mem_inst__abc_19396_new_n4113_; 
wire w_mem_inst__abc_19396_new_n4115_; 
wire w_mem_inst__abc_19396_new_n4116_; 
wire w_mem_inst__abc_19396_new_n4117_; 
wire w_mem_inst__abc_19396_new_n4119_; 
wire w_mem_inst__abc_19396_new_n4120_; 
wire w_mem_inst__abc_19396_new_n4121_; 
wire w_mem_inst__abc_19396_new_n4123_; 
wire w_mem_inst__abc_19396_new_n4124_; 
wire w_mem_inst__abc_19396_new_n4125_; 
wire w_mem_inst__abc_19396_new_n4127_; 
wire w_mem_inst__abc_19396_new_n4128_; 
wire w_mem_inst__abc_19396_new_n4129_; 
wire w_mem_inst__abc_19396_new_n4131_; 
wire w_mem_inst__abc_19396_new_n4132_; 
wire w_mem_inst__abc_19396_new_n4133_; 
wire w_mem_inst__abc_19396_new_n4135_; 
wire w_mem_inst__abc_19396_new_n4136_; 
wire w_mem_inst__abc_19396_new_n4137_; 
wire w_mem_inst__abc_19396_new_n4139_; 
wire w_mem_inst__abc_19396_new_n4140_; 
wire w_mem_inst__abc_19396_new_n4141_; 
wire w_mem_inst__abc_19396_new_n4143_; 
wire w_mem_inst__abc_19396_new_n4144_; 
wire w_mem_inst__abc_19396_new_n4145_; 
wire w_mem_inst__abc_19396_new_n4147_; 
wire w_mem_inst__abc_19396_new_n4148_; 
wire w_mem_inst__abc_19396_new_n4149_; 
wire w_mem_inst__abc_19396_new_n4151_; 
wire w_mem_inst__abc_19396_new_n4152_; 
wire w_mem_inst__abc_19396_new_n4153_; 
wire w_mem_inst__abc_19396_new_n4154_; 
wire w_mem_inst__abc_19396_new_n4156_; 
wire w_mem_inst__abc_19396_new_n4157_; 
wire w_mem_inst__abc_19396_new_n4158_; 
wire w_mem_inst__abc_19396_new_n4159_; 
wire w_mem_inst__abc_19396_new_n4161_; 
wire w_mem_inst__abc_19396_new_n4162_; 
wire w_mem_inst__abc_19396_new_n4163_; 
wire w_mem_inst__abc_19396_new_n4164_; 
wire w_mem_inst__abc_19396_new_n4166_; 
wire w_mem_inst__abc_19396_new_n4167_; 
wire w_mem_inst__abc_19396_new_n4168_; 
wire w_mem_inst__abc_19396_new_n4169_; 
wire w_mem_inst__abc_19396_new_n4171_; 
wire w_mem_inst__abc_19396_new_n4172_; 
wire w_mem_inst__abc_19396_new_n4173_; 
wire w_mem_inst__abc_19396_new_n4174_; 
wire w_mem_inst__abc_19396_new_n4176_; 
wire w_mem_inst__abc_19396_new_n4177_; 
wire w_mem_inst__abc_19396_new_n4178_; 
wire w_mem_inst__abc_19396_new_n4179_; 
wire w_mem_inst__abc_19396_new_n4181_; 
wire w_mem_inst__abc_19396_new_n4182_; 
wire w_mem_inst__abc_19396_new_n4183_; 
wire w_mem_inst__abc_19396_new_n4184_; 
wire w_mem_inst__abc_19396_new_n4186_; 
wire w_mem_inst__abc_19396_new_n4187_; 
wire w_mem_inst__abc_19396_new_n4188_; 
wire w_mem_inst__abc_19396_new_n4189_; 
wire w_mem_inst__abc_19396_new_n4191_; 
wire w_mem_inst__abc_19396_new_n4192_; 
wire w_mem_inst__abc_19396_new_n4193_; 
wire w_mem_inst__abc_19396_new_n4194_; 
wire w_mem_inst__abc_19396_new_n4196_; 
wire w_mem_inst__abc_19396_new_n4197_; 
wire w_mem_inst__abc_19396_new_n4198_; 
wire w_mem_inst__abc_19396_new_n4199_; 
wire w_mem_inst__abc_19396_new_n4201_; 
wire w_mem_inst__abc_19396_new_n4202_; 
wire w_mem_inst__abc_19396_new_n4203_; 
wire w_mem_inst__abc_19396_new_n4204_; 
wire w_mem_inst__abc_19396_new_n4206_; 
wire w_mem_inst__abc_19396_new_n4207_; 
wire w_mem_inst__abc_19396_new_n4208_; 
wire w_mem_inst__abc_19396_new_n4209_; 
wire w_mem_inst__abc_19396_new_n4211_; 
wire w_mem_inst__abc_19396_new_n4212_; 
wire w_mem_inst__abc_19396_new_n4213_; 
wire w_mem_inst__abc_19396_new_n4214_; 
wire w_mem_inst__abc_19396_new_n4216_; 
wire w_mem_inst__abc_19396_new_n4217_; 
wire w_mem_inst__abc_19396_new_n4218_; 
wire w_mem_inst__abc_19396_new_n4219_; 
wire w_mem_inst__abc_19396_new_n4221_; 
wire w_mem_inst__abc_19396_new_n4222_; 
wire w_mem_inst__abc_19396_new_n4223_; 
wire w_mem_inst__abc_19396_new_n4224_; 
wire w_mem_inst__abc_19396_new_n4226_; 
wire w_mem_inst__abc_19396_new_n4227_; 
wire w_mem_inst__abc_19396_new_n4228_; 
wire w_mem_inst__abc_19396_new_n4229_; 
wire w_mem_inst__abc_19396_new_n4231_; 
wire w_mem_inst__abc_19396_new_n4232_; 
wire w_mem_inst__abc_19396_new_n4233_; 
wire w_mem_inst__abc_19396_new_n4234_; 
wire w_mem_inst__abc_19396_new_n4236_; 
wire w_mem_inst__abc_19396_new_n4237_; 
wire w_mem_inst__abc_19396_new_n4238_; 
wire w_mem_inst__abc_19396_new_n4239_; 
wire w_mem_inst__abc_19396_new_n4241_; 
wire w_mem_inst__abc_19396_new_n4242_; 
wire w_mem_inst__abc_19396_new_n4243_; 
wire w_mem_inst__abc_19396_new_n4244_; 
wire w_mem_inst__abc_19396_new_n4246_; 
wire w_mem_inst__abc_19396_new_n4247_; 
wire w_mem_inst__abc_19396_new_n4248_; 
wire w_mem_inst__abc_19396_new_n4249_; 
wire w_mem_inst__abc_19396_new_n4251_; 
wire w_mem_inst__abc_19396_new_n4252_; 
wire w_mem_inst__abc_19396_new_n4253_; 
wire w_mem_inst__abc_19396_new_n4254_; 
wire w_mem_inst__abc_19396_new_n4256_; 
wire w_mem_inst__abc_19396_new_n4257_; 
wire w_mem_inst__abc_19396_new_n4258_; 
wire w_mem_inst__abc_19396_new_n4259_; 
wire w_mem_inst__abc_19396_new_n4261_; 
wire w_mem_inst__abc_19396_new_n4262_; 
wire w_mem_inst__abc_19396_new_n4263_; 
wire w_mem_inst__abc_19396_new_n4264_; 
wire w_mem_inst__abc_19396_new_n4266_; 
wire w_mem_inst__abc_19396_new_n4267_; 
wire w_mem_inst__abc_19396_new_n4268_; 
wire w_mem_inst__abc_19396_new_n4269_; 
wire w_mem_inst__abc_19396_new_n4271_; 
wire w_mem_inst__abc_19396_new_n4272_; 
wire w_mem_inst__abc_19396_new_n4273_; 
wire w_mem_inst__abc_19396_new_n4274_; 
wire w_mem_inst__abc_19396_new_n4276_; 
wire w_mem_inst__abc_19396_new_n4277_; 
wire w_mem_inst__abc_19396_new_n4278_; 
wire w_mem_inst__abc_19396_new_n4279_; 
wire w_mem_inst__abc_19396_new_n4281_; 
wire w_mem_inst__abc_19396_new_n4282_; 
wire w_mem_inst__abc_19396_new_n4283_; 
wire w_mem_inst__abc_19396_new_n4284_; 
wire w_mem_inst__abc_19396_new_n4286_; 
wire w_mem_inst__abc_19396_new_n4287_; 
wire w_mem_inst__abc_19396_new_n4288_; 
wire w_mem_inst__abc_19396_new_n4289_; 
wire w_mem_inst__abc_19396_new_n4291_; 
wire w_mem_inst__abc_19396_new_n4292_; 
wire w_mem_inst__abc_19396_new_n4293_; 
wire w_mem_inst__abc_19396_new_n4294_; 
wire w_mem_inst__abc_19396_new_n4296_; 
wire w_mem_inst__abc_19396_new_n4297_; 
wire w_mem_inst__abc_19396_new_n4298_; 
wire w_mem_inst__abc_19396_new_n4299_; 
wire w_mem_inst__abc_19396_new_n4301_; 
wire w_mem_inst__abc_19396_new_n4302_; 
wire w_mem_inst__abc_19396_new_n4303_; 
wire w_mem_inst__abc_19396_new_n4304_; 
wire w_mem_inst__abc_19396_new_n4306_; 
wire w_mem_inst__abc_19396_new_n4307_; 
wire w_mem_inst__abc_19396_new_n4308_; 
wire w_mem_inst__abc_19396_new_n4309_; 
wire w_mem_inst__abc_19396_new_n4311_; 
wire w_mem_inst__abc_19396_new_n4312_; 
wire w_mem_inst__abc_19396_new_n4313_; 
wire w_mem_inst__abc_19396_new_n4314_; 
wire w_mem_inst__abc_19396_new_n4316_; 
wire w_mem_inst__abc_19396_new_n4317_; 
wire w_mem_inst__abc_19396_new_n4318_; 
wire w_mem_inst__abc_19396_new_n4319_; 
wire w_mem_inst__abc_19396_new_n4321_; 
wire w_mem_inst__abc_19396_new_n4322_; 
wire w_mem_inst__abc_19396_new_n4323_; 
wire w_mem_inst__abc_19396_new_n4324_; 
wire w_mem_inst__abc_19396_new_n4326_; 
wire w_mem_inst__abc_19396_new_n4327_; 
wire w_mem_inst__abc_19396_new_n4328_; 
wire w_mem_inst__abc_19396_new_n4329_; 
wire w_mem_inst__abc_19396_new_n4331_; 
wire w_mem_inst__abc_19396_new_n4332_; 
wire w_mem_inst__abc_19396_new_n4333_; 
wire w_mem_inst__abc_19396_new_n4334_; 
wire w_mem_inst__abc_19396_new_n4336_; 
wire w_mem_inst__abc_19396_new_n4337_; 
wire w_mem_inst__abc_19396_new_n4338_; 
wire w_mem_inst__abc_19396_new_n4339_; 
wire w_mem_inst__abc_19396_new_n4341_; 
wire w_mem_inst__abc_19396_new_n4342_; 
wire w_mem_inst__abc_19396_new_n4343_; 
wire w_mem_inst__abc_19396_new_n4344_; 
wire w_mem_inst__abc_19396_new_n4346_; 
wire w_mem_inst__abc_19396_new_n4347_; 
wire w_mem_inst__abc_19396_new_n4348_; 
wire w_mem_inst__abc_19396_new_n4349_; 
wire w_mem_inst__abc_19396_new_n4351_; 
wire w_mem_inst__abc_19396_new_n4352_; 
wire w_mem_inst__abc_19396_new_n4353_; 
wire w_mem_inst__abc_19396_new_n4354_; 
wire w_mem_inst__abc_19396_new_n4356_; 
wire w_mem_inst__abc_19396_new_n4357_; 
wire w_mem_inst__abc_19396_new_n4358_; 
wire w_mem_inst__abc_19396_new_n4359_; 
wire w_mem_inst__abc_19396_new_n4361_; 
wire w_mem_inst__abc_19396_new_n4362_; 
wire w_mem_inst__abc_19396_new_n4363_; 
wire w_mem_inst__abc_19396_new_n4364_; 
wire w_mem_inst__abc_19396_new_n4366_; 
wire w_mem_inst__abc_19396_new_n4367_; 
wire w_mem_inst__abc_19396_new_n4368_; 
wire w_mem_inst__abc_19396_new_n4369_; 
wire w_mem_inst__abc_19396_new_n4371_; 
wire w_mem_inst__abc_19396_new_n4372_; 
wire w_mem_inst__abc_19396_new_n4373_; 
wire w_mem_inst__abc_19396_new_n4374_; 
wire w_mem_inst__abc_19396_new_n4376_; 
wire w_mem_inst__abc_19396_new_n4377_; 
wire w_mem_inst__abc_19396_new_n4378_; 
wire w_mem_inst__abc_19396_new_n4379_; 
wire w_mem_inst__abc_19396_new_n4381_; 
wire w_mem_inst__abc_19396_new_n4382_; 
wire w_mem_inst__abc_19396_new_n4383_; 
wire w_mem_inst__abc_19396_new_n4384_; 
wire w_mem_inst__abc_19396_new_n4386_; 
wire w_mem_inst__abc_19396_new_n4387_; 
wire w_mem_inst__abc_19396_new_n4388_; 
wire w_mem_inst__abc_19396_new_n4389_; 
wire w_mem_inst__abc_19396_new_n4391_; 
wire w_mem_inst__abc_19396_new_n4392_; 
wire w_mem_inst__abc_19396_new_n4393_; 
wire w_mem_inst__abc_19396_new_n4394_; 
wire w_mem_inst__abc_19396_new_n4396_; 
wire w_mem_inst__abc_19396_new_n4397_; 
wire w_mem_inst__abc_19396_new_n4398_; 
wire w_mem_inst__abc_19396_new_n4399_; 
wire w_mem_inst__abc_19396_new_n4401_; 
wire w_mem_inst__abc_19396_new_n4402_; 
wire w_mem_inst__abc_19396_new_n4403_; 
wire w_mem_inst__abc_19396_new_n4404_; 
wire w_mem_inst__abc_19396_new_n4406_; 
wire w_mem_inst__abc_19396_new_n4407_; 
wire w_mem_inst__abc_19396_new_n4408_; 
wire w_mem_inst__abc_19396_new_n4409_; 
wire w_mem_inst__abc_19396_new_n4411_; 
wire w_mem_inst__abc_19396_new_n4412_; 
wire w_mem_inst__abc_19396_new_n4413_; 
wire w_mem_inst__abc_19396_new_n4414_; 
wire w_mem_inst__abc_19396_new_n4416_; 
wire w_mem_inst__abc_19396_new_n4417_; 
wire w_mem_inst__abc_19396_new_n4418_; 
wire w_mem_inst__abc_19396_new_n4419_; 
wire w_mem_inst__abc_19396_new_n4421_; 
wire w_mem_inst__abc_19396_new_n4422_; 
wire w_mem_inst__abc_19396_new_n4423_; 
wire w_mem_inst__abc_19396_new_n4424_; 
wire w_mem_inst__abc_19396_new_n4426_; 
wire w_mem_inst__abc_19396_new_n4427_; 
wire w_mem_inst__abc_19396_new_n4428_; 
wire w_mem_inst__abc_19396_new_n4429_; 
wire w_mem_inst__abc_19396_new_n4431_; 
wire w_mem_inst__abc_19396_new_n4432_; 
wire w_mem_inst__abc_19396_new_n4433_; 
wire w_mem_inst__abc_19396_new_n4434_; 
wire w_mem_inst__abc_19396_new_n4436_; 
wire w_mem_inst__abc_19396_new_n4437_; 
wire w_mem_inst__abc_19396_new_n4438_; 
wire w_mem_inst__abc_19396_new_n4439_; 
wire w_mem_inst__abc_19396_new_n4441_; 
wire w_mem_inst__abc_19396_new_n4442_; 
wire w_mem_inst__abc_19396_new_n4443_; 
wire w_mem_inst__abc_19396_new_n4444_; 
wire w_mem_inst__abc_19396_new_n4446_; 
wire w_mem_inst__abc_19396_new_n4447_; 
wire w_mem_inst__abc_19396_new_n4448_; 
wire w_mem_inst__abc_19396_new_n4449_; 
wire w_mem_inst__abc_19396_new_n4451_; 
wire w_mem_inst__abc_19396_new_n4452_; 
wire w_mem_inst__abc_19396_new_n4453_; 
wire w_mem_inst__abc_19396_new_n4454_; 
wire w_mem_inst__abc_19396_new_n4456_; 
wire w_mem_inst__abc_19396_new_n4457_; 
wire w_mem_inst__abc_19396_new_n4458_; 
wire w_mem_inst__abc_19396_new_n4459_; 
wire w_mem_inst__abc_19396_new_n4461_; 
wire w_mem_inst__abc_19396_new_n4462_; 
wire w_mem_inst__abc_19396_new_n4463_; 
wire w_mem_inst__abc_19396_new_n4464_; 
wire w_mem_inst__abc_19396_new_n4466_; 
wire w_mem_inst__abc_19396_new_n4467_; 
wire w_mem_inst__abc_19396_new_n4468_; 
wire w_mem_inst__abc_19396_new_n4469_; 
wire w_mem_inst__abc_19396_new_n4471_; 
wire w_mem_inst__abc_19396_new_n4472_; 
wire w_mem_inst__abc_19396_new_n4473_; 
wire w_mem_inst__abc_19396_new_n4474_; 
wire w_mem_inst__abc_19396_new_n4476_; 
wire w_mem_inst__abc_19396_new_n4477_; 
wire w_mem_inst__abc_19396_new_n4478_; 
wire w_mem_inst__abc_19396_new_n4479_; 
wire w_mem_inst__abc_19396_new_n4481_; 
wire w_mem_inst__abc_19396_new_n4482_; 
wire w_mem_inst__abc_19396_new_n4483_; 
wire w_mem_inst__abc_19396_new_n4484_; 
wire w_mem_inst__abc_19396_new_n4486_; 
wire w_mem_inst__abc_19396_new_n4487_; 
wire w_mem_inst__abc_19396_new_n4488_; 
wire w_mem_inst__abc_19396_new_n4489_; 
wire w_mem_inst__abc_19396_new_n4491_; 
wire w_mem_inst__abc_19396_new_n4492_; 
wire w_mem_inst__abc_19396_new_n4493_; 
wire w_mem_inst__abc_19396_new_n4494_; 
wire w_mem_inst__abc_19396_new_n4496_; 
wire w_mem_inst__abc_19396_new_n4497_; 
wire w_mem_inst__abc_19396_new_n4498_; 
wire w_mem_inst__abc_19396_new_n4499_; 
wire w_mem_inst__abc_19396_new_n4501_; 
wire w_mem_inst__abc_19396_new_n4502_; 
wire w_mem_inst__abc_19396_new_n4503_; 
wire w_mem_inst__abc_19396_new_n4504_; 
wire w_mem_inst__abc_19396_new_n4506_; 
wire w_mem_inst__abc_19396_new_n4507_; 
wire w_mem_inst__abc_19396_new_n4508_; 
wire w_mem_inst__abc_19396_new_n4509_; 
wire w_mem_inst__abc_19396_new_n4511_; 
wire w_mem_inst__abc_19396_new_n4512_; 
wire w_mem_inst__abc_19396_new_n4513_; 
wire w_mem_inst__abc_19396_new_n4514_; 
wire w_mem_inst__abc_19396_new_n4516_; 
wire w_mem_inst__abc_19396_new_n4517_; 
wire w_mem_inst__abc_19396_new_n4518_; 
wire w_mem_inst__abc_19396_new_n4519_; 
wire w_mem_inst__abc_19396_new_n4521_; 
wire w_mem_inst__abc_19396_new_n4522_; 
wire w_mem_inst__abc_19396_new_n4523_; 
wire w_mem_inst__abc_19396_new_n4524_; 
wire w_mem_inst__abc_19396_new_n4526_; 
wire w_mem_inst__abc_19396_new_n4527_; 
wire w_mem_inst__abc_19396_new_n4528_; 
wire w_mem_inst__abc_19396_new_n4529_; 
wire w_mem_inst__abc_19396_new_n4531_; 
wire w_mem_inst__abc_19396_new_n4532_; 
wire w_mem_inst__abc_19396_new_n4533_; 
wire w_mem_inst__abc_19396_new_n4534_; 
wire w_mem_inst__abc_19396_new_n4536_; 
wire w_mem_inst__abc_19396_new_n4537_; 
wire w_mem_inst__abc_19396_new_n4538_; 
wire w_mem_inst__abc_19396_new_n4539_; 
wire w_mem_inst__abc_19396_new_n4541_; 
wire w_mem_inst__abc_19396_new_n4542_; 
wire w_mem_inst__abc_19396_new_n4543_; 
wire w_mem_inst__abc_19396_new_n4544_; 
wire w_mem_inst__abc_19396_new_n4546_; 
wire w_mem_inst__abc_19396_new_n4547_; 
wire w_mem_inst__abc_19396_new_n4548_; 
wire w_mem_inst__abc_19396_new_n4549_; 
wire w_mem_inst__abc_19396_new_n4551_; 
wire w_mem_inst__abc_19396_new_n4552_; 
wire w_mem_inst__abc_19396_new_n4553_; 
wire w_mem_inst__abc_19396_new_n4554_; 
wire w_mem_inst__abc_19396_new_n4556_; 
wire w_mem_inst__abc_19396_new_n4557_; 
wire w_mem_inst__abc_19396_new_n4558_; 
wire w_mem_inst__abc_19396_new_n4559_; 
wire w_mem_inst__abc_19396_new_n4561_; 
wire w_mem_inst__abc_19396_new_n4562_; 
wire w_mem_inst__abc_19396_new_n4563_; 
wire w_mem_inst__abc_19396_new_n4564_; 
wire w_mem_inst__abc_19396_new_n4566_; 
wire w_mem_inst__abc_19396_new_n4567_; 
wire w_mem_inst__abc_19396_new_n4568_; 
wire w_mem_inst__abc_19396_new_n4569_; 
wire w_mem_inst__abc_19396_new_n4571_; 
wire w_mem_inst__abc_19396_new_n4572_; 
wire w_mem_inst__abc_19396_new_n4573_; 
wire w_mem_inst__abc_19396_new_n4574_; 
wire w_mem_inst__abc_19396_new_n4576_; 
wire w_mem_inst__abc_19396_new_n4577_; 
wire w_mem_inst__abc_19396_new_n4578_; 
wire w_mem_inst__abc_19396_new_n4579_; 
wire w_mem_inst__abc_19396_new_n4581_; 
wire w_mem_inst__abc_19396_new_n4582_; 
wire w_mem_inst__abc_19396_new_n4583_; 
wire w_mem_inst__abc_19396_new_n4584_; 
wire w_mem_inst__abc_19396_new_n4586_; 
wire w_mem_inst__abc_19396_new_n4587_; 
wire w_mem_inst__abc_19396_new_n4588_; 
wire w_mem_inst__abc_19396_new_n4589_; 
wire w_mem_inst__abc_19396_new_n4591_; 
wire w_mem_inst__abc_19396_new_n4592_; 
wire w_mem_inst__abc_19396_new_n4593_; 
wire w_mem_inst__abc_19396_new_n4594_; 
wire w_mem_inst__abc_19396_new_n4596_; 
wire w_mem_inst__abc_19396_new_n4597_; 
wire w_mem_inst__abc_19396_new_n4598_; 
wire w_mem_inst__abc_19396_new_n4599_; 
wire w_mem_inst__abc_19396_new_n4601_; 
wire w_mem_inst__abc_19396_new_n4602_; 
wire w_mem_inst__abc_19396_new_n4603_; 
wire w_mem_inst__abc_19396_new_n4604_; 
wire w_mem_inst__abc_19396_new_n4606_; 
wire w_mem_inst__abc_19396_new_n4607_; 
wire w_mem_inst__abc_19396_new_n4608_; 
wire w_mem_inst__abc_19396_new_n4609_; 
wire w_mem_inst__abc_19396_new_n4611_; 
wire w_mem_inst__abc_19396_new_n4612_; 
wire w_mem_inst__abc_19396_new_n4613_; 
wire w_mem_inst__abc_19396_new_n4614_; 
wire w_mem_inst__abc_19396_new_n4616_; 
wire w_mem_inst__abc_19396_new_n4617_; 
wire w_mem_inst__abc_19396_new_n4618_; 
wire w_mem_inst__abc_19396_new_n4619_; 
wire w_mem_inst__abc_19396_new_n4621_; 
wire w_mem_inst__abc_19396_new_n4622_; 
wire w_mem_inst__abc_19396_new_n4623_; 
wire w_mem_inst__abc_19396_new_n4624_; 
wire w_mem_inst__abc_19396_new_n4626_; 
wire w_mem_inst__abc_19396_new_n4627_; 
wire w_mem_inst__abc_19396_new_n4628_; 
wire w_mem_inst__abc_19396_new_n4629_; 
wire w_mem_inst__abc_19396_new_n4631_; 
wire w_mem_inst__abc_19396_new_n4632_; 
wire w_mem_inst__abc_19396_new_n4633_; 
wire w_mem_inst__abc_19396_new_n4634_; 
wire w_mem_inst__abc_19396_new_n4636_; 
wire w_mem_inst__abc_19396_new_n4637_; 
wire w_mem_inst__abc_19396_new_n4638_; 
wire w_mem_inst__abc_19396_new_n4639_; 
wire w_mem_inst__abc_19396_new_n4641_; 
wire w_mem_inst__abc_19396_new_n4642_; 
wire w_mem_inst__abc_19396_new_n4643_; 
wire w_mem_inst__abc_19396_new_n4644_; 
wire w_mem_inst__abc_19396_new_n4646_; 
wire w_mem_inst__abc_19396_new_n4647_; 
wire w_mem_inst__abc_19396_new_n4648_; 
wire w_mem_inst__abc_19396_new_n4649_; 
wire w_mem_inst__abc_19396_new_n4651_; 
wire w_mem_inst__abc_19396_new_n4652_; 
wire w_mem_inst__abc_19396_new_n4653_; 
wire w_mem_inst__abc_19396_new_n4654_; 
wire w_mem_inst__abc_19396_new_n4656_; 
wire w_mem_inst__abc_19396_new_n4657_; 
wire w_mem_inst__abc_19396_new_n4658_; 
wire w_mem_inst__abc_19396_new_n4659_; 
wire w_mem_inst__abc_19396_new_n4661_; 
wire w_mem_inst__abc_19396_new_n4662_; 
wire w_mem_inst__abc_19396_new_n4663_; 
wire w_mem_inst__abc_19396_new_n4664_; 
wire w_mem_inst__abc_19396_new_n4666_; 
wire w_mem_inst__abc_19396_new_n4667_; 
wire w_mem_inst__abc_19396_new_n4668_; 
wire w_mem_inst__abc_19396_new_n4669_; 
wire w_mem_inst__abc_19396_new_n4671_; 
wire w_mem_inst__abc_19396_new_n4672_; 
wire w_mem_inst__abc_19396_new_n4673_; 
wire w_mem_inst__abc_19396_new_n4674_; 
wire w_mem_inst__abc_19396_new_n4676_; 
wire w_mem_inst__abc_19396_new_n4677_; 
wire w_mem_inst__abc_19396_new_n4678_; 
wire w_mem_inst__abc_19396_new_n4679_; 
wire w_mem_inst__abc_19396_new_n4681_; 
wire w_mem_inst__abc_19396_new_n4682_; 
wire w_mem_inst__abc_19396_new_n4683_; 
wire w_mem_inst__abc_19396_new_n4684_; 
wire w_mem_inst__abc_19396_new_n4686_; 
wire w_mem_inst__abc_19396_new_n4687_; 
wire w_mem_inst__abc_19396_new_n4688_; 
wire w_mem_inst__abc_19396_new_n4689_; 
wire w_mem_inst__abc_19396_new_n4691_; 
wire w_mem_inst__abc_19396_new_n4692_; 
wire w_mem_inst__abc_19396_new_n4693_; 
wire w_mem_inst__abc_19396_new_n4694_; 
wire w_mem_inst__abc_19396_new_n4696_; 
wire w_mem_inst__abc_19396_new_n4697_; 
wire w_mem_inst__abc_19396_new_n4698_; 
wire w_mem_inst__abc_19396_new_n4699_; 
wire w_mem_inst__abc_19396_new_n4701_; 
wire w_mem_inst__abc_19396_new_n4702_; 
wire w_mem_inst__abc_19396_new_n4703_; 
wire w_mem_inst__abc_19396_new_n4704_; 
wire w_mem_inst__abc_19396_new_n4706_; 
wire w_mem_inst__abc_19396_new_n4707_; 
wire w_mem_inst__abc_19396_new_n4708_; 
wire w_mem_inst__abc_19396_new_n4709_; 
wire w_mem_inst__abc_19396_new_n4711_; 
wire w_mem_inst__abc_19396_new_n4712_; 
wire w_mem_inst__abc_19396_new_n4713_; 
wire w_mem_inst__abc_19396_new_n4714_; 
wire w_mem_inst__abc_19396_new_n4716_; 
wire w_mem_inst__abc_19396_new_n4717_; 
wire w_mem_inst__abc_19396_new_n4718_; 
wire w_mem_inst__abc_19396_new_n4719_; 
wire w_mem_inst__abc_19396_new_n4721_; 
wire w_mem_inst__abc_19396_new_n4722_; 
wire w_mem_inst__abc_19396_new_n4723_; 
wire w_mem_inst__abc_19396_new_n4724_; 
wire w_mem_inst__abc_19396_new_n4726_; 
wire w_mem_inst__abc_19396_new_n4727_; 
wire w_mem_inst__abc_19396_new_n4728_; 
wire w_mem_inst__abc_19396_new_n4729_; 
wire w_mem_inst__abc_19396_new_n4731_; 
wire w_mem_inst__abc_19396_new_n4732_; 
wire w_mem_inst__abc_19396_new_n4733_; 
wire w_mem_inst__abc_19396_new_n4734_; 
wire w_mem_inst__abc_19396_new_n4736_; 
wire w_mem_inst__abc_19396_new_n4737_; 
wire w_mem_inst__abc_19396_new_n4738_; 
wire w_mem_inst__abc_19396_new_n4739_; 
wire w_mem_inst__abc_19396_new_n4741_; 
wire w_mem_inst__abc_19396_new_n4742_; 
wire w_mem_inst__abc_19396_new_n4743_; 
wire w_mem_inst__abc_19396_new_n4744_; 
wire w_mem_inst__abc_19396_new_n4746_; 
wire w_mem_inst__abc_19396_new_n4747_; 
wire w_mem_inst__abc_19396_new_n4748_; 
wire w_mem_inst__abc_19396_new_n4749_; 
wire w_mem_inst__abc_19396_new_n4751_; 
wire w_mem_inst__abc_19396_new_n4752_; 
wire w_mem_inst__abc_19396_new_n4753_; 
wire w_mem_inst__abc_19396_new_n4754_; 
wire w_mem_inst__abc_19396_new_n4756_; 
wire w_mem_inst__abc_19396_new_n4757_; 
wire w_mem_inst__abc_19396_new_n4758_; 
wire w_mem_inst__abc_19396_new_n4759_; 
wire w_mem_inst__abc_19396_new_n4761_; 
wire w_mem_inst__abc_19396_new_n4762_; 
wire w_mem_inst__abc_19396_new_n4763_; 
wire w_mem_inst__abc_19396_new_n4764_; 
wire w_mem_inst__abc_19396_new_n4766_; 
wire w_mem_inst__abc_19396_new_n4767_; 
wire w_mem_inst__abc_19396_new_n4768_; 
wire w_mem_inst__abc_19396_new_n4769_; 
wire w_mem_inst__abc_19396_new_n4771_; 
wire w_mem_inst__abc_19396_new_n4772_; 
wire w_mem_inst__abc_19396_new_n4773_; 
wire w_mem_inst__abc_19396_new_n4774_; 
wire w_mem_inst__abc_19396_new_n4776_; 
wire w_mem_inst__abc_19396_new_n4777_; 
wire w_mem_inst__abc_19396_new_n4778_; 
wire w_mem_inst__abc_19396_new_n4779_; 
wire w_mem_inst__abc_19396_new_n4781_; 
wire w_mem_inst__abc_19396_new_n4782_; 
wire w_mem_inst__abc_19396_new_n4783_; 
wire w_mem_inst__abc_19396_new_n4784_; 
wire w_mem_inst__abc_19396_new_n4786_; 
wire w_mem_inst__abc_19396_new_n4787_; 
wire w_mem_inst__abc_19396_new_n4788_; 
wire w_mem_inst__abc_19396_new_n4789_; 
wire w_mem_inst__abc_19396_new_n4791_; 
wire w_mem_inst__abc_19396_new_n4792_; 
wire w_mem_inst__abc_19396_new_n4794_; 
wire w_mem_inst__abc_19396_new_n4796_; 
wire w_mem_inst__abc_19396_new_n4797_; 
wire w_mem_inst__abc_19396_new_n4799_; 
wire w_mem_inst__abc_19396_new_n4800_; 
wire w_mem_inst__abc_19396_new_n4801_; 
wire w_mem_inst__abc_19396_new_n4803_; 
wire w_mem_inst__abc_19396_new_n4804_; 
wire w_mem_inst__abc_19396_new_n4805_; 
wire w_mem_inst__abc_19396_new_n4807_; 
wire w_mem_inst__abc_19396_new_n4808_; 
wire w_mem_inst__abc_19396_new_n4809_; 
wire w_mem_inst__abc_19396_new_n4811_; 
wire w_mem_inst_w_ctr_reg_0_; 
wire w_mem_inst_w_ctr_reg_1_; 
wire w_mem_inst_w_ctr_reg_2_; 
wire w_mem_inst_w_ctr_reg_3_; 
wire w_mem_inst_w_ctr_reg_4_; 
wire w_mem_inst_w_ctr_reg_5_; 
wire w_mem_inst_w_ctr_reg_6_; 
wire w_mem_inst_w_mem_0__0_; 
wire w_mem_inst_w_mem_0__10_; 
wire w_mem_inst_w_mem_0__11_; 
wire w_mem_inst_w_mem_0__12_; 
wire w_mem_inst_w_mem_0__13_; 
wire w_mem_inst_w_mem_0__14_; 
wire w_mem_inst_w_mem_0__15_; 
wire w_mem_inst_w_mem_0__16_; 
wire w_mem_inst_w_mem_0__17_; 
wire w_mem_inst_w_mem_0__18_; 
wire w_mem_inst_w_mem_0__19_; 
wire w_mem_inst_w_mem_0__1_; 
wire w_mem_inst_w_mem_0__20_; 
wire w_mem_inst_w_mem_0__21_; 
wire w_mem_inst_w_mem_0__22_; 
wire w_mem_inst_w_mem_0__23_; 
wire w_mem_inst_w_mem_0__24_; 
wire w_mem_inst_w_mem_0__25_; 
wire w_mem_inst_w_mem_0__26_; 
wire w_mem_inst_w_mem_0__27_; 
wire w_mem_inst_w_mem_0__28_; 
wire w_mem_inst_w_mem_0__29_; 
wire w_mem_inst_w_mem_0__2_; 
wire w_mem_inst_w_mem_0__30_; 
wire w_mem_inst_w_mem_0__31_; 
wire w_mem_inst_w_mem_0__3_; 
wire w_mem_inst_w_mem_0__4_; 
wire w_mem_inst_w_mem_0__5_; 
wire w_mem_inst_w_mem_0__6_; 
wire w_mem_inst_w_mem_0__7_; 
wire w_mem_inst_w_mem_0__8_; 
wire w_mem_inst_w_mem_0__9_; 
wire w_mem_inst_w_mem_10__0_; 
wire w_mem_inst_w_mem_10__10_; 
wire w_mem_inst_w_mem_10__11_; 
wire w_mem_inst_w_mem_10__12_; 
wire w_mem_inst_w_mem_10__13_; 
wire w_mem_inst_w_mem_10__14_; 
wire w_mem_inst_w_mem_10__15_; 
wire w_mem_inst_w_mem_10__16_; 
wire w_mem_inst_w_mem_10__17_; 
wire w_mem_inst_w_mem_10__18_; 
wire w_mem_inst_w_mem_10__19_; 
wire w_mem_inst_w_mem_10__1_; 
wire w_mem_inst_w_mem_10__20_; 
wire w_mem_inst_w_mem_10__21_; 
wire w_mem_inst_w_mem_10__22_; 
wire w_mem_inst_w_mem_10__23_; 
wire w_mem_inst_w_mem_10__24_; 
wire w_mem_inst_w_mem_10__25_; 
wire w_mem_inst_w_mem_10__26_; 
wire w_mem_inst_w_mem_10__27_; 
wire w_mem_inst_w_mem_10__28_; 
wire w_mem_inst_w_mem_10__29_; 
wire w_mem_inst_w_mem_10__2_; 
wire w_mem_inst_w_mem_10__30_; 
wire w_mem_inst_w_mem_10__31_; 
wire w_mem_inst_w_mem_10__3_; 
wire w_mem_inst_w_mem_10__4_; 
wire w_mem_inst_w_mem_10__5_; 
wire w_mem_inst_w_mem_10__6_; 
wire w_mem_inst_w_mem_10__7_; 
wire w_mem_inst_w_mem_10__8_; 
wire w_mem_inst_w_mem_10__9_; 
wire w_mem_inst_w_mem_11__0_; 
wire w_mem_inst_w_mem_11__10_; 
wire w_mem_inst_w_mem_11__11_; 
wire w_mem_inst_w_mem_11__12_; 
wire w_mem_inst_w_mem_11__13_; 
wire w_mem_inst_w_mem_11__14_; 
wire w_mem_inst_w_mem_11__15_; 
wire w_mem_inst_w_mem_11__16_; 
wire w_mem_inst_w_mem_11__17_; 
wire w_mem_inst_w_mem_11__18_; 
wire w_mem_inst_w_mem_11__19_; 
wire w_mem_inst_w_mem_11__1_; 
wire w_mem_inst_w_mem_11__20_; 
wire w_mem_inst_w_mem_11__21_; 
wire w_mem_inst_w_mem_11__22_; 
wire w_mem_inst_w_mem_11__23_; 
wire w_mem_inst_w_mem_11__24_; 
wire w_mem_inst_w_mem_11__25_; 
wire w_mem_inst_w_mem_11__26_; 
wire w_mem_inst_w_mem_11__27_; 
wire w_mem_inst_w_mem_11__28_; 
wire w_mem_inst_w_mem_11__29_; 
wire w_mem_inst_w_mem_11__2_; 
wire w_mem_inst_w_mem_11__30_; 
wire w_mem_inst_w_mem_11__31_; 
wire w_mem_inst_w_mem_11__3_; 
wire w_mem_inst_w_mem_11__4_; 
wire w_mem_inst_w_mem_11__5_; 
wire w_mem_inst_w_mem_11__6_; 
wire w_mem_inst_w_mem_11__7_; 
wire w_mem_inst_w_mem_11__8_; 
wire w_mem_inst_w_mem_11__9_; 
wire w_mem_inst_w_mem_12__0_; 
wire w_mem_inst_w_mem_12__10_; 
wire w_mem_inst_w_mem_12__11_; 
wire w_mem_inst_w_mem_12__12_; 
wire w_mem_inst_w_mem_12__13_; 
wire w_mem_inst_w_mem_12__14_; 
wire w_mem_inst_w_mem_12__15_; 
wire w_mem_inst_w_mem_12__16_; 
wire w_mem_inst_w_mem_12__17_; 
wire w_mem_inst_w_mem_12__18_; 
wire w_mem_inst_w_mem_12__19_; 
wire w_mem_inst_w_mem_12__1_; 
wire w_mem_inst_w_mem_12__20_; 
wire w_mem_inst_w_mem_12__21_; 
wire w_mem_inst_w_mem_12__22_; 
wire w_mem_inst_w_mem_12__23_; 
wire w_mem_inst_w_mem_12__24_; 
wire w_mem_inst_w_mem_12__25_; 
wire w_mem_inst_w_mem_12__26_; 
wire w_mem_inst_w_mem_12__27_; 
wire w_mem_inst_w_mem_12__28_; 
wire w_mem_inst_w_mem_12__29_; 
wire w_mem_inst_w_mem_12__2_; 
wire w_mem_inst_w_mem_12__30_; 
wire w_mem_inst_w_mem_12__31_; 
wire w_mem_inst_w_mem_12__3_; 
wire w_mem_inst_w_mem_12__4_; 
wire w_mem_inst_w_mem_12__5_; 
wire w_mem_inst_w_mem_12__6_; 
wire w_mem_inst_w_mem_12__7_; 
wire w_mem_inst_w_mem_12__8_; 
wire w_mem_inst_w_mem_12__9_; 
wire w_mem_inst_w_mem_13__0_; 
wire w_mem_inst_w_mem_13__10_; 
wire w_mem_inst_w_mem_13__11_; 
wire w_mem_inst_w_mem_13__12_; 
wire w_mem_inst_w_mem_13__13_; 
wire w_mem_inst_w_mem_13__14_; 
wire w_mem_inst_w_mem_13__15_; 
wire w_mem_inst_w_mem_13__16_; 
wire w_mem_inst_w_mem_13__17_; 
wire w_mem_inst_w_mem_13__18_; 
wire w_mem_inst_w_mem_13__19_; 
wire w_mem_inst_w_mem_13__1_; 
wire w_mem_inst_w_mem_13__20_; 
wire w_mem_inst_w_mem_13__21_; 
wire w_mem_inst_w_mem_13__22_; 
wire w_mem_inst_w_mem_13__23_; 
wire w_mem_inst_w_mem_13__24_; 
wire w_mem_inst_w_mem_13__25_; 
wire w_mem_inst_w_mem_13__26_; 
wire w_mem_inst_w_mem_13__27_; 
wire w_mem_inst_w_mem_13__28_; 
wire w_mem_inst_w_mem_13__29_; 
wire w_mem_inst_w_mem_13__2_; 
wire w_mem_inst_w_mem_13__30_; 
wire w_mem_inst_w_mem_13__31_; 
wire w_mem_inst_w_mem_13__3_; 
wire w_mem_inst_w_mem_13__4_; 
wire w_mem_inst_w_mem_13__5_; 
wire w_mem_inst_w_mem_13__6_; 
wire w_mem_inst_w_mem_13__7_; 
wire w_mem_inst_w_mem_13__8_; 
wire w_mem_inst_w_mem_13__9_; 
wire w_mem_inst_w_mem_14__0_; 
wire w_mem_inst_w_mem_14__10_; 
wire w_mem_inst_w_mem_14__11_; 
wire w_mem_inst_w_mem_14__12_; 
wire w_mem_inst_w_mem_14__13_; 
wire w_mem_inst_w_mem_14__14_; 
wire w_mem_inst_w_mem_14__15_; 
wire w_mem_inst_w_mem_14__16_; 
wire w_mem_inst_w_mem_14__17_; 
wire w_mem_inst_w_mem_14__18_; 
wire w_mem_inst_w_mem_14__19_; 
wire w_mem_inst_w_mem_14__1_; 
wire w_mem_inst_w_mem_14__20_; 
wire w_mem_inst_w_mem_14__21_; 
wire w_mem_inst_w_mem_14__22_; 
wire w_mem_inst_w_mem_14__23_; 
wire w_mem_inst_w_mem_14__24_; 
wire w_mem_inst_w_mem_14__25_; 
wire w_mem_inst_w_mem_14__26_; 
wire w_mem_inst_w_mem_14__27_; 
wire w_mem_inst_w_mem_14__28_; 
wire w_mem_inst_w_mem_14__29_; 
wire w_mem_inst_w_mem_14__2_; 
wire w_mem_inst_w_mem_14__30_; 
wire w_mem_inst_w_mem_14__31_; 
wire w_mem_inst_w_mem_14__3_; 
wire w_mem_inst_w_mem_14__4_; 
wire w_mem_inst_w_mem_14__5_; 
wire w_mem_inst_w_mem_14__6_; 
wire w_mem_inst_w_mem_14__7_; 
wire w_mem_inst_w_mem_14__8_; 
wire w_mem_inst_w_mem_14__9_; 
wire w_mem_inst_w_mem_15__0_; 
wire w_mem_inst_w_mem_15__10_; 
wire w_mem_inst_w_mem_15__11_; 
wire w_mem_inst_w_mem_15__12_; 
wire w_mem_inst_w_mem_15__13_; 
wire w_mem_inst_w_mem_15__14_; 
wire w_mem_inst_w_mem_15__15_; 
wire w_mem_inst_w_mem_15__16_; 
wire w_mem_inst_w_mem_15__17_; 
wire w_mem_inst_w_mem_15__18_; 
wire w_mem_inst_w_mem_15__19_; 
wire w_mem_inst_w_mem_15__1_; 
wire w_mem_inst_w_mem_15__20_; 
wire w_mem_inst_w_mem_15__21_; 
wire w_mem_inst_w_mem_15__22_; 
wire w_mem_inst_w_mem_15__23_; 
wire w_mem_inst_w_mem_15__24_; 
wire w_mem_inst_w_mem_15__25_; 
wire w_mem_inst_w_mem_15__26_; 
wire w_mem_inst_w_mem_15__27_; 
wire w_mem_inst_w_mem_15__28_; 
wire w_mem_inst_w_mem_15__29_; 
wire w_mem_inst_w_mem_15__2_; 
wire w_mem_inst_w_mem_15__30_; 
wire w_mem_inst_w_mem_15__31_; 
wire w_mem_inst_w_mem_15__3_; 
wire w_mem_inst_w_mem_15__4_; 
wire w_mem_inst_w_mem_15__5_; 
wire w_mem_inst_w_mem_15__6_; 
wire w_mem_inst_w_mem_15__7_; 
wire w_mem_inst_w_mem_15__8_; 
wire w_mem_inst_w_mem_15__9_; 
wire w_mem_inst_w_mem_1__0_; 
wire w_mem_inst_w_mem_1__10_; 
wire w_mem_inst_w_mem_1__11_; 
wire w_mem_inst_w_mem_1__12_; 
wire w_mem_inst_w_mem_1__13_; 
wire w_mem_inst_w_mem_1__14_; 
wire w_mem_inst_w_mem_1__15_; 
wire w_mem_inst_w_mem_1__16_; 
wire w_mem_inst_w_mem_1__17_; 
wire w_mem_inst_w_mem_1__18_; 
wire w_mem_inst_w_mem_1__19_; 
wire w_mem_inst_w_mem_1__1_; 
wire w_mem_inst_w_mem_1__20_; 
wire w_mem_inst_w_mem_1__21_; 
wire w_mem_inst_w_mem_1__22_; 
wire w_mem_inst_w_mem_1__23_; 
wire w_mem_inst_w_mem_1__24_; 
wire w_mem_inst_w_mem_1__25_; 
wire w_mem_inst_w_mem_1__26_; 
wire w_mem_inst_w_mem_1__27_; 
wire w_mem_inst_w_mem_1__28_; 
wire w_mem_inst_w_mem_1__29_; 
wire w_mem_inst_w_mem_1__2_; 
wire w_mem_inst_w_mem_1__30_; 
wire w_mem_inst_w_mem_1__31_; 
wire w_mem_inst_w_mem_1__3_; 
wire w_mem_inst_w_mem_1__4_; 
wire w_mem_inst_w_mem_1__5_; 
wire w_mem_inst_w_mem_1__6_; 
wire w_mem_inst_w_mem_1__7_; 
wire w_mem_inst_w_mem_1__8_; 
wire w_mem_inst_w_mem_1__9_; 
wire w_mem_inst_w_mem_2__0_; 
wire w_mem_inst_w_mem_2__10_; 
wire w_mem_inst_w_mem_2__11_; 
wire w_mem_inst_w_mem_2__12_; 
wire w_mem_inst_w_mem_2__13_; 
wire w_mem_inst_w_mem_2__14_; 
wire w_mem_inst_w_mem_2__15_; 
wire w_mem_inst_w_mem_2__16_; 
wire w_mem_inst_w_mem_2__17_; 
wire w_mem_inst_w_mem_2__18_; 
wire w_mem_inst_w_mem_2__19_; 
wire w_mem_inst_w_mem_2__1_; 
wire w_mem_inst_w_mem_2__20_; 
wire w_mem_inst_w_mem_2__21_; 
wire w_mem_inst_w_mem_2__22_; 
wire w_mem_inst_w_mem_2__23_; 
wire w_mem_inst_w_mem_2__24_; 
wire w_mem_inst_w_mem_2__25_; 
wire w_mem_inst_w_mem_2__26_; 
wire w_mem_inst_w_mem_2__27_; 
wire w_mem_inst_w_mem_2__28_; 
wire w_mem_inst_w_mem_2__29_; 
wire w_mem_inst_w_mem_2__2_; 
wire w_mem_inst_w_mem_2__30_; 
wire w_mem_inst_w_mem_2__31_; 
wire w_mem_inst_w_mem_2__3_; 
wire w_mem_inst_w_mem_2__4_; 
wire w_mem_inst_w_mem_2__5_; 
wire w_mem_inst_w_mem_2__6_; 
wire w_mem_inst_w_mem_2__7_; 
wire w_mem_inst_w_mem_2__8_; 
wire w_mem_inst_w_mem_2__9_; 
wire w_mem_inst_w_mem_3__0_; 
wire w_mem_inst_w_mem_3__10_; 
wire w_mem_inst_w_mem_3__11_; 
wire w_mem_inst_w_mem_3__12_; 
wire w_mem_inst_w_mem_3__13_; 
wire w_mem_inst_w_mem_3__14_; 
wire w_mem_inst_w_mem_3__15_; 
wire w_mem_inst_w_mem_3__16_; 
wire w_mem_inst_w_mem_3__17_; 
wire w_mem_inst_w_mem_3__18_; 
wire w_mem_inst_w_mem_3__19_; 
wire w_mem_inst_w_mem_3__1_; 
wire w_mem_inst_w_mem_3__20_; 
wire w_mem_inst_w_mem_3__21_; 
wire w_mem_inst_w_mem_3__22_; 
wire w_mem_inst_w_mem_3__23_; 
wire w_mem_inst_w_mem_3__24_; 
wire w_mem_inst_w_mem_3__25_; 
wire w_mem_inst_w_mem_3__26_; 
wire w_mem_inst_w_mem_3__27_; 
wire w_mem_inst_w_mem_3__28_; 
wire w_mem_inst_w_mem_3__29_; 
wire w_mem_inst_w_mem_3__2_; 
wire w_mem_inst_w_mem_3__30_; 
wire w_mem_inst_w_mem_3__31_; 
wire w_mem_inst_w_mem_3__3_; 
wire w_mem_inst_w_mem_3__4_; 
wire w_mem_inst_w_mem_3__5_; 
wire w_mem_inst_w_mem_3__6_; 
wire w_mem_inst_w_mem_3__7_; 
wire w_mem_inst_w_mem_3__8_; 
wire w_mem_inst_w_mem_3__9_; 
wire w_mem_inst_w_mem_4__0_; 
wire w_mem_inst_w_mem_4__10_; 
wire w_mem_inst_w_mem_4__11_; 
wire w_mem_inst_w_mem_4__12_; 
wire w_mem_inst_w_mem_4__13_; 
wire w_mem_inst_w_mem_4__14_; 
wire w_mem_inst_w_mem_4__15_; 
wire w_mem_inst_w_mem_4__16_; 
wire w_mem_inst_w_mem_4__17_; 
wire w_mem_inst_w_mem_4__18_; 
wire w_mem_inst_w_mem_4__19_; 
wire w_mem_inst_w_mem_4__1_; 
wire w_mem_inst_w_mem_4__20_; 
wire w_mem_inst_w_mem_4__21_; 
wire w_mem_inst_w_mem_4__22_; 
wire w_mem_inst_w_mem_4__23_; 
wire w_mem_inst_w_mem_4__24_; 
wire w_mem_inst_w_mem_4__25_; 
wire w_mem_inst_w_mem_4__26_; 
wire w_mem_inst_w_mem_4__27_; 
wire w_mem_inst_w_mem_4__28_; 
wire w_mem_inst_w_mem_4__29_; 
wire w_mem_inst_w_mem_4__2_; 
wire w_mem_inst_w_mem_4__30_; 
wire w_mem_inst_w_mem_4__31_; 
wire w_mem_inst_w_mem_4__3_; 
wire w_mem_inst_w_mem_4__4_; 
wire w_mem_inst_w_mem_4__5_; 
wire w_mem_inst_w_mem_4__6_; 
wire w_mem_inst_w_mem_4__7_; 
wire w_mem_inst_w_mem_4__8_; 
wire w_mem_inst_w_mem_4__9_; 
wire w_mem_inst_w_mem_5__0_; 
wire w_mem_inst_w_mem_5__10_; 
wire w_mem_inst_w_mem_5__11_; 
wire w_mem_inst_w_mem_5__12_; 
wire w_mem_inst_w_mem_5__13_; 
wire w_mem_inst_w_mem_5__14_; 
wire w_mem_inst_w_mem_5__15_; 
wire w_mem_inst_w_mem_5__16_; 
wire w_mem_inst_w_mem_5__17_; 
wire w_mem_inst_w_mem_5__18_; 
wire w_mem_inst_w_mem_5__19_; 
wire w_mem_inst_w_mem_5__1_; 
wire w_mem_inst_w_mem_5__20_; 
wire w_mem_inst_w_mem_5__21_; 
wire w_mem_inst_w_mem_5__22_; 
wire w_mem_inst_w_mem_5__23_; 
wire w_mem_inst_w_mem_5__24_; 
wire w_mem_inst_w_mem_5__25_; 
wire w_mem_inst_w_mem_5__26_; 
wire w_mem_inst_w_mem_5__27_; 
wire w_mem_inst_w_mem_5__28_; 
wire w_mem_inst_w_mem_5__29_; 
wire w_mem_inst_w_mem_5__2_; 
wire w_mem_inst_w_mem_5__30_; 
wire w_mem_inst_w_mem_5__31_; 
wire w_mem_inst_w_mem_5__3_; 
wire w_mem_inst_w_mem_5__4_; 
wire w_mem_inst_w_mem_5__5_; 
wire w_mem_inst_w_mem_5__6_; 
wire w_mem_inst_w_mem_5__7_; 
wire w_mem_inst_w_mem_5__8_; 
wire w_mem_inst_w_mem_5__9_; 
wire w_mem_inst_w_mem_6__0_; 
wire w_mem_inst_w_mem_6__10_; 
wire w_mem_inst_w_mem_6__11_; 
wire w_mem_inst_w_mem_6__12_; 
wire w_mem_inst_w_mem_6__13_; 
wire w_mem_inst_w_mem_6__14_; 
wire w_mem_inst_w_mem_6__15_; 
wire w_mem_inst_w_mem_6__16_; 
wire w_mem_inst_w_mem_6__17_; 
wire w_mem_inst_w_mem_6__18_; 
wire w_mem_inst_w_mem_6__19_; 
wire w_mem_inst_w_mem_6__1_; 
wire w_mem_inst_w_mem_6__20_; 
wire w_mem_inst_w_mem_6__21_; 
wire w_mem_inst_w_mem_6__22_; 
wire w_mem_inst_w_mem_6__23_; 
wire w_mem_inst_w_mem_6__24_; 
wire w_mem_inst_w_mem_6__25_; 
wire w_mem_inst_w_mem_6__26_; 
wire w_mem_inst_w_mem_6__27_; 
wire w_mem_inst_w_mem_6__28_; 
wire w_mem_inst_w_mem_6__29_; 
wire w_mem_inst_w_mem_6__2_; 
wire w_mem_inst_w_mem_6__30_; 
wire w_mem_inst_w_mem_6__31_; 
wire w_mem_inst_w_mem_6__3_; 
wire w_mem_inst_w_mem_6__4_; 
wire w_mem_inst_w_mem_6__5_; 
wire w_mem_inst_w_mem_6__6_; 
wire w_mem_inst_w_mem_6__7_; 
wire w_mem_inst_w_mem_6__8_; 
wire w_mem_inst_w_mem_6__9_; 
wire w_mem_inst_w_mem_7__0_; 
wire w_mem_inst_w_mem_7__10_; 
wire w_mem_inst_w_mem_7__11_; 
wire w_mem_inst_w_mem_7__12_; 
wire w_mem_inst_w_mem_7__13_; 
wire w_mem_inst_w_mem_7__14_; 
wire w_mem_inst_w_mem_7__15_; 
wire w_mem_inst_w_mem_7__16_; 
wire w_mem_inst_w_mem_7__17_; 
wire w_mem_inst_w_mem_7__18_; 
wire w_mem_inst_w_mem_7__19_; 
wire w_mem_inst_w_mem_7__1_; 
wire w_mem_inst_w_mem_7__20_; 
wire w_mem_inst_w_mem_7__21_; 
wire w_mem_inst_w_mem_7__22_; 
wire w_mem_inst_w_mem_7__23_; 
wire w_mem_inst_w_mem_7__24_; 
wire w_mem_inst_w_mem_7__25_; 
wire w_mem_inst_w_mem_7__26_; 
wire w_mem_inst_w_mem_7__27_; 
wire w_mem_inst_w_mem_7__28_; 
wire w_mem_inst_w_mem_7__29_; 
wire w_mem_inst_w_mem_7__2_; 
wire w_mem_inst_w_mem_7__30_; 
wire w_mem_inst_w_mem_7__31_; 
wire w_mem_inst_w_mem_7__3_; 
wire w_mem_inst_w_mem_7__4_; 
wire w_mem_inst_w_mem_7__5_; 
wire w_mem_inst_w_mem_7__6_; 
wire w_mem_inst_w_mem_7__7_; 
wire w_mem_inst_w_mem_7__8_; 
wire w_mem_inst_w_mem_7__9_; 
wire w_mem_inst_w_mem_8__0_; 
wire w_mem_inst_w_mem_8__10_; 
wire w_mem_inst_w_mem_8__11_; 
wire w_mem_inst_w_mem_8__12_; 
wire w_mem_inst_w_mem_8__13_; 
wire w_mem_inst_w_mem_8__14_; 
wire w_mem_inst_w_mem_8__15_; 
wire w_mem_inst_w_mem_8__16_; 
wire w_mem_inst_w_mem_8__17_; 
wire w_mem_inst_w_mem_8__18_; 
wire w_mem_inst_w_mem_8__19_; 
wire w_mem_inst_w_mem_8__1_; 
wire w_mem_inst_w_mem_8__20_; 
wire w_mem_inst_w_mem_8__21_; 
wire w_mem_inst_w_mem_8__22_; 
wire w_mem_inst_w_mem_8__23_; 
wire w_mem_inst_w_mem_8__24_; 
wire w_mem_inst_w_mem_8__25_; 
wire w_mem_inst_w_mem_8__26_; 
wire w_mem_inst_w_mem_8__27_; 
wire w_mem_inst_w_mem_8__28_; 
wire w_mem_inst_w_mem_8__29_; 
wire w_mem_inst_w_mem_8__2_; 
wire w_mem_inst_w_mem_8__30_; 
wire w_mem_inst_w_mem_8__31_; 
wire w_mem_inst_w_mem_8__3_; 
wire w_mem_inst_w_mem_8__4_; 
wire w_mem_inst_w_mem_8__5_; 
wire w_mem_inst_w_mem_8__6_; 
wire w_mem_inst_w_mem_8__7_; 
wire w_mem_inst_w_mem_8__8_; 
wire w_mem_inst_w_mem_8__9_; 
wire w_mem_inst_w_mem_9__0_; 
wire w_mem_inst_w_mem_9__10_; 
wire w_mem_inst_w_mem_9__11_; 
wire w_mem_inst_w_mem_9__12_; 
wire w_mem_inst_w_mem_9__13_; 
wire w_mem_inst_w_mem_9__14_; 
wire w_mem_inst_w_mem_9__15_; 
wire w_mem_inst_w_mem_9__16_; 
wire w_mem_inst_w_mem_9__17_; 
wire w_mem_inst_w_mem_9__18_; 
wire w_mem_inst_w_mem_9__19_; 
wire w_mem_inst_w_mem_9__1_; 
wire w_mem_inst_w_mem_9__20_; 
wire w_mem_inst_w_mem_9__21_; 
wire w_mem_inst_w_mem_9__22_; 
wire w_mem_inst_w_mem_9__23_; 
wire w_mem_inst_w_mem_9__24_; 
wire w_mem_inst_w_mem_9__25_; 
wire w_mem_inst_w_mem_9__26_; 
wire w_mem_inst_w_mem_9__27_; 
wire w_mem_inst_w_mem_9__28_; 
wire w_mem_inst_w_mem_9__29_; 
wire w_mem_inst_w_mem_9__2_; 
wire w_mem_inst_w_mem_9__30_; 
wire w_mem_inst_w_mem_9__31_; 
wire w_mem_inst_w_mem_9__3_; 
wire w_mem_inst_w_mem_9__4_; 
wire w_mem_inst_w_mem_9__5_; 
wire w_mem_inst_w_mem_9__6_; 
wire w_mem_inst_w_mem_9__7_; 
wire w_mem_inst_w_mem_9__8_; 
wire w_mem_inst_w_mem_9__9_; 
AND2X2 AND2X2_1 ( .A(c_reg_15_), .B(_auto_iopadmap_cc_368_execute_22625_79_), .Y(_abc_15497_new_n699_));
AND2X2 AND2X2_10 ( .A(c_reg_17_), .B(_auto_iopadmap_cc_368_execute_22625_81_), .Y(_abc_15497_new_n829_));
AND2X2 AND2X2_100 ( .A(_abc_15497_new_n3712_), .B(_abc_15497_new_n3710_), .Y(_abc_15497_new_n3713_));
AND2X2 AND2X2_101 ( .A(_abc_15497_new_n3717_), .B(_abc_15497_new_n3718_), .Y(_abc_15497_new_n3719_));
AND2X2 AND2X2_102 ( .A(_abc_15497_new_n3695_), .B(_abc_15497_new_n3694_), .Y(_abc_15497_new_n3723_));
AND2X2 AND2X2_103 ( .A(_abc_15497_new_n3743_), .B(_abc_15497_new_n3741_), .Y(_abc_15497_new_n3744_));
AND2X2 AND2X2_104 ( .A(_abc_15497_new_n3745_), .B(_abc_15497_new_n3748_), .Y(_abc_15497_new_n3749_));
AND2X2 AND2X2_105 ( .A(_abc_15497_new_n3808_), .B(_abc_15497_new_n3803_), .Y(_abc_15497_new_n3809_));
AND2X2 AND2X2_106 ( .A(_abc_15497_new_n3781_), .B(_abc_15497_new_n3819_), .Y(_abc_15497_new_n3820_));
AND2X2 AND2X2_107 ( .A(_abc_15497_new_n3826_), .B(_abc_15497_new_n3864_), .Y(_abc_15497_new_n3865_));
AND2X2 AND2X2_108 ( .A(_abc_15497_new_n3894_), .B(c_reg_20_), .Y(_abc_15497_new_n3895_));
AND2X2 AND2X2_109 ( .A(_abc_15497_new_n3944_), .B(c_reg_21_), .Y(_abc_15497_new_n3945_));
AND2X2 AND2X2_11 ( .A(_abc_15497_new_n819_), .B(_abc_15497_new_n846_), .Y(_abc_15497_new_n847_));
AND2X2 AND2X2_110 ( .A(_abc_15497_new_n3936_), .B(_abc_15497_new_n3980_), .Y(_abc_15497_new_n3981_));
AND2X2 AND2X2_111 ( .A(_abc_15497_new_n3987_), .B(_abc_15497_new_n3990_), .Y(_abc_15497_new_n3991_));
AND2X2 AND2X2_112 ( .A(_abc_15497_new_n3999_), .B(c_reg_22_), .Y(_abc_15497_new_n4000_));
AND2X2 AND2X2_113 ( .A(_abc_15497_new_n3991_), .B(_abc_15497_new_n4035_), .Y(_abc_15497_new_n4036_));
AND2X2 AND2X2_114 ( .A(_abc_15497_new_n4043_), .B(_abc_15497_new_n4090_), .Y(_abc_15497_new_n4091_));
AND2X2 AND2X2_115 ( .A(_abc_15497_new_n4097_), .B(_abc_15497_new_n3986_), .Y(_abc_15497_new_n4098_));
AND2X2 AND2X2_116 ( .A(_abc_15497_new_n4145_), .B(_abc_15497_new_n4146_), .Y(_abc_15497_new_n4147_));
AND2X2 AND2X2_117 ( .A(_abc_15497_new_n4177_), .B(_abc_15497_new_n4178_), .Y(_abc_15497_new_n4182_));
AND2X2 AND2X2_118 ( .A(_abc_15497_new_n4201_), .B(_abc_15497_new_n4195_), .Y(_abc_15497_new_n4202_));
AND2X2 AND2X2_119 ( .A(_abc_15497_new_n4215_), .B(_abc_15497_new_n4193_), .Y(_abc_15497_new_n4217_));
AND2X2 AND2X2_12 ( .A(_abc_15497_new_n868_), .B(_abc_15497_new_n881_), .Y(_abc_15497_new_n886_));
AND2X2 AND2X2_120 ( .A(_abc_15497_new_n4218_), .B(_abc_15497_new_n3678_), .Y(_abc_15497_new_n4219_));
AND2X2 AND2X2_121 ( .A(_abc_15497_new_n4227_), .B(_abc_15497_new_n4228_), .Y(_abc_15497_new_n4229_));
AND2X2 AND2X2_122 ( .A(_abc_15497_new_n4235_), .B(_abc_15497_new_n4260_), .Y(_abc_15497_new_n4262_));
AND2X2 AND2X2_123 ( .A(_abc_15497_new_n4233_), .B(_abc_15497_new_n4263_), .Y(_abc_15497_new_n4264_));
AND2X2 AND2X2_124 ( .A(_abc_15497_new_n4301_), .B(_abc_15497_new_n4277_), .Y(_abc_15497_new_n4303_));
AND2X2 AND2X2_125 ( .A(_abc_15497_new_n4358_), .B(_abc_15497_new_n4357_), .Y(_abc_15497_new_n4359_));
AND2X2 AND2X2_126 ( .A(_abc_15497_new_n4325_), .B(_abc_15497_new_n4359_), .Y(_abc_15497_new_n4360_));
AND2X2 AND2X2_127 ( .A(_abc_15497_new_n4391_), .B(_abc_15497_new_n4392_), .Y(_abc_15497_new_n4393_));
AND2X2 AND2X2_128 ( .A(_abc_15497_new_n4359_), .B(_abc_15497_new_n4318_), .Y(_abc_15497_new_n4407_));
AND2X2 AND2X2_129 ( .A(c_reg_31_), .B(b_reg_31_), .Y(_abc_15497_new_n4418_));
AND2X2 AND2X2_13 ( .A(_abc_15497_new_n902_), .B(_abc_15497_new_n907_), .Y(_abc_15497_new_n908_));
AND2X2 AND2X2_130 ( .A(_abc_15497_new_n781_), .B(_abc_15497_new_n4493_), .Y(_abc_15497_new_n4494_));
AND2X2 AND2X2_131 ( .A(_abc_15497_new_n4515_), .B(_abc_15497_new_n784_), .Y(_abc_15497_new_n4516_));
AND2X2 AND2X2_132 ( .A(_abc_15497_new_n4535_), .B(_abc_15497_new_n718_), .Y(_abc_15497_new_n4536_));
AND2X2 AND2X2_133 ( .A(_abc_15497_new_n792_), .B(_abc_15497_new_n846_), .Y(_abc_15497_new_n4564_));
AND2X2 AND2X2_134 ( .A(_abc_15497_new_n4571_), .B(_abc_15497_new_n809_), .Y(_abc_15497_new_n4572_));
AND2X2 AND2X2_135 ( .A(_abc_15497_new_n848_), .B(_abc_15497_new_n860_), .Y(_abc_15497_new_n4588_));
AND2X2 AND2X2_136 ( .A(_abc_15497_new_n4592_), .B(_abc_15497_new_n854_), .Y(_abc_15497_new_n4593_));
AND2X2 AND2X2_137 ( .A(w_mem_inst__abc_19396_new_n1619__bF_buf4), .B(w_mem_inst__abc_19396_new_n1620__bF_buf7), .Y(w_mem_inst__abc_19396_new_n1621_));
AND2X2 AND2X2_138 ( .A(w_mem_inst__abc_19396_new_n4800_), .B(w_mem_inst__abc_19396_new_n4801_), .Y(w_mem_inst__0w_ctr_reg_6_0__3_));
AND2X2 AND2X2_139 ( .A(w_mem_inst__abc_19396_new_n4805_), .B(w_mem_inst_w_ctr_reg_5_), .Y(w_mem_inst__abc_19396_new_n4809_));
AND2X2 AND2X2_14 ( .A(_abc_15497_new_n906_), .B(_abc_15497_new_n896_), .Y(_abc_15497_new_n918_));
AND2X2 AND2X2_15 ( .A(_abc_15497_new_n892_), .B(_abc_15497_new_n918_), .Y(_abc_15497_new_n927_));
AND2X2 AND2X2_16 ( .A(e_reg_5_), .B(_auto_iopadmap_cc_368_execute_22625_5_), .Y(_abc_15497_new_n978_));
AND2X2 AND2X2_17 ( .A(_abc_15497_new_n976_), .B(_abc_15497_new_n979_), .Y(_abc_15497_new_n980_));
AND2X2 AND2X2_18 ( .A(_abc_15497_new_n985_), .B(_abc_15497_new_n986_), .Y(_abc_15497_new_n987_));
AND2X2 AND2X2_19 ( .A(e_reg_6_), .B(_auto_iopadmap_cc_368_execute_22625_6_), .Y(_abc_15497_new_n991_));
AND2X2 AND2X2_2 ( .A(c_reg_12_), .B(_auto_iopadmap_cc_368_execute_22625_76_), .Y(_abc_15497_new_n711_));
AND2X2 AND2X2_20 ( .A(_abc_15497_new_n1138_), .B(_abc_15497_new_n1133_), .Y(_abc_15497_new_n1139_));
AND2X2 AND2X2_21 ( .A(_abc_15497_new_n1110_), .B(_abc_15497_new_n1157_), .Y(_abc_15497_new_n1158_));
AND2X2 AND2X2_22 ( .A(_abc_15497_new_n1183_), .B(_abc_15497_new_n1188_), .Y(_abc_15497_new_n1189_));
AND2X2 AND2X2_23 ( .A(_abc_15497_new_n1237_), .B(_abc_15497_new_n1259_), .Y(_abc_15497_new_n1260_));
AND2X2 AND2X2_24 ( .A(_abc_15497_new_n1266_), .B(_abc_15497_new_n1270_), .Y(_abc_15497_new_n1271_));
AND2X2 AND2X2_25 ( .A(_abc_15497_new_n1276_), .B(_abc_15497_new_n1264_), .Y(_abc_15497_new_n1284_));
AND2X2 AND2X2_26 ( .A(_abc_15497_new_n1285_), .B(_abc_15497_new_n1281_), .Y(_abc_15497_new_n1286_));
AND2X2 AND2X2_27 ( .A(_abc_15497_new_n1291_), .B(_abc_15497_new_n1292_), .Y(_abc_15497_new_n1294_));
AND2X2 AND2X2_28 ( .A(_auto_iopadmap_cc_368_execute_22625_34_), .B(d_reg_2_), .Y(_abc_15497_new_n1312_));
AND2X2 AND2X2_29 ( .A(_abc_15497_new_n1318_), .B(_abc_15497_new_n1322_), .Y(_abc_15497_new_n1323_));
AND2X2 AND2X2_3 ( .A(c_reg_11_), .B(_auto_iopadmap_cc_368_execute_22625_75_), .Y(_abc_15497_new_n726_));
AND2X2 AND2X2_30 ( .A(_abc_15497_new_n1362_), .B(_abc_15497_new_n1367_), .Y(_abc_15497_new_n1368_));
AND2X2 AND2X2_31 ( .A(_abc_15497_new_n1385_), .B(_abc_15497_new_n1389_), .Y(_abc_15497_new_n1390_));
AND2X2 AND2X2_32 ( .A(_abc_15497_new_n1396_), .B(_abc_15497_new_n1401_), .Y(_abc_15497_new_n1402_));
AND2X2 AND2X2_33 ( .A(_abc_15497_new_n1434_), .B(_abc_15497_new_n1439_), .Y(_abc_15497_new_n1440_));
AND2X2 AND2X2_34 ( .A(_abc_15497_new_n1467_), .B(_abc_15497_new_n1471_), .Y(_abc_15497_new_n1472_));
AND2X2 AND2X2_35 ( .A(_abc_15497_new_n1493_), .B(_abc_15497_new_n1498_), .Y(_abc_15497_new_n1499_));
AND2X2 AND2X2_36 ( .A(_abc_15497_new_n1536_), .B(_abc_15497_new_n1533_), .Y(_abc_15497_new_n1537_));
AND2X2 AND2X2_37 ( .A(_abc_15497_new_n1542_), .B(_abc_15497_new_n1546_), .Y(_abc_15497_new_n1547_));
AND2X2 AND2X2_38 ( .A(_abc_15497_new_n1584_), .B(_abc_15497_new_n1589_), .Y(_abc_15497_new_n1590_));
AND2X2 AND2X2_39 ( .A(_abc_15497_new_n1613_), .B(_abc_15497_new_n1618_), .Y(_abc_15497_new_n1619_));
AND2X2 AND2X2_4 ( .A(c_reg_7_), .B(_auto_iopadmap_cc_368_execute_22625_71_), .Y(_abc_15497_new_n747_));
AND2X2 AND2X2_40 ( .A(_abc_15497_new_n1624_), .B(_abc_15497_new_n1611_), .Y(_abc_15497_new_n1633_));
AND2X2 AND2X2_41 ( .A(_abc_15497_new_n1639_), .B(_abc_15497_new_n1640_), .Y(_abc_15497_new_n1641_));
AND2X2 AND2X2_42 ( .A(_auto_iopadmap_cc_368_execute_22625_99_), .B(b_reg_3_), .Y(_abc_15497_new_n1774_));
AND2X2 AND2X2_43 ( .A(_auto_iopadmap_cc_368_execute_22625_105_), .B(b_reg_9_), .Y(_abc_15497_new_n1831_));
AND2X2 AND2X2_44 ( .A(_abc_15497_new_n1885_), .B(_abc_15497_new_n1883_), .Y(_abc_15497_new_n1886_));
AND2X2 AND2X2_45 ( .A(_abc_15497_new_n1886_), .B(_abc_15497_new_n1879_), .Y(_abc_15497_new_n1887_));
AND2X2 AND2X2_46 ( .A(_abc_15497_new_n1956_), .B(_abc_15497_new_n1961_), .Y(_abc_15497_new_n1962_));
AND2X2 AND2X2_47 ( .A(_abc_15497_new_n1995_), .B(_abc_15497_new_n1955_), .Y(_abc_15497_new_n2002_));
AND2X2 AND2X2_48 ( .A(_abc_15497_new_n2003_), .B(_abc_15497_new_n2009_), .Y(_abc_15497_new_n2010_));
AND2X2 AND2X2_49 ( .A(_abc_15497_new_n2033_), .B(_abc_15497_new_n2043_), .Y(_abc_15497_new_n2048_));
AND2X2 AND2X2_5 ( .A(c_reg_2_), .B(_auto_iopadmap_cc_368_execute_22625_66_), .Y(_abc_15497_new_n767_));
AND2X2 AND2X2_50 ( .A(_abc_15497_new_n2193_), .B(_abc_15497_new_n2185_), .Y(_abc_15497_new_n2194_));
AND2X2 AND2X2_51 ( .A(_auto_iopadmap_cc_368_execute_22625_141_), .B(a_reg_13_), .Y(_abc_15497_new_n2223_));
AND2X2 AND2X2_52 ( .A(_abc_15497_new_n2281_), .B(_abc_15497_new_n2286_), .Y(_abc_15497_new_n2287_));
AND2X2 AND2X2_53 ( .A(_abc_15497_new_n2294_), .B(_abc_15497_new_n2299_), .Y(_abc_15497_new_n2300_));
AND2X2 AND2X2_54 ( .A(_abc_15497_new_n2308_), .B(_abc_15497_new_n2313_), .Y(_abc_15497_new_n2314_));
AND2X2 AND2X2_55 ( .A(_abc_15497_new_n2338_), .B(_abc_15497_new_n2339_), .Y(_abc_15497_new_n2340_));
AND2X2 AND2X2_56 ( .A(_abc_15497_new_n2357_), .B(_abc_15497_new_n2363_), .Y(_abc_15497_new_n2364_));
AND2X2 AND2X2_57 ( .A(_abc_15497_new_n2387_), .B(_abc_15497_new_n2397_), .Y(_abc_15497_new_n2402_));
AND2X2 AND2X2_58 ( .A(_abc_15497_new_n2415_), .B(_abc_15497_new_n2420_), .Y(_abc_15497_new_n2421_));
AND2X2 AND2X2_59 ( .A(_abc_15497_new_n2420_), .B(_abc_15497_new_n2409_), .Y(_abc_15497_new_n2432_));
AND2X2 AND2X2_6 ( .A(_abc_15497_new_n780_), .B(_abc_15497_new_n764_), .Y(_abc_15497_new_n781_));
AND2X2 AND2X2_60 ( .A(_abc_15497_new_n2433_), .B(_abc_15497_new_n2429_), .Y(_abc_15497_new_n2434_));
AND2X2 AND2X2_61 ( .A(_abc_15497_new_n2439_), .B(_abc_15497_new_n2440_), .Y(_abc_15497_new_n2441_));
AND2X2 AND2X2_62 ( .A(_abc_15497_new_n2741_), .B(_abc_15497_new_n2740_), .Y(_abc_15497_new_n2751_));
AND2X2 AND2X2_63 ( .A(_abc_15497_new_n2776_), .B(_abc_15497_new_n2777_), .Y(_abc_15497_new_n2778_));
AND2X2 AND2X2_64 ( .A(_abc_15497_new_n2787_), .B(_abc_15497_new_n2789_), .Y(_abc_15497_new_n2806_));
AND2X2 AND2X2_65 ( .A(_abc_15497_new_n2803_), .B(_abc_15497_new_n2799_), .Y(_abc_15497_new_n2807_));
AND2X2 AND2X2_66 ( .A(_abc_15497_new_n2850_), .B(_abc_15497_new_n2847_), .Y(_abc_15497_new_n2851_));
AND2X2 AND2X2_67 ( .A(_abc_15497_new_n2835_), .B(_abc_15497_new_n2837_), .Y(_abc_15497_new_n2853_));
AND2X2 AND2X2_68 ( .A(_abc_15497_new_n2894_), .B(_abc_15497_new_n2896_), .Y(_abc_15497_new_n2912_));
AND2X2 AND2X2_69 ( .A(_abc_15497_new_n2968_), .B(_abc_15497_new_n2964_), .Y(_abc_15497_new_n2971_));
AND2X2 AND2X2_7 ( .A(c_reg_21_), .B(_auto_iopadmap_cc_368_execute_22625_85_), .Y(_abc_15497_new_n806_));
AND2X2 AND2X2_70 ( .A(_abc_15497_new_n2950_), .B(_abc_15497_new_n2947_), .Y(_abc_15497_new_n2976_));
AND2X2 AND2X2_71 ( .A(_abc_15497_new_n2993_), .B(_abc_15497_new_n2989_), .Y(_abc_15497_new_n2994_));
AND2X2 AND2X2_72 ( .A(_abc_15497_new_n3002_), .B(_abc_15497_new_n2993_), .Y(_abc_15497_new_n3003_));
AND2X2 AND2X2_73 ( .A(_abc_15497_new_n3029_), .B(_abc_15497_new_n3025_), .Y(_abc_15497_new_n3030_));
AND2X2 AND2X2_74 ( .A(_abc_15497_new_n3013_), .B(_abc_15497_new_n3015_), .Y(_abc_15497_new_n3032_));
AND2X2 AND2X2_75 ( .A(_abc_15497_new_n3003_), .B(_abc_15497_new_n3052_), .Y(_abc_15497_new_n3053_));
AND2X2 AND2X2_76 ( .A(_abc_15497_new_n3087_), .B(_abc_15497_new_n3083_), .Y(_abc_15497_new_n3088_));
AND2X2 AND2X2_77 ( .A(_abc_15497_new_n3071_), .B(_abc_15497_new_n3073_), .Y(_abc_15497_new_n3090_));
AND2X2 AND2X2_78 ( .A(_abc_15497_new_n3152_), .B(_abc_15497_new_n3157_), .Y(_abc_15497_new_n3158_));
AND2X2 AND2X2_79 ( .A(_abc_15497_new_n3175_), .B(_abc_15497_new_n3177_), .Y(_abc_15497_new_n3199_));
AND2X2 AND2X2_8 ( .A(c_reg_20_), .B(_auto_iopadmap_cc_368_execute_22625_84_), .Y(_abc_15497_new_n807_));
AND2X2 AND2X2_80 ( .A(_abc_15497_new_n3051_), .B(_abc_15497_new_n3045_), .Y(_abc_15497_new_n3212_));
AND2X2 AND2X2_81 ( .A(_abc_15497_new_n3217_), .B(_abc_15497_new_n3211_), .Y(_abc_15497_new_n3218_));
AND2X2 AND2X2_82 ( .A(_abc_15497_new_n3220_), .B(_abc_15497_new_n3221_), .Y(_abc_15497_new_n3222_));
AND2X2 AND2X2_83 ( .A(b_reg_9_), .B(c_reg_9_), .Y(_abc_15497_new_n3231_));
AND2X2 AND2X2_84 ( .A(_abc_15497_new_n3278_), .B(_abc_15497_new_n3274_), .Y(_abc_15497_new_n3279_));
AND2X2 AND2X2_85 ( .A(_abc_15497_new_n3287_), .B(_abc_15497_new_n3342_), .Y(_abc_15497_new_n3343_));
AND2X2 AND2X2_86 ( .A(e_reg_11_), .B(a_reg_6_), .Y(_abc_15497_new_n3363_));
AND2X2 AND2X2_87 ( .A(round_ctr_reg_3_), .B(round_ctr_reg_2_), .Y(_abc_15497_new_n3392_));
AND2X2 AND2X2_88 ( .A(_abc_15497_new_n3396_), .B(_abc_15497_new_n3390_), .Y(_abc_15497_new_n3397_));
AND2X2 AND2X2_89 ( .A(_abc_15497_new_n3349_), .B(_abc_15497_new_n3397_), .Y(_abc_15497_new_n3398_));
AND2X2 AND2X2_9 ( .A(c_reg_19_), .B(_auto_iopadmap_cc_368_execute_22625_83_), .Y(_abc_15497_new_n820_));
AND2X2 AND2X2_90 ( .A(b_reg_12_), .B(c_reg_12_), .Y(_abc_15497_new_n3422_));
AND2X2 AND2X2_91 ( .A(_abc_15497_new_n3470_), .B(_abc_15497_new_n3463_), .Y(_abc_15497_new_n3471_));
AND2X2 AND2X2_92 ( .A(b_reg_13_), .B(c_reg_13_), .Y(_abc_15497_new_n3482_));
AND2X2 AND2X2_93 ( .A(e_reg_13_), .B(a_reg_8_), .Y(_abc_15497_new_n3496_));
AND2X2 AND2X2_94 ( .A(_abc_15497_new_n3486_), .B(_abc_15497_new_n3483_), .Y(_abc_15497_new_n3506_));
AND2X2 AND2X2_95 ( .A(b_reg_14_), .B(c_reg_14_), .Y(_abc_15497_new_n3545_));
AND2X2 AND2X2_96 ( .A(e_reg_14_), .B(a_reg_9_), .Y(_abc_15497_new_n3561_));
AND2X2 AND2X2_97 ( .A(_abc_15497_new_n3549_), .B(_abc_15497_new_n3546_), .Y(_abc_15497_new_n3572_));
AND2X2 AND2X2_98 ( .A(b_reg_15_), .B(c_reg_15_), .Y(_abc_15497_new_n3607_));
AND2X2 AND2X2_99 ( .A(_abc_15497_new_n3682_), .B(c_reg_16_), .Y(_abc_15497_new_n3683_));
AOI21X1 AOI21X1_1 ( .A(_abc_15497_new_n713_), .B(_abc_15497_new_n711_), .C(_abc_15497_new_n710_), .Y(_abc_15497_new_n714_));
AOI21X1 AOI21X1_10 ( .A(_abc_15497_new_n796_), .B(_abc_15497_new_n800_), .C(_abc_15497_new_n795_), .Y(_abc_15497_new_n811_));
AOI21X1 AOI21X1_100 ( .A(_abc_15497_new_n1308_), .B(_abc_15497_new_n2783_), .C(_abc_15497_new_n2782_), .Y(_abc_15497_new_n2784_));
AOI21X1 AOI21X1_101 ( .A(_abc_15497_new_n2797_), .B(_abc_15497_new_n2794_), .C(w_1_), .Y(_abc_15497_new_n2801_));
AOI21X1 AOI21X1_102 ( .A(_abc_15497_new_n2808_), .B(_abc_15497_new_n2805_), .C(_abc_15497_new_n2771_), .Y(_abc_15497_new_n2809_));
AOI21X1 AOI21X1_103 ( .A(_abc_15497_new_n2811_), .B(_abc_15497_new_n2810_), .C(_abc_15497_new_n2771_), .Y(_abc_15497_new_n2814_));
AOI21X1 AOI21X1_104 ( .A(_abc_15497_new_n2826_), .B(_abc_15497_new_n2780__bF_buf0), .C(_abc_15497_new_n2809_), .Y(_abc_15497_new_n2827_));
AOI21X1 AOI21X1_105 ( .A(_abc_15497_new_n2829_), .B(_abc_15497_new_n2831_), .C(_abc_15497_new_n2830_), .Y(_abc_15497_new_n2832_));
AOI21X1 AOI21X1_106 ( .A(_abc_15497_new_n2790_), .B(_abc_15497_new_n2803_), .C(_abc_15497_new_n2857_), .Y(_abc_15497_new_n2858_));
AOI21X1 AOI21X1_107 ( .A(_abc_15497_new_n2856_), .B(_abc_15497_new_n2861_), .C(_abc_15497_new_n2738_), .Y(_abc_15497_new_n2862_));
AOI21X1 AOI21X1_108 ( .A(round_ctr_reg_5_), .B(round_ctr_reg_3_), .C(round_ctr_reg_6_), .Y(_abc_15497_new_n2863_));
AOI21X1 AOI21X1_109 ( .A(_abc_15497_new_n2870_), .B(_abc_15497_new_n2871_), .C(_abc_15497_new_n2869_), .Y(_abc_15497_new_n2872_));
AOI21X1 AOI21X1_11 ( .A(_abc_15497_new_n831_), .B(_abc_15497_new_n834_), .C(_abc_15497_new_n829_), .Y(_abc_15497_new_n835_));
AOI21X1 AOI21X1_110 ( .A(_abc_15497_new_n2813_), .B(_abc_15497_new_n2816_), .C(_abc_15497_new_n2874_), .Y(_abc_15497_new_n2875_));
AOI21X1 AOI21X1_111 ( .A(_abc_15497_new_n2860_), .B(_abc_15497_new_n2859_), .C(_abc_15497_new_n2858_), .Y(_abc_15497_new_n2884_));
AOI21X1 AOI21X1_112 ( .A(_abc_15497_new_n2861_), .B(_abc_15497_new_n2738_), .C(_abc_15497_new_n2884_), .Y(_abc_15497_new_n2885_));
AOI21X1 AOI21X1_113 ( .A(_abc_15497_new_n2838_), .B(_abc_15497_new_n2850_), .C(_abc_15497_new_n2887_), .Y(_abc_15497_new_n2888_));
AOI21X1 AOI21X1_114 ( .A(_abc_15497_new_n1320_), .B(_abc_15497_new_n2890_), .C(_abc_15497_new_n2889_), .Y(_abc_15497_new_n2891_));
AOI21X1 AOI21X1_115 ( .A(_abc_15497_new_n2899_), .B(_abc_15497_new_n2900_), .C(w_3_), .Y(_abc_15497_new_n2901_));
AOI21X1 AOI21X1_116 ( .A(_abc_15497_new_n2916_), .B(_abc_15497_new_n2911_), .C(_abc_15497_new_n2888_), .Y(_abc_15497_new_n2917_));
AOI21X1 AOI21X1_117 ( .A(_abc_15497_new_n2920_), .B(_abc_15497_new_n2919_), .C(_abc_15497_new_n2918_), .Y(_abc_15497_new_n2921_));
AOI21X1 AOI21X1_118 ( .A(round_ctr_reg_4_), .B(round_ctr_reg_2_), .C(round_ctr_reg_6_), .Y(_abc_15497_new_n2923_));
AOI21X1 AOI21X1_119 ( .A(_abc_15497_new_n2926_), .B(_abc_15497_new_n2927_), .C(_abc_15497_new_n2925__bF_buf2), .Y(_abc_15497_new_n2930_));
AOI21X1 AOI21X1_12 ( .A(_abc_15497_new_n822_), .B(_abc_15497_new_n825_), .C(_abc_15497_new_n820_), .Y(_abc_15497_new_n836_));
AOI21X1 AOI21X1_120 ( .A(_abc_15497_new_n2931_), .B(_abc_15497_new_n2932_), .C(_abc_15497_new_n2756__bF_buf1), .Y(_abc_15497_new_n2933_));
AOI21X1 AOI21X1_121 ( .A(_abc_15497_new_n2867_), .B(_abc_15497_new_n2934_), .C(_abc_15497_new_n2940_), .Y(_abc_15497_new_n2941_));
AOI21X1 AOI21X1_122 ( .A(_abc_15497_new_n2927_), .B(_abc_15497_new_n2925__bF_buf1), .C(_abc_15497_new_n2917_), .Y(_abc_15497_new_n2943_));
AOI21X1 AOI21X1_123 ( .A(_abc_15497_new_n1333_), .B(_abc_15497_new_n2948_), .C(_abc_15497_new_n2946_), .Y(_abc_15497_new_n2949_));
AOI21X1 AOI21X1_124 ( .A(_abc_15497_new_n2899_), .B(w_3_), .C(_abc_15497_new_n2965_), .Y(_abc_15497_new_n2966_));
AOI21X1 AOI21X1_125 ( .A(_abc_15497_new_n2897_), .B(_abc_15497_new_n2909_), .C(_abc_15497_new_n2974_), .Y(_abc_15497_new_n2975_));
AOI21X1 AOI21X1_126 ( .A(_abc_15497_new_n2976_), .B(_abc_15497_new_n2756__bF_buf0), .C(_abc_15497_new_n2979_), .Y(_abc_15497_new_n2980_));
AOI21X1 AOI21X1_127 ( .A(_abc_15497_new_n2883_), .B(_abc_15497_new_n2934_), .C(_abc_15497_new_n2940_), .Y(_abc_15497_new_n2996_));
AOI21X1 AOI21X1_128 ( .A(_abc_15497_new_n2969_), .B(_abc_15497_new_n3004_), .C(_abc_15497_new_n2945_), .Y(_abc_15497_new_n3005_));
AOI21X1 AOI21X1_129 ( .A(_abc_15497_new_n1343_), .B(_abc_15497_new_n3009_), .C(_abc_15497_new_n3008_), .Y(_abc_15497_new_n3010_));
AOI21X1 AOI21X1_13 ( .A(_abc_15497_new_n819_), .B(_abc_15497_new_n837_), .C(_abc_15497_new_n812_), .Y(_abc_15497_new_n838_));
AOI21X1 AOI21X1_130 ( .A(_abc_15497_new_n3023_), .B(_abc_15497_new_n3020_), .C(w_5_), .Y(_abc_15497_new_n3027_));
AOI21X1 AOI21X1_131 ( .A(_abc_15497_new_n3031_), .B(_abc_15497_new_n3034_), .C(_abc_15497_new_n3007_), .Y(_abc_15497_new_n3035_));
AOI21X1 AOI21X1_132 ( .A(_abc_15497_new_n2954_), .B(_abc_15497_new_n2968_), .C(_abc_15497_new_n3036_), .Y(_abc_15497_new_n3037_));
AOI21X1 AOI21X1_133 ( .A(_abc_15497_new_n3039_), .B(_abc_15497_new_n3038_), .C(_abc_15497_new_n3037_), .Y(_abc_15497_new_n3040_));
AOI21X1 AOI21X1_134 ( .A(_abc_15497_new_n2987_), .B(_abc_15497_new_n2944_), .C(_abc_15497_new_n3047_), .Y(_abc_15497_new_n3048_));
AOI21X1 AOI21X1_135 ( .A(_abc_15497_new_n3043_), .B(_abc_15497_new_n3042_), .C(_abc_15497_new_n2781__bF_buf0), .Y(_abc_15497_new_n3049_));
AOI21X1 AOI21X1_136 ( .A(_abc_15497_new_n3041_), .B(_abc_15497_new_n3044_), .C(_abc_15497_new_n3006_), .Y(_abc_15497_new_n3060_));
AOI21X1 AOI21X1_137 ( .A(_abc_15497_new_n3042_), .B(_abc_15497_new_n2781__bF_buf3), .C(_abc_15497_new_n3040_), .Y(_abc_15497_new_n3064_));
AOI21X1 AOI21X1_138 ( .A(_abc_15497_new_n1357_), .B(_abc_15497_new_n3067_), .C(_abc_15497_new_n3066_), .Y(_abc_15497_new_n3068_));
AOI21X1 AOI21X1_139 ( .A(_abc_15497_new_n3081_), .B(_abc_15497_new_n3078_), .C(w_6_), .Y(_abc_15497_new_n3085_));
AOI21X1 AOI21X1_14 ( .A(_abc_15497_new_n792_), .B(_abc_15497_new_n847_), .C(_abc_15497_new_n839_), .Y(_abc_15497_new_n848_));
AOI21X1 AOI21X1_140 ( .A(_abc_15497_new_n3089_), .B(_abc_15497_new_n3092_), .C(_abc_15497_new_n3065_), .Y(_abc_15497_new_n3093_));
AOI21X1 AOI21X1_141 ( .A(_abc_15497_new_n3016_), .B(_abc_15497_new_n3029_), .C(_abc_15497_new_n3094_), .Y(_abc_15497_new_n3095_));
AOI21X1 AOI21X1_142 ( .A(_abc_15497_new_n3097_), .B(_abc_15497_new_n3096_), .C(_abc_15497_new_n3095_), .Y(_abc_15497_new_n3098_));
AOI21X1 AOI21X1_143 ( .A(_abc_15497_new_n3101_), .B(_abc_15497_new_n3100_), .C(_abc_15497_new_n2738_), .Y(_abc_15497_new_n3105_));
AOI21X1 AOI21X1_144 ( .A(_abc_15497_new_n1353_), .B(_abc_15497_new_n3121_), .C(_abc_15497_new_n3120_), .Y(_abc_15497_new_n3122_));
AOI21X1 AOI21X1_145 ( .A(_abc_15497_new_n2756__bF_buf3), .B(_abc_15497_new_n3124_), .C(_abc_15497_new_n3128_), .Y(_abc_15497_new_n3129_));
AOI21X1 AOI21X1_146 ( .A(_abc_15497_new_n3136_), .B(_abc_15497_new_n3133_), .C(w_7_), .Y(_abc_15497_new_n3140_));
AOI21X1 AOI21X1_147 ( .A(_abc_15497_new_n3074_), .B(_abc_15497_new_n3087_), .C(_abc_15497_new_n3153_), .Y(_abc_15497_new_n3154_));
AOI21X1 AOI21X1_148 ( .A(_abc_15497_new_n1364_), .B(_abc_15497_new_n3171_), .C(_abc_15497_new_n3170_), .Y(_abc_15497_new_n3172_));
AOI21X1 AOI21X1_149 ( .A(_abc_15497_new_n3191_), .B(_abc_15497_new_n3193_), .C(_abc_15497_new_n3190_), .Y(_abc_15497_new_n3194_));
AOI21X1 AOI21X1_15 ( .A(_abc_15497_new_n853_), .B(_abc_15497_new_n857_), .C(_abc_15497_new_n851_), .Y(_abc_15497_new_n863_));
AOI21X1 AOI21X1_150 ( .A(_abc_15497_new_n3147_), .B(_abc_15497_new_n3142_), .C(_abc_15497_new_n3196_), .Y(_abc_15497_new_n3197_));
AOI21X1 AOI21X1_151 ( .A(_abc_15497_new_n3205_), .B(_abc_15497_new_n3204_), .C(_abc_15497_new_n2924__bF_buf0), .Y(_abc_15497_new_n3208_));
AOI21X1 AOI21X1_152 ( .A(_abc_15497_new_n3195_), .B(_abc_15497_new_n3202_), .C(_abc_15497_new_n2759__bF_buf1), .Y(_abc_15497_new_n3209_));
AOI21X1 AOI21X1_153 ( .A(_abc_15497_new_n3103_), .B(_abc_15497_new_n3107_), .C(_abc_15497_new_n3162_), .Y(_abc_15497_new_n3213_));
AOI21X1 AOI21X1_154 ( .A(_abc_15497_new_n3213_), .B(_abc_15497_new_n3061_), .C(_abc_15497_new_n3215_), .Y(_abc_15497_new_n3216_));
AOI21X1 AOI21X1_155 ( .A(_abc_15497_new_n3201_), .B(_abc_15497_new_n3198_), .C(_abc_15497_new_n3169_), .Y(_abc_15497_new_n3228_));
AOI21X1 AOI21X1_156 ( .A(_abc_15497_new_n2944_), .B(_abc_15497_new_n2755_), .C(_abc_15497_new_n3237_), .Y(_abc_15497_new_n3238_));
AOI21X1 AOI21X1_157 ( .A(d_reg_9_), .B(_abc_15497_new_n3232_), .C(_abc_15497_new_n3231_), .Y(_abc_15497_new_n3239_));
AOI21X1 AOI21X1_158 ( .A(_abc_15497_new_n3248_), .B(_abc_15497_new_n3246_), .C(_abc_15497_new_n3251_), .Y(_abc_15497_new_n3252_));
AOI21X1 AOI21X1_159 ( .A(_abc_15497_new_n1374_), .B(_abc_15497_new_n3254_), .C(_abc_15497_new_n3235_), .Y(_abc_15497_new_n3255_));
AOI21X1 AOI21X1_16 ( .A(_abc_15497_new_n888_), .B(_abc_15497_new_n886_), .C(_abc_15497_new_n890_), .Y(_abc_15497_new_n891_));
AOI21X1 AOI21X1_160 ( .A(_abc_15497_new_n2756__bF_buf2), .B(_abc_15497_new_n3257_), .C(_abc_15497_new_n3240_), .Y(_abc_15497_new_n3258_));
AOI21X1 AOI21X1_161 ( .A(_abc_15497_new_n3247_), .B(_abc_15497_new_n3244_), .C(w_9_), .Y(_abc_15497_new_n3260_));
AOI21X1 AOI21X1_162 ( .A(_abc_15497_new_n3253_), .B(_abc_15497_new_n3264_), .C(_abc_15497_new_n3230_), .Y(_abc_15497_new_n3265_));
AOI21X1 AOI21X1_163 ( .A(_abc_15497_new_n3271_), .B(_abc_15497_new_n3272_), .C(_abc_15497_new_n2781__bF_buf2), .Y(_abc_15497_new_n3276_));
AOI21X1 AOI21X1_164 ( .A(_abc_15497_new_n3269_), .B(_abc_15497_new_n3273_), .C(_abc_15497_new_n3229_), .Y(_abc_15497_new_n3283_));
AOI21X1 AOI21X1_165 ( .A(_abc_15497_new_n3217_), .B(_abc_15497_new_n3286_), .C(_abc_15497_new_n3284_), .Y(_abc_15497_new_n3287_));
AOI21X1 AOI21X1_166 ( .A(_abc_15497_new_n3271_), .B(_abc_15497_new_n2781__bF_buf1), .C(_abc_15497_new_n3268_), .Y(_abc_15497_new_n3288_));
AOI21X1 AOI21X1_167 ( .A(_abc_15497_new_n3290_), .B(_abc_15497_new_n3292_), .C(_abc_15497_new_n3291_), .Y(_abc_15497_new_n3293_));
AOI21X1 AOI21X1_168 ( .A(_abc_15497_new_n3307_), .B(_abc_15497_new_n3304_), .C(w_10_), .Y(_abc_15497_new_n3310_));
AOI21X1 AOI21X1_169 ( .A(_abc_15497_new_n2756__bF_buf1), .B(_abc_15497_new_n3295_), .C(_abc_15497_new_n3317_), .Y(_abc_15497_new_n3318_));
AOI21X1 AOI21X1_17 ( .A(_abc_15497_new_n892_), .B(_abc_15497_new_n896_), .C(_abc_15497_new_n870__bF_buf8), .Y(_abc_15497_new_n897_));
AOI21X1 AOI21X1_170 ( .A(_abc_15497_new_n3314_), .B(_abc_15497_new_n3322_), .C(_abc_15497_new_n3289_), .Y(_abc_15497_new_n3323_));
AOI21X1 AOI21X1_171 ( .A(_abc_15497_new_n2759__bF_buf4), .B(_abc_15497_new_n3255_), .C(_abc_15497_new_n3328_), .Y(_abc_15497_new_n3329_));
AOI21X1 AOI21X1_172 ( .A(_abc_15497_new_n3330_), .B(_abc_15497_new_n3262_), .C(_abc_15497_new_n3331_), .Y(_abc_15497_new_n3332_));
AOI21X1 AOI21X1_173 ( .A(_abc_15497_new_n3333_), .B(_abc_15497_new_n3334_), .C(_abc_15497_new_n2759__bF_buf2), .Y(_abc_15497_new_n3338_));
AOI21X1 AOI21X1_174 ( .A(_abc_15497_new_n1398_), .B(_abc_15497_new_n3353_), .C(_abc_15497_new_n3352_), .Y(_abc_15497_new_n3354_));
AOI21X1 AOI21X1_175 ( .A(_abc_15497_new_n3365_), .B(_abc_15497_new_n3366_), .C(w_11_), .Y(_abc_15497_new_n3370_));
AOI21X1 AOI21X1_176 ( .A(_abc_15497_new_n3357_), .B(_abc_15497_new_n3359_), .C(_abc_15497_new_n3373_), .Y(_abc_15497_new_n3374_));
AOI21X1 AOI21X1_177 ( .A(_abc_15497_new_n3299_), .B(_abc_15497_new_n3313_), .C(_abc_15497_new_n3381_), .Y(_abc_15497_new_n3382_));
AOI21X1 AOI21X1_178 ( .A(_abc_15497_new_n3357_), .B(_abc_15497_new_n3359_), .C(_abc_15497_new_n3378_), .Y(_abc_15497_new_n3383_));
AOI21X1 AOI21X1_179 ( .A(_abc_15497_new_n3376_), .B(_abc_15497_new_n3377_), .C(_abc_15497_new_n3375_), .Y(_abc_15497_new_n3384_));
AOI21X1 AOI21X1_18 ( .A(_abc_15497_new_n892_), .B(_abc_15497_new_n896_), .C(_abc_15497_new_n895_), .Y(_abc_15497_new_n902_));
AOI21X1 AOI21X1_180 ( .A(_abc_15497_new_n3333_), .B(_abc_15497_new_n2759__bF_buf0), .C(_abc_15497_new_n3326_), .Y(_abc_15497_new_n3391_));
AOI21X1 AOI21X1_181 ( .A(_abc_15497_new_n3336_), .B(_abc_15497_new_n3340_), .C(_abc_15497_new_n3404_), .Y(_abc_15497_new_n3405_));
AOI21X1 AOI21X1_182 ( .A(_abc_15497_new_n3405_), .B(_abc_15497_new_n3284_), .C(_abc_15497_new_n3406_), .Y(_abc_15497_new_n3407_));
AOI21X1 AOI21X1_183 ( .A(_abc_15497_new_n2756__bF_buf0), .B(_abc_15497_new_n3356_), .C(_abc_15497_new_n3413_), .Y(_abc_15497_new_n3414_));
AOI21X1 AOI21X1_184 ( .A(_abc_15497_new_n3415_), .B(_abc_15497_new_n3410_), .C(_abc_15497_new_n3382_), .Y(_abc_15497_new_n3416_));
AOI21X1 AOI21X1_185 ( .A(_abc_15497_new_n3388_), .B(_abc_15497_new_n2755_), .C(_abc_15497_new_n3416_), .Y(_abc_15497_new_n3417_));
AOI21X1 AOI21X1_186 ( .A(_abc_15497_new_n1414_), .B(_abc_15497_new_n3420_), .C(_abc_15497_new_n3419_), .Y(_abc_15497_new_n3421_));
AOI21X1 AOI21X1_187 ( .A(_abc_15497_new_n3436_), .B(_abc_15497_new_n3433_), .C(w_12_), .Y(_abc_15497_new_n3439_));
AOI21X1 AOI21X1_188 ( .A(_abc_15497_new_n2756__bF_buf4), .B(_abc_15497_new_n3424_), .C(_abc_15497_new_n3447_), .Y(_abc_15497_new_n3448_));
AOI21X1 AOI21X1_189 ( .A(_abc_15497_new_n3443_), .B(_abc_15497_new_n3452_), .C(_abc_15497_new_n3418_), .Y(_abc_15497_new_n3453_));
AOI21X1 AOI21X1_19 ( .A(_abc_15497_new_n942_), .B(_abc_15497_new_n938_), .C(_abc_15497_new_n870__bF_buf4), .Y(_abc_15497_new_n943_));
AOI21X1 AOI21X1_190 ( .A(_abc_15497_new_n3375_), .B(_abc_15497_new_n3372_), .C(_abc_15497_new_n3454_), .Y(_abc_15497_new_n3455_));
AOI21X1 AOI21X1_191 ( .A(_abc_15497_new_n3456_), .B(_abc_15497_new_n3457_), .C(_abc_15497_new_n3455_), .Y(_abc_15497_new_n3458_));
AOI21X1 AOI21X1_192 ( .A(_abc_15497_new_n3464_), .B(_abc_15497_new_n3465_), .C(_abc_15497_new_n3351_), .Y(_abc_15497_new_n3466_));
AOI21X1 AOI21X1_193 ( .A(_abc_15497_new_n2944_), .B(_abc_15497_new_n2755_), .C(_abc_15497_new_n3487_), .Y(_abc_15497_new_n3488_));
AOI21X1 AOI21X1_194 ( .A(_abc_15497_new_n3497_), .B(_abc_15497_new_n3500_), .C(_abc_15497_new_n3503_), .Y(_abc_15497_new_n3504_));
AOI21X1 AOI21X1_195 ( .A(_abc_15497_new_n2756__bF_buf0), .B(_abc_15497_new_n3506_), .C(_abc_15497_new_n3492_), .Y(_abc_15497_new_n3507_));
AOI21X1 AOI21X1_196 ( .A(_abc_15497_new_n3505_), .B(_abc_15497_new_n3511_), .C(_abc_15497_new_n3480_), .Y(_abc_15497_new_n3512_));
AOI21X1 AOI21X1_197 ( .A(_abc_15497_new_n3428_), .B(_abc_15497_new_n3442_), .C(_abc_15497_new_n3517_), .Y(_abc_15497_new_n3518_));
AOI21X1 AOI21X1_198 ( .A(_abc_15497_new_n3460_), .B(_abc_15497_new_n2925__bF_buf0), .C(_abc_15497_new_n3458_), .Y(_abc_15497_new_n3523_));
AOI21X1 AOI21X1_199 ( .A(_abc_15497_new_n3520_), .B(_abc_15497_new_n3519_), .C(_abc_15497_new_n2755_), .Y(_abc_15497_new_n3524_));
AOI21X1 AOI21X1_2 ( .A(_abc_15497_new_n701_), .B(_abc_15497_new_n704_), .C(_abc_15497_new_n699_), .Y(_abc_15497_new_n715_));
AOI21X1 AOI21X1_20 ( .A(_abc_15497_new_n957_), .B(_abc_15497_new_n959_), .C(_abc_15497_new_n961_), .Y(_abc_15497_new_n969_));
AOI21X1 AOI21X1_200 ( .A(_abc_15497_new_n3478_), .B(_abc_15497_new_n3528_), .C(_abc_15497_new_n3529_), .Y(_abc_15497_new_n3530_));
AOI21X1 AOI21X1_201 ( .A(_abc_15497_new_n3459_), .B(_abc_15497_new_n3462_), .C(_abc_15497_new_n3417_), .Y(_abc_15497_new_n3535_));
AOI21X1 AOI21X1_202 ( .A(_abc_15497_new_n3519_), .B(_abc_15497_new_n2755_), .C(_abc_15497_new_n3515_), .Y(_abc_15497_new_n3541_));
AOI21X1 AOI21X1_203 ( .A(_abc_15497_new_n2944_), .B(_abc_15497_new_n2755_), .C(_abc_15497_new_n3550_), .Y(_abc_15497_new_n3551_));
AOI21X1 AOI21X1_204 ( .A(_abc_15497_new_n3543_), .B(_abc_15497_new_n3548_), .C(_abc_15497_new_n3544_), .Y(_abc_15497_new_n3552_));
AOI21X1 AOI21X1_205 ( .A(_abc_15497_new_n3563_), .B(_abc_15497_new_n3564_), .C(w_14_), .Y(_abc_15497_new_n3567_));
AOI21X1 AOI21X1_206 ( .A(_abc_15497_new_n2756__bF_buf4), .B(_abc_15497_new_n3572_), .C(_abc_15497_new_n3556_), .Y(_abc_15497_new_n3573_));
AOI21X1 AOI21X1_207 ( .A(_abc_15497_new_n3571_), .B(_abc_15497_new_n3577_), .C(_abc_15497_new_n3542_), .Y(_abc_15497_new_n3578_));
AOI21X1 AOI21X1_208 ( .A(_abc_15497_new_n1425_), .B(_abc_15497_new_n3485_), .C(_abc_15497_new_n3481_), .Y(_abc_15497_new_n3583_));
AOI21X1 AOI21X1_209 ( .A(_abc_15497_new_n3585_), .B(_abc_15497_new_n3509_), .C(_abc_15497_new_n3586_), .Y(_abc_15497_new_n3587_));
AOI21X1 AOI21X1_21 ( .A(_abc_15497_new_n971_), .B(_abc_15497_new_n972_), .C(_abc_15497_new_n870__bF_buf2), .Y(_abc_15497_new_n973_));
AOI21X1 AOI21X1_210 ( .A(_abc_15497_new_n3588_), .B(_abc_15497_new_n3589_), .C(_abc_15497_new_n2924__bF_buf4), .Y(_abc_15497_new_n3593_));
AOI21X1 AOI21X1_211 ( .A(_abc_15497_new_n3627_), .B(_abc_15497_new_n3624_), .C(w_15_), .Y(_abc_15497_new_n3630_));
AOI21X1 AOI21X1_212 ( .A(_abc_15497_new_n1447_), .B(_abc_15497_new_n3616_), .C(_abc_15497_new_n3612_), .Y(_abc_15497_new_n3635_));
AOI21X1 AOI21X1_213 ( .A(_abc_15497_new_n3634_), .B(_abc_15497_new_n3642_), .C(_abc_15497_new_n3606_), .Y(_abc_15497_new_n3643_));
AOI21X1 AOI21X1_214 ( .A(_abc_15497_new_n3649_), .B(_abc_15497_new_n3575_), .C(_abc_15497_new_n3650_), .Y(_abc_15497_new_n3651_));
AOI21X1 AOI21X1_215 ( .A(_abc_15497_new_n3588_), .B(_abc_15497_new_n2924__bF_buf2), .C(_abc_15497_new_n3581_), .Y(_abc_15497_new_n3656_));
AOI21X1 AOI21X1_216 ( .A(_abc_15497_new_n3653_), .B(_abc_15497_new_n3652_), .C(_abc_15497_new_n2742__bF_buf2), .Y(_abc_15497_new_n3657_));
AOI21X1 AOI21X1_217 ( .A(_abc_15497_new_n3598_), .B(_abc_15497_new_n3604_), .C(_abc_15497_new_n3660_), .Y(_abc_15497_new_n3661_));
AOI21X1 AOI21X1_218 ( .A(_abc_15497_new_n3591_), .B(_abc_15497_new_n3595_), .C(_abc_15497_new_n3660_), .Y(_abc_15497_new_n3668_));
AOI21X1 AOI21X1_219 ( .A(_abc_15497_new_n3668_), .B(_abc_15497_new_n3670_), .C(_abc_15497_new_n3671_), .Y(_abc_15497_new_n3672_));
AOI21X1 AOI21X1_22 ( .A(_abc_15497_new_n870__bF_buf1), .B(_abc_15497_new_n974_), .C(_abc_15497_new_n973_), .Y(_0H4_reg_31_0__4_));
AOI21X1 AOI21X1_220 ( .A(_abc_15497_new_n3217_), .B(_abc_15497_new_n3674_), .C(_abc_15497_new_n3673_), .Y(_abc_15497_new_n3675_));
AOI21X1 AOI21X1_221 ( .A(_abc_15497_new_n3704_), .B(_abc_15497_new_n3703_), .C(_abc_15497_new_n3680_), .Y(_abc_15497_new_n3707_));
AOI21X1 AOI21X1_222 ( .A(_abc_15497_new_n3701_), .B(_abc_15497_new_n3698_), .C(_abc_15497_new_n3681_), .Y(_abc_15497_new_n3708_));
AOI21X1 AOI21X1_223 ( .A(_abc_15497_new_n3709_), .B(_abc_15497_new_n3706_), .C(_abc_15497_new_n3677_), .Y(_abc_15497_new_n3711_));
AOI21X1 AOI21X1_224 ( .A(_abc_15497_new_n3726_), .B(_abc_15497_new_n3729_), .C(_abc_15497_new_n3727_), .Y(_abc_15497_new_n3730_));
AOI21X1 AOI21X1_225 ( .A(_abc_15497_new_n3750_), .B(_abc_15497_new_n3753_), .C(_abc_15497_new_n3725_), .Y(_abc_15497_new_n3754_));
AOI21X1 AOI21X1_226 ( .A(_abc_15497_new_n3700_), .B(_abc_15497_new_n3690_), .C(_abc_15497_new_n3755_), .Y(_abc_15497_new_n3756_));
AOI21X1 AOI21X1_227 ( .A(_abc_15497_new_n3721_), .B(_abc_15497_new_n3770_), .C(_abc_15497_new_n3771_), .Y(_abc_15497_new_n3772_));
AOI21X1 AOI21X1_228 ( .A(_abc_15497_new_n1650__bF_buf0), .B(_abc_15497_new_n3773_), .C(_abc_15497_new_n3772_), .Y(_abc_15497_new_n3774_));
AOI21X1 AOI21X1_229 ( .A(_abc_15497_new_n3764_), .B(_abc_15497_new_n3768_), .C(_abc_15497_new_n3714_), .Y(_abc_15497_new_n3776_));
AOI21X1 AOI21X1_23 ( .A(e_reg_4_), .B(_auto_iopadmap_cc_368_execute_22625_4_), .C(_abc_15497_new_n970_), .Y(_abc_15497_new_n976_));
AOI21X1 AOI21X1_230 ( .A(_abc_15497_new_n3760_), .B(_abc_15497_new_n3763_), .C(_abc_15497_new_n3765_), .Y(_abc_15497_new_n3777_));
AOI21X1 AOI21X1_231 ( .A(_abc_15497_new_n3711_), .B(_abc_15497_new_n3778_), .C(_abc_15497_new_n3777_), .Y(_abc_15497_new_n3779_));
AOI21X1 AOI21X1_232 ( .A(_abc_15497_new_n3676_), .B(_abc_15497_new_n3776_), .C(_abc_15497_new_n3780_), .Y(_abc_15497_new_n3781_));
AOI21X1 AOI21X1_233 ( .A(_abc_15497_new_n3761_), .B(_abc_15497_new_n2944_), .C(_abc_15497_new_n3759_), .Y(_abc_15497_new_n3816_));
AOI21X1 AOI21X1_234 ( .A(_abc_15497_new_n3804_), .B(_abc_15497_new_n3807_), .C(_abc_15497_new_n3828_), .Y(_abc_15497_new_n3829_));
AOI21X1 AOI21X1_235 ( .A(_abc_15497_new_n3853_), .B(_abc_15497_new_n3854_), .C(_abc_15497_new_n3852_), .Y(_abc_15497_new_n3857_));
AOI21X1 AOI21X1_236 ( .A(_abc_15497_new_n3847_), .B(_abc_15497_new_n3850_), .C(_abc_15497_new_n3829_), .Y(_abc_15497_new_n3858_));
AOI21X1 AOI21X1_237 ( .A(_abc_15497_new_n3810_), .B(_abc_15497_new_n3813_), .C(_abc_15497_new_n3816_), .Y(_abc_15497_new_n3870_));
AOI21X1 AOI21X1_238 ( .A(_abc_15497_new_n3871_), .B(_abc_15497_new_n3872_), .C(_abc_15497_new_n3782_), .Y(_abc_15497_new_n3873_));
AOI21X1 AOI21X1_239 ( .A(_abc_15497_new_n3862_), .B(_abc_15497_new_n3861_), .C(_abc_15497_new_n3810_), .Y(_abc_15497_new_n3874_));
AOI21X1 AOI21X1_24 ( .A(_abc_15497_new_n1025_), .B(_abc_15497_new_n1008_), .C(_abc_15497_new_n870__bF_buf7), .Y(_abc_15497_new_n1030_));
AOI21X1 AOI21X1_240 ( .A(_abc_15497_new_n3859_), .B(_abc_15497_new_n3856_), .C(_abc_15497_new_n3827_), .Y(_abc_15497_new_n3875_));
AOI21X1 AOI21X1_241 ( .A(_abc_15497_new_n3859_), .B(_abc_15497_new_n3856_), .C(_abc_15497_new_n3810_), .Y(_abc_15497_new_n3877_));
AOI21X1 AOI21X1_242 ( .A(_abc_15497_new_n3849_), .B(_abc_15497_new_n3887_), .C(_abc_15497_new_n3892_), .Y(_abc_15497_new_n3893_));
AOI21X1 AOI21X1_243 ( .A(_abc_15497_new_n3916_), .B(_abc_15497_new_n3917_), .C(_abc_15497_new_n3915_), .Y(_abc_15497_new_n3920_));
AOI21X1 AOI21X1_244 ( .A(_abc_15497_new_n3913_), .B(_abc_15497_new_n3910_), .C(_abc_15497_new_n3893_), .Y(_abc_15497_new_n3921_));
AOI21X1 AOI21X1_245 ( .A(_abc_15497_new_n3851_), .B(_abc_15497_new_n3678_), .C(_abc_15497_new_n3858_), .Y(_abc_15497_new_n3924_));
AOI21X1 AOI21X1_246 ( .A(_abc_15497_new_n3922_), .B(_abc_15497_new_n3919_), .C(_abc_15497_new_n3924_), .Y(_abc_15497_new_n3935_));
AOI21X1 AOI21X1_247 ( .A(_abc_15497_new_n3885_), .B(_abc_15497_new_n3928_), .C(_abc_15497_new_n3935_), .Y(_abc_15497_new_n3936_));
AOI21X1 AOI21X1_248 ( .A(_abc_15497_new_n3912_), .B(_abc_15497_new_n3902_), .C(_abc_15497_new_n3942_), .Y(_abc_15497_new_n3943_));
AOI21X1 AOI21X1_249 ( .A(_abc_15497_new_n3967_), .B(_abc_15497_new_n3968_), .C(_abc_15497_new_n3966_), .Y(_abc_15497_new_n3971_));
AOI21X1 AOI21X1_25 ( .A(_abc_15497_new_n1036_), .B(_abc_15497_new_n1058_), .C(_abc_15497_new_n1060_), .Y(_abc_15497_new_n1061_));
AOI21X1 AOI21X1_250 ( .A(_abc_15497_new_n3961_), .B(_abc_15497_new_n3964_), .C(_abc_15497_new_n3943_), .Y(_abc_15497_new_n3972_));
AOI21X1 AOI21X1_251 ( .A(_abc_15497_new_n3914_), .B(_abc_15497_new_n3678_), .C(_abc_15497_new_n3921_), .Y(_abc_15497_new_n3975_));
AOI21X1 AOI21X1_252 ( .A(_abc_15497_new_n3973_), .B(_abc_15497_new_n3970_), .C(_abc_15497_new_n3975_), .Y(_abc_15497_new_n3988_));
AOI21X1 AOI21X1_253 ( .A(_abc_15497_new_n3935_), .B(_abc_15497_new_n3989_), .C(_abc_15497_new_n3988_), .Y(_abc_15497_new_n3990_));
AOI21X1 AOI21X1_254 ( .A(_abc_15497_new_n3963_), .B(_abc_15497_new_n3953_), .C(_abc_15497_new_n3997_), .Y(_abc_15497_new_n3998_));
AOI21X1 AOI21X1_255 ( .A(_abc_15497_new_n4022_), .B(_abc_15497_new_n4023_), .C(_abc_15497_new_n4021_), .Y(_abc_15497_new_n4026_));
AOI21X1 AOI21X1_256 ( .A(_abc_15497_new_n4016_), .B(_abc_15497_new_n4019_), .C(_abc_15497_new_n3998_), .Y(_abc_15497_new_n4027_));
AOI21X1 AOI21X1_257 ( .A(_abc_15497_new_n3965_), .B(_abc_15497_new_n2780__bF_buf0), .C(_abc_15497_new_n3972_), .Y(_abc_15497_new_n4030_));
AOI21X1 AOI21X1_258 ( .A(_abc_15497_new_n4028_), .B(_abc_15497_new_n4025_), .C(_abc_15497_new_n4030_), .Y(_abc_15497_new_n4041_));
AOI21X1 AOI21X1_259 ( .A(_abc_15497_new_n3987_), .B(_abc_15497_new_n3990_), .C(_abc_15497_new_n4035_), .Y(_abc_15497_new_n4042_));
AOI21X1 AOI21X1_26 ( .A(_abc_15497_new_n1075_), .B(_abc_15497_new_n1065_), .C(_abc_15497_new_n1074_), .Y(_abc_15497_new_n1085_));
AOI21X1 AOI21X1_260 ( .A(_abc_15497_new_n1543_), .B(_abc_15497_new_n4052_), .C(_abc_15497_new_n4050_), .Y(_abc_15497_new_n4053_));
AOI21X1 AOI21X1_261 ( .A(_abc_15497_new_n4072_), .B(_abc_15497_new_n4073_), .C(_abc_15497_new_n4049_), .Y(_abc_15497_new_n4074_));
AOI21X1 AOI21X1_262 ( .A(_abc_15497_new_n4018_), .B(_abc_15497_new_n4008_), .C(_abc_15497_new_n4075_), .Y(_abc_15497_new_n4076_));
AOI21X1 AOI21X1_263 ( .A(_abc_15497_new_n4078_), .B(_abc_15497_new_n4077_), .C(_abc_15497_new_n4076_), .Y(_abc_15497_new_n4079_));
AOI21X1 AOI21X1_264 ( .A(_abc_15497_new_n4020_), .B(_abc_15497_new_n2756__bF_buf1), .C(_abc_15497_new_n4027_), .Y(_abc_15497_new_n4085_));
AOI21X1 AOI21X1_265 ( .A(_abc_15497_new_n4080_), .B(_abc_15497_new_n4083_), .C(_abc_15497_new_n4085_), .Y(_abc_15497_new_n4100_));
AOI21X1 AOI21X1_266 ( .A(_abc_15497_new_n4041_), .B(_abc_15497_new_n4101_), .C(_abc_15497_new_n4100_), .Y(_abc_15497_new_n4102_));
AOI21X1 AOI21X1_267 ( .A(_abc_15497_new_n3881_), .B(_abc_15497_new_n4098_), .C(_abc_15497_new_n4103_), .Y(_abc_15497_new_n4104_));
AOI21X1 AOI21X1_268 ( .A(_abc_15497_new_n1562_), .B(_abc_15497_new_n4110_), .C(_abc_15497_new_n4109_), .Y(_abc_15497_new_n4111_));
AOI21X1 AOI21X1_269 ( .A(_abc_15497_new_n4106_), .B(_abc_15497_new_n4143_), .C(_abc_15497_new_n1646_), .Y(_abc_15497_new_n4144_));
AOI21X1 AOI21X1_27 ( .A(_abc_15497_new_n1097_), .B(_abc_15497_new_n1082_), .C(_abc_15497_new_n1096_), .Y(_abc_15497_new_n1105_));
AOI21X1 AOI21X1_270 ( .A(_abc_15497_new_n1572_), .B(_abc_15497_new_n4156_), .C(_abc_15497_new_n4154_), .Y(_abc_15497_new_n4157_));
AOI21X1 AOI21X1_271 ( .A(_abc_15497_new_n4126_), .B(w_24_), .C(_abc_15497_new_n4124_), .Y(_abc_15497_new_n4163_));
AOI21X1 AOI21X1_272 ( .A(_abc_15497_new_n4150_), .B(_abc_15497_new_n4149_), .C(_abc_15497_new_n4179_), .Y(_abc_15497_new_n4180_));
AOI21X1 AOI21X1_273 ( .A(_abc_15497_new_n4140_), .B(_abc_15497_new_n4142_), .C(_abc_15497_new_n4179_), .Y(_abc_15497_new_n4189_));
AOI21X1 AOI21X1_274 ( .A(_abc_15497_new_n4195_), .B(_abc_15497_new_n4194_), .C(_abc_15497_new_n1586_), .Y(_abc_15497_new_n4196_));
AOI21X1 AOI21X1_275 ( .A(_abc_15497_new_n4191_), .B(_abc_15497_new_n4225_), .C(_abc_15497_new_n1646_), .Y(_abc_15497_new_n4226_));
AOI21X1 AOI21X1_276 ( .A(_abc_15497_new_n4211_), .B(w_26_), .C(_abc_15497_new_n4209_), .Y(_abc_15497_new_n4250_));
AOI21X1 AOI21X1_277 ( .A(_abc_15497_new_n4263_), .B(_abc_15497_new_n4272_), .C(_abc_15497_new_n4262_), .Y(_abc_15497_new_n4273_));
AOI21X1 AOI21X1_278 ( .A(_abc_15497_new_n4106_), .B(_abc_15497_new_n4271_), .C(_abc_15497_new_n4274_), .Y(_abc_15497_new_n4275_));
AOI21X1 AOI21X1_279 ( .A(b_reg_28_), .B(_abc_15497_new_n4280_), .C(_abc_15497_new_n4285_), .Y(_abc_15497_new_n4286_));
AOI21X1 AOI21X1_28 ( .A(_abc_15497_new_n1102_), .B(_abc_15497_new_n1104_), .C(_abc_15497_new_n1106_), .Y(_abc_15497_new_n1107_));
AOI21X1 AOI21X1_280 ( .A(_abc_15497_new_n4305_), .B(_abc_15497_new_n3216_), .C(_abc_15497_new_n4311_), .Y(_abc_15497_new_n4312_));
AOI21X1 AOI21X1_281 ( .A(_abc_15497_new_n4315_), .B(_abc_15497_new_n4104_), .C(_abc_15497_new_n4316_), .Y(_abc_15497_new_n4317_));
AOI21X1 AOI21X1_282 ( .A(_abc_15497_new_n4256_), .B(_abc_15497_new_n4278_), .C(_abc_15497_new_n4299_), .Y(_abc_15497_new_n4326_));
AOI21X1 AOI21X1_283 ( .A(_abc_15497_new_n4300_), .B(_abc_15497_new_n2743__bF_buf4), .C(_abc_15497_new_n4326_), .Y(_abc_15497_new_n4327_));
AOI21X1 AOI21X1_284 ( .A(d_reg_29_), .B(_abc_15497_new_n4330_), .C(_abc_15497_new_n4331_), .Y(_abc_15497_new_n4332_));
AOI21X1 AOI21X1_285 ( .A(_abc_15497_new_n4336_), .B(_abc_15497_new_n4337_), .C(_abc_15497_new_n2925__bF_buf3), .Y(_abc_15497_new_n4338_));
AOI21X1 AOI21X1_286 ( .A(_abc_15497_new_n4294_), .B(w_28_), .C(_abc_15497_new_n4293_), .Y(_abc_15497_new_n4343_));
AOI21X1 AOI21X1_287 ( .A(_abc_15497_new_n4303_), .B(_abc_15497_new_n4357_), .C(_abc_15497_new_n4366_), .Y(_abc_15497_new_n4367_));
AOI21X1 AOI21X1_288 ( .A(d_reg_30_), .B(_abc_15497_new_n4372_), .C(_abc_15497_new_n4373_), .Y(_abc_15497_new_n4374_));
AOI21X1 AOI21X1_289 ( .A(_abc_15497_new_n4378_), .B(_abc_15497_new_n4379_), .C(_abc_15497_new_n2925__bF_buf2), .Y(_abc_15497_new_n4380_));
AOI21X1 AOI21X1_29 ( .A(_abc_15497_new_n1148_), .B(_abc_15497_new_n1131_), .C(_abc_15497_new_n1147_), .Y(_abc_15497_new_n1152_));
AOI21X1 AOI21X1_290 ( .A(_abc_15497_new_n4369_), .B(_abc_15497_new_n4355_), .C(_abc_15497_new_n4400_), .Y(_abc_15497_new_n4406_));
AOI21X1 AOI21X1_291 ( .A(_abc_15497_new_n4408_), .B(_abc_15497_new_n4367_), .C(_abc_15497_new_n4409_), .Y(_abc_15497_new_n4410_));
AOI21X1 AOI21X1_292 ( .A(_abc_15497_new_n4368_), .B(_abc_15497_new_n4401_), .C(_abc_15497_new_n4406_), .Y(_abc_15497_new_n4435_));
AOI21X1 AOI21X1_293 ( .A(_abc_15497_new_n4447_), .B(round_ctr_inc_bF_buf10), .C(_abc_15497_new_n1647_), .Y(_abc_15497_new_n4449_));
AOI21X1 AOI21X1_294 ( .A(_abc_15497_new_n4463_), .B(_abc_15497_new_n4462_), .C(_abc_15497_new_n4464_), .Y(_0round_ctr_reg_6_0__3_));
AOI21X1 AOI21X1_295 ( .A(_abc_15497_new_n4468_), .B(_abc_15497_new_n4469_), .C(_abc_15497_new_n4470_), .Y(_0round_ctr_reg_6_0__5_));
AOI21X1 AOI21X1_296 ( .A(_abc_15497_new_n4500_), .B(_abc_15497_new_n4499_), .C(_abc_15497_new_n761_), .Y(_abc_15497_new_n4501_));
AOI21X1 AOI21X1_297 ( .A(_abc_15497_new_n4511_), .B(_abc_15497_new_n786_), .C(_abc_15497_new_n743_), .Y(_abc_15497_new_n4515_));
AOI21X1 AOI21X1_298 ( .A(_abc_15497_new_n4511_), .B(_abc_15497_new_n788_), .C(_abc_15497_new_n4519_), .Y(_abc_15497_new_n4520_));
AOI21X1 AOI21X1_299 ( .A(_abc_15497_new_n4530_), .B(_abc_15497_new_n720_), .C(_abc_15497_new_n711_), .Y(_abc_15497_new_n4535_));
AOI21X1 AOI21X1_3 ( .A(_abc_15497_new_n731_), .B(_abc_15497_new_n729_), .C(_abc_15497_new_n726_), .Y(_abc_15497_new_n732_));
AOI21X1 AOI21X1_30 ( .A(_abc_15497_new_n1160_), .B(_abc_15497_new_n1180_), .C(_abc_15497_new_n1182_), .Y(_abc_15497_new_n1183_));
AOI21X1 AOI21X1_300 ( .A(_abc_15497_new_n4530_), .B(_abc_15497_new_n724_), .C(_abc_15497_new_n716_), .Y(_abc_15497_new_n4550_));
AOI21X1 AOI21X1_301 ( .A(_abc_15497_new_n792_), .B(_abc_15497_new_n842_), .C(_abc_15497_new_n834_), .Y(_abc_15497_new_n4553_));
AOI21X1 AOI21X1_302 ( .A(_abc_15497_new_n4557_), .B(_abc_15497_new_n827_), .C(_abc_15497_new_n825_), .Y(_abc_15497_new_n4560_));
AOI21X1 AOI21X1_303 ( .A(_abc_15497_new_n4565_), .B(_abc_15497_new_n815_), .C(_abc_15497_new_n807_), .Y(_abc_15497_new_n4571_));
AOI21X1 AOI21X1_304 ( .A(_abc_15497_new_n4584_), .B(_abc_15497_new_n797_), .C(_abc_15497_new_n870__bF_buf9), .Y(_abc_15497_new_n4586_));
AOI21X1 AOI21X1_305 ( .A(w_mem_inst__abc_19396_new_n4801_), .B(w_mem_inst__abc_19396_new_n4803_), .C(w_mem_inst__abc_19396_new_n4805_), .Y(w_mem_inst__0w_ctr_reg_6_0__4_));
AOI21X1 AOI21X1_306 ( .A(w_mem_inst_w_ctr_reg_5_), .B(w_mem_inst__abc_19396_new_n4807_), .C(w_mem_inst__abc_19396_new_n4805_), .Y(w_mem_inst__abc_19396_new_n4808_));
AOI21X1 AOI21X1_307 ( .A(w_mem_inst_w_ctr_reg_6_), .B(w_mem_inst__abc_19396_new_n4807_), .C(w_mem_inst__abc_19396_new_n4809_), .Y(w_mem_inst__abc_19396_new_n4811_));
AOI21X1 AOI21X1_308 ( .A(w_mem_inst__abc_19396_new_n4809_), .B(w_mem_inst_w_ctr_reg_6_), .C(w_mem_inst__abc_19396_new_n4811_), .Y(w_mem_inst__0w_ctr_reg_6_0__6_));
AOI21X1 AOI21X1_31 ( .A(_abc_15497_new_n1175_), .B(_abc_15497_new_n1164_), .C(_abc_15497_new_n1174_), .Y(_abc_15497_new_n1205_));
AOI21X1 AOI21X1_32 ( .A(_abc_15497_new_n1197_), .B(_abc_15497_new_n1186_), .C(_abc_15497_new_n1196_), .Y(_abc_15497_new_n1206_));
AOI21X1 AOI21X1_33 ( .A(_abc_15497_new_n1158_), .B(_abc_15497_new_n1202_), .C(_abc_15497_new_n1209_), .Y(_abc_15497_new_n1210_));
AOI21X1 AOI21X1_34 ( .A(_abc_15497_new_n1271_), .B(_abc_15497_new_n1276_), .C(_abc_15497_new_n1277_), .Y(_abc_15497_new_n1278_));
AOI21X1 AOI21X1_35 ( .A(_abc_15497_new_n870__bF_buf0), .B(_abc_15497_new_n1269_), .C(_abc_15497_new_n1278_), .Y(_0H4_reg_31_0__29_));
AOI21X1 AOI21X1_36 ( .A(_abc_15497_new_n1263_), .B(_abc_15497_new_n1284_), .C(_abc_15497_new_n1283_), .Y(_abc_15497_new_n1285_));
AOI21X1 AOI21X1_37 ( .A(_abc_15497_new_n1310_), .B(_abc_15497_new_n1313_), .C(_abc_15497_new_n1312_), .Y(_abc_15497_new_n1318_));
AOI21X1 AOI21X1_38 ( .A(_abc_15497_new_n1358_), .B(_abc_15497_new_n1355_), .C(_abc_15497_new_n1354_), .Y(_abc_15497_new_n1362_));
AOI21X1 AOI21X1_39 ( .A(_abc_15497_new_n1376_), .B(_abc_15497_new_n1365_), .C(_abc_15497_new_n1375_), .Y(_abc_15497_new_n1384_));
AOI21X1 AOI21X1_4 ( .A(_abc_15497_new_n745_), .B(_abc_15497_new_n743_), .C(_abc_15497_new_n740_), .Y(_abc_15497_new_n746_));
AOI21X1 AOI21X1_40 ( .A(_abc_15497_new_n1400_), .B(_abc_15497_new_n1388_), .C(_abc_15497_new_n1399_), .Y(_abc_15497_new_n1408_));
AOI21X1 AOI21X1_41 ( .A(_abc_15497_new_n1427_), .B(_abc_15497_new_n1415_), .C(_abc_15497_new_n1426_), .Y(_abc_15497_new_n1432_));
AOI21X1 AOI21X1_42 ( .A(_abc_15497_new_n1423_), .B(_abc_15497_new_n1427_), .C(_abc_15497_new_n1433_), .Y(_abc_15497_new_n1434_));
AOI21X1 AOI21X1_43 ( .A(_abc_15497_new_n1449_), .B(_abc_15497_new_n1437_), .C(_abc_15497_new_n1448_), .Y(_abc_15497_new_n1454_));
AOI21X1 AOI21X1_44 ( .A(_abc_15497_new_n1409_), .B(_abc_15497_new_n1457_), .C(_abc_15497_new_n1455_), .Y(_abc_15497_new_n1458_));
AOI21X1 AOI21X1_45 ( .A(_abc_15497_new_n1460_), .B(_abc_15497_new_n1464_), .C(_abc_15497_new_n1463_), .Y(_abc_15497_new_n1467_));
AOI21X1 AOI21X1_46 ( .A(_abc_15497_new_n1471_), .B(_abc_15497_new_n1463_), .C(_abc_15497_new_n1470_), .Y(_abc_15497_new_n1478_));
AOI21X1 AOI21X1_47 ( .A(_abc_15497_new_n1460_), .B(_abc_15497_new_n1481_), .C(_abc_15497_new_n1479_), .Y(_abc_15497_new_n1482_));
AOI21X1 AOI21X1_48 ( .A(_abc_15497_new_n1483_), .B(_abc_15497_new_n1487_), .C(_abc_15497_new_n1486_), .Y(_abc_15497_new_n1493_));
AOI21X1 AOI21X1_49 ( .A(_abc_15497_new_n1497_), .B(_abc_15497_new_n1486_), .C(_abc_15497_new_n1496_), .Y(_abc_15497_new_n1505_));
AOI21X1 AOI21X1_5 ( .A(_abc_15497_new_n752_), .B(_abc_15497_new_n750_), .C(_abc_15497_new_n747_), .Y(_abc_15497_new_n753_));
AOI21X1 AOI21X1_50 ( .A(_abc_15497_new_n1460_), .B(_abc_15497_new_n1504_), .C(_abc_15497_new_n1506_), .Y(_abc_15497_new_n1507_));
AOI21X1 AOI21X1_51 ( .A(_abc_15497_new_n1508_), .B(_abc_15497_new_n1535_), .C(_abc_15497_new_n1534_), .Y(_abc_15497_new_n1536_));
AOI21X1 AOI21X1_52 ( .A(_abc_15497_new_n1460_), .B(_abc_15497_new_n1558_), .C(_abc_15497_new_n1556_), .Y(_abc_15497_new_n1559_));
AOI21X1 AOI21X1_53 ( .A(_abc_15497_new_n1574_), .B(_abc_15497_new_n1563_), .C(_abc_15497_new_n1573_), .Y(_abc_15497_new_n1582_));
AOI21X1 AOI21X1_54 ( .A(_abc_15497_new_n1560_), .B(_abc_15497_new_n1581_), .C(_abc_15497_new_n1583_), .Y(_abc_15497_new_n1584_));
AOI21X1 AOI21X1_55 ( .A(_abc_15497_new_n1598_), .B(_abc_15497_new_n1587_), .C(_abc_15497_new_n1597_), .Y(_abc_15497_new_n1607_));
AOI21X1 AOI21X1_56 ( .A(_abc_15497_new_n1619_), .B(_abc_15497_new_n1624_), .C(_abc_15497_new_n1625_), .Y(_abc_15497_new_n1626_));
AOI21X1 AOI21X1_57 ( .A(_abc_15497_new_n870__bF_buf3), .B(_abc_15497_new_n1617_), .C(_abc_15497_new_n1626_), .Y(_0H3_reg_31_0__29_));
AOI21X1 AOI21X1_58 ( .A(_abc_15497_new_n1610_), .B(_abc_15497_new_n1633_), .C(_abc_15497_new_n1632_), .Y(_abc_15497_new_n1634_));
AOI21X1 AOI21X1_59 ( .A(_abc_15497_new_n1758_), .B(_abc_15497_new_n1757_), .C(_abc_15497_new_n870__bF_buf0), .Y(_abc_15497_new_n1759_));
AOI21X1 AOI21X1_6 ( .A(_abc_15497_new_n774_), .B(_abc_15497_new_n776_), .C(_abc_15497_new_n767_), .Y(_abc_15497_new_n777_));
AOI21X1 AOI21X1_60 ( .A(_abc_15497_new_n1772_), .B(_abc_15497_new_n1781_), .C(_abc_15497_new_n1774_), .Y(_abc_15497_new_n1782_));
AOI21X1 AOI21X1_61 ( .A(_abc_15497_new_n1800_), .B(_abc_15497_new_n1804_), .C(_abc_15497_new_n1803_), .Y(_abc_15497_new_n1807_));
AOI21X1 AOI21X1_62 ( .A(_abc_15497_new_n1825_), .B(_abc_15497_new_n1822_), .C(_abc_15497_new_n1821_), .Y(_abc_15497_new_n1829_));
AOI21X1 AOI21X1_63 ( .A(_abc_15497_new_n1832_), .B(_abc_15497_new_n1821_), .C(_abc_15497_new_n1831_), .Y(_abc_15497_new_n1838_));
AOI21X1 AOI21X1_64 ( .A(_abc_15497_new_n1852_), .B(_abc_15497_new_n1842_), .C(_abc_15497_new_n1851_), .Y(_abc_15497_new_n1861_));
AOI21X1 AOI21X1_65 ( .A(_abc_15497_new_n1825_), .B(_abc_15497_new_n1864_), .C(_abc_15497_new_n1863_), .Y(_abc_15497_new_n1865_));
AOI21X1 AOI21X1_66 ( .A(_abc_15497_new_n1895_), .B(_abc_15497_new_n1877_), .C(_abc_15497_new_n1894_), .Y(_abc_15497_new_n1899_));
AOI21X1 AOI21X1_67 ( .A(_abc_15497_new_n1863_), .B(_abc_15497_new_n1902_), .C(_abc_15497_new_n1901_), .Y(_abc_15497_new_n1903_));
AOI21X1 AOI21X1_68 ( .A(_abc_15497_new_n1934_), .B(_abc_15497_new_n1930_), .C(_abc_15497_new_n1942_), .Y(_abc_15497_new_n1945_));
AOI21X1 AOI21X1_69 ( .A(_abc_15497_new_n1920_), .B(_abc_15497_new_n1909_), .C(_abc_15497_new_n1919_), .Y(_abc_15497_new_n1950_));
AOI21X1 AOI21X1_7 ( .A(_abc_15497_new_n782_), .B(_abc_15497_new_n758_), .C(_abc_15497_new_n754_), .Y(_abc_15497_new_n783_));
AOI21X1 AOI21X1_70 ( .A(_abc_15497_new_n1942_), .B(_abc_15497_new_n1931_), .C(_abc_15497_new_n1941_), .Y(_abc_15497_new_n1952_));
AOI21X1 AOI21X1_71 ( .A(_abc_15497_new_n1905_), .B(_abc_15497_new_n1955_), .C(_abc_15497_new_n1953_), .Y(_abc_15497_new_n1956_));
AOI21X1 AOI21X1_72 ( .A(_abc_15497_new_n1969_), .B(_abc_15497_new_n1959_), .C(_abc_15497_new_n1968_), .Y(_abc_15497_new_n1977_));
AOI21X1 AOI21X1_73 ( .A(_abc_15497_new_n1978_), .B(_abc_15497_new_n1982_), .C(_abc_15497_new_n1981_), .Y(_abc_15497_new_n1986_));
AOI21X1 AOI21X1_74 ( .A(_abc_15497_new_n1990_), .B(_abc_15497_new_n1981_), .C(_abc_15497_new_n1989_), .Y(_abc_15497_new_n1998_));
AOI21X1 AOI21X1_75 ( .A(_abc_15497_new_n1905_), .B(_abc_15497_new_n2002_), .C(_abc_15497_new_n2001_), .Y(_abc_15497_new_n2003_));
AOI21X1 AOI21X1_76 ( .A(_abc_15497_new_n2048_), .B(_abc_15497_new_n2026_), .C(_abc_15497_new_n2051_), .Y(_abc_15497_new_n2052_));
AOI21X1 AOI21X1_77 ( .A(_abc_15497_new_n2055_), .B(_abc_15497_new_n2056_), .C(_abc_15497_new_n2053_), .Y(_abc_15497_new_n2057_));
AOI21X1 AOI21X1_78 ( .A(_abc_15497_new_n2063_), .B(_abc_15497_new_n2068_), .C(_abc_15497_new_n870__bF_buf4), .Y(_abc_15497_new_n2070_));
AOI21X1 AOI21X1_79 ( .A(_abc_15497_new_n2053_), .B(_abc_15497_new_n2075_), .C(_abc_15497_new_n2074_), .Y(_abc_15497_new_n2076_));
AOI21X1 AOI21X1_8 ( .A(_abc_15497_new_n790_), .B(_abc_15497_new_n737_), .C(_abc_15497_new_n733_), .Y(_abc_15497_new_n791_));
AOI21X1 AOI21X1_80 ( .A(_abc_15497_new_n2099_), .B(_abc_15497_new_n2098_), .C(_abc_15497_new_n870__bF_buf10), .Y(_abc_15497_new_n2100_));
AOI21X1 AOI21X1_81 ( .A(_abc_15497_new_n2114_), .B(_abc_15497_new_n2116_), .C(_abc_15497_new_n2117_), .Y(_abc_15497_new_n2124_));
AOI21X1 AOI21X1_82 ( .A(_abc_15497_new_n2152_), .B(_abc_15497_new_n2145_), .C(_abc_15497_new_n870__bF_buf7), .Y(_abc_15497_new_n2156_));
AOI21X1 AOI21X1_83 ( .A(_abc_15497_new_n2163_), .B(_abc_15497_new_n2192_), .C(_abc_15497_new_n2190_), .Y(_abc_15497_new_n2193_));
AOI21X1 AOI21X1_84 ( .A(_abc_15497_new_n2163_), .B(_abc_15497_new_n2205_), .C(_abc_15497_new_n2210_), .Y(_abc_15497_new_n2233_));
AOI21X1 AOI21X1_85 ( .A(_abc_15497_new_n2224_), .B(_abc_15497_new_n2215_), .C(_abc_15497_new_n2223_), .Y(_abc_15497_new_n2234_));
AOI21X1 AOI21X1_86 ( .A(_abc_15497_new_n2246_), .B(_abc_15497_new_n2231_), .C(_abc_15497_new_n2245_), .Y(_abc_15497_new_n2249_));
AOI21X1 AOI21X1_87 ( .A(_abc_15497_new_n2210_), .B(_abc_15497_new_n2252_), .C(_abc_15497_new_n2251_), .Y(_abc_15497_new_n2253_));
AOI21X1 AOI21X1_88 ( .A(_abc_15497_new_n2272_), .B(_abc_15497_new_n2259_), .C(_abc_15497_new_n2271_), .Y(_abc_15497_new_n2280_));
AOI21X1 AOI21X1_89 ( .A(_abc_15497_new_n2298_), .B(_abc_15497_new_n2285_), .C(_abc_15497_new_n2297_), .Y(_abc_15497_new_n2306_));
AOI21X1 AOI21X1_9 ( .A(_abc_15497_new_n809_), .B(_abc_15497_new_n807_), .C(_abc_15497_new_n806_), .Y(_abc_15497_new_n810_));
AOI21X1 AOI21X1_90 ( .A(_abc_15497_new_n2255_), .B(_abc_15497_new_n2305_), .C(_abc_15497_new_n2307_), .Y(_abc_15497_new_n2308_));
AOI21X1 AOI21X1_91 ( .A(_abc_15497_new_n2329_), .B(_abc_15497_new_n2334_), .C(_abc_15497_new_n2333_), .Y(_abc_15497_new_n2338_));
AOI21X1 AOI21X1_92 ( .A(_abc_15497_new_n2348_), .B(_abc_15497_new_n2346_), .C(_abc_15497_new_n2351_), .Y(_abc_15497_new_n2352_));
AOI21X1 AOI21X1_93 ( .A(_abc_15497_new_n2255_), .B(_abc_15497_new_n2356_), .C(_abc_15497_new_n2354_), .Y(_abc_15497_new_n2357_));
AOI21X1 AOI21X1_94 ( .A(_abc_15497_new_n2374_), .B(_abc_15497_new_n2361_), .C(_abc_15497_new_n2373_), .Y(_abc_15497_new_n2381_));
AOI21X1 AOI21X1_95 ( .A(_abc_15497_new_n2397_), .B(_abc_15497_new_n2386_), .C(_abc_15497_new_n2396_), .Y(_abc_15497_new_n2405_));
AOI21X1 AOI21X1_96 ( .A(_abc_15497_new_n2404_), .B(_abc_15497_new_n2402_), .C(_abc_15497_new_n2406_), .Y(_abc_15497_new_n2407_));
AOI21X1 AOI21X1_97 ( .A(_abc_15497_new_n2408_), .B(_abc_15497_new_n2432_), .C(_abc_15497_new_n2431_), .Y(_abc_15497_new_n2433_));
AOI21X1 AOI21X1_98 ( .A(_abc_15497_new_n2759__bF_buf5), .B(_abc_15497_new_n2749_), .C(_abc_15497_new_n2743__bF_buf5), .Y(_abc_15497_new_n2760_));
AOI21X1 AOI21X1_99 ( .A(_abc_15497_new_n2740_), .B(_abc_15497_new_n2741_), .C(_abc_15497_new_n2738_), .Y(_abc_15497_new_n2781_));
AOI22X1 AOI22X1_1 ( .A(_abc_15497_new_n913_), .B(_abc_15497_new_n914_), .C(_abc_15497_new_n917_), .D(_abc_15497_new_n919_), .Y(_abc_15497_new_n920_));
AOI22X1 AOI22X1_10 ( .A(d_reg_7_), .B(round_ctr_inc_bF_buf1), .C(e_reg_7_), .D(_abc_15497_new_n1663__bF_buf4), .Y(_abc_15497_new_n1673_));
AOI22X1 AOI22X1_100 ( .A(round_ctr_inc_bF_buf8), .B(b_reg_4_), .C(c_reg_2_), .D(_abc_15497_new_n1663__bF_buf6), .Y(_abc_15497_new_n2646_));
AOI22X1 AOI22X1_101 ( .A(round_ctr_inc_bF_buf6), .B(b_reg_5_), .C(c_reg_3_), .D(_abc_15497_new_n1663__bF_buf5), .Y(_abc_15497_new_n2649_));
AOI22X1 AOI22X1_102 ( .A(round_ctr_inc_bF_buf4), .B(b_reg_6_), .C(c_reg_4_), .D(_abc_15497_new_n1663__bF_buf4), .Y(_abc_15497_new_n2652_));
AOI22X1 AOI22X1_103 ( .A(round_ctr_inc_bF_buf2), .B(b_reg_7_), .C(_abc_15497_new_n2654_), .D(_abc_15497_new_n1650__bF_buf2), .Y(_abc_15497_new_n2655_));
AOI22X1 AOI22X1_104 ( .A(round_ctr_inc_bF_buf1), .B(b_reg_8_), .C(_abc_15497_new_n2657_), .D(_abc_15497_new_n1650__bF_buf1), .Y(_abc_15497_new_n2658_));
AOI22X1 AOI22X1_105 ( .A(round_ctr_inc_bF_buf0), .B(b_reg_9_), .C(c_reg_7_), .D(_abc_15497_new_n1663__bF_buf3), .Y(_abc_15497_new_n2661_));
AOI22X1 AOI22X1_106 ( .A(round_ctr_inc_bF_buf12), .B(b_reg_10_), .C(_abc_15497_new_n1650__bF_buf0), .D(_abc_15497_new_n2663_), .Y(_abc_15497_new_n2664_));
AOI22X1 AOI22X1_107 ( .A(round_ctr_inc_bF_buf11), .B(b_reg_11_), .C(_abc_15497_new_n1650__bF_buf9), .D(_abc_15497_new_n2666_), .Y(_abc_15497_new_n2667_));
AOI22X1 AOI22X1_108 ( .A(round_ctr_inc_bF_buf10), .B(b_reg_12_), .C(_abc_15497_new_n2669_), .D(_abc_15497_new_n1650__bF_buf8), .Y(_abc_15497_new_n2670_));
AOI22X1 AOI22X1_109 ( .A(round_ctr_inc_bF_buf9), .B(b_reg_13_), .C(c_reg_11_), .D(_abc_15497_new_n1663__bF_buf2), .Y(_abc_15497_new_n2673_));
AOI22X1 AOI22X1_11 ( .A(d_reg_8_), .B(round_ctr_inc_bF_buf13), .C(_abc_15497_new_n1675_), .D(_abc_15497_new_n1650__bF_buf5), .Y(_abc_15497_new_n1676_));
AOI22X1 AOI22X1_110 ( .A(round_ctr_inc_bF_buf7), .B(b_reg_14_), .C(c_reg_12_), .D(_abc_15497_new_n1663__bF_buf1), .Y(_abc_15497_new_n2676_));
AOI22X1 AOI22X1_111 ( .A(round_ctr_inc_bF_buf5), .B(b_reg_15_), .C(_abc_15497_new_n1650__bF_buf7), .D(_abc_15497_new_n2678_), .Y(_abc_15497_new_n2679_));
AOI22X1 AOI22X1_112 ( .A(round_ctr_inc_bF_buf4), .B(b_reg_16_), .C(_abc_15497_new_n2681_), .D(_abc_15497_new_n1650__bF_buf6), .Y(_abc_15497_new_n2682_));
AOI22X1 AOI22X1_113 ( .A(round_ctr_inc_bF_buf3), .B(b_reg_17_), .C(c_reg_15_), .D(_abc_15497_new_n1663__bF_buf0), .Y(_abc_15497_new_n2685_));
AOI22X1 AOI22X1_114 ( .A(round_ctr_inc_bF_buf1), .B(b_reg_18_), .C(_abc_15497_new_n1650__bF_buf5), .D(_abc_15497_new_n2687_), .Y(_abc_15497_new_n2688_));
AOI22X1 AOI22X1_115 ( .A(round_ctr_inc_bF_buf0), .B(b_reg_19_), .C(c_reg_17_), .D(_abc_15497_new_n1663__bF_buf7), .Y(_abc_15497_new_n2691_));
AOI22X1 AOI22X1_116 ( .A(round_ctr_inc_bF_buf12), .B(b_reg_20_), .C(_abc_15497_new_n1650__bF_buf4), .D(_abc_15497_new_n2693_), .Y(_abc_15497_new_n2694_));
AOI22X1 AOI22X1_117 ( .A(round_ctr_inc_bF_buf11), .B(b_reg_21_), .C(c_reg_19_), .D(_abc_15497_new_n1663__bF_buf6), .Y(_abc_15497_new_n2697_));
AOI22X1 AOI22X1_118 ( .A(round_ctr_inc_bF_buf9), .B(b_reg_22_), .C(c_reg_20_), .D(_abc_15497_new_n1663__bF_buf5), .Y(_abc_15497_new_n2700_));
AOI22X1 AOI22X1_119 ( .A(round_ctr_inc_bF_buf7), .B(b_reg_23_), .C(c_reg_21_), .D(_abc_15497_new_n1663__bF_buf4), .Y(_abc_15497_new_n2703_));
AOI22X1 AOI22X1_12 ( .A(d_reg_9_), .B(round_ctr_inc_bF_buf12), .C(_abc_15497_new_n1650__bF_buf4), .D(_abc_15497_new_n1678_), .Y(_abc_15497_new_n1679_));
AOI22X1 AOI22X1_120 ( .A(round_ctr_inc_bF_buf5), .B(b_reg_24_), .C(_abc_15497_new_n1650__bF_buf3), .D(_abc_15497_new_n2705_), .Y(_abc_15497_new_n2706_));
AOI22X1 AOI22X1_121 ( .A(round_ctr_inc_bF_buf4), .B(b_reg_25_), .C(c_reg_23_), .D(_abc_15497_new_n1663__bF_buf3), .Y(_abc_15497_new_n2709_));
AOI22X1 AOI22X1_122 ( .A(round_ctr_inc_bF_buf2), .B(b_reg_26_), .C(_abc_15497_new_n1650__bF_buf2), .D(_abc_15497_new_n2711_), .Y(_abc_15497_new_n2712_));
AOI22X1 AOI22X1_123 ( .A(round_ctr_inc_bF_buf1), .B(b_reg_27_), .C(_abc_15497_new_n1650__bF_buf1), .D(_abc_15497_new_n2714_), .Y(_abc_15497_new_n2715_));
AOI22X1 AOI22X1_124 ( .A(round_ctr_inc_bF_buf0), .B(b_reg_28_), .C(_abc_15497_new_n1650__bF_buf0), .D(_abc_15497_new_n2717_), .Y(_abc_15497_new_n2718_));
AOI22X1 AOI22X1_125 ( .A(round_ctr_inc_bF_buf13), .B(b_reg_29_), .C(c_reg_27_), .D(_abc_15497_new_n1663__bF_buf2), .Y(_abc_15497_new_n2721_));
AOI22X1 AOI22X1_126 ( .A(round_ctr_inc_bF_buf11), .B(b_reg_30_), .C(c_reg_28_), .D(_abc_15497_new_n1663__bF_buf1), .Y(_abc_15497_new_n2724_));
AOI22X1 AOI22X1_127 ( .A(round_ctr_inc_bF_buf9), .B(b_reg_31_), .C(_abc_15497_new_n1650__bF_buf9), .D(_abc_15497_new_n2726_), .Y(_abc_15497_new_n2727_));
AOI22X1 AOI22X1_128 ( .A(round_ctr_inc_bF_buf8), .B(b_reg_0_), .C(_abc_15497_new_n1650__bF_buf8), .D(_abc_15497_new_n2729_), .Y(_abc_15497_new_n2730_));
AOI22X1 AOI22X1_129 ( .A(round_ctr_inc_bF_buf7), .B(b_reg_1_), .C(c_reg_31_), .D(_abc_15497_new_n1663__bF_buf0), .Y(_abc_15497_new_n2733_));
AOI22X1 AOI22X1_13 ( .A(d_reg_10_), .B(round_ctr_inc_bF_buf11), .C(_abc_15497_new_n1650__bF_buf3), .D(_abc_15497_new_n1681_), .Y(_abc_15497_new_n1682_));
AOI22X1 AOI22X1_130 ( .A(_abc_15497_new_n2735_), .B(_abc_15497_new_n2758_), .C(_abc_15497_new_n2752_), .D(_abc_15497_new_n2754_), .Y(_abc_15497_new_n2759_));
AOI22X1 AOI22X1_131 ( .A(_abc_15497_new_n2743__bF_buf4), .B(_abc_15497_new_n2745_), .C(_abc_15497_new_n2760_), .D(_abc_15497_new_n2757_), .Y(_abc_15497_new_n2761_));
AOI22X1 AOI22X1_132 ( .A(_abc_15497_new_n1308_), .B(_abc_15497_new_n2782_), .C(_abc_15497_new_n2784_), .D(_abc_15497_new_n2785_), .Y(_abc_15497_new_n2786_));
AOI22X1 AOI22X1_133 ( .A(_abc_15497_new_n2759__bF_buf4), .B(_abc_15497_new_n2784_), .C(_abc_15497_new_n2743__bF_buf2), .D(_abc_15497_new_n2788_), .Y(_abc_15497_new_n2789_));
AOI22X1 AOI22X1_134 ( .A(_abc_15497_new_n2761_), .B(_abc_15497_new_n2767_), .C(_abc_15497_new_n2810_), .D(_abc_15497_new_n2811_), .Y(_abc_15497_new_n2812_));
AOI22X1 AOI22X1_135 ( .A(_abc_15497_new_n2761_), .B(_abc_15497_new_n2767_), .C(_abc_15497_new_n2805_), .D(_abc_15497_new_n2808_), .Y(_abc_15497_new_n2815_));
AOI22X1 AOI22X1_136 ( .A(_abc_15497_new_n2823_), .B(_abc_15497_new_n1650__bF_buf6), .C(a_reg_1_), .D(_abc_15497_new_n1663__bF_buf7), .Y(_abc_15497_new_n2824_));
AOI22X1 AOI22X1_137 ( .A(_abc_15497_new_n2829_), .B(_abc_15497_new_n2830_), .C(_abc_15497_new_n2832_), .D(_abc_15497_new_n2833_), .Y(_abc_15497_new_n2834_));
AOI22X1 AOI22X1_138 ( .A(_abc_15497_new_n2759__bF_buf3), .B(_abc_15497_new_n2832_), .C(_abc_15497_new_n2743__bF_buf1), .D(_abc_15497_new_n2836_), .Y(_abc_15497_new_n2837_));
AOI22X1 AOI22X1_139 ( .A(_abc_15497_new_n2736_), .B(_abc_15497_new_n2863_), .C(_abc_15497_new_n2865_), .D(_abc_15497_new_n2864_), .Y(_abc_15497_new_n2866_));
AOI22X1 AOI22X1_14 ( .A(d_reg_11_), .B(round_ctr_inc_bF_buf10), .C(_abc_15497_new_n1650__bF_buf2), .D(_abc_15497_new_n1685_), .Y(_abc_15497_new_n1686_));
AOI22X1 AOI22X1_140 ( .A(_abc_15497_new_n2880_), .B(_abc_15497_new_n1650__bF_buf5), .C(a_reg_2_), .D(_abc_15497_new_n1663__bF_buf6), .Y(_abc_15497_new_n2881_));
AOI22X1 AOI22X1_141 ( .A(_abc_15497_new_n2759__bF_buf2), .B(_abc_15497_new_n2891_), .C(_abc_15497_new_n2743__bF_buf0), .D(_abc_15497_new_n2895_), .Y(_abc_15497_new_n2896_));
AOI22X1 AOI22X1_142 ( .A(_abc_15497_new_n2937_), .B(_abc_15497_new_n1650__bF_buf4), .C(a_reg_3_), .D(_abc_15497_new_n1663__bF_buf5), .Y(_abc_15497_new_n2938_));
AOI22X1 AOI22X1_143 ( .A(_abc_15497_new_n2759__bF_buf1), .B(_abc_15497_new_n2949_), .C(_abc_15497_new_n2743__bF_buf5), .D(_abc_15497_new_n2952_), .Y(_abc_15497_new_n2953_));
AOI22X1 AOI22X1_144 ( .A(_abc_15497_new_n2999_), .B(_abc_15497_new_n1650__bF_buf3), .C(a_reg_4_), .D(_abc_15497_new_n1663__bF_buf4), .Y(_abc_15497_new_n3000_));
AOI22X1 AOI22X1_145 ( .A(_abc_15497_new_n1343_), .B(_abc_15497_new_n3008_), .C(_abc_15497_new_n3010_), .D(_abc_15497_new_n3011_), .Y(_abc_15497_new_n3012_));
AOI22X1 AOI22X1_146 ( .A(_abc_15497_new_n2759__bF_buf0), .B(_abc_15497_new_n3010_), .C(_abc_15497_new_n2743__bF_buf4), .D(_abc_15497_new_n3014_), .Y(_abc_15497_new_n3015_));
AOI22X1 AOI22X1_147 ( .A(_abc_15497_new_n3055_), .B(_abc_15497_new_n1650__bF_buf2), .C(a_reg_5_), .D(_abc_15497_new_n1663__bF_buf3), .Y(_abc_15497_new_n3056_));
AOI22X1 AOI22X1_148 ( .A(_abc_15497_new_n1357_), .B(_abc_15497_new_n3066_), .C(_abc_15497_new_n3068_), .D(_abc_15497_new_n3069_), .Y(_abc_15497_new_n3070_));
AOI22X1 AOI22X1_149 ( .A(_abc_15497_new_n2759__bF_buf5), .B(_abc_15497_new_n3068_), .C(_abc_15497_new_n2743__bF_buf3), .D(_abc_15497_new_n3072_), .Y(_abc_15497_new_n3073_));
AOI22X1 AOI22X1_15 ( .A(d_reg_12_), .B(round_ctr_inc_bF_buf9), .C(_abc_15497_new_n1650__bF_buf1), .D(_abc_15497_new_n1688_), .Y(_abc_15497_new_n1689_));
AOI22X1 AOI22X1_150 ( .A(_abc_15497_new_n3113_), .B(_abc_15497_new_n1650__bF_buf1), .C(a_reg_6_), .D(_abc_15497_new_n1663__bF_buf2), .Y(_abc_15497_new_n3114_));
AOI22X1 AOI22X1_151 ( .A(_abc_15497_new_n1353_), .B(_abc_15497_new_n3120_), .C(_abc_15497_new_n3123_), .D(_abc_15497_new_n3122_), .Y(_abc_15497_new_n3124_));
AOI22X1 AOI22X1_152 ( .A(_abc_15497_new_n2759__bF_buf4), .B(_abc_15497_new_n3122_), .C(_abc_15497_new_n2743__bF_buf2), .D(_abc_15497_new_n3126_), .Y(_abc_15497_new_n3146_));
AOI22X1 AOI22X1_153 ( .A(_abc_15497_new_n1650__bF_buf0), .B(_abc_15497_new_n3164_), .C(round_ctr_inc_bF_buf1), .D(_abc_15497_new_n3163_), .Y(_abc_15497_new_n3165_));
AOI22X1 AOI22X1_154 ( .A(_abc_15497_new_n1364_), .B(_abc_15497_new_n3170_), .C(_abc_15497_new_n3172_), .D(_abc_15497_new_n3173_), .Y(_abc_15497_new_n3174_));
AOI22X1 AOI22X1_155 ( .A(_abc_15497_new_n2759__bF_buf3), .B(_abc_15497_new_n3172_), .C(_abc_15497_new_n2743__bF_buf1), .D(_abc_15497_new_n3176_), .Y(_abc_15497_new_n3177_));
AOI22X1 AOI22X1_156 ( .A(_abc_15497_new_n3175_), .B(_abc_15497_new_n3177_), .C(_abc_15497_new_n3188_), .D(_abc_15497_new_n3187_), .Y(_abc_15497_new_n3189_));
AOI22X1 AOI22X1_157 ( .A(_abc_15497_new_n1374_), .B(_abc_15497_new_n3235_), .C(_abc_15497_new_n3256_), .D(_abc_15497_new_n3255_), .Y(_abc_15497_new_n3257_));
AOI22X1 AOI22X1_158 ( .A(_abc_15497_new_n3267_), .B(_abc_15497_new_n3266_), .C(_abc_15497_new_n3191_), .D(_abc_15497_new_n3198_), .Y(_abc_15497_new_n3268_));
AOI22X1 AOI22X1_159 ( .A(_abc_15497_new_n1650__bF_buf8), .B(_abc_15497_new_n3224_), .C(round_ctr_inc_bF_buf0), .D(_abc_15497_new_n3280_), .Y(_abc_15497_new_n3281_));
AOI22X1 AOI22X1_16 ( .A(d_reg_13_), .B(round_ctr_inc_bF_buf8), .C(e_reg_13_), .D(_abc_15497_new_n1663__bF_buf3), .Y(_abc_15497_new_n1692_));
AOI22X1 AOI22X1_160 ( .A(_abc_15497_new_n3290_), .B(_abc_15497_new_n3291_), .C(_abc_15497_new_n3293_), .D(_abc_15497_new_n3294_), .Y(_abc_15497_new_n3295_));
AOI22X1 AOI22X1_161 ( .A(_abc_15497_new_n2759__bF_buf5), .B(_abc_15497_new_n3293_), .C(_abc_15497_new_n2743__bF_buf0), .D(_abc_15497_new_n3297_), .Y(_abc_15497_new_n3298_));
AOI22X1 AOI22X1_162 ( .A(_abc_15497_new_n3253_), .B(_abc_15497_new_n3259_), .C(_abc_15497_new_n3324_), .D(_abc_15497_new_n3325_), .Y(_abc_15497_new_n3326_));
AOI22X1 AOI22X1_163 ( .A(_abc_15497_new_n3345_), .B(_abc_15497_new_n1650__bF_buf7), .C(a_reg_10_), .D(_abc_15497_new_n1663__bF_buf1), .Y(_abc_15497_new_n3346_));
AOI22X1 AOI22X1_164 ( .A(_abc_15497_new_n1398_), .B(_abc_15497_new_n3352_), .C(_abc_15497_new_n3355_), .D(_abc_15497_new_n3354_), .Y(_abc_15497_new_n3356_));
AOI22X1 AOI22X1_165 ( .A(_abc_15497_new_n2759__bF_buf1), .B(_abc_15497_new_n3354_), .C(_abc_15497_new_n2743__bF_buf5), .D(_abc_15497_new_n3358_), .Y(_abc_15497_new_n3359_));
AOI22X1 AOI22X1_166 ( .A(_abc_15497_new_n2735_), .B(_abc_15497_new_n3393_), .C(_abc_15497_new_n3387_), .D(_abc_15497_new_n3388_), .Y(_abc_15497_new_n3394_));
AOI22X1 AOI22X1_167 ( .A(_abc_15497_new_n2752_), .B(_abc_15497_new_n2754_), .C(_abc_15497_new_n3385_), .D(_abc_15497_new_n3380_), .Y(_abc_15497_new_n3395_));
AOI22X1 AOI22X1_168 ( .A(_abc_15497_new_n3400_), .B(_abc_15497_new_n1650__bF_buf6), .C(a_reg_11_), .D(_abc_15497_new_n1663__bF_buf0), .Y(_abc_15497_new_n3401_));
AOI22X1 AOI22X1_169 ( .A(_abc_15497_new_n1414_), .B(_abc_15497_new_n3419_), .C(_abc_15497_new_n3423_), .D(_abc_15497_new_n3421_), .Y(_abc_15497_new_n3424_));
AOI22X1 AOI22X1_17 ( .A(d_reg_14_), .B(round_ctr_inc_bF_buf6), .C(_abc_15497_new_n1694_), .D(_abc_15497_new_n1650__bF_buf0), .Y(_abc_15497_new_n1695_));
AOI22X1 AOI22X1_170 ( .A(_abc_15497_new_n2759__bF_buf5), .B(_abc_15497_new_n3421_), .C(_abc_15497_new_n2743__bF_buf4), .D(_abc_15497_new_n3426_), .Y(_abc_15497_new_n3427_));
AOI22X1 AOI22X1_171 ( .A(_abc_15497_new_n3475_), .B(_abc_15497_new_n1650__bF_buf5), .C(a_reg_12_), .D(_abc_15497_new_n1663__bF_buf7), .Y(_abc_15497_new_n3476_));
AOI22X1 AOI22X1_172 ( .A(_abc_15497_new_n3443_), .B(_abc_15497_new_n3449_), .C(_abc_15497_new_n3514_), .D(_abc_15497_new_n3513_), .Y(_abc_15497_new_n3515_));
AOI22X1 AOI22X1_173 ( .A(_abc_15497_new_n3508_), .B(_abc_15497_new_n3505_), .C(_abc_15497_new_n3579_), .D(_abc_15497_new_n3580_), .Y(_abc_15497_new_n3581_));
AOI22X1 AOI22X1_174 ( .A(_abc_15497_new_n2759__bF_buf3), .B(_abc_15497_new_n3583_), .C(_abc_15497_new_n2743__bF_buf3), .D(_abc_15497_new_n3490_), .Y(_abc_15497_new_n3584_));
AOI22X1 AOI22X1_175 ( .A(_abc_15497_new_n3600_), .B(_abc_15497_new_n1650__bF_buf3), .C(a_reg_14_), .D(_abc_15497_new_n1663__bF_buf6), .Y(_abc_15497_new_n3601_));
AOI22X1 AOI22X1_176 ( .A(_abc_15497_new_n2759__bF_buf0), .B(_abc_15497_new_n3635_), .C(_abc_15497_new_n2743__bF_buf1), .D(_abc_15497_new_n3617_), .Y(_abc_15497_new_n3638_));
AOI22X1 AOI22X1_177 ( .A(_abc_15497_new_n3574_), .B(_abc_15497_new_n3571_), .C(_abc_15497_new_n3645_), .D(_abc_15497_new_n3644_), .Y(_abc_15497_new_n3646_));
AOI22X1 AOI22X1_178 ( .A(_abc_15497_new_n2759__bF_buf5), .B(_abc_15497_new_n3552_), .C(_abc_15497_new_n2743__bF_buf5), .D(_abc_15497_new_n3554_), .Y(_abc_15497_new_n3648_));
AOI22X1 AOI22X1_179 ( .A(_abc_15497_new_n3665_), .B(_abc_15497_new_n1650__bF_buf2), .C(a_reg_15_), .D(_abc_15497_new_n1663__bF_buf5), .Y(_abc_15497_new_n3666_));
AOI22X1 AOI22X1_18 ( .A(d_reg_15_), .B(round_ctr_inc_bF_buf5), .C(e_reg_15_), .D(_abc_15497_new_n1663__bF_buf2), .Y(_abc_15497_new_n1698_));
AOI22X1 AOI22X1_180 ( .A(_abc_15497_new_n2759__bF_buf4), .B(_abc_15497_new_n3688_), .C(_abc_15497_new_n2743__bF_buf3), .D(_abc_15497_new_n3687_), .Y(_abc_15497_new_n3689_));
AOI22X1 AOI22X1_181 ( .A(_abc_15497_new_n2759__bF_buf3), .B(_abc_15497_new_n3730_), .C(_abc_15497_new_n2743__bF_buf2), .D(_abc_15497_new_n3733_), .Y(_abc_15497_new_n3734_));
AOI22X1 AOI22X1_182 ( .A(_abc_15497_new_n1650__bF_buf9), .B(_abc_15497_new_n2290_), .C(a_reg_18_), .D(_abc_15497_new_n1663__bF_buf4), .Y(_abc_15497_new_n3822_));
AOI22X1 AOI22X1_183 ( .A(_abc_15497_new_n3867_), .B(_abc_15497_new_n1650__bF_buf8), .C(a_reg_19_), .D(_abc_15497_new_n1663__bF_buf3), .Y(_abc_15497_new_n3868_));
AOI22X1 AOI22X1_184 ( .A(_abc_15497_new_n3860_), .B(_abc_15497_new_n3863_), .C(_abc_15497_new_n3815_), .D(_abc_15497_new_n3817_), .Y(_abc_15497_new_n3883_));
AOI22X1 AOI22X1_185 ( .A(_abc_15497_new_n2759__bF_buf0), .B(_abc_15497_new_n3900_), .C(_abc_15497_new_n2743__bF_buf1), .D(_abc_15497_new_n3899_), .Y(_abc_15497_new_n3901_));
AOI22X1 AOI22X1_186 ( .A(_abc_15497_new_n3932_), .B(_abc_15497_new_n1650__bF_buf7), .C(a_reg_20_), .D(_abc_15497_new_n1663__bF_buf2), .Y(_abc_15497_new_n3933_));
AOI22X1 AOI22X1_187 ( .A(_abc_15497_new_n2759__bF_buf5), .B(_abc_15497_new_n3951_), .C(_abc_15497_new_n2743__bF_buf0), .D(_abc_15497_new_n3950_), .Y(_abc_15497_new_n3952_));
AOI22X1 AOI22X1_188 ( .A(_abc_15497_new_n3983_), .B(_abc_15497_new_n1650__bF_buf6), .C(a_reg_21_), .D(_abc_15497_new_n1663__bF_buf1), .Y(_abc_15497_new_n3984_));
AOI22X1 AOI22X1_189 ( .A(_abc_15497_new_n3923_), .B(_abc_15497_new_n3927_), .C(_abc_15497_new_n3974_), .D(_abc_15497_new_n3978_), .Y(_abc_15497_new_n3986_));
AOI22X1 AOI22X1_19 ( .A(d_reg_16_), .B(round_ctr_inc_bF_buf3), .C(_abc_15497_new_n1650__bF_buf9), .D(_abc_15497_new_n1700_), .Y(_abc_15497_new_n1701_));
AOI22X1 AOI22X1_190 ( .A(_abc_15497_new_n2759__bF_buf4), .B(_abc_15497_new_n4006_), .C(_abc_15497_new_n2743__bF_buf5), .D(_abc_15497_new_n4004_), .Y(_abc_15497_new_n4007_));
AOI22X1 AOI22X1_191 ( .A(_abc_15497_new_n1650__bF_buf5), .B(_abc_15497_new_n4038_), .C(a_reg_22_), .D(_abc_15497_new_n1663__bF_buf0), .Y(_abc_15497_new_n4039_));
AOI22X1 AOI22X1_192 ( .A(_abc_15497_new_n2759__bF_buf3), .B(_abc_15497_new_n4053_), .C(_abc_15497_new_n2743__bF_buf4), .D(_abc_15497_new_n4056_), .Y(_abc_15497_new_n4057_));
AOI22X1 AOI22X1_193 ( .A(_abc_15497_new_n4094_), .B(_abc_15497_new_n1650__bF_buf4), .C(a_reg_23_), .D(_abc_15497_new_n1663__bF_buf7), .Y(_abc_15497_new_n4095_));
AOI22X1 AOI22X1_194 ( .A(_abc_15497_new_n4033_), .B(_abc_15497_new_n4029_), .C(_abc_15497_new_n4084_), .D(_abc_15497_new_n4088_), .Y(_abc_15497_new_n4097_));
AOI22X1 AOI22X1_195 ( .A(_abc_15497_new_n2759__bF_buf2), .B(_abc_15497_new_n4111_), .C(_abc_15497_new_n2743__bF_buf3), .D(_abc_15497_new_n4115_), .Y(_abc_15497_new_n4116_));
AOI22X1 AOI22X1_196 ( .A(_abc_15497_new_n2759__bF_buf0), .B(_abc_15497_new_n4157_), .C(_abc_15497_new_n2743__bF_buf2), .D(_abc_15497_new_n4160_), .Y(_abc_15497_new_n4161_));
AOI22X1 AOI22X1_197 ( .A(_abc_15497_new_n1650__bF_buf2), .B(_abc_15497_new_n4184_), .C(a_reg_25_), .D(_abc_15497_new_n1663__bF_buf6), .Y(_abc_15497_new_n4185_));
AOI22X1 AOI22X1_198 ( .A(_abc_15497_new_n2743__bF_buf1), .B(_abc_15497_new_n4200_), .C(_abc_15497_new_n2759__bF_buf5), .D(_abc_15497_new_n4202_), .Y(_abc_15497_new_n4203_));
AOI22X1 AOI22X1_199 ( .A(_abc_15497_new_n2743__bF_buf0), .B(_abc_15497_new_n4247_), .C(_abc_15497_new_n2756__bF_buf3), .D(_abc_15497_new_n4246_), .Y(_abc_15497_new_n4248_));
AOI22X1 AOI22X1_2 ( .A(_abc_15497_new_n1544_), .B(_abc_15497_new_n1552_), .C(_abc_15497_new_n1534_), .D(_abc_15497_new_n1553_), .Y(_abc_15497_new_n1554_));
AOI22X1 AOI22X1_20 ( .A(d_reg_17_), .B(round_ctr_inc_bF_buf2), .C(_abc_15497_new_n1703_), .D(_abc_15497_new_n1650__bF_buf8), .Y(_abc_15497_new_n1704_));
AOI22X1 AOI22X1_200 ( .A(_abc_15497_new_n4266_), .B(_abc_15497_new_n1650__bF_buf0), .C(a_reg_27_), .D(_abc_15497_new_n1663__bF_buf5), .Y(_abc_15497_new_n4267_));
AOI22X1 AOI22X1_201 ( .A(_abc_15497_new_n4286_), .B(_abc_15497_new_n2743__bF_buf5), .C(_abc_15497_new_n2759__bF_buf3), .D(_abc_15497_new_n4287_), .Y(_abc_15497_new_n4288_));
AOI22X1 AOI22X1_202 ( .A(_abc_15497_new_n4321_), .B(_abc_15497_new_n1650__bF_buf9), .C(a_reg_28_), .D(_abc_15497_new_n1663__bF_buf4), .Y(_abc_15497_new_n4322_));
AOI22X1 AOI22X1_203 ( .A(_abc_15497_new_n1650__bF_buf8), .B(_abc_15497_new_n4362_), .C(a_reg_29_), .D(_abc_15497_new_n1663__bF_buf3), .Y(_abc_15497_new_n4363_));
AOI22X1 AOI22X1_204 ( .A(_abc_15497_new_n1650__bF_buf7), .B(_abc_15497_new_n4403_), .C(a_reg_30_), .D(_abc_15497_new_n1663__bF_buf2), .Y(_abc_15497_new_n4404_));
AOI22X1 AOI22X1_205 ( .A(_abc_15497_new_n4438_), .B(_abc_15497_new_n1650__bF_buf6), .C(a_reg_31_), .D(_abc_15497_new_n1663__bF_buf1), .Y(_abc_15497_new_n4439_));
AOI22X1 AOI22X1_206 ( .A(_abc_15497_new_n4442_), .B(_abc_15497_new_n4443_), .C(_abc_15497_new_n4456_), .D(_abc_15497_new_n4455_), .Y(_0round_ctr_reg_6_0__1_));
AOI22X1 AOI22X1_207 ( .A(round_ctr_inc_bF_buf7), .B(_abc_15497_new_n4459_), .C(round_ctr_reg_2_), .D(_abc_15497_new_n1663__bF_buf7), .Y(_abc_15497_new_n4460_));
AOI22X1 AOI22X1_208 ( .A(_abc_15497_new_n870__bF_buf8), .B(_abc_15497_new_n4582_), .C(_abc_15497_new_n4586_), .D(_abc_15497_new_n4585_), .Y(_0H2_reg_31_0__23_));
AOI22X1 AOI22X1_209 ( .A(w_mem_inst__abc_19396_new_n1625__bF_buf4), .B(w_mem_inst_w_mem_9__0_), .C(w_mem_inst_w_mem_10__0_), .D(w_mem_inst__abc_19396_new_n1628__bF_buf4), .Y(w_mem_inst__abc_19396_new_n1629_));
AOI22X1 AOI22X1_21 ( .A(d_reg_18_), .B(round_ctr_inc_bF_buf1), .C(_abc_15497_new_n1650__bF_buf7), .D(_abc_15497_new_n1706_), .Y(_abc_15497_new_n1707_));
AOI22X1 AOI22X1_210 ( .A(w_mem_inst__abc_19396_new_n1630__bF_buf4), .B(w_mem_inst_w_mem_4__0_), .C(w_mem_inst_w_mem_6__0_), .D(w_mem_inst__abc_19396_new_n1631__bF_buf4), .Y(w_mem_inst__abc_19396_new_n1632_));
AOI22X1 AOI22X1_211 ( .A(w_mem_inst__abc_19396_new_n1637__bF_buf4), .B(w_mem_inst_w_mem_3__0_), .C(w_mem_inst_w_mem_14__0_), .D(w_mem_inst__abc_19396_new_n1638__bF_buf4), .Y(w_mem_inst__abc_19396_new_n1639_));
AOI22X1 AOI22X1_212 ( .A(w_mem_inst__abc_19396_new_n1587__bF_buf4), .B(w_mem_inst__abc_19396_new_n1590_), .C(w_mem_inst__abc_19396_new_n1616_), .D(w_mem_inst__abc_19396_new_n1641_), .Y(w_0_));
AOI22X1 AOI22X1_213 ( .A(w_mem_inst__abc_19396_new_n1625__bF_buf3), .B(w_mem_inst_w_mem_9__1_), .C(w_mem_inst_w_mem_10__1_), .D(w_mem_inst__abc_19396_new_n1628__bF_buf3), .Y(w_mem_inst__abc_19396_new_n1659_));
AOI22X1 AOI22X1_214 ( .A(w_mem_inst__abc_19396_new_n1630__bF_buf3), .B(w_mem_inst_w_mem_4__1_), .C(w_mem_inst_w_mem_6__1_), .D(w_mem_inst__abc_19396_new_n1631__bF_buf3), .Y(w_mem_inst__abc_19396_new_n1660_));
AOI22X1 AOI22X1_215 ( .A(w_mem_inst__abc_19396_new_n1637__bF_buf3), .B(w_mem_inst_w_mem_3__1_), .C(w_mem_inst_w_mem_14__1_), .D(w_mem_inst__abc_19396_new_n1638__bF_buf3), .Y(w_mem_inst__abc_19396_new_n1664_));
AOI22X1 AOI22X1_216 ( .A(w_mem_inst__abc_19396_new_n1587__bF_buf3), .B(w_mem_inst__abc_19396_new_n1645_), .C(w_mem_inst__abc_19396_new_n1654_), .D(w_mem_inst__abc_19396_new_n1666_), .Y(w_1_));
AOI22X1 AOI22X1_217 ( .A(w_mem_inst__abc_19396_new_n1625__bF_buf2), .B(w_mem_inst_w_mem_9__2_), .C(w_mem_inst_w_mem_10__2_), .D(w_mem_inst__abc_19396_new_n1628__bF_buf2), .Y(w_mem_inst__abc_19396_new_n1684_));
AOI22X1 AOI22X1_218 ( .A(w_mem_inst__abc_19396_new_n1630__bF_buf2), .B(w_mem_inst_w_mem_4__2_), .C(w_mem_inst_w_mem_6__2_), .D(w_mem_inst__abc_19396_new_n1631__bF_buf2), .Y(w_mem_inst__abc_19396_new_n1685_));
AOI22X1 AOI22X1_219 ( .A(w_mem_inst__abc_19396_new_n1637__bF_buf2), .B(w_mem_inst_w_mem_3__2_), .C(w_mem_inst_w_mem_14__2_), .D(w_mem_inst__abc_19396_new_n1638__bF_buf2), .Y(w_mem_inst__abc_19396_new_n1689_));
AOI22X1 AOI22X1_22 ( .A(d_reg_19_), .B(round_ctr_inc_bF_buf0), .C(_abc_15497_new_n1650__bF_buf6), .D(_abc_15497_new_n1709_), .Y(_abc_15497_new_n1710_));
AOI22X1 AOI22X1_220 ( .A(w_mem_inst__abc_19396_new_n1587__bF_buf2), .B(w_mem_inst__abc_19396_new_n1670_), .C(w_mem_inst__abc_19396_new_n1679_), .D(w_mem_inst__abc_19396_new_n1691_), .Y(w_2_));
AOI22X1 AOI22X1_221 ( .A(w_mem_inst__abc_19396_new_n1625__bF_buf1), .B(w_mem_inst_w_mem_9__3_), .C(w_mem_inst_w_mem_10__3_), .D(w_mem_inst__abc_19396_new_n1628__bF_buf1), .Y(w_mem_inst__abc_19396_new_n1709_));
AOI22X1 AOI22X1_222 ( .A(w_mem_inst__abc_19396_new_n1630__bF_buf1), .B(w_mem_inst_w_mem_4__3_), .C(w_mem_inst_w_mem_6__3_), .D(w_mem_inst__abc_19396_new_n1631__bF_buf1), .Y(w_mem_inst__abc_19396_new_n1710_));
AOI22X1 AOI22X1_223 ( .A(w_mem_inst__abc_19396_new_n1637__bF_buf1), .B(w_mem_inst_w_mem_3__3_), .C(w_mem_inst_w_mem_14__3_), .D(w_mem_inst__abc_19396_new_n1638__bF_buf1), .Y(w_mem_inst__abc_19396_new_n1714_));
AOI22X1 AOI22X1_224 ( .A(w_mem_inst__abc_19396_new_n1587__bF_buf1), .B(w_mem_inst__abc_19396_new_n1695_), .C(w_mem_inst__abc_19396_new_n1704_), .D(w_mem_inst__abc_19396_new_n1716_), .Y(w_3_));
AOI22X1 AOI22X1_225 ( .A(w_mem_inst__abc_19396_new_n1625__bF_buf0), .B(w_mem_inst_w_mem_9__4_), .C(w_mem_inst_w_mem_10__4_), .D(w_mem_inst__abc_19396_new_n1628__bF_buf0), .Y(w_mem_inst__abc_19396_new_n1734_));
AOI22X1 AOI22X1_226 ( .A(w_mem_inst__abc_19396_new_n1630__bF_buf0), .B(w_mem_inst_w_mem_4__4_), .C(w_mem_inst_w_mem_6__4_), .D(w_mem_inst__abc_19396_new_n1631__bF_buf0), .Y(w_mem_inst__abc_19396_new_n1735_));
AOI22X1 AOI22X1_227 ( .A(w_mem_inst__abc_19396_new_n1637__bF_buf0), .B(w_mem_inst_w_mem_3__4_), .C(w_mem_inst_w_mem_14__4_), .D(w_mem_inst__abc_19396_new_n1638__bF_buf0), .Y(w_mem_inst__abc_19396_new_n1739_));
AOI22X1 AOI22X1_228 ( .A(w_mem_inst__abc_19396_new_n1587__bF_buf0), .B(w_mem_inst__abc_19396_new_n1720_), .C(w_mem_inst__abc_19396_new_n1729_), .D(w_mem_inst__abc_19396_new_n1741_), .Y(w_4_));
AOI22X1 AOI22X1_229 ( .A(w_mem_inst__abc_19396_new_n1625__bF_buf4), .B(w_mem_inst_w_mem_9__5_), .C(w_mem_inst_w_mem_10__5_), .D(w_mem_inst__abc_19396_new_n1628__bF_buf4), .Y(w_mem_inst__abc_19396_new_n1759_));
AOI22X1 AOI22X1_23 ( .A(d_reg_20_), .B(round_ctr_inc_bF_buf13), .C(_abc_15497_new_n1712_), .D(_abc_15497_new_n1650__bF_buf5), .Y(_abc_15497_new_n1713_));
AOI22X1 AOI22X1_230 ( .A(w_mem_inst__abc_19396_new_n1630__bF_buf4), .B(w_mem_inst_w_mem_4__5_), .C(w_mem_inst_w_mem_6__5_), .D(w_mem_inst__abc_19396_new_n1631__bF_buf4), .Y(w_mem_inst__abc_19396_new_n1760_));
AOI22X1 AOI22X1_231 ( .A(w_mem_inst__abc_19396_new_n1637__bF_buf4), .B(w_mem_inst_w_mem_3__5_), .C(w_mem_inst_w_mem_14__5_), .D(w_mem_inst__abc_19396_new_n1638__bF_buf4), .Y(w_mem_inst__abc_19396_new_n1764_));
AOI22X1 AOI22X1_232 ( .A(w_mem_inst__abc_19396_new_n1587__bF_buf4), .B(w_mem_inst__abc_19396_new_n1745_), .C(w_mem_inst__abc_19396_new_n1754_), .D(w_mem_inst__abc_19396_new_n1766_), .Y(w_5_));
AOI22X1 AOI22X1_233 ( .A(w_mem_inst__abc_19396_new_n1625__bF_buf3), .B(w_mem_inst_w_mem_9__6_), .C(w_mem_inst_w_mem_10__6_), .D(w_mem_inst__abc_19396_new_n1628__bF_buf3), .Y(w_mem_inst__abc_19396_new_n1784_));
AOI22X1 AOI22X1_234 ( .A(w_mem_inst__abc_19396_new_n1630__bF_buf3), .B(w_mem_inst_w_mem_4__6_), .C(w_mem_inst_w_mem_6__6_), .D(w_mem_inst__abc_19396_new_n1631__bF_buf3), .Y(w_mem_inst__abc_19396_new_n1785_));
AOI22X1 AOI22X1_235 ( .A(w_mem_inst__abc_19396_new_n1637__bF_buf3), .B(w_mem_inst_w_mem_3__6_), .C(w_mem_inst_w_mem_14__6_), .D(w_mem_inst__abc_19396_new_n1638__bF_buf3), .Y(w_mem_inst__abc_19396_new_n1789_));
AOI22X1 AOI22X1_236 ( .A(w_mem_inst__abc_19396_new_n1587__bF_buf3), .B(w_mem_inst__abc_19396_new_n1770_), .C(w_mem_inst__abc_19396_new_n1779_), .D(w_mem_inst__abc_19396_new_n1791_), .Y(w_6_));
AOI22X1 AOI22X1_237 ( .A(w_mem_inst__abc_19396_new_n1625__bF_buf2), .B(w_mem_inst_w_mem_9__7_), .C(w_mem_inst_w_mem_10__7_), .D(w_mem_inst__abc_19396_new_n1628__bF_buf2), .Y(w_mem_inst__abc_19396_new_n1809_));
AOI22X1 AOI22X1_238 ( .A(w_mem_inst__abc_19396_new_n1630__bF_buf2), .B(w_mem_inst_w_mem_4__7_), .C(w_mem_inst_w_mem_6__7_), .D(w_mem_inst__abc_19396_new_n1631__bF_buf2), .Y(w_mem_inst__abc_19396_new_n1810_));
AOI22X1 AOI22X1_239 ( .A(w_mem_inst__abc_19396_new_n1637__bF_buf2), .B(w_mem_inst_w_mem_3__7_), .C(w_mem_inst_w_mem_14__7_), .D(w_mem_inst__abc_19396_new_n1638__bF_buf2), .Y(w_mem_inst__abc_19396_new_n1814_));
AOI22X1 AOI22X1_24 ( .A(d_reg_21_), .B(round_ctr_inc_bF_buf12), .C(_abc_15497_new_n1650__bF_buf4), .D(_abc_15497_new_n1715_), .Y(_abc_15497_new_n1716_));
AOI22X1 AOI22X1_240 ( .A(w_mem_inst__abc_19396_new_n1587__bF_buf2), .B(w_mem_inst__abc_19396_new_n1795_), .C(w_mem_inst__abc_19396_new_n1804_), .D(w_mem_inst__abc_19396_new_n1816_), .Y(w_7_));
AOI22X1 AOI22X1_241 ( .A(w_mem_inst__abc_19396_new_n1625__bF_buf1), .B(w_mem_inst_w_mem_9__8_), .C(w_mem_inst_w_mem_10__8_), .D(w_mem_inst__abc_19396_new_n1628__bF_buf1), .Y(w_mem_inst__abc_19396_new_n1834_));
AOI22X1 AOI22X1_242 ( .A(w_mem_inst__abc_19396_new_n1630__bF_buf1), .B(w_mem_inst_w_mem_4__8_), .C(w_mem_inst_w_mem_6__8_), .D(w_mem_inst__abc_19396_new_n1631__bF_buf1), .Y(w_mem_inst__abc_19396_new_n1835_));
AOI22X1 AOI22X1_243 ( .A(w_mem_inst__abc_19396_new_n1637__bF_buf1), .B(w_mem_inst_w_mem_3__8_), .C(w_mem_inst_w_mem_14__8_), .D(w_mem_inst__abc_19396_new_n1638__bF_buf1), .Y(w_mem_inst__abc_19396_new_n1839_));
AOI22X1 AOI22X1_244 ( .A(w_mem_inst__abc_19396_new_n1587__bF_buf1), .B(w_mem_inst__abc_19396_new_n1820_), .C(w_mem_inst__abc_19396_new_n1829_), .D(w_mem_inst__abc_19396_new_n1841_), .Y(w_8_));
AOI22X1 AOI22X1_245 ( .A(w_mem_inst__abc_19396_new_n1625__bF_buf0), .B(w_mem_inst_w_mem_9__9_), .C(w_mem_inst_w_mem_10__9_), .D(w_mem_inst__abc_19396_new_n1628__bF_buf0), .Y(w_mem_inst__abc_19396_new_n1859_));
AOI22X1 AOI22X1_246 ( .A(w_mem_inst__abc_19396_new_n1630__bF_buf0), .B(w_mem_inst_w_mem_4__9_), .C(w_mem_inst_w_mem_6__9_), .D(w_mem_inst__abc_19396_new_n1631__bF_buf0), .Y(w_mem_inst__abc_19396_new_n1860_));
AOI22X1 AOI22X1_247 ( .A(w_mem_inst__abc_19396_new_n1637__bF_buf0), .B(w_mem_inst_w_mem_3__9_), .C(w_mem_inst_w_mem_14__9_), .D(w_mem_inst__abc_19396_new_n1638__bF_buf0), .Y(w_mem_inst__abc_19396_new_n1864_));
AOI22X1 AOI22X1_248 ( .A(w_mem_inst__abc_19396_new_n1587__bF_buf0), .B(w_mem_inst__abc_19396_new_n1845_), .C(w_mem_inst__abc_19396_new_n1854_), .D(w_mem_inst__abc_19396_new_n1866_), .Y(w_9_));
AOI22X1 AOI22X1_249 ( .A(w_mem_inst__abc_19396_new_n1625__bF_buf4), .B(w_mem_inst_w_mem_9__10_), .C(w_mem_inst_w_mem_10__10_), .D(w_mem_inst__abc_19396_new_n1628__bF_buf4), .Y(w_mem_inst__abc_19396_new_n1884_));
AOI22X1 AOI22X1_25 ( .A(d_reg_22_), .B(round_ctr_inc_bF_buf11), .C(e_reg_22_), .D(_abc_15497_new_n1663__bF_buf1), .Y(_abc_15497_new_n1719_));
AOI22X1 AOI22X1_250 ( .A(w_mem_inst__abc_19396_new_n1630__bF_buf4), .B(w_mem_inst_w_mem_4__10_), .C(w_mem_inst_w_mem_6__10_), .D(w_mem_inst__abc_19396_new_n1631__bF_buf4), .Y(w_mem_inst__abc_19396_new_n1885_));
AOI22X1 AOI22X1_251 ( .A(w_mem_inst__abc_19396_new_n1637__bF_buf4), .B(w_mem_inst_w_mem_3__10_), .C(w_mem_inst_w_mem_14__10_), .D(w_mem_inst__abc_19396_new_n1638__bF_buf4), .Y(w_mem_inst__abc_19396_new_n1889_));
AOI22X1 AOI22X1_252 ( .A(w_mem_inst__abc_19396_new_n1587__bF_buf4), .B(w_mem_inst__abc_19396_new_n1870_), .C(w_mem_inst__abc_19396_new_n1879_), .D(w_mem_inst__abc_19396_new_n1891_), .Y(w_10_));
AOI22X1 AOI22X1_253 ( .A(w_mem_inst__abc_19396_new_n1625__bF_buf3), .B(w_mem_inst_w_mem_9__11_), .C(w_mem_inst_w_mem_10__11_), .D(w_mem_inst__abc_19396_new_n1628__bF_buf3), .Y(w_mem_inst__abc_19396_new_n1909_));
AOI22X1 AOI22X1_254 ( .A(w_mem_inst__abc_19396_new_n1630__bF_buf3), .B(w_mem_inst_w_mem_4__11_), .C(w_mem_inst_w_mem_6__11_), .D(w_mem_inst__abc_19396_new_n1631__bF_buf3), .Y(w_mem_inst__abc_19396_new_n1910_));
AOI22X1 AOI22X1_255 ( .A(w_mem_inst__abc_19396_new_n1637__bF_buf3), .B(w_mem_inst_w_mem_3__11_), .C(w_mem_inst_w_mem_14__11_), .D(w_mem_inst__abc_19396_new_n1638__bF_buf3), .Y(w_mem_inst__abc_19396_new_n1914_));
AOI22X1 AOI22X1_256 ( .A(w_mem_inst__abc_19396_new_n1587__bF_buf3), .B(w_mem_inst__abc_19396_new_n1895_), .C(w_mem_inst__abc_19396_new_n1904_), .D(w_mem_inst__abc_19396_new_n1916_), .Y(w_11_));
AOI22X1 AOI22X1_257 ( .A(w_mem_inst__abc_19396_new_n1625__bF_buf2), .B(w_mem_inst_w_mem_9__12_), .C(w_mem_inst_w_mem_10__12_), .D(w_mem_inst__abc_19396_new_n1628__bF_buf2), .Y(w_mem_inst__abc_19396_new_n1934_));
AOI22X1 AOI22X1_258 ( .A(w_mem_inst__abc_19396_new_n1630__bF_buf2), .B(w_mem_inst_w_mem_4__12_), .C(w_mem_inst_w_mem_6__12_), .D(w_mem_inst__abc_19396_new_n1631__bF_buf2), .Y(w_mem_inst__abc_19396_new_n1935_));
AOI22X1 AOI22X1_259 ( .A(w_mem_inst__abc_19396_new_n1637__bF_buf2), .B(w_mem_inst_w_mem_3__12_), .C(w_mem_inst_w_mem_14__12_), .D(w_mem_inst__abc_19396_new_n1638__bF_buf2), .Y(w_mem_inst__abc_19396_new_n1939_));
AOI22X1 AOI22X1_26 ( .A(d_reg_23_), .B(round_ctr_inc_bF_buf9), .C(e_reg_23_), .D(_abc_15497_new_n1663__bF_buf0), .Y(_abc_15497_new_n1722_));
AOI22X1 AOI22X1_260 ( .A(w_mem_inst__abc_19396_new_n1587__bF_buf2), .B(w_mem_inst__abc_19396_new_n1920_), .C(w_mem_inst__abc_19396_new_n1929_), .D(w_mem_inst__abc_19396_new_n1941_), .Y(w_12_));
AOI22X1 AOI22X1_261 ( .A(w_mem_inst__abc_19396_new_n1625__bF_buf1), .B(w_mem_inst_w_mem_9__13_), .C(w_mem_inst_w_mem_10__13_), .D(w_mem_inst__abc_19396_new_n1628__bF_buf1), .Y(w_mem_inst__abc_19396_new_n1959_));
AOI22X1 AOI22X1_262 ( .A(w_mem_inst__abc_19396_new_n1630__bF_buf1), .B(w_mem_inst_w_mem_4__13_), .C(w_mem_inst_w_mem_6__13_), .D(w_mem_inst__abc_19396_new_n1631__bF_buf1), .Y(w_mem_inst__abc_19396_new_n1960_));
AOI22X1 AOI22X1_263 ( .A(w_mem_inst__abc_19396_new_n1637__bF_buf1), .B(w_mem_inst_w_mem_3__13_), .C(w_mem_inst_w_mem_14__13_), .D(w_mem_inst__abc_19396_new_n1638__bF_buf1), .Y(w_mem_inst__abc_19396_new_n1964_));
AOI22X1 AOI22X1_264 ( .A(w_mem_inst__abc_19396_new_n1587__bF_buf1), .B(w_mem_inst__abc_19396_new_n1945_), .C(w_mem_inst__abc_19396_new_n1954_), .D(w_mem_inst__abc_19396_new_n1966_), .Y(w_13_));
AOI22X1 AOI22X1_265 ( .A(w_mem_inst__abc_19396_new_n1625__bF_buf0), .B(w_mem_inst_w_mem_9__14_), .C(w_mem_inst_w_mem_10__14_), .D(w_mem_inst__abc_19396_new_n1628__bF_buf0), .Y(w_mem_inst__abc_19396_new_n1984_));
AOI22X1 AOI22X1_266 ( .A(w_mem_inst__abc_19396_new_n1630__bF_buf0), .B(w_mem_inst_w_mem_4__14_), .C(w_mem_inst_w_mem_6__14_), .D(w_mem_inst__abc_19396_new_n1631__bF_buf0), .Y(w_mem_inst__abc_19396_new_n1985_));
AOI22X1 AOI22X1_267 ( .A(w_mem_inst__abc_19396_new_n1637__bF_buf0), .B(w_mem_inst_w_mem_3__14_), .C(w_mem_inst_w_mem_14__14_), .D(w_mem_inst__abc_19396_new_n1638__bF_buf0), .Y(w_mem_inst__abc_19396_new_n1989_));
AOI22X1 AOI22X1_268 ( .A(w_mem_inst__abc_19396_new_n1587__bF_buf0), .B(w_mem_inst__abc_19396_new_n1970_), .C(w_mem_inst__abc_19396_new_n1979_), .D(w_mem_inst__abc_19396_new_n1991_), .Y(w_14_));
AOI22X1 AOI22X1_269 ( .A(w_mem_inst__abc_19396_new_n1625__bF_buf4), .B(w_mem_inst_w_mem_9__15_), .C(w_mem_inst_w_mem_10__15_), .D(w_mem_inst__abc_19396_new_n1628__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2009_));
AOI22X1 AOI22X1_27 ( .A(d_reg_24_), .B(round_ctr_inc_bF_buf7), .C(_abc_15497_new_n1724_), .D(_abc_15497_new_n1650__bF_buf3), .Y(_abc_15497_new_n1725_));
AOI22X1 AOI22X1_270 ( .A(w_mem_inst__abc_19396_new_n1630__bF_buf4), .B(w_mem_inst_w_mem_4__15_), .C(w_mem_inst_w_mem_6__15_), .D(w_mem_inst__abc_19396_new_n1631__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2010_));
AOI22X1 AOI22X1_271 ( .A(w_mem_inst__abc_19396_new_n1637__bF_buf4), .B(w_mem_inst_w_mem_3__15_), .C(w_mem_inst_w_mem_14__15_), .D(w_mem_inst__abc_19396_new_n1638__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2014_));
AOI22X1 AOI22X1_272 ( .A(w_mem_inst__abc_19396_new_n1587__bF_buf4), .B(w_mem_inst__abc_19396_new_n1995_), .C(w_mem_inst__abc_19396_new_n2004_), .D(w_mem_inst__abc_19396_new_n2016_), .Y(w_15_));
AOI22X1 AOI22X1_273 ( .A(w_mem_inst__abc_19396_new_n1625__bF_buf3), .B(w_mem_inst_w_mem_9__16_), .C(w_mem_inst_w_mem_10__16_), .D(w_mem_inst__abc_19396_new_n1628__bF_buf3), .Y(w_mem_inst__abc_19396_new_n2034_));
AOI22X1 AOI22X1_274 ( .A(w_mem_inst__abc_19396_new_n1630__bF_buf3), .B(w_mem_inst_w_mem_4__16_), .C(w_mem_inst_w_mem_6__16_), .D(w_mem_inst__abc_19396_new_n1631__bF_buf3), .Y(w_mem_inst__abc_19396_new_n2035_));
AOI22X1 AOI22X1_275 ( .A(w_mem_inst__abc_19396_new_n1637__bF_buf3), .B(w_mem_inst_w_mem_3__16_), .C(w_mem_inst_w_mem_14__16_), .D(w_mem_inst__abc_19396_new_n1638__bF_buf3), .Y(w_mem_inst__abc_19396_new_n2039_));
AOI22X1 AOI22X1_276 ( .A(w_mem_inst__abc_19396_new_n1587__bF_buf3), .B(w_mem_inst__abc_19396_new_n2020_), .C(w_mem_inst__abc_19396_new_n2029_), .D(w_mem_inst__abc_19396_new_n2041_), .Y(w_16_));
AOI22X1 AOI22X1_277 ( .A(w_mem_inst__abc_19396_new_n1625__bF_buf2), .B(w_mem_inst_w_mem_9__17_), .C(w_mem_inst_w_mem_10__17_), .D(w_mem_inst__abc_19396_new_n1628__bF_buf2), .Y(w_mem_inst__abc_19396_new_n2059_));
AOI22X1 AOI22X1_278 ( .A(w_mem_inst__abc_19396_new_n1630__bF_buf2), .B(w_mem_inst_w_mem_4__17_), .C(w_mem_inst_w_mem_6__17_), .D(w_mem_inst__abc_19396_new_n1631__bF_buf2), .Y(w_mem_inst__abc_19396_new_n2060_));
AOI22X1 AOI22X1_279 ( .A(w_mem_inst__abc_19396_new_n1637__bF_buf2), .B(w_mem_inst_w_mem_3__17_), .C(w_mem_inst_w_mem_14__17_), .D(w_mem_inst__abc_19396_new_n1638__bF_buf2), .Y(w_mem_inst__abc_19396_new_n2064_));
AOI22X1 AOI22X1_28 ( .A(d_reg_25_), .B(round_ctr_inc_bF_buf6), .C(e_reg_25_), .D(_abc_15497_new_n1663__bF_buf7), .Y(_abc_15497_new_n1728_));
AOI22X1 AOI22X1_280 ( .A(w_mem_inst__abc_19396_new_n1587__bF_buf2), .B(w_mem_inst__abc_19396_new_n2045_), .C(w_mem_inst__abc_19396_new_n2054_), .D(w_mem_inst__abc_19396_new_n2066_), .Y(w_17_));
AOI22X1 AOI22X1_281 ( .A(w_mem_inst__abc_19396_new_n1625__bF_buf1), .B(w_mem_inst_w_mem_9__18_), .C(w_mem_inst_w_mem_10__18_), .D(w_mem_inst__abc_19396_new_n1628__bF_buf1), .Y(w_mem_inst__abc_19396_new_n2084_));
AOI22X1 AOI22X1_282 ( .A(w_mem_inst__abc_19396_new_n1630__bF_buf1), .B(w_mem_inst_w_mem_4__18_), .C(w_mem_inst_w_mem_6__18_), .D(w_mem_inst__abc_19396_new_n1631__bF_buf1), .Y(w_mem_inst__abc_19396_new_n2085_));
AOI22X1 AOI22X1_283 ( .A(w_mem_inst__abc_19396_new_n1637__bF_buf1), .B(w_mem_inst_w_mem_3__18_), .C(w_mem_inst_w_mem_14__18_), .D(w_mem_inst__abc_19396_new_n1638__bF_buf1), .Y(w_mem_inst__abc_19396_new_n2089_));
AOI22X1 AOI22X1_284 ( .A(w_mem_inst__abc_19396_new_n1587__bF_buf1), .B(w_mem_inst__abc_19396_new_n2070_), .C(w_mem_inst__abc_19396_new_n2079_), .D(w_mem_inst__abc_19396_new_n2091_), .Y(w_18_));
AOI22X1 AOI22X1_285 ( .A(w_mem_inst__abc_19396_new_n1625__bF_buf0), .B(w_mem_inst_w_mem_9__19_), .C(w_mem_inst_w_mem_10__19_), .D(w_mem_inst__abc_19396_new_n1628__bF_buf0), .Y(w_mem_inst__abc_19396_new_n2109_));
AOI22X1 AOI22X1_286 ( .A(w_mem_inst__abc_19396_new_n1630__bF_buf0), .B(w_mem_inst_w_mem_4__19_), .C(w_mem_inst_w_mem_6__19_), .D(w_mem_inst__abc_19396_new_n1631__bF_buf0), .Y(w_mem_inst__abc_19396_new_n2110_));
AOI22X1 AOI22X1_287 ( .A(w_mem_inst__abc_19396_new_n1637__bF_buf0), .B(w_mem_inst_w_mem_3__19_), .C(w_mem_inst_w_mem_14__19_), .D(w_mem_inst__abc_19396_new_n1638__bF_buf0), .Y(w_mem_inst__abc_19396_new_n2114_));
AOI22X1 AOI22X1_288 ( .A(w_mem_inst__abc_19396_new_n1587__bF_buf0), .B(w_mem_inst__abc_19396_new_n2095_), .C(w_mem_inst__abc_19396_new_n2104_), .D(w_mem_inst__abc_19396_new_n2116_), .Y(w_19_));
AOI22X1 AOI22X1_289 ( .A(w_mem_inst__abc_19396_new_n1625__bF_buf4), .B(w_mem_inst_w_mem_9__20_), .C(w_mem_inst_w_mem_10__20_), .D(w_mem_inst__abc_19396_new_n1628__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2134_));
AOI22X1 AOI22X1_29 ( .A(d_reg_26_), .B(round_ctr_inc_bF_buf4), .C(_abc_15497_new_n1650__bF_buf2), .D(_abc_15497_new_n1730_), .Y(_abc_15497_new_n1731_));
AOI22X1 AOI22X1_290 ( .A(w_mem_inst__abc_19396_new_n1630__bF_buf4), .B(w_mem_inst_w_mem_4__20_), .C(w_mem_inst_w_mem_6__20_), .D(w_mem_inst__abc_19396_new_n1631__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2135_));
AOI22X1 AOI22X1_291 ( .A(w_mem_inst__abc_19396_new_n1637__bF_buf4), .B(w_mem_inst_w_mem_3__20_), .C(w_mem_inst_w_mem_14__20_), .D(w_mem_inst__abc_19396_new_n1638__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2139_));
AOI22X1 AOI22X1_292 ( .A(w_mem_inst__abc_19396_new_n1587__bF_buf4), .B(w_mem_inst__abc_19396_new_n2120_), .C(w_mem_inst__abc_19396_new_n2129_), .D(w_mem_inst__abc_19396_new_n2141_), .Y(w_20_));
AOI22X1 AOI22X1_293 ( .A(w_mem_inst__abc_19396_new_n1625__bF_buf3), .B(w_mem_inst_w_mem_9__21_), .C(w_mem_inst_w_mem_10__21_), .D(w_mem_inst__abc_19396_new_n1628__bF_buf3), .Y(w_mem_inst__abc_19396_new_n2159_));
AOI22X1 AOI22X1_294 ( .A(w_mem_inst__abc_19396_new_n1630__bF_buf3), .B(w_mem_inst_w_mem_4__21_), .C(w_mem_inst_w_mem_6__21_), .D(w_mem_inst__abc_19396_new_n1631__bF_buf3), .Y(w_mem_inst__abc_19396_new_n2160_));
AOI22X1 AOI22X1_295 ( .A(w_mem_inst__abc_19396_new_n1637__bF_buf3), .B(w_mem_inst_w_mem_3__21_), .C(w_mem_inst_w_mem_14__21_), .D(w_mem_inst__abc_19396_new_n1638__bF_buf3), .Y(w_mem_inst__abc_19396_new_n2164_));
AOI22X1 AOI22X1_296 ( .A(w_mem_inst__abc_19396_new_n1587__bF_buf3), .B(w_mem_inst__abc_19396_new_n2145_), .C(w_mem_inst__abc_19396_new_n2154_), .D(w_mem_inst__abc_19396_new_n2166_), .Y(w_21_));
AOI22X1 AOI22X1_297 ( .A(w_mem_inst__abc_19396_new_n1625__bF_buf2), .B(w_mem_inst_w_mem_9__22_), .C(w_mem_inst_w_mem_10__22_), .D(w_mem_inst__abc_19396_new_n1628__bF_buf2), .Y(w_mem_inst__abc_19396_new_n2184_));
AOI22X1 AOI22X1_298 ( .A(w_mem_inst__abc_19396_new_n1630__bF_buf2), .B(w_mem_inst_w_mem_4__22_), .C(w_mem_inst_w_mem_6__22_), .D(w_mem_inst__abc_19396_new_n1631__bF_buf2), .Y(w_mem_inst__abc_19396_new_n2185_));
AOI22X1 AOI22X1_299 ( .A(w_mem_inst__abc_19396_new_n1637__bF_buf2), .B(w_mem_inst_w_mem_3__22_), .C(w_mem_inst_w_mem_14__22_), .D(w_mem_inst__abc_19396_new_n1638__bF_buf2), .Y(w_mem_inst__abc_19396_new_n2189_));
AOI22X1 AOI22X1_3 ( .A(d_reg_0_), .B(round_ctr_inc_bF_buf11), .C(_abc_15497_new_n1650__bF_buf9), .D(_abc_15497_new_n1649_), .Y(_abc_15497_new_n1651_));
AOI22X1 AOI22X1_30 ( .A(d_reg_27_), .B(round_ctr_inc_bF_buf3), .C(_abc_15497_new_n1650__bF_buf1), .D(_abc_15497_new_n1733_), .Y(_abc_15497_new_n1734_));
AOI22X1 AOI22X1_300 ( .A(w_mem_inst__abc_19396_new_n1587__bF_buf2), .B(w_mem_inst__abc_19396_new_n2170_), .C(w_mem_inst__abc_19396_new_n2179_), .D(w_mem_inst__abc_19396_new_n2191_), .Y(w_22_));
AOI22X1 AOI22X1_301 ( .A(w_mem_inst__abc_19396_new_n1625__bF_buf1), .B(w_mem_inst_w_mem_9__23_), .C(w_mem_inst_w_mem_10__23_), .D(w_mem_inst__abc_19396_new_n1628__bF_buf1), .Y(w_mem_inst__abc_19396_new_n2209_));
AOI22X1 AOI22X1_302 ( .A(w_mem_inst__abc_19396_new_n1630__bF_buf1), .B(w_mem_inst_w_mem_4__23_), .C(w_mem_inst_w_mem_6__23_), .D(w_mem_inst__abc_19396_new_n1631__bF_buf1), .Y(w_mem_inst__abc_19396_new_n2210_));
AOI22X1 AOI22X1_303 ( .A(w_mem_inst__abc_19396_new_n1637__bF_buf1), .B(w_mem_inst_w_mem_3__23_), .C(w_mem_inst_w_mem_14__23_), .D(w_mem_inst__abc_19396_new_n1638__bF_buf1), .Y(w_mem_inst__abc_19396_new_n2214_));
AOI22X1 AOI22X1_304 ( .A(w_mem_inst__abc_19396_new_n1587__bF_buf1), .B(w_mem_inst__abc_19396_new_n2195_), .C(w_mem_inst__abc_19396_new_n2204_), .D(w_mem_inst__abc_19396_new_n2216_), .Y(w_23_));
AOI22X1 AOI22X1_305 ( .A(w_mem_inst__abc_19396_new_n1625__bF_buf0), .B(w_mem_inst_w_mem_9__24_), .C(w_mem_inst_w_mem_10__24_), .D(w_mem_inst__abc_19396_new_n1628__bF_buf0), .Y(w_mem_inst__abc_19396_new_n2234_));
AOI22X1 AOI22X1_306 ( .A(w_mem_inst__abc_19396_new_n1630__bF_buf0), .B(w_mem_inst_w_mem_4__24_), .C(w_mem_inst_w_mem_6__24_), .D(w_mem_inst__abc_19396_new_n1631__bF_buf0), .Y(w_mem_inst__abc_19396_new_n2235_));
AOI22X1 AOI22X1_307 ( .A(w_mem_inst__abc_19396_new_n1637__bF_buf0), .B(w_mem_inst_w_mem_3__24_), .C(w_mem_inst_w_mem_14__24_), .D(w_mem_inst__abc_19396_new_n1638__bF_buf0), .Y(w_mem_inst__abc_19396_new_n2239_));
AOI22X1 AOI22X1_308 ( .A(w_mem_inst__abc_19396_new_n1587__bF_buf0), .B(w_mem_inst__abc_19396_new_n2220_), .C(w_mem_inst__abc_19396_new_n2229_), .D(w_mem_inst__abc_19396_new_n2241_), .Y(w_24_));
AOI22X1 AOI22X1_309 ( .A(w_mem_inst__abc_19396_new_n1625__bF_buf4), .B(w_mem_inst_w_mem_9__25_), .C(w_mem_inst_w_mem_10__25_), .D(w_mem_inst__abc_19396_new_n1628__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2259_));
AOI22X1 AOI22X1_31 ( .A(d_reg_28_), .B(round_ctr_inc_bF_buf2), .C(_abc_15497_new_n1650__bF_buf0), .D(_abc_15497_new_n1737_), .Y(_abc_15497_new_n1738_));
AOI22X1 AOI22X1_310 ( .A(w_mem_inst__abc_19396_new_n1630__bF_buf4), .B(w_mem_inst_w_mem_4__25_), .C(w_mem_inst_w_mem_6__25_), .D(w_mem_inst__abc_19396_new_n1631__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2260_));
AOI22X1 AOI22X1_311 ( .A(w_mem_inst__abc_19396_new_n1637__bF_buf4), .B(w_mem_inst_w_mem_3__25_), .C(w_mem_inst_w_mem_14__25_), .D(w_mem_inst__abc_19396_new_n1638__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2264_));
AOI22X1 AOI22X1_312 ( .A(w_mem_inst__abc_19396_new_n1587__bF_buf4), .B(w_mem_inst__abc_19396_new_n2245_), .C(w_mem_inst__abc_19396_new_n2254_), .D(w_mem_inst__abc_19396_new_n2266_), .Y(w_25_));
AOI22X1 AOI22X1_313 ( .A(w_mem_inst__abc_19396_new_n1625__bF_buf3), .B(w_mem_inst_w_mem_9__26_), .C(w_mem_inst_w_mem_10__26_), .D(w_mem_inst__abc_19396_new_n1628__bF_buf3), .Y(w_mem_inst__abc_19396_new_n2284_));
AOI22X1 AOI22X1_314 ( .A(w_mem_inst__abc_19396_new_n1630__bF_buf3), .B(w_mem_inst_w_mem_4__26_), .C(w_mem_inst_w_mem_6__26_), .D(w_mem_inst__abc_19396_new_n1631__bF_buf3), .Y(w_mem_inst__abc_19396_new_n2285_));
AOI22X1 AOI22X1_315 ( .A(w_mem_inst__abc_19396_new_n1637__bF_buf3), .B(w_mem_inst_w_mem_3__26_), .C(w_mem_inst_w_mem_14__26_), .D(w_mem_inst__abc_19396_new_n1638__bF_buf3), .Y(w_mem_inst__abc_19396_new_n2289_));
AOI22X1 AOI22X1_316 ( .A(w_mem_inst__abc_19396_new_n1587__bF_buf3), .B(w_mem_inst__abc_19396_new_n2270_), .C(w_mem_inst__abc_19396_new_n2279_), .D(w_mem_inst__abc_19396_new_n2291_), .Y(w_26_));
AOI22X1 AOI22X1_317 ( .A(w_mem_inst__abc_19396_new_n1625__bF_buf2), .B(w_mem_inst_w_mem_9__27_), .C(w_mem_inst_w_mem_10__27_), .D(w_mem_inst__abc_19396_new_n1628__bF_buf2), .Y(w_mem_inst__abc_19396_new_n2309_));
AOI22X1 AOI22X1_318 ( .A(w_mem_inst__abc_19396_new_n1630__bF_buf2), .B(w_mem_inst_w_mem_4__27_), .C(w_mem_inst_w_mem_6__27_), .D(w_mem_inst__abc_19396_new_n1631__bF_buf2), .Y(w_mem_inst__abc_19396_new_n2310_));
AOI22X1 AOI22X1_319 ( .A(w_mem_inst__abc_19396_new_n1637__bF_buf2), .B(w_mem_inst_w_mem_3__27_), .C(w_mem_inst_w_mem_14__27_), .D(w_mem_inst__abc_19396_new_n1638__bF_buf2), .Y(w_mem_inst__abc_19396_new_n2314_));
AOI22X1 AOI22X1_32 ( .A(d_reg_29_), .B(round_ctr_inc_bF_buf1), .C(_abc_15497_new_n1650__bF_buf9), .D(_abc_15497_new_n1740_), .Y(_abc_15497_new_n1741_));
AOI22X1 AOI22X1_320 ( .A(w_mem_inst__abc_19396_new_n1587__bF_buf2), .B(w_mem_inst__abc_19396_new_n2295_), .C(w_mem_inst__abc_19396_new_n2304_), .D(w_mem_inst__abc_19396_new_n2316_), .Y(w_27_));
AOI22X1 AOI22X1_321 ( .A(w_mem_inst__abc_19396_new_n1625__bF_buf1), .B(w_mem_inst_w_mem_9__28_), .C(w_mem_inst_w_mem_10__28_), .D(w_mem_inst__abc_19396_new_n1628__bF_buf1), .Y(w_mem_inst__abc_19396_new_n2334_));
AOI22X1 AOI22X1_322 ( .A(w_mem_inst__abc_19396_new_n1630__bF_buf1), .B(w_mem_inst_w_mem_4__28_), .C(w_mem_inst_w_mem_6__28_), .D(w_mem_inst__abc_19396_new_n1631__bF_buf1), .Y(w_mem_inst__abc_19396_new_n2335_));
AOI22X1 AOI22X1_323 ( .A(w_mem_inst__abc_19396_new_n1637__bF_buf1), .B(w_mem_inst_w_mem_3__28_), .C(w_mem_inst_w_mem_14__28_), .D(w_mem_inst__abc_19396_new_n1638__bF_buf1), .Y(w_mem_inst__abc_19396_new_n2339_));
AOI22X1 AOI22X1_324 ( .A(w_mem_inst__abc_19396_new_n1587__bF_buf1), .B(w_mem_inst__abc_19396_new_n2320_), .C(w_mem_inst__abc_19396_new_n2329_), .D(w_mem_inst__abc_19396_new_n2341_), .Y(w_28_));
AOI22X1 AOI22X1_325 ( .A(w_mem_inst__abc_19396_new_n1625__bF_buf0), .B(w_mem_inst_w_mem_9__29_), .C(w_mem_inst_w_mem_10__29_), .D(w_mem_inst__abc_19396_new_n1628__bF_buf0), .Y(w_mem_inst__abc_19396_new_n2359_));
AOI22X1 AOI22X1_326 ( .A(w_mem_inst__abc_19396_new_n1630__bF_buf0), .B(w_mem_inst_w_mem_4__29_), .C(w_mem_inst_w_mem_6__29_), .D(w_mem_inst__abc_19396_new_n1631__bF_buf0), .Y(w_mem_inst__abc_19396_new_n2360_));
AOI22X1 AOI22X1_327 ( .A(w_mem_inst__abc_19396_new_n1637__bF_buf0), .B(w_mem_inst_w_mem_3__29_), .C(w_mem_inst_w_mem_14__29_), .D(w_mem_inst__abc_19396_new_n1638__bF_buf0), .Y(w_mem_inst__abc_19396_new_n2364_));
AOI22X1 AOI22X1_328 ( .A(w_mem_inst__abc_19396_new_n1587__bF_buf0), .B(w_mem_inst__abc_19396_new_n2345_), .C(w_mem_inst__abc_19396_new_n2354_), .D(w_mem_inst__abc_19396_new_n2366_), .Y(w_29_));
AOI22X1 AOI22X1_329 ( .A(w_mem_inst__abc_19396_new_n1625__bF_buf4), .B(w_mem_inst_w_mem_9__30_), .C(w_mem_inst_w_mem_10__30_), .D(w_mem_inst__abc_19396_new_n1628__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2384_));
AOI22X1 AOI22X1_33 ( .A(d_reg_30_), .B(round_ctr_inc_bF_buf0), .C(e_reg_30_), .D(_abc_15497_new_n1663__bF_buf6), .Y(_abc_15497_new_n1744_));
AOI22X1 AOI22X1_330 ( .A(w_mem_inst__abc_19396_new_n1630__bF_buf4), .B(w_mem_inst_w_mem_4__30_), .C(w_mem_inst_w_mem_6__30_), .D(w_mem_inst__abc_19396_new_n1631__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2385_));
AOI22X1 AOI22X1_331 ( .A(w_mem_inst__abc_19396_new_n1637__bF_buf4), .B(w_mem_inst_w_mem_3__30_), .C(w_mem_inst_w_mem_14__30_), .D(w_mem_inst__abc_19396_new_n1638__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2389_));
AOI22X1 AOI22X1_332 ( .A(w_mem_inst__abc_19396_new_n1587__bF_buf4), .B(w_mem_inst__abc_19396_new_n2370_), .C(w_mem_inst__abc_19396_new_n2379_), .D(w_mem_inst__abc_19396_new_n2391_), .Y(w_30_));
AOI22X1 AOI22X1_333 ( .A(w_mem_inst__abc_19396_new_n1625__bF_buf3), .B(w_mem_inst_w_mem_9__31_), .C(w_mem_inst_w_mem_10__31_), .D(w_mem_inst__abc_19396_new_n1628__bF_buf3), .Y(w_mem_inst__abc_19396_new_n2409_));
AOI22X1 AOI22X1_334 ( .A(w_mem_inst__abc_19396_new_n1630__bF_buf3), .B(w_mem_inst_w_mem_4__31_), .C(w_mem_inst_w_mem_6__31_), .D(w_mem_inst__abc_19396_new_n1631__bF_buf3), .Y(w_mem_inst__abc_19396_new_n2410_));
AOI22X1 AOI22X1_335 ( .A(w_mem_inst__abc_19396_new_n1637__bF_buf3), .B(w_mem_inst_w_mem_3__31_), .C(w_mem_inst_w_mem_14__31_), .D(w_mem_inst__abc_19396_new_n1638__bF_buf3), .Y(w_mem_inst__abc_19396_new_n2414_));
AOI22X1 AOI22X1_336 ( .A(w_mem_inst__abc_19396_new_n1587__bF_buf3), .B(w_mem_inst__abc_19396_new_n2395_), .C(w_mem_inst__abc_19396_new_n2404_), .D(w_mem_inst__abc_19396_new_n2416_), .Y(w_31_));
AOI22X1 AOI22X1_34 ( .A(_abc_15497_new_n870__bF_buf3), .B(_abc_15497_new_n2062_), .C(_abc_15497_new_n2070_), .D(_abc_15497_new_n2069_), .Y(_0H1_reg_31_0__29_));
AOI22X1 AOI22X1_35 ( .A(round_ctr_inc_bF_buf11), .B(a_reg_0_), .C(_abc_15497_new_n2444_), .D(_abc_15497_new_n1650__bF_buf7), .Y(_abc_15497_new_n2445_));
AOI22X1 AOI22X1_36 ( .A(round_ctr_inc_bF_buf10), .B(a_reg_1_), .C(_abc_15497_new_n1650__bF_buf6), .D(_abc_15497_new_n2447_), .Y(_abc_15497_new_n2448_));
AOI22X1 AOI22X1_37 ( .A(round_ctr_inc_bF_buf9), .B(a_reg_2_), .C(_abc_15497_new_n1650__bF_buf5), .D(_abc_15497_new_n2450_), .Y(_abc_15497_new_n2451_));
AOI22X1 AOI22X1_38 ( .A(round_ctr_inc_bF_buf8), .B(a_reg_3_), .C(b_reg_3_), .D(_abc_15497_new_n1663__bF_buf4), .Y(_abc_15497_new_n2454_));
AOI22X1 AOI22X1_39 ( .A(round_ctr_inc_bF_buf6), .B(a_reg_4_), .C(_abc_15497_new_n1650__bF_buf4), .D(_abc_15497_new_n2456_), .Y(_abc_15497_new_n2457_));
AOI22X1 AOI22X1_4 ( .A(d_reg_1_), .B(round_ctr_inc_bF_buf10), .C(_abc_15497_new_n1650__bF_buf8), .D(_abc_15497_new_n1653_), .Y(_abc_15497_new_n1654_));
AOI22X1 AOI22X1_40 ( .A(round_ctr_inc_bF_buf5), .B(a_reg_5_), .C(_abc_15497_new_n1650__bF_buf3), .D(_abc_15497_new_n2459_), .Y(_abc_15497_new_n2460_));
AOI22X1 AOI22X1_41 ( .A(round_ctr_inc_bF_buf4), .B(a_reg_6_), .C(_abc_15497_new_n1650__bF_buf2), .D(_abc_15497_new_n2462_), .Y(_abc_15497_new_n2463_));
AOI22X1 AOI22X1_42 ( .A(round_ctr_inc_bF_buf3), .B(a_reg_7_), .C(b_reg_7_), .D(_abc_15497_new_n1663__bF_buf3), .Y(_abc_15497_new_n2466_));
AOI22X1 AOI22X1_43 ( .A(round_ctr_inc_bF_buf1), .B(a_reg_8_), .C(_abc_15497_new_n2468_), .D(_abc_15497_new_n1650__bF_buf1), .Y(_abc_15497_new_n2469_));
AOI22X1 AOI22X1_44 ( .A(round_ctr_inc_bF_buf0), .B(a_reg_9_), .C(b_reg_9_), .D(_abc_15497_new_n1663__bF_buf2), .Y(_abc_15497_new_n2472_));
AOI22X1 AOI22X1_45 ( .A(round_ctr_inc_bF_buf12), .B(a_reg_10_), .C(_abc_15497_new_n1650__bF_buf0), .D(_abc_15497_new_n2474_), .Y(_abc_15497_new_n2475_));
AOI22X1 AOI22X1_46 ( .A(round_ctr_inc_bF_buf11), .B(a_reg_11_), .C(b_reg_11_), .D(_abc_15497_new_n1663__bF_buf1), .Y(_abc_15497_new_n2478_));
AOI22X1 AOI22X1_47 ( .A(round_ctr_inc_bF_buf9), .B(a_reg_12_), .C(_abc_15497_new_n1650__bF_buf9), .D(_abc_15497_new_n2480_), .Y(_abc_15497_new_n2481_));
AOI22X1 AOI22X1_48 ( .A(round_ctr_inc_bF_buf8), .B(a_reg_13_), .C(_abc_15497_new_n2483_), .D(_abc_15497_new_n1650__bF_buf8), .Y(_abc_15497_new_n2484_));
AOI22X1 AOI22X1_49 ( .A(round_ctr_inc_bF_buf7), .B(a_reg_14_), .C(_abc_15497_new_n1650__bF_buf7), .D(_abc_15497_new_n2486_), .Y(_abc_15497_new_n2487_));
AOI22X1 AOI22X1_5 ( .A(d_reg_2_), .B(round_ctr_inc_bF_buf9), .C(_abc_15497_new_n1650__bF_buf7), .D(_abc_15497_new_n1656_), .Y(_abc_15497_new_n1657_));
AOI22X1 AOI22X1_50 ( .A(round_ctr_inc_bF_buf6), .B(a_reg_15_), .C(b_reg_15_), .D(_abc_15497_new_n1663__bF_buf0), .Y(_abc_15497_new_n2490_));
AOI22X1 AOI22X1_51 ( .A(round_ctr_inc_bF_buf4), .B(a_reg_16_), .C(_abc_15497_new_n2492_), .D(_abc_15497_new_n1650__bF_buf6), .Y(_abc_15497_new_n2493_));
AOI22X1 AOI22X1_52 ( .A(round_ctr_inc_bF_buf3), .B(a_reg_17_), .C(_abc_15497_new_n1650__bF_buf5), .D(_abc_15497_new_n2495_), .Y(_abc_15497_new_n2496_));
AOI22X1 AOI22X1_53 ( .A(round_ctr_inc_bF_buf2), .B(a_reg_18_), .C(b_reg_18_), .D(_abc_15497_new_n1663__bF_buf7), .Y(_abc_15497_new_n2499_));
AOI22X1 AOI22X1_54 ( .A(round_ctr_inc_bF_buf0), .B(a_reg_19_), .C(b_reg_19_), .D(_abc_15497_new_n1663__bF_buf6), .Y(_abc_15497_new_n2502_));
AOI22X1 AOI22X1_55 ( .A(round_ctr_inc_bF_buf12), .B(a_reg_20_), .C(_abc_15497_new_n1650__bF_buf4), .D(_abc_15497_new_n2504_), .Y(_abc_15497_new_n2505_));
AOI22X1 AOI22X1_56 ( .A(round_ctr_inc_bF_buf11), .B(a_reg_21_), .C(_abc_15497_new_n1650__bF_buf3), .D(_abc_15497_new_n2507_), .Y(_abc_15497_new_n2508_));
AOI22X1 AOI22X1_57 ( .A(round_ctr_inc_bF_buf10), .B(a_reg_22_), .C(b_reg_22_), .D(_abc_15497_new_n1663__bF_buf5), .Y(_abc_15497_new_n2511_));
AOI22X1 AOI22X1_58 ( .A(round_ctr_inc_bF_buf8), .B(a_reg_23_), .C(b_reg_23_), .D(_abc_15497_new_n1663__bF_buf4), .Y(_abc_15497_new_n2514_));
AOI22X1 AOI22X1_59 ( .A(round_ctr_inc_bF_buf6), .B(a_reg_24_), .C(_abc_15497_new_n2516_), .D(_abc_15497_new_n1650__bF_buf2), .Y(_abc_15497_new_n2517_));
AOI22X1 AOI22X1_6 ( .A(d_reg_3_), .B(round_ctr_inc_bF_buf8), .C(_abc_15497_new_n1650__bF_buf6), .D(_abc_15497_new_n1659_), .Y(_abc_15497_new_n1660_));
AOI22X1 AOI22X1_60 ( .A(round_ctr_inc_bF_buf5), .B(a_reg_25_), .C(b_reg_25_), .D(_abc_15497_new_n1663__bF_buf3), .Y(_abc_15497_new_n2520_));
AOI22X1 AOI22X1_61 ( .A(round_ctr_inc_bF_buf3), .B(a_reg_26_), .C(_abc_15497_new_n2522_), .D(_abc_15497_new_n1650__bF_buf1), .Y(_abc_15497_new_n2523_));
AOI22X1 AOI22X1_62 ( .A(round_ctr_inc_bF_buf2), .B(a_reg_27_), .C(b_reg_27_), .D(_abc_15497_new_n1663__bF_buf2), .Y(_abc_15497_new_n2526_));
AOI22X1 AOI22X1_63 ( .A(round_ctr_inc_bF_buf0), .B(a_reg_28_), .C(_abc_15497_new_n1650__bF_buf0), .D(_abc_15497_new_n2528_), .Y(_abc_15497_new_n2529_));
AOI22X1 AOI22X1_64 ( .A(round_ctr_inc_bF_buf13), .B(a_reg_29_), .C(b_reg_29_), .D(_abc_15497_new_n1663__bF_buf1), .Y(_abc_15497_new_n2532_));
AOI22X1 AOI22X1_65 ( .A(round_ctr_inc_bF_buf11), .B(a_reg_30_), .C(b_reg_30_), .D(_abc_15497_new_n1663__bF_buf0), .Y(_abc_15497_new_n2535_));
AOI22X1 AOI22X1_66 ( .A(round_ctr_inc_bF_buf9), .B(a_reg_31_), .C(b_reg_31_), .D(_abc_15497_new_n1663__bF_buf7), .Y(_abc_15497_new_n2538_));
AOI22X1 AOI22X1_67 ( .A(round_ctr_inc_bF_buf7), .B(c_reg_0_), .C(_abc_15497_new_n1650__bF_buf9), .D(_abc_15497_new_n2540_), .Y(_abc_15497_new_n2541_));
AOI22X1 AOI22X1_68 ( .A(round_ctr_inc_bF_buf6), .B(c_reg_1_), .C(_abc_15497_new_n2543_), .D(_abc_15497_new_n1650__bF_buf8), .Y(_abc_15497_new_n2544_));
AOI22X1 AOI22X1_69 ( .A(round_ctr_inc_bF_buf5), .B(c_reg_2_), .C(d_reg_2_), .D(_abc_15497_new_n1663__bF_buf6), .Y(_abc_15497_new_n2547_));
AOI22X1 AOI22X1_7 ( .A(d_reg_4_), .B(round_ctr_inc_bF_buf7), .C(e_reg_4_), .D(_abc_15497_new_n1663__bF_buf7), .Y(_abc_15497_new_n1664_));
AOI22X1 AOI22X1_70 ( .A(round_ctr_inc_bF_buf3), .B(c_reg_3_), .C(_abc_15497_new_n1650__bF_buf7), .D(_abc_15497_new_n2549_), .Y(_abc_15497_new_n2550_));
AOI22X1 AOI22X1_71 ( .A(round_ctr_inc_bF_buf2), .B(c_reg_4_), .C(_abc_15497_new_n2552_), .D(_abc_15497_new_n1650__bF_buf6), .Y(_abc_15497_new_n2553_));
AOI22X1 AOI22X1_72 ( .A(round_ctr_inc_bF_buf1), .B(c_reg_5_), .C(_abc_15497_new_n2555_), .D(_abc_15497_new_n1650__bF_buf5), .Y(_abc_15497_new_n2556_));
AOI22X1 AOI22X1_73 ( .A(round_ctr_inc_bF_buf0), .B(c_reg_6_), .C(_abc_15497_new_n2558_), .D(_abc_15497_new_n1650__bF_buf4), .Y(_abc_15497_new_n2559_));
AOI22X1 AOI22X1_74 ( .A(round_ctr_inc_bF_buf13), .B(c_reg_7_), .C(_abc_15497_new_n1650__bF_buf3), .D(_abc_15497_new_n2561_), .Y(_abc_15497_new_n2562_));
AOI22X1 AOI22X1_75 ( .A(round_ctr_inc_bF_buf12), .B(c_reg_8_), .C(_abc_15497_new_n1650__bF_buf2), .D(_abc_15497_new_n2564_), .Y(_abc_15497_new_n2565_));
AOI22X1 AOI22X1_76 ( .A(round_ctr_inc_bF_buf11), .B(c_reg_9_), .C(_abc_15497_new_n1650__bF_buf1), .D(_abc_15497_new_n2567_), .Y(_abc_15497_new_n2568_));
AOI22X1 AOI22X1_77 ( .A(round_ctr_inc_bF_buf10), .B(c_reg_10_), .C(d_reg_10_), .D(_abc_15497_new_n1663__bF_buf5), .Y(_abc_15497_new_n2571_));
AOI22X1 AOI22X1_78 ( .A(round_ctr_inc_bF_buf8), .B(c_reg_11_), .C(_abc_15497_new_n1650__bF_buf0), .D(_abc_15497_new_n2573_), .Y(_abc_15497_new_n2574_));
AOI22X1 AOI22X1_79 ( .A(round_ctr_inc_bF_buf7), .B(c_reg_12_), .C(_abc_15497_new_n2576_), .D(_abc_15497_new_n1650__bF_buf9), .Y(_abc_15497_new_n2577_));
AOI22X1 AOI22X1_8 ( .A(d_reg_5_), .B(round_ctr_inc_bF_buf5), .C(e_reg_5_), .D(_abc_15497_new_n1663__bF_buf6), .Y(_abc_15497_new_n1667_));
AOI22X1 AOI22X1_80 ( .A(round_ctr_inc_bF_buf6), .B(c_reg_13_), .C(_abc_15497_new_n1650__bF_buf8), .D(_abc_15497_new_n2579_), .Y(_abc_15497_new_n2580_));
AOI22X1 AOI22X1_81 ( .A(round_ctr_inc_bF_buf5), .B(c_reg_14_), .C(d_reg_14_), .D(_abc_15497_new_n1663__bF_buf4), .Y(_abc_15497_new_n2583_));
AOI22X1 AOI22X1_82 ( .A(round_ctr_inc_bF_buf3), .B(c_reg_15_), .C(_abc_15497_new_n1650__bF_buf7), .D(_abc_15497_new_n2585_), .Y(_abc_15497_new_n2586_));
AOI22X1 AOI22X1_83 ( .A(round_ctr_inc_bF_buf2), .B(c_reg_16_), .C(_abc_15497_new_n1650__bF_buf6), .D(_abc_15497_new_n2588_), .Y(_abc_15497_new_n2589_));
AOI22X1 AOI22X1_84 ( .A(round_ctr_inc_bF_buf1), .B(c_reg_17_), .C(d_reg_17_), .D(_abc_15497_new_n1663__bF_buf3), .Y(_abc_15497_new_n2592_));
AOI22X1 AOI22X1_85 ( .A(round_ctr_inc_bF_buf13), .B(c_reg_18_), .C(_abc_15497_new_n1650__bF_buf5), .D(_abc_15497_new_n2594_), .Y(_abc_15497_new_n2595_));
AOI22X1 AOI22X1_86 ( .A(round_ctr_inc_bF_buf12), .B(c_reg_19_), .C(_abc_15497_new_n1650__bF_buf4), .D(_abc_15497_new_n2597_), .Y(_abc_15497_new_n2598_));
AOI22X1 AOI22X1_87 ( .A(round_ctr_inc_bF_buf11), .B(c_reg_20_), .C(_abc_15497_new_n2600_), .D(_abc_15497_new_n1650__bF_buf3), .Y(_abc_15497_new_n2601_));
AOI22X1 AOI22X1_88 ( .A(round_ctr_inc_bF_buf10), .B(c_reg_21_), .C(d_reg_21_), .D(_abc_15497_new_n1663__bF_buf2), .Y(_abc_15497_new_n2604_));
AOI22X1 AOI22X1_89 ( .A(round_ctr_inc_bF_buf8), .B(c_reg_22_), .C(_abc_15497_new_n1650__bF_buf2), .D(_abc_15497_new_n2606_), .Y(_abc_15497_new_n2607_));
AOI22X1 AOI22X1_9 ( .A(d_reg_6_), .B(round_ctr_inc_bF_buf3), .C(e_reg_6_), .D(_abc_15497_new_n1663__bF_buf5), .Y(_abc_15497_new_n1670_));
AOI22X1 AOI22X1_90 ( .A(round_ctr_inc_bF_buf7), .B(c_reg_23_), .C(_abc_15497_new_n1650__bF_buf1), .D(_abc_15497_new_n2609_), .Y(_abc_15497_new_n2610_));
AOI22X1 AOI22X1_91 ( .A(round_ctr_inc_bF_buf6), .B(c_reg_24_), .C(_abc_15497_new_n1650__bF_buf0), .D(_abc_15497_new_n2612_), .Y(_abc_15497_new_n2613_));
AOI22X1 AOI22X1_92 ( .A(round_ctr_inc_bF_buf5), .B(c_reg_25_), .C(_abc_15497_new_n1650__bF_buf9), .D(_abc_15497_new_n2615_), .Y(_abc_15497_new_n2616_));
AOI22X1 AOI22X1_93 ( .A(c_reg_26_), .B(round_ctr_inc_bF_buf4), .C(_abc_15497_new_n1650__bF_buf8), .D(_abc_15497_new_n2618_), .Y(_abc_15497_new_n2619_));
AOI22X1 AOI22X1_94 ( .A(c_reg_27_), .B(round_ctr_inc_bF_buf3), .C(_abc_15497_new_n1650__bF_buf7), .D(_abc_15497_new_n2621_), .Y(_abc_15497_new_n2622_));
AOI22X1 AOI22X1_95 ( .A(c_reg_28_), .B(round_ctr_inc_bF_buf2), .C(d_reg_28_), .D(_abc_15497_new_n1663__bF_buf1), .Y(_abc_15497_new_n2625_));
AOI22X1 AOI22X1_96 ( .A(c_reg_29_), .B(round_ctr_inc_bF_buf0), .C(_abc_15497_new_n1650__bF_buf6), .D(_abc_15497_new_n2627_), .Y(_abc_15497_new_n2628_));
AOI22X1 AOI22X1_97 ( .A(c_reg_30_), .B(round_ctr_inc_bF_buf13), .C(_abc_15497_new_n1650__bF_buf5), .D(_abc_15497_new_n2631_), .Y(_abc_15497_new_n2632_));
AOI22X1 AOI22X1_98 ( .A(round_ctr_inc_bF_buf11), .B(b_reg_2_), .C(_abc_15497_new_n1650__bF_buf3), .D(_abc_15497_new_n2639_), .Y(_abc_15497_new_n2640_));
AOI22X1 AOI22X1_99 ( .A(round_ctr_inc_bF_buf10), .B(b_reg_3_), .C(c_reg_1_), .D(_abc_15497_new_n1663__bF_buf7), .Y(_abc_15497_new_n2643_));
BUFX2 BUFX2_1 ( .A(_auto_iopadmap_cc_368_execute_22625_0_), .Y(\digest[0] ));
BUFX2 BUFX2_10 ( .A(_auto_iopadmap_cc_368_execute_22625_9_), .Y(\digest[9] ));
BUFX2 BUFX2_100 ( .A(_auto_iopadmap_cc_368_execute_22625_99_), .Y(\digest[99] ));
BUFX2 BUFX2_101 ( .A(_auto_iopadmap_cc_368_execute_22625_100_), .Y(\digest[100] ));
BUFX2 BUFX2_102 ( .A(_auto_iopadmap_cc_368_execute_22625_101_), .Y(\digest[101] ));
BUFX2 BUFX2_103 ( .A(_auto_iopadmap_cc_368_execute_22625_102_), .Y(\digest[102] ));
BUFX2 BUFX2_104 ( .A(_auto_iopadmap_cc_368_execute_22625_103_), .Y(\digest[103] ));
BUFX2 BUFX2_105 ( .A(_auto_iopadmap_cc_368_execute_22625_104_), .Y(\digest[104] ));
BUFX2 BUFX2_106 ( .A(_auto_iopadmap_cc_368_execute_22625_105_), .Y(\digest[105] ));
BUFX2 BUFX2_107 ( .A(_auto_iopadmap_cc_368_execute_22625_106_), .Y(\digest[106] ));
BUFX2 BUFX2_108 ( .A(_auto_iopadmap_cc_368_execute_22625_107_), .Y(\digest[107] ));
BUFX2 BUFX2_109 ( .A(_auto_iopadmap_cc_368_execute_22625_108_), .Y(\digest[108] ));
BUFX2 BUFX2_11 ( .A(_auto_iopadmap_cc_368_execute_22625_10_), .Y(\digest[10] ));
BUFX2 BUFX2_110 ( .A(_auto_iopadmap_cc_368_execute_22625_109_), .Y(\digest[109] ));
BUFX2 BUFX2_111 ( .A(_auto_iopadmap_cc_368_execute_22625_110_), .Y(\digest[110] ));
BUFX2 BUFX2_112 ( .A(_auto_iopadmap_cc_368_execute_22625_111_), .Y(\digest[111] ));
BUFX2 BUFX2_113 ( .A(_auto_iopadmap_cc_368_execute_22625_112_), .Y(\digest[112] ));
BUFX2 BUFX2_114 ( .A(_auto_iopadmap_cc_368_execute_22625_113_), .Y(\digest[113] ));
BUFX2 BUFX2_115 ( .A(_auto_iopadmap_cc_368_execute_22625_114_), .Y(\digest[114] ));
BUFX2 BUFX2_116 ( .A(_auto_iopadmap_cc_368_execute_22625_115_), .Y(\digest[115] ));
BUFX2 BUFX2_117 ( .A(_auto_iopadmap_cc_368_execute_22625_116_), .Y(\digest[116] ));
BUFX2 BUFX2_118 ( .A(_auto_iopadmap_cc_368_execute_22625_117_), .Y(\digest[117] ));
BUFX2 BUFX2_119 ( .A(_auto_iopadmap_cc_368_execute_22625_118_), .Y(\digest[118] ));
BUFX2 BUFX2_12 ( .A(_auto_iopadmap_cc_368_execute_22625_11_), .Y(\digest[11] ));
BUFX2 BUFX2_120 ( .A(_auto_iopadmap_cc_368_execute_22625_119_), .Y(\digest[119] ));
BUFX2 BUFX2_121 ( .A(_auto_iopadmap_cc_368_execute_22625_120_), .Y(\digest[120] ));
BUFX2 BUFX2_122 ( .A(_auto_iopadmap_cc_368_execute_22625_121_), .Y(\digest[121] ));
BUFX2 BUFX2_123 ( .A(_auto_iopadmap_cc_368_execute_22625_122_), .Y(\digest[122] ));
BUFX2 BUFX2_124 ( .A(_auto_iopadmap_cc_368_execute_22625_123_), .Y(\digest[123] ));
BUFX2 BUFX2_125 ( .A(_auto_iopadmap_cc_368_execute_22625_124_), .Y(\digest[124] ));
BUFX2 BUFX2_126 ( .A(_auto_iopadmap_cc_368_execute_22625_125_), .Y(\digest[125] ));
BUFX2 BUFX2_127 ( .A(_auto_iopadmap_cc_368_execute_22625_126_), .Y(\digest[126] ));
BUFX2 BUFX2_128 ( .A(_auto_iopadmap_cc_368_execute_22625_127_), .Y(\digest[127] ));
BUFX2 BUFX2_129 ( .A(_auto_iopadmap_cc_368_execute_22625_128_), .Y(\digest[128] ));
BUFX2 BUFX2_13 ( .A(_auto_iopadmap_cc_368_execute_22625_12_), .Y(\digest[12] ));
BUFX2 BUFX2_130 ( .A(_auto_iopadmap_cc_368_execute_22625_129_), .Y(\digest[129] ));
BUFX2 BUFX2_131 ( .A(_auto_iopadmap_cc_368_execute_22625_130_), .Y(\digest[130] ));
BUFX2 BUFX2_132 ( .A(_auto_iopadmap_cc_368_execute_22625_131_), .Y(\digest[131] ));
BUFX2 BUFX2_133 ( .A(_auto_iopadmap_cc_368_execute_22625_132_), .Y(\digest[132] ));
BUFX2 BUFX2_134 ( .A(_auto_iopadmap_cc_368_execute_22625_133_), .Y(\digest[133] ));
BUFX2 BUFX2_135 ( .A(_auto_iopadmap_cc_368_execute_22625_134_), .Y(\digest[134] ));
BUFX2 BUFX2_136 ( .A(_auto_iopadmap_cc_368_execute_22625_135_), .Y(\digest[135] ));
BUFX2 BUFX2_137 ( .A(_auto_iopadmap_cc_368_execute_22625_136_), .Y(\digest[136] ));
BUFX2 BUFX2_138 ( .A(_auto_iopadmap_cc_368_execute_22625_137_), .Y(\digest[137] ));
BUFX2 BUFX2_139 ( .A(_auto_iopadmap_cc_368_execute_22625_138_), .Y(\digest[138] ));
BUFX2 BUFX2_14 ( .A(_auto_iopadmap_cc_368_execute_22625_13_), .Y(\digest[13] ));
BUFX2 BUFX2_140 ( .A(_auto_iopadmap_cc_368_execute_22625_139_), .Y(\digest[139] ));
BUFX2 BUFX2_141 ( .A(_auto_iopadmap_cc_368_execute_22625_140_), .Y(\digest[140] ));
BUFX2 BUFX2_142 ( .A(_auto_iopadmap_cc_368_execute_22625_141_), .Y(\digest[141] ));
BUFX2 BUFX2_143 ( .A(_auto_iopadmap_cc_368_execute_22625_142_), .Y(\digest[142] ));
BUFX2 BUFX2_144 ( .A(_auto_iopadmap_cc_368_execute_22625_143_), .Y(\digest[143] ));
BUFX2 BUFX2_145 ( .A(_auto_iopadmap_cc_368_execute_22625_144_), .Y(\digest[144] ));
BUFX2 BUFX2_146 ( .A(_auto_iopadmap_cc_368_execute_22625_145_), .Y(\digest[145] ));
BUFX2 BUFX2_147 ( .A(_auto_iopadmap_cc_368_execute_22625_146_), .Y(\digest[146] ));
BUFX2 BUFX2_148 ( .A(_auto_iopadmap_cc_368_execute_22625_147_), .Y(\digest[147] ));
BUFX2 BUFX2_149 ( .A(_auto_iopadmap_cc_368_execute_22625_148_), .Y(\digest[148] ));
BUFX2 BUFX2_15 ( .A(_auto_iopadmap_cc_368_execute_22625_14_), .Y(\digest[14] ));
BUFX2 BUFX2_150 ( .A(_auto_iopadmap_cc_368_execute_22625_149_), .Y(\digest[149] ));
BUFX2 BUFX2_151 ( .A(_auto_iopadmap_cc_368_execute_22625_150_), .Y(\digest[150] ));
BUFX2 BUFX2_152 ( .A(_auto_iopadmap_cc_368_execute_22625_151_), .Y(\digest[151] ));
BUFX2 BUFX2_153 ( .A(_auto_iopadmap_cc_368_execute_22625_152_), .Y(\digest[152] ));
BUFX2 BUFX2_154 ( .A(_auto_iopadmap_cc_368_execute_22625_153_), .Y(\digest[153] ));
BUFX2 BUFX2_155 ( .A(_auto_iopadmap_cc_368_execute_22625_154_), .Y(\digest[154] ));
BUFX2 BUFX2_156 ( .A(_auto_iopadmap_cc_368_execute_22625_155_), .Y(\digest[155] ));
BUFX2 BUFX2_157 ( .A(_auto_iopadmap_cc_368_execute_22625_156_), .Y(\digest[156] ));
BUFX2 BUFX2_158 ( .A(_auto_iopadmap_cc_368_execute_22625_157_), .Y(\digest[157] ));
BUFX2 BUFX2_159 ( .A(_auto_iopadmap_cc_368_execute_22625_158_), .Y(\digest[158] ));
BUFX2 BUFX2_16 ( .A(_auto_iopadmap_cc_368_execute_22625_15_), .Y(\digest[15] ));
BUFX2 BUFX2_160 ( .A(_auto_iopadmap_cc_368_execute_22625_159_), .Y(\digest[159] ));
BUFX2 BUFX2_161 ( .A(_auto_iopadmap_cc_368_execute_22786), .Y(digest_valid));
BUFX2 BUFX2_162 ( .A(_auto_iopadmap_cc_368_execute_22788), .Y(ready));
BUFX2 BUFX2_17 ( .A(_auto_iopadmap_cc_368_execute_22625_16_), .Y(\digest[16] ));
BUFX2 BUFX2_18 ( .A(_auto_iopadmap_cc_368_execute_22625_17_), .Y(\digest[17] ));
BUFX2 BUFX2_19 ( .A(_auto_iopadmap_cc_368_execute_22625_18_), .Y(\digest[18] ));
BUFX2 BUFX2_2 ( .A(_auto_iopadmap_cc_368_execute_22625_1_), .Y(\digest[1] ));
BUFX2 BUFX2_20 ( .A(_auto_iopadmap_cc_368_execute_22625_19_), .Y(\digest[19] ));
BUFX2 BUFX2_21 ( .A(_auto_iopadmap_cc_368_execute_22625_20_), .Y(\digest[20] ));
BUFX2 BUFX2_22 ( .A(_auto_iopadmap_cc_368_execute_22625_21_), .Y(\digest[21] ));
BUFX2 BUFX2_23 ( .A(_auto_iopadmap_cc_368_execute_22625_22_), .Y(\digest[22] ));
BUFX2 BUFX2_24 ( .A(_auto_iopadmap_cc_368_execute_22625_23_), .Y(\digest[23] ));
BUFX2 BUFX2_25 ( .A(_auto_iopadmap_cc_368_execute_22625_24_), .Y(\digest[24] ));
BUFX2 BUFX2_26 ( .A(_auto_iopadmap_cc_368_execute_22625_25_), .Y(\digest[25] ));
BUFX2 BUFX2_27 ( .A(_auto_iopadmap_cc_368_execute_22625_26_), .Y(\digest[26] ));
BUFX2 BUFX2_28 ( .A(_auto_iopadmap_cc_368_execute_22625_27_), .Y(\digest[27] ));
BUFX2 BUFX2_29 ( .A(_auto_iopadmap_cc_368_execute_22625_28_), .Y(\digest[28] ));
BUFX2 BUFX2_3 ( .A(_auto_iopadmap_cc_368_execute_22625_2_), .Y(\digest[2] ));
BUFX2 BUFX2_30 ( .A(_auto_iopadmap_cc_368_execute_22625_29_), .Y(\digest[29] ));
BUFX2 BUFX2_31 ( .A(_auto_iopadmap_cc_368_execute_22625_30_), .Y(\digest[30] ));
BUFX2 BUFX2_32 ( .A(_auto_iopadmap_cc_368_execute_22625_31_), .Y(\digest[31] ));
BUFX2 BUFX2_33 ( .A(_auto_iopadmap_cc_368_execute_22625_32_), .Y(\digest[32] ));
BUFX2 BUFX2_34 ( .A(_auto_iopadmap_cc_368_execute_22625_33_), .Y(\digest[33] ));
BUFX2 BUFX2_35 ( .A(_auto_iopadmap_cc_368_execute_22625_34_), .Y(\digest[34] ));
BUFX2 BUFX2_36 ( .A(_auto_iopadmap_cc_368_execute_22625_35_), .Y(\digest[35] ));
BUFX2 BUFX2_37 ( .A(_auto_iopadmap_cc_368_execute_22625_36_), .Y(\digest[36] ));
BUFX2 BUFX2_38 ( .A(_auto_iopadmap_cc_368_execute_22625_37_), .Y(\digest[37] ));
BUFX2 BUFX2_39 ( .A(_auto_iopadmap_cc_368_execute_22625_38_), .Y(\digest[38] ));
BUFX2 BUFX2_4 ( .A(_auto_iopadmap_cc_368_execute_22625_3_), .Y(\digest[3] ));
BUFX2 BUFX2_40 ( .A(_auto_iopadmap_cc_368_execute_22625_39_), .Y(\digest[39] ));
BUFX2 BUFX2_41 ( .A(_auto_iopadmap_cc_368_execute_22625_40_), .Y(\digest[40] ));
BUFX2 BUFX2_42 ( .A(_auto_iopadmap_cc_368_execute_22625_41_), .Y(\digest[41] ));
BUFX2 BUFX2_43 ( .A(_auto_iopadmap_cc_368_execute_22625_42_), .Y(\digest[42] ));
BUFX2 BUFX2_44 ( .A(_auto_iopadmap_cc_368_execute_22625_43_), .Y(\digest[43] ));
BUFX2 BUFX2_45 ( .A(_auto_iopadmap_cc_368_execute_22625_44_), .Y(\digest[44] ));
BUFX2 BUFX2_46 ( .A(_auto_iopadmap_cc_368_execute_22625_45_), .Y(\digest[45] ));
BUFX2 BUFX2_47 ( .A(_auto_iopadmap_cc_368_execute_22625_46_), .Y(\digest[46] ));
BUFX2 BUFX2_48 ( .A(_auto_iopadmap_cc_368_execute_22625_47_), .Y(\digest[47] ));
BUFX2 BUFX2_49 ( .A(_auto_iopadmap_cc_368_execute_22625_48_), .Y(\digest[48] ));
BUFX2 BUFX2_5 ( .A(_auto_iopadmap_cc_368_execute_22625_4_), .Y(\digest[4] ));
BUFX2 BUFX2_50 ( .A(_auto_iopadmap_cc_368_execute_22625_49_), .Y(\digest[49] ));
BUFX2 BUFX2_51 ( .A(_auto_iopadmap_cc_368_execute_22625_50_), .Y(\digest[50] ));
BUFX2 BUFX2_52 ( .A(_auto_iopadmap_cc_368_execute_22625_51_), .Y(\digest[51] ));
BUFX2 BUFX2_53 ( .A(_auto_iopadmap_cc_368_execute_22625_52_), .Y(\digest[52] ));
BUFX2 BUFX2_54 ( .A(_auto_iopadmap_cc_368_execute_22625_53_), .Y(\digest[53] ));
BUFX2 BUFX2_55 ( .A(_auto_iopadmap_cc_368_execute_22625_54_), .Y(\digest[54] ));
BUFX2 BUFX2_56 ( .A(_auto_iopadmap_cc_368_execute_22625_55_), .Y(\digest[55] ));
BUFX2 BUFX2_57 ( .A(_auto_iopadmap_cc_368_execute_22625_56_), .Y(\digest[56] ));
BUFX2 BUFX2_58 ( .A(_auto_iopadmap_cc_368_execute_22625_57_), .Y(\digest[57] ));
BUFX2 BUFX2_59 ( .A(_auto_iopadmap_cc_368_execute_22625_58_), .Y(\digest[58] ));
BUFX2 BUFX2_6 ( .A(_auto_iopadmap_cc_368_execute_22625_5_), .Y(\digest[5] ));
BUFX2 BUFX2_60 ( .A(_auto_iopadmap_cc_368_execute_22625_59_), .Y(\digest[59] ));
BUFX2 BUFX2_61 ( .A(_auto_iopadmap_cc_368_execute_22625_60_), .Y(\digest[60] ));
BUFX2 BUFX2_62 ( .A(_auto_iopadmap_cc_368_execute_22625_61_), .Y(\digest[61] ));
BUFX2 BUFX2_63 ( .A(_auto_iopadmap_cc_368_execute_22625_62_), .Y(\digest[62] ));
BUFX2 BUFX2_64 ( .A(_auto_iopadmap_cc_368_execute_22625_63_), .Y(\digest[63] ));
BUFX2 BUFX2_65 ( .A(_auto_iopadmap_cc_368_execute_22625_64_), .Y(\digest[64] ));
BUFX2 BUFX2_66 ( .A(_auto_iopadmap_cc_368_execute_22625_65_), .Y(\digest[65] ));
BUFX2 BUFX2_67 ( .A(_auto_iopadmap_cc_368_execute_22625_66_), .Y(\digest[66] ));
BUFX2 BUFX2_68 ( .A(_auto_iopadmap_cc_368_execute_22625_67_), .Y(\digest[67] ));
BUFX2 BUFX2_69 ( .A(_auto_iopadmap_cc_368_execute_22625_68_), .Y(\digest[68] ));
BUFX2 BUFX2_7 ( .A(_auto_iopadmap_cc_368_execute_22625_6_), .Y(\digest[6] ));
BUFX2 BUFX2_70 ( .A(_auto_iopadmap_cc_368_execute_22625_69_), .Y(\digest[69] ));
BUFX2 BUFX2_71 ( .A(_auto_iopadmap_cc_368_execute_22625_70_), .Y(\digest[70] ));
BUFX2 BUFX2_72 ( .A(_auto_iopadmap_cc_368_execute_22625_71_), .Y(\digest[71] ));
BUFX2 BUFX2_73 ( .A(_auto_iopadmap_cc_368_execute_22625_72_), .Y(\digest[72] ));
BUFX2 BUFX2_74 ( .A(_auto_iopadmap_cc_368_execute_22625_73_), .Y(\digest[73] ));
BUFX2 BUFX2_75 ( .A(_auto_iopadmap_cc_368_execute_22625_74_), .Y(\digest[74] ));
BUFX2 BUFX2_76 ( .A(_auto_iopadmap_cc_368_execute_22625_75_), .Y(\digest[75] ));
BUFX2 BUFX2_77 ( .A(_auto_iopadmap_cc_368_execute_22625_76_), .Y(\digest[76] ));
BUFX2 BUFX2_78 ( .A(_auto_iopadmap_cc_368_execute_22625_77_), .Y(\digest[77] ));
BUFX2 BUFX2_79 ( .A(_auto_iopadmap_cc_368_execute_22625_78_), .Y(\digest[78] ));
BUFX2 BUFX2_8 ( .A(_auto_iopadmap_cc_368_execute_22625_7_), .Y(\digest[7] ));
BUFX2 BUFX2_80 ( .A(_auto_iopadmap_cc_368_execute_22625_79_), .Y(\digest[79] ));
BUFX2 BUFX2_81 ( .A(_auto_iopadmap_cc_368_execute_22625_80_), .Y(\digest[80] ));
BUFX2 BUFX2_82 ( .A(_auto_iopadmap_cc_368_execute_22625_81_), .Y(\digest[81] ));
BUFX2 BUFX2_83 ( .A(_auto_iopadmap_cc_368_execute_22625_82_), .Y(\digest[82] ));
BUFX2 BUFX2_84 ( .A(_auto_iopadmap_cc_368_execute_22625_83_), .Y(\digest[83] ));
BUFX2 BUFX2_85 ( .A(_auto_iopadmap_cc_368_execute_22625_84_), .Y(\digest[84] ));
BUFX2 BUFX2_86 ( .A(_auto_iopadmap_cc_368_execute_22625_85_), .Y(\digest[85] ));
BUFX2 BUFX2_87 ( .A(_auto_iopadmap_cc_368_execute_22625_86_), .Y(\digest[86] ));
BUFX2 BUFX2_88 ( .A(_auto_iopadmap_cc_368_execute_22625_87_), .Y(\digest[87] ));
BUFX2 BUFX2_89 ( .A(_auto_iopadmap_cc_368_execute_22625_88_), .Y(\digest[88] ));
BUFX2 BUFX2_9 ( .A(_auto_iopadmap_cc_368_execute_22625_8_), .Y(\digest[8] ));
BUFX2 BUFX2_90 ( .A(_auto_iopadmap_cc_368_execute_22625_89_), .Y(\digest[89] ));
BUFX2 BUFX2_91 ( .A(_auto_iopadmap_cc_368_execute_22625_90_), .Y(\digest[90] ));
BUFX2 BUFX2_92 ( .A(_auto_iopadmap_cc_368_execute_22625_91_), .Y(\digest[91] ));
BUFX2 BUFX2_93 ( .A(_auto_iopadmap_cc_368_execute_22625_92_), .Y(\digest[92] ));
BUFX2 BUFX2_94 ( .A(_auto_iopadmap_cc_368_execute_22625_93_), .Y(\digest[93] ));
BUFX2 BUFX2_95 ( .A(_auto_iopadmap_cc_368_execute_22625_94_), .Y(\digest[94] ));
BUFX2 BUFX2_96 ( .A(_auto_iopadmap_cc_368_execute_22625_95_), .Y(\digest[95] ));
BUFX2 BUFX2_97 ( .A(_auto_iopadmap_cc_368_execute_22625_96_), .Y(\digest[96] ));
BUFX2 BUFX2_98 ( .A(_auto_iopadmap_cc_368_execute_22625_97_), .Y(\digest[97] ));
BUFX2 BUFX2_99 ( .A(_auto_iopadmap_cc_368_execute_22625_98_), .Y(\digest[98] ));
BUFX4 BUFX4_1 ( .A(clk), .Y(clk_hier0_bF_buf8));
BUFX4 BUFX4_10 ( .A(w_mem_inst__abc_19396_new_n2422_), .Y(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf8));
BUFX4 BUFX4_100 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf75));
BUFX4 BUFX4_101 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf74));
BUFX4 BUFX4_102 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf73));
BUFX4 BUFX4_103 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf72));
BUFX4 BUFX4_104 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf71));
BUFX4 BUFX4_105 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf70));
BUFX4 BUFX4_106 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf69));
BUFX4 BUFX4_107 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf68));
BUFX4 BUFX4_108 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf67));
BUFX4 BUFX4_109 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf66));
BUFX4 BUFX4_11 ( .A(w_mem_inst__abc_19396_new_n2422_), .Y(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf7));
BUFX4 BUFX4_110 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf65));
BUFX4 BUFX4_111 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf64));
BUFX4 BUFX4_112 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf63));
BUFX4 BUFX4_113 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf62));
BUFX4 BUFX4_114 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf61));
BUFX4 BUFX4_115 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf60));
BUFX4 BUFX4_116 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf59));
BUFX4 BUFX4_117 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf58));
BUFX4 BUFX4_118 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf57));
BUFX4 BUFX4_119 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf56));
BUFX4 BUFX4_12 ( .A(w_mem_inst__abc_19396_new_n2422_), .Y(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf6));
BUFX4 BUFX4_120 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf55));
BUFX4 BUFX4_121 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf54));
BUFX4 BUFX4_122 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf53));
BUFX4 BUFX4_123 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf52));
BUFX4 BUFX4_124 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf51));
BUFX4 BUFX4_125 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf50));
BUFX4 BUFX4_126 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf49));
BUFX4 BUFX4_127 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf48));
BUFX4 BUFX4_128 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf47));
BUFX4 BUFX4_129 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf46));
BUFX4 BUFX4_13 ( .A(w_mem_inst__abc_19396_new_n2422_), .Y(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf5));
BUFX4 BUFX4_130 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf45));
BUFX4 BUFX4_131 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf44));
BUFX4 BUFX4_132 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf43));
BUFX4 BUFX4_133 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf42));
BUFX4 BUFX4_134 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf41));
BUFX4 BUFX4_135 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf40));
BUFX4 BUFX4_136 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf39));
BUFX4 BUFX4_137 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf38));
BUFX4 BUFX4_138 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf37));
BUFX4 BUFX4_139 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf36));
BUFX4 BUFX4_14 ( .A(w_mem_inst__abc_19396_new_n2422_), .Y(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf4));
BUFX4 BUFX4_140 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf35));
BUFX4 BUFX4_141 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf34));
BUFX4 BUFX4_142 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf33));
BUFX4 BUFX4_143 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf32));
BUFX4 BUFX4_144 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf31));
BUFX4 BUFX4_145 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf30));
BUFX4 BUFX4_146 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf29));
BUFX4 BUFX4_147 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf28));
BUFX4 BUFX4_148 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf27));
BUFX4 BUFX4_149 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf26));
BUFX4 BUFX4_15 ( .A(w_mem_inst__abc_19396_new_n2422_), .Y(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf3));
BUFX4 BUFX4_150 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf25));
BUFX4 BUFX4_151 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf24));
BUFX4 BUFX4_152 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf23));
BUFX4 BUFX4_153 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf22));
BUFX4 BUFX4_154 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf21));
BUFX4 BUFX4_155 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf20));
BUFX4 BUFX4_156 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf19));
BUFX4 BUFX4_157 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf18));
BUFX4 BUFX4_158 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf17));
BUFX4 BUFX4_159 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf16));
BUFX4 BUFX4_16 ( .A(w_mem_inst__abc_19396_new_n2422_), .Y(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf2));
BUFX4 BUFX4_160 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf15));
BUFX4 BUFX4_161 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf14));
BUFX4 BUFX4_162 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf13));
BUFX4 BUFX4_163 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf12));
BUFX4 BUFX4_164 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf11));
BUFX4 BUFX4_165 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf10));
BUFX4 BUFX4_166 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf9));
BUFX4 BUFX4_167 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf8));
BUFX4 BUFX4_168 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf7));
BUFX4 BUFX4_169 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf6));
BUFX4 BUFX4_17 ( .A(w_mem_inst__abc_19396_new_n2422_), .Y(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf1));
BUFX4 BUFX4_170 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf5));
BUFX4 BUFX4_171 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf4));
BUFX4 BUFX4_172 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf3));
BUFX4 BUFX4_173 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf2));
BUFX4 BUFX4_174 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf1));
BUFX4 BUFX4_175 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf0));
BUFX4 BUFX4_176 ( .A(_abc_15497_new_n1650_), .Y(_abc_15497_new_n1650__bF_buf9));
BUFX4 BUFX4_177 ( .A(_abc_15497_new_n1650_), .Y(_abc_15497_new_n1650__bF_buf8));
BUFX4 BUFX4_178 ( .A(_abc_15497_new_n1650_), .Y(_abc_15497_new_n1650__bF_buf7));
BUFX4 BUFX4_179 ( .A(_abc_15497_new_n1650_), .Y(_abc_15497_new_n1650__bF_buf6));
BUFX4 BUFX4_18 ( .A(w_mem_inst__abc_19396_new_n2422_), .Y(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf0));
BUFX4 BUFX4_180 ( .A(_abc_15497_new_n1650_), .Y(_abc_15497_new_n1650__bF_buf5));
BUFX4 BUFX4_181 ( .A(_abc_15497_new_n1650_), .Y(_abc_15497_new_n1650__bF_buf4));
BUFX4 BUFX4_182 ( .A(_abc_15497_new_n1650_), .Y(_abc_15497_new_n1650__bF_buf3));
BUFX4 BUFX4_183 ( .A(_abc_15497_new_n1650_), .Y(_abc_15497_new_n1650__bF_buf2));
BUFX4 BUFX4_184 ( .A(_abc_15497_new_n1650_), .Y(_abc_15497_new_n1650__bF_buf1));
BUFX4 BUFX4_185 ( .A(_abc_15497_new_n1650_), .Y(_abc_15497_new_n1650__bF_buf0));
BUFX4 BUFX4_186 ( .A(w_mem_inst__abc_19396_new_n1637_), .Y(w_mem_inst__abc_19396_new_n1637__bF_buf4));
BUFX4 BUFX4_187 ( .A(w_mem_inst__abc_19396_new_n1637_), .Y(w_mem_inst__abc_19396_new_n1637__bF_buf3));
BUFX4 BUFX4_188 ( .A(w_mem_inst__abc_19396_new_n1637_), .Y(w_mem_inst__abc_19396_new_n1637__bF_buf2));
BUFX4 BUFX4_189 ( .A(w_mem_inst__abc_19396_new_n1637_), .Y(w_mem_inst__abc_19396_new_n1637__bF_buf1));
BUFX4 BUFX4_19 ( .A(w_mem_inst__abc_19396_new_n2421_), .Y(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf6));
BUFX4 BUFX4_190 ( .A(w_mem_inst__abc_19396_new_n1637_), .Y(w_mem_inst__abc_19396_new_n1637__bF_buf0));
BUFX4 BUFX4_191 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf8), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf96));
BUFX4 BUFX4_192 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf7), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf95));
BUFX4 BUFX4_193 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf6), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf94));
BUFX4 BUFX4_194 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf5), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf93));
BUFX4 BUFX4_195 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf4), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf92));
BUFX4 BUFX4_196 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf3), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf91));
BUFX4 BUFX4_197 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf2), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf90));
BUFX4 BUFX4_198 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf1), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf89));
BUFX4 BUFX4_199 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf0), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf88));
BUFX4 BUFX4_2 ( .A(clk), .Y(clk_hier0_bF_buf7));
BUFX4 BUFX4_20 ( .A(w_mem_inst__abc_19396_new_n2421_), .Y(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf5));
BUFX4 BUFX4_200 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf8), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf87));
BUFX4 BUFX4_201 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf7), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf86));
BUFX4 BUFX4_202 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf6), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf85));
BUFX4 BUFX4_203 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf5), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf84));
BUFX4 BUFX4_204 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf4), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf83));
BUFX4 BUFX4_205 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf3), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf82));
BUFX4 BUFX4_206 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf2), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf81));
BUFX4 BUFX4_207 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf1), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf80));
BUFX4 BUFX4_208 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf0), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf79));
BUFX4 BUFX4_209 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf8), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf78));
BUFX4 BUFX4_21 ( .A(w_mem_inst__abc_19396_new_n2421_), .Y(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf4));
BUFX4 BUFX4_210 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf7), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf77));
BUFX4 BUFX4_211 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf6), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf76));
BUFX4 BUFX4_212 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf5), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf75));
BUFX4 BUFX4_213 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf4), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf74));
BUFX4 BUFX4_214 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf3), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf73));
BUFX4 BUFX4_215 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf2), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf72));
BUFX4 BUFX4_216 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf1), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf71));
BUFX4 BUFX4_217 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf0), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf70));
BUFX4 BUFX4_218 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf8), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf69));
BUFX4 BUFX4_219 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf7), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf68));
BUFX4 BUFX4_22 ( .A(w_mem_inst__abc_19396_new_n2421_), .Y(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf3));
BUFX4 BUFX4_220 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf6), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf67));
BUFX4 BUFX4_221 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf5), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf66));
BUFX4 BUFX4_222 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf4), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf65));
BUFX4 BUFX4_223 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf3), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf64));
BUFX4 BUFX4_224 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf2), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf63));
BUFX4 BUFX4_225 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf1), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf62));
BUFX4 BUFX4_226 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf0), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf61));
BUFX4 BUFX4_227 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf8), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf60));
BUFX4 BUFX4_228 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf7), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf59));
BUFX4 BUFX4_229 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf6), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf58));
BUFX4 BUFX4_23 ( .A(w_mem_inst__abc_19396_new_n2421_), .Y(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf2));
BUFX4 BUFX4_230 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf5), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf57));
BUFX4 BUFX4_231 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf4), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf56));
BUFX4 BUFX4_232 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf3), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf55));
BUFX4 BUFX4_233 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf2), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf54));
BUFX4 BUFX4_234 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf1), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf53));
BUFX4 BUFX4_235 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf0), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf52));
BUFX4 BUFX4_236 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf8), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf51));
BUFX4 BUFX4_237 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf7), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf50));
BUFX4 BUFX4_238 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf6), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf49));
BUFX4 BUFX4_239 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf5), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf48));
BUFX4 BUFX4_24 ( .A(w_mem_inst__abc_19396_new_n2421_), .Y(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf1));
BUFX4 BUFX4_240 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf4), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf47));
BUFX4 BUFX4_241 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf3), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf46));
BUFX4 BUFX4_242 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf2), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf45));
BUFX4 BUFX4_243 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf1), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf44));
BUFX4 BUFX4_244 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf0), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf43));
BUFX4 BUFX4_245 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf8), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf42));
BUFX4 BUFX4_246 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf7), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf41));
BUFX4 BUFX4_247 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf6), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf40));
BUFX4 BUFX4_248 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf5), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf39));
BUFX4 BUFX4_249 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf4), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf38));
BUFX4 BUFX4_25 ( .A(w_mem_inst__abc_19396_new_n2421_), .Y(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf0));
BUFX4 BUFX4_250 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf3), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf37));
BUFX4 BUFX4_251 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf2), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf36));
BUFX4 BUFX4_252 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf1), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf35));
BUFX4 BUFX4_253 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf0), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf34));
BUFX4 BUFX4_254 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf8), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf33));
BUFX4 BUFX4_255 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf7), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf32));
BUFX4 BUFX4_256 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf6), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf31));
BUFX4 BUFX4_257 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf5), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf30));
BUFX4 BUFX4_258 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf4), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf29));
BUFX4 BUFX4_259 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf3), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf28));
BUFX4 BUFX4_26 ( .A(reset_n), .Y(reset_n_hier0_bF_buf8));
BUFX4 BUFX4_260 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf2), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf27));
BUFX4 BUFX4_261 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf1), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf26));
BUFX4 BUFX4_262 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf0), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf25));
BUFX4 BUFX4_263 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf8), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf24));
BUFX4 BUFX4_264 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf7), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf23));
BUFX4 BUFX4_265 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf6), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf22));
BUFX4 BUFX4_266 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf5), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf21));
BUFX4 BUFX4_267 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf4), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf20));
BUFX4 BUFX4_268 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf3), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf19));
BUFX4 BUFX4_269 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf2), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf18));
BUFX4 BUFX4_27 ( .A(reset_n), .Y(reset_n_hier0_bF_buf7));
BUFX4 BUFX4_270 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf1), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf17));
BUFX4 BUFX4_271 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf0), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf16));
BUFX4 BUFX4_272 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf8), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf15));
BUFX4 BUFX4_273 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf7), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf14));
BUFX4 BUFX4_274 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf6), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf13));
BUFX4 BUFX4_275 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf5), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf12));
BUFX4 BUFX4_276 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf4), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf11));
BUFX4 BUFX4_277 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf3), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf10));
BUFX4 BUFX4_278 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf2), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf9));
BUFX4 BUFX4_279 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf1), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf8));
BUFX4 BUFX4_28 ( .A(reset_n), .Y(reset_n_hier0_bF_buf6));
BUFX4 BUFX4_280 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf0), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf7));
BUFX4 BUFX4_281 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf8), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf6));
BUFX4 BUFX4_282 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf7), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf5));
BUFX4 BUFX4_283 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf6), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf4));
BUFX4 BUFX4_284 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf5), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf3));
BUFX4 BUFX4_285 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf4), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf2));
BUFX4 BUFX4_286 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf3), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf1));
BUFX4 BUFX4_287 ( .A(w_mem_inst__abc_19396_new_n2422__hier0_bF_buf2), .Y(w_mem_inst__abc_19396_new_n2422__bF_buf0));
BUFX4 BUFX4_288 ( .A(_abc_15497_new_n883_), .Y(_abc_15497_new_n883__bF_buf13));
BUFX4 BUFX4_289 ( .A(_abc_15497_new_n883_), .Y(_abc_15497_new_n883__bF_buf12));
BUFX4 BUFX4_29 ( .A(reset_n), .Y(reset_n_hier0_bF_buf5));
BUFX4 BUFX4_290 ( .A(_abc_15497_new_n883_), .Y(_abc_15497_new_n883__bF_buf11));
BUFX4 BUFX4_291 ( .A(_abc_15497_new_n883_), .Y(_abc_15497_new_n883__bF_buf10));
BUFX4 BUFX4_292 ( .A(_abc_15497_new_n883_), .Y(_abc_15497_new_n883__bF_buf9));
BUFX4 BUFX4_293 ( .A(_abc_15497_new_n883_), .Y(_abc_15497_new_n883__bF_buf8));
BUFX4 BUFX4_294 ( .A(_abc_15497_new_n883_), .Y(_abc_15497_new_n883__bF_buf7));
BUFX4 BUFX4_295 ( .A(_abc_15497_new_n883_), .Y(_abc_15497_new_n883__bF_buf6));
BUFX4 BUFX4_296 ( .A(_abc_15497_new_n883_), .Y(_abc_15497_new_n883__bF_buf5));
BUFX4 BUFX4_297 ( .A(_abc_15497_new_n883_), .Y(_abc_15497_new_n883__bF_buf4));
BUFX4 BUFX4_298 ( .A(_abc_15497_new_n883_), .Y(_abc_15497_new_n883__bF_buf3));
BUFX4 BUFX4_299 ( .A(_abc_15497_new_n883_), .Y(_abc_15497_new_n883__bF_buf2));
BUFX4 BUFX4_3 ( .A(clk), .Y(clk_hier0_bF_buf6));
BUFX4 BUFX4_30 ( .A(reset_n), .Y(reset_n_hier0_bF_buf4));
BUFX4 BUFX4_300 ( .A(_abc_15497_new_n883_), .Y(_abc_15497_new_n883__bF_buf1));
BUFX4 BUFX4_301 ( .A(_abc_15497_new_n883_), .Y(_abc_15497_new_n883__bF_buf0));
BUFX4 BUFX4_302 ( .A(w_mem_inst__abc_19396_new_n1631_), .Y(w_mem_inst__abc_19396_new_n1631__bF_buf4));
BUFX4 BUFX4_303 ( .A(w_mem_inst__abc_19396_new_n1631_), .Y(w_mem_inst__abc_19396_new_n1631__bF_buf3));
BUFX4 BUFX4_304 ( .A(w_mem_inst__abc_19396_new_n1631_), .Y(w_mem_inst__abc_19396_new_n1631__bF_buf2));
BUFX4 BUFX4_305 ( .A(w_mem_inst__abc_19396_new_n1631_), .Y(w_mem_inst__abc_19396_new_n1631__bF_buf1));
BUFX4 BUFX4_306 ( .A(w_mem_inst__abc_19396_new_n1631_), .Y(w_mem_inst__abc_19396_new_n1631__bF_buf0));
BUFX4 BUFX4_307 ( .A(w_mem_inst__abc_19396_new_n1628_), .Y(w_mem_inst__abc_19396_new_n1628__bF_buf4));
BUFX4 BUFX4_308 ( .A(w_mem_inst__abc_19396_new_n1628_), .Y(w_mem_inst__abc_19396_new_n1628__bF_buf3));
BUFX4 BUFX4_309 ( .A(w_mem_inst__abc_19396_new_n1628_), .Y(w_mem_inst__abc_19396_new_n1628__bF_buf2));
BUFX4 BUFX4_31 ( .A(reset_n), .Y(reset_n_hier0_bF_buf3));
BUFX4 BUFX4_310 ( .A(w_mem_inst__abc_19396_new_n1628_), .Y(w_mem_inst__abc_19396_new_n1628__bF_buf1));
BUFX4 BUFX4_311 ( .A(w_mem_inst__abc_19396_new_n1628_), .Y(w_mem_inst__abc_19396_new_n1628__bF_buf0));
BUFX4 BUFX4_312 ( .A(w_mem_inst__abc_19396_new_n1625_), .Y(w_mem_inst__abc_19396_new_n1625__bF_buf4));
BUFX4 BUFX4_313 ( .A(w_mem_inst__abc_19396_new_n1625_), .Y(w_mem_inst__abc_19396_new_n1625__bF_buf3));
BUFX4 BUFX4_314 ( .A(w_mem_inst__abc_19396_new_n1625_), .Y(w_mem_inst__abc_19396_new_n1625__bF_buf2));
BUFX4 BUFX4_315 ( .A(w_mem_inst__abc_19396_new_n1625_), .Y(w_mem_inst__abc_19396_new_n1625__bF_buf1));
BUFX4 BUFX4_316 ( .A(w_mem_inst__abc_19396_new_n1625_), .Y(w_mem_inst__abc_19396_new_n1625__bF_buf0));
BUFX4 BUFX4_317 ( .A(_abc_15497_new_n2743_), .Y(_abc_15497_new_n2743__bF_buf5));
BUFX4 BUFX4_318 ( .A(_abc_15497_new_n2743_), .Y(_abc_15497_new_n2743__bF_buf4));
BUFX4 BUFX4_319 ( .A(_abc_15497_new_n2743_), .Y(_abc_15497_new_n2743__bF_buf3));
BUFX4 BUFX4_32 ( .A(reset_n), .Y(reset_n_hier0_bF_buf2));
BUFX4 BUFX4_320 ( .A(_abc_15497_new_n2743_), .Y(_abc_15497_new_n2743__bF_buf2));
BUFX4 BUFX4_321 ( .A(_abc_15497_new_n2743_), .Y(_abc_15497_new_n2743__bF_buf1));
BUFX4 BUFX4_322 ( .A(_abc_15497_new_n2743_), .Y(_abc_15497_new_n2743__bF_buf0));
BUFX4 BUFX4_323 ( .A(_abc_15497_new_n2781_), .Y(_abc_15497_new_n2781__bF_buf3));
BUFX4 BUFX4_324 ( .A(_abc_15497_new_n2781_), .Y(_abc_15497_new_n2781__bF_buf2));
BUFX4 BUFX4_325 ( .A(_abc_15497_new_n2781_), .Y(_abc_15497_new_n2781__bF_buf1));
BUFX4 BUFX4_326 ( .A(_abc_15497_new_n2781_), .Y(_abc_15497_new_n2781__bF_buf0));
BUFX4 BUFX4_327 ( .A(_abc_15497_new_n871_), .Y(_abc_15497_new_n871__bF_buf4));
BUFX4 BUFX4_328 ( .A(_abc_15497_new_n871_), .Y(_abc_15497_new_n871__bF_buf3));
BUFX4 BUFX4_329 ( .A(_abc_15497_new_n871_), .Y(_abc_15497_new_n871__bF_buf2));
BUFX4 BUFX4_33 ( .A(reset_n), .Y(reset_n_hier0_bF_buf1));
BUFX4 BUFX4_330 ( .A(_abc_15497_new_n871_), .Y(_abc_15497_new_n871__bF_buf1));
BUFX4 BUFX4_331 ( .A(_abc_15497_new_n871_), .Y(_abc_15497_new_n871__bF_buf0));
BUFX4 BUFX4_332 ( .A(w_mem_inst__abc_19396_new_n1619_), .Y(w_mem_inst__abc_19396_new_n1619__bF_buf4));
BUFX4 BUFX4_333 ( .A(w_mem_inst__abc_19396_new_n1619_), .Y(w_mem_inst__abc_19396_new_n1619__bF_buf3));
BUFX4 BUFX4_334 ( .A(w_mem_inst__abc_19396_new_n1619_), .Y(w_mem_inst__abc_19396_new_n1619__bF_buf2));
BUFX4 BUFX4_335 ( .A(w_mem_inst__abc_19396_new_n1619_), .Y(w_mem_inst__abc_19396_new_n1619__bF_buf1));
BUFX4 BUFX4_336 ( .A(w_mem_inst__abc_19396_new_n1619_), .Y(w_mem_inst__abc_19396_new_n1619__bF_buf0));
BUFX4 BUFX4_337 ( .A(w_mem_inst__abc_19396_new_n1598_), .Y(w_mem_inst__abc_19396_new_n1598__bF_buf4));
BUFX4 BUFX4_338 ( .A(w_mem_inst__abc_19396_new_n1598_), .Y(w_mem_inst__abc_19396_new_n1598__bF_buf3));
BUFX4 BUFX4_339 ( .A(w_mem_inst__abc_19396_new_n1598_), .Y(w_mem_inst__abc_19396_new_n1598__bF_buf2));
BUFX4 BUFX4_34 ( .A(reset_n), .Y(reset_n_hier0_bF_buf0));
BUFX4 BUFX4_340 ( .A(w_mem_inst__abc_19396_new_n1598_), .Y(w_mem_inst__abc_19396_new_n1598__bF_buf1));
BUFX4 BUFX4_341 ( .A(w_mem_inst__abc_19396_new_n1598_), .Y(w_mem_inst__abc_19396_new_n1598__bF_buf0));
BUFX4 BUFX4_342 ( .A(_abc_15497_new_n2925_), .Y(_abc_15497_new_n2925__bF_buf3));
BUFX4 BUFX4_343 ( .A(_abc_15497_new_n2925_), .Y(_abc_15497_new_n2925__bF_buf2));
BUFX4 BUFX4_344 ( .A(_abc_15497_new_n2925_), .Y(_abc_15497_new_n2925__bF_buf1));
BUFX4 BUFX4_345 ( .A(_abc_15497_new_n2925_), .Y(_abc_15497_new_n2925__bF_buf0));
BUFX4 BUFX4_346 ( .A(w_mem_inst__abc_19396_new_n1613_), .Y(w_mem_inst__abc_19396_new_n1613__bF_buf4));
BUFX4 BUFX4_347 ( .A(w_mem_inst__abc_19396_new_n1613_), .Y(w_mem_inst__abc_19396_new_n1613__bF_buf3));
BUFX4 BUFX4_348 ( .A(w_mem_inst__abc_19396_new_n1613_), .Y(w_mem_inst__abc_19396_new_n1613__bF_buf2));
BUFX4 BUFX4_349 ( .A(w_mem_inst__abc_19396_new_n1613_), .Y(w_mem_inst__abc_19396_new_n1613__bF_buf1));
BUFX4 BUFX4_35 ( .A(w_mem_inst__abc_19396_new_n2420_), .Y(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf6));
BUFX4 BUFX4_350 ( .A(w_mem_inst__abc_19396_new_n1613_), .Y(w_mem_inst__abc_19396_new_n1613__bF_buf0));
BUFX4 BUFX4_351 ( .A(w_mem_inst__abc_19396_new_n1586_), .Y(w_mem_inst__abc_19396_new_n1586__bF_buf4));
BUFX4 BUFX4_352 ( .A(w_mem_inst__abc_19396_new_n1586_), .Y(w_mem_inst__abc_19396_new_n1586__bF_buf3));
BUFX4 BUFX4_353 ( .A(w_mem_inst__abc_19396_new_n1586_), .Y(w_mem_inst__abc_19396_new_n1586__bF_buf2));
BUFX4 BUFX4_354 ( .A(w_mem_inst__abc_19396_new_n1586_), .Y(w_mem_inst__abc_19396_new_n1586__bF_buf1));
BUFX4 BUFX4_355 ( .A(w_mem_inst__abc_19396_new_n1586_), .Y(w_mem_inst__abc_19396_new_n1586__bF_buf0));
BUFX4 BUFX4_356 ( .A(w_mem_inst__abc_19396_new_n1604_), .Y(w_mem_inst__abc_19396_new_n1604__bF_buf4));
BUFX4 BUFX4_357 ( .A(w_mem_inst__abc_19396_new_n1604_), .Y(w_mem_inst__abc_19396_new_n1604__bF_buf3));
BUFX4 BUFX4_358 ( .A(w_mem_inst__abc_19396_new_n1604_), .Y(w_mem_inst__abc_19396_new_n1604__bF_buf2));
BUFX4 BUFX4_359 ( .A(w_mem_inst__abc_19396_new_n1604_), .Y(w_mem_inst__abc_19396_new_n1604__bF_buf1));
BUFX4 BUFX4_36 ( .A(w_mem_inst__abc_19396_new_n2420_), .Y(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf5));
BUFX4 BUFX4_360 ( .A(w_mem_inst__abc_19396_new_n1604_), .Y(w_mem_inst__abc_19396_new_n1604__bF_buf0));
BUFX4 BUFX4_361 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf6), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf60));
BUFX4 BUFX4_362 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf5), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf59));
BUFX4 BUFX4_363 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf4), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf58));
BUFX4 BUFX4_364 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf3), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf57));
BUFX4 BUFX4_365 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf2), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf56));
BUFX4 BUFX4_366 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf1), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf55));
BUFX4 BUFX4_367 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf0), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf54));
BUFX4 BUFX4_368 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf6), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf53));
BUFX4 BUFX4_369 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf5), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf52));
BUFX4 BUFX4_37 ( .A(w_mem_inst__abc_19396_new_n2420_), .Y(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf4));
BUFX4 BUFX4_370 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf4), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf51));
BUFX4 BUFX4_371 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf3), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf50));
BUFX4 BUFX4_372 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf2), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf49));
BUFX4 BUFX4_373 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf1), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf48));
BUFX4 BUFX4_374 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf0), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf47));
BUFX4 BUFX4_375 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf6), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf46));
BUFX4 BUFX4_376 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf5), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf45));
BUFX4 BUFX4_377 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf4), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf44));
BUFX4 BUFX4_378 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf3), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf43));
BUFX4 BUFX4_379 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf2), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf42));
BUFX4 BUFX4_38 ( .A(w_mem_inst__abc_19396_new_n2420_), .Y(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf3));
BUFX4 BUFX4_380 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf1), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf41));
BUFX4 BUFX4_381 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf0), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf40));
BUFX4 BUFX4_382 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf6), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf39));
BUFX4 BUFX4_383 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf5), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf38));
BUFX4 BUFX4_384 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf4), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf37));
BUFX4 BUFX4_385 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf3), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf36));
BUFX4 BUFX4_386 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf2), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf35));
BUFX4 BUFX4_387 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf1), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf34));
BUFX4 BUFX4_388 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf0), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf33));
BUFX4 BUFX4_389 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf6), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf32));
BUFX4 BUFX4_39 ( .A(w_mem_inst__abc_19396_new_n2420_), .Y(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf2));
BUFX4 BUFX4_390 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf5), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf31));
BUFX4 BUFX4_391 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf4), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf30));
BUFX4 BUFX4_392 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf3), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf29));
BUFX4 BUFX4_393 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf2), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf28));
BUFX4 BUFX4_394 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf1), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf27));
BUFX4 BUFX4_395 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf0), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf26));
BUFX4 BUFX4_396 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf6), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf25));
BUFX4 BUFX4_397 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf5), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf24));
BUFX4 BUFX4_398 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf4), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf23));
BUFX4 BUFX4_399 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf3), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf22));
BUFX4 BUFX4_4 ( .A(clk), .Y(clk_hier0_bF_buf5));
BUFX4 BUFX4_40 ( .A(w_mem_inst__abc_19396_new_n2420_), .Y(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf1));
BUFX4 BUFX4_400 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf2), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf21));
BUFX4 BUFX4_401 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf1), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf20));
BUFX4 BUFX4_402 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf0), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf19));
BUFX4 BUFX4_403 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf6), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf18));
BUFX4 BUFX4_404 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf5), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf17));
BUFX4 BUFX4_405 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf4), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf16));
BUFX4 BUFX4_406 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf3), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf15));
BUFX4 BUFX4_407 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf2), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf14));
BUFX4 BUFX4_408 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf1), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf13));
BUFX4 BUFX4_409 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf0), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf12));
BUFX4 BUFX4_41 ( .A(w_mem_inst__abc_19396_new_n2420_), .Y(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf0));
BUFX4 BUFX4_410 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf6), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf11));
BUFX4 BUFX4_411 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf5), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf10));
BUFX4 BUFX4_412 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf4), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf9));
BUFX4 BUFX4_413 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf3), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf8));
BUFX4 BUFX4_414 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf2), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf7));
BUFX4 BUFX4_415 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf1), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf6));
BUFX4 BUFX4_416 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf0), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf5));
BUFX4 BUFX4_417 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf6), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf4));
BUFX4 BUFX4_418 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf5), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf3));
BUFX4 BUFX4_419 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf4), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf2));
BUFX4 BUFX4_42 ( .A(_abc_15497_new_n872_), .Y(_abc_15497_new_n872__bF_buf4));
BUFX4 BUFX4_420 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf3), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf1));
BUFX4 BUFX4_421 ( .A(w_mem_inst__abc_19396_new_n2421__hier0_bF_buf2), .Y(w_mem_inst__abc_19396_new_n2421__bF_buf0));
BUFX4 BUFX4_422 ( .A(round_ctr_rst), .Y(round_ctr_rst_bF_buf8));
BUFX4 BUFX4_423 ( .A(round_ctr_rst), .Y(round_ctr_rst_bF_buf7));
BUFX4 BUFX4_424 ( .A(round_ctr_rst), .Y(round_ctr_rst_bF_buf6));
BUFX4 BUFX4_425 ( .A(round_ctr_rst), .Y(round_ctr_rst_bF_buf5));
BUFX4 BUFX4_426 ( .A(round_ctr_rst), .Y(round_ctr_rst_bF_buf4));
BUFX4 BUFX4_427 ( .A(round_ctr_rst), .Y(round_ctr_rst_bF_buf3));
BUFX4 BUFX4_428 ( .A(round_ctr_rst), .Y(round_ctr_rst_bF_buf2));
BUFX4 BUFX4_429 ( .A(round_ctr_rst), .Y(round_ctr_rst_bF_buf1));
BUFX4 BUFX4_43 ( .A(_abc_15497_new_n872_), .Y(_abc_15497_new_n872__bF_buf3));
BUFX4 BUFX4_430 ( .A(round_ctr_rst), .Y(round_ctr_rst_bF_buf0));
BUFX4 BUFX4_431 ( .A(w_mem_inst__abc_19396_new_n1630_), .Y(w_mem_inst__abc_19396_new_n1630__bF_buf4));
BUFX4 BUFX4_432 ( .A(w_mem_inst__abc_19396_new_n1630_), .Y(w_mem_inst__abc_19396_new_n1630__bF_buf3));
BUFX4 BUFX4_433 ( .A(w_mem_inst__abc_19396_new_n1630_), .Y(w_mem_inst__abc_19396_new_n1630__bF_buf2));
BUFX4 BUFX4_434 ( .A(w_mem_inst__abc_19396_new_n1630_), .Y(w_mem_inst__abc_19396_new_n1630__bF_buf1));
BUFX4 BUFX4_435 ( .A(w_mem_inst__abc_19396_new_n1630_), .Y(w_mem_inst__abc_19396_new_n1630__bF_buf0));
BUFX4 BUFX4_436 ( .A(w_mem_inst__abc_19396_new_n2582_), .Y(w_mem_inst__abc_19396_new_n2582__bF_buf4));
BUFX4 BUFX4_437 ( .A(w_mem_inst__abc_19396_new_n2582_), .Y(w_mem_inst__abc_19396_new_n2582__bF_buf3));
BUFX4 BUFX4_438 ( .A(w_mem_inst__abc_19396_new_n2582_), .Y(w_mem_inst__abc_19396_new_n2582__bF_buf2));
BUFX4 BUFX4_439 ( .A(w_mem_inst__abc_19396_new_n2582_), .Y(w_mem_inst__abc_19396_new_n2582__bF_buf1));
BUFX4 BUFX4_44 ( .A(_abc_15497_new_n872_), .Y(_abc_15497_new_n872__bF_buf2));
BUFX4 BUFX4_440 ( .A(w_mem_inst__abc_19396_new_n2582_), .Y(w_mem_inst__abc_19396_new_n2582__bF_buf0));
BUFX4 BUFX4_441 ( .A(_abc_15497_new_n873_), .Y(_abc_15497_new_n873__bF_buf7));
BUFX4 BUFX4_442 ( .A(_abc_15497_new_n873_), .Y(_abc_15497_new_n873__bF_buf6));
BUFX4 BUFX4_443 ( .A(_abc_15497_new_n873_), .Y(_abc_15497_new_n873__bF_buf5));
BUFX4 BUFX4_444 ( .A(_abc_15497_new_n873_), .Y(_abc_15497_new_n873__bF_buf4));
BUFX4 BUFX4_445 ( .A(_abc_15497_new_n873_), .Y(_abc_15497_new_n873__bF_buf3));
BUFX4 BUFX4_446 ( .A(_abc_15497_new_n873_), .Y(_abc_15497_new_n873__bF_buf2));
BUFX4 BUFX4_447 ( .A(_abc_15497_new_n873_), .Y(_abc_15497_new_n873__bF_buf1));
BUFX4 BUFX4_448 ( .A(_abc_15497_new_n873_), .Y(_abc_15497_new_n873__bF_buf0));
BUFX4 BUFX4_449 ( .A(_abc_15497_new_n2742_), .Y(_abc_15497_new_n2742__bF_buf3));
BUFX4 BUFX4_45 ( .A(_abc_15497_new_n872_), .Y(_abc_15497_new_n872__bF_buf1));
BUFX4 BUFX4_450 ( .A(_abc_15497_new_n2742_), .Y(_abc_15497_new_n2742__bF_buf2));
BUFX4 BUFX4_451 ( .A(_abc_15497_new_n2742_), .Y(_abc_15497_new_n2742__bF_buf1));
BUFX4 BUFX4_452 ( .A(_abc_15497_new_n2742_), .Y(_abc_15497_new_n2742__bF_buf0));
BUFX4 BUFX4_453 ( .A(_abc_15497_new_n2780_), .Y(_abc_15497_new_n2780__bF_buf3));
BUFX4 BUFX4_454 ( .A(_abc_15497_new_n2780_), .Y(_abc_15497_new_n2780__bF_buf2));
BUFX4 BUFX4_455 ( .A(_abc_15497_new_n2780_), .Y(_abc_15497_new_n2780__bF_buf1));
BUFX4 BUFX4_456 ( .A(_abc_15497_new_n2780_), .Y(_abc_15497_new_n2780__bF_buf0));
BUFX4 BUFX4_457 ( .A(w_mem_inst__abc_19396_new_n1621_), .Y(w_mem_inst__abc_19396_new_n1621__bF_buf4));
BUFX4 BUFX4_458 ( .A(w_mem_inst__abc_19396_new_n1621_), .Y(w_mem_inst__abc_19396_new_n1621__bF_buf3));
BUFX4 BUFX4_459 ( .A(w_mem_inst__abc_19396_new_n1621_), .Y(w_mem_inst__abc_19396_new_n1621__bF_buf2));
BUFX4 BUFX4_46 ( .A(_abc_15497_new_n872_), .Y(_abc_15497_new_n872__bF_buf0));
BUFX4 BUFX4_460 ( .A(w_mem_inst__abc_19396_new_n1621_), .Y(w_mem_inst__abc_19396_new_n1621__bF_buf1));
BUFX4 BUFX4_461 ( .A(w_mem_inst__abc_19396_new_n1621_), .Y(w_mem_inst__abc_19396_new_n1621__bF_buf0));
BUFX4 BUFX4_462 ( .A(_abc_15497_new_n870_), .Y(_abc_15497_new_n870__bF_buf11));
BUFX4 BUFX4_463 ( .A(_abc_15497_new_n870_), .Y(_abc_15497_new_n870__bF_buf10));
BUFX4 BUFX4_464 ( .A(_abc_15497_new_n870_), .Y(_abc_15497_new_n870__bF_buf9));
BUFX4 BUFX4_465 ( .A(_abc_15497_new_n870_), .Y(_abc_15497_new_n870__bF_buf8));
BUFX4 BUFX4_466 ( .A(_abc_15497_new_n870_), .Y(_abc_15497_new_n870__bF_buf7));
BUFX4 BUFX4_467 ( .A(_abc_15497_new_n870_), .Y(_abc_15497_new_n870__bF_buf6));
BUFX4 BUFX4_468 ( .A(_abc_15497_new_n870_), .Y(_abc_15497_new_n870__bF_buf5));
BUFX4 BUFX4_469 ( .A(_abc_15497_new_n870_), .Y(_abc_15497_new_n870__bF_buf4));
BUFX4 BUFX4_47 ( .A(w_mem_inst__abc_19396_new_n1620_), .Y(w_mem_inst__abc_19396_new_n1620__bF_buf7));
BUFX4 BUFX4_470 ( .A(_abc_15497_new_n870_), .Y(_abc_15497_new_n870__bF_buf3));
BUFX4 BUFX4_471 ( .A(_abc_15497_new_n870_), .Y(_abc_15497_new_n870__bF_buf2));
BUFX4 BUFX4_472 ( .A(_abc_15497_new_n870_), .Y(_abc_15497_new_n870__bF_buf1));
BUFX4 BUFX4_473 ( .A(_abc_15497_new_n870_), .Y(_abc_15497_new_n870__bF_buf0));
BUFX4 BUFX4_474 ( .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf88));
BUFX4 BUFX4_475 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf87));
BUFX4 BUFX4_476 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf86));
BUFX4 BUFX4_477 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf85));
BUFX4 BUFX4_478 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf84));
BUFX4 BUFX4_479 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf83));
BUFX4 BUFX4_48 ( .A(w_mem_inst__abc_19396_new_n1620_), .Y(w_mem_inst__abc_19396_new_n1620__bF_buf6));
BUFX4 BUFX4_480 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf82));
BUFX4 BUFX4_481 ( .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf81));
BUFX4 BUFX4_482 ( .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf80));
BUFX4 BUFX4_483 ( .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf79));
BUFX4 BUFX4_484 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf78));
BUFX4 BUFX4_485 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf77));
BUFX4 BUFX4_486 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf76));
BUFX4 BUFX4_487 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf75));
BUFX4 BUFX4_488 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf74));
BUFX4 BUFX4_489 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf73));
BUFX4 BUFX4_49 ( .A(w_mem_inst__abc_19396_new_n1620_), .Y(w_mem_inst__abc_19396_new_n1620__bF_buf5));
BUFX4 BUFX4_490 ( .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf72));
BUFX4 BUFX4_491 ( .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf71));
BUFX4 BUFX4_492 ( .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf70));
BUFX4 BUFX4_493 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf69));
BUFX4 BUFX4_494 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf68));
BUFX4 BUFX4_495 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf67));
BUFX4 BUFX4_496 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf66));
BUFX4 BUFX4_497 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf65));
BUFX4 BUFX4_498 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf64));
BUFX4 BUFX4_499 ( .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf63));
BUFX4 BUFX4_5 ( .A(clk), .Y(clk_hier0_bF_buf4));
BUFX4 BUFX4_50 ( .A(w_mem_inst__abc_19396_new_n1620_), .Y(w_mem_inst__abc_19396_new_n1620__bF_buf4));
BUFX4 BUFX4_500 ( .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf62));
BUFX4 BUFX4_501 ( .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf61));
BUFX4 BUFX4_502 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf60));
BUFX4 BUFX4_503 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf59));
BUFX4 BUFX4_504 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf58));
BUFX4 BUFX4_505 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf57));
BUFX4 BUFX4_506 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf56));
BUFX4 BUFX4_507 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf55));
BUFX4 BUFX4_508 ( .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf54));
BUFX4 BUFX4_509 ( .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf53));
BUFX4 BUFX4_51 ( .A(w_mem_inst__abc_19396_new_n1620_), .Y(w_mem_inst__abc_19396_new_n1620__bF_buf3));
BUFX4 BUFX4_510 ( .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf52));
BUFX4 BUFX4_511 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf51));
BUFX4 BUFX4_512 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf50));
BUFX4 BUFX4_513 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf49));
BUFX4 BUFX4_514 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf48));
BUFX4 BUFX4_515 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf47));
BUFX4 BUFX4_516 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf46));
BUFX4 BUFX4_517 ( .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf45));
BUFX4 BUFX4_518 ( .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf44));
BUFX4 BUFX4_519 ( .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf43));
BUFX4 BUFX4_52 ( .A(w_mem_inst__abc_19396_new_n1620_), .Y(w_mem_inst__abc_19396_new_n1620__bF_buf2));
BUFX4 BUFX4_520 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf42));
BUFX4 BUFX4_521 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf41));
BUFX4 BUFX4_522 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf40));
BUFX4 BUFX4_523 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf39));
BUFX4 BUFX4_524 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf38));
BUFX4 BUFX4_525 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf37));
BUFX4 BUFX4_526 ( .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf36));
BUFX4 BUFX4_527 ( .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf35));
BUFX4 BUFX4_528 ( .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf34));
BUFX4 BUFX4_529 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf33));
BUFX4 BUFX4_53 ( .A(w_mem_inst__abc_19396_new_n1620_), .Y(w_mem_inst__abc_19396_new_n1620__bF_buf1));
BUFX4 BUFX4_530 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf32));
BUFX4 BUFX4_531 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf31));
BUFX4 BUFX4_532 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf30));
BUFX4 BUFX4_533 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf29));
BUFX4 BUFX4_534 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf28));
BUFX4 BUFX4_535 ( .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf27));
BUFX4 BUFX4_536 ( .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf26));
BUFX4 BUFX4_537 ( .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf25));
BUFX4 BUFX4_538 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf24));
BUFX4 BUFX4_539 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf23));
BUFX4 BUFX4_54 ( .A(w_mem_inst__abc_19396_new_n1620_), .Y(w_mem_inst__abc_19396_new_n1620__bF_buf0));
BUFX4 BUFX4_540 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf22));
BUFX4 BUFX4_541 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf21));
BUFX4 BUFX4_542 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf20));
BUFX4 BUFX4_543 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf19));
BUFX4 BUFX4_544 ( .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf18));
BUFX4 BUFX4_545 ( .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf17));
BUFX4 BUFX4_546 ( .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf16));
BUFX4 BUFX4_547 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf15));
BUFX4 BUFX4_548 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf14));
BUFX4 BUFX4_549 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf13));
BUFX4 BUFX4_55 ( .A(w_mem_inst__abc_19396_new_n1617_), .Y(w_mem_inst__abc_19396_new_n1617__bF_buf7));
BUFX4 BUFX4_550 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf12));
BUFX4 BUFX4_551 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf11));
BUFX4 BUFX4_552 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf10));
BUFX4 BUFX4_553 ( .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf9));
BUFX4 BUFX4_554 ( .A(reset_n_hier0_bF_buf0), .Y(reset_n_bF_buf8));
BUFX4 BUFX4_555 ( .A(reset_n_hier0_bF_buf8), .Y(reset_n_bF_buf7));
BUFX4 BUFX4_556 ( .A(reset_n_hier0_bF_buf7), .Y(reset_n_bF_buf6));
BUFX4 BUFX4_557 ( .A(reset_n_hier0_bF_buf6), .Y(reset_n_bF_buf5));
BUFX4 BUFX4_558 ( .A(reset_n_hier0_bF_buf5), .Y(reset_n_bF_buf4));
BUFX4 BUFX4_559 ( .A(reset_n_hier0_bF_buf4), .Y(reset_n_bF_buf3));
BUFX4 BUFX4_56 ( .A(w_mem_inst__abc_19396_new_n1617_), .Y(w_mem_inst__abc_19396_new_n1617__bF_buf6));
BUFX4 BUFX4_560 ( .A(reset_n_hier0_bF_buf3), .Y(reset_n_bF_buf2));
BUFX4 BUFX4_561 ( .A(reset_n_hier0_bF_buf2), .Y(reset_n_bF_buf1));
BUFX4 BUFX4_562 ( .A(reset_n_hier0_bF_buf1), .Y(reset_n_bF_buf0));
BUFX4 BUFX4_563 ( .A(_abc_15497_new_n1663_), .Y(_abc_15497_new_n1663__bF_buf7));
BUFX4 BUFX4_564 ( .A(_abc_15497_new_n1663_), .Y(_abc_15497_new_n1663__bF_buf6));
BUFX4 BUFX4_565 ( .A(_abc_15497_new_n1663_), .Y(_abc_15497_new_n1663__bF_buf5));
BUFX4 BUFX4_566 ( .A(_abc_15497_new_n1663_), .Y(_abc_15497_new_n1663__bF_buf4));
BUFX4 BUFX4_567 ( .A(_abc_15497_new_n1663_), .Y(_abc_15497_new_n1663__bF_buf3));
BUFX4 BUFX4_568 ( .A(_abc_15497_new_n1663_), .Y(_abc_15497_new_n1663__bF_buf2));
BUFX4 BUFX4_569 ( .A(_abc_15497_new_n1663_), .Y(_abc_15497_new_n1663__bF_buf1));
BUFX4 BUFX4_57 ( .A(w_mem_inst__abc_19396_new_n1617_), .Y(w_mem_inst__abc_19396_new_n1617__bF_buf5));
BUFX4 BUFX4_570 ( .A(_abc_15497_new_n1663_), .Y(_abc_15497_new_n1663__bF_buf0));
BUFX4 BUFX4_571 ( .A(_abc_15497_new_n2924_), .Y(_abc_15497_new_n2924__bF_buf4));
BUFX4 BUFX4_572 ( .A(_abc_15497_new_n2924_), .Y(_abc_15497_new_n2924__bF_buf3));
BUFX4 BUFX4_573 ( .A(_abc_15497_new_n2924_), .Y(_abc_15497_new_n2924__bF_buf2));
BUFX4 BUFX4_574 ( .A(_abc_15497_new_n2924_), .Y(_abc_15497_new_n2924__bF_buf1));
BUFX4 BUFX4_575 ( .A(_abc_15497_new_n2924_), .Y(_abc_15497_new_n2924__bF_buf0));
BUFX4 BUFX4_576 ( .A(w_mem_inst__abc_19396_new_n1594_), .Y(w_mem_inst__abc_19396_new_n1594__bF_buf7));
BUFX4 BUFX4_577 ( .A(w_mem_inst__abc_19396_new_n1594_), .Y(w_mem_inst__abc_19396_new_n1594__bF_buf6));
BUFX4 BUFX4_578 ( .A(w_mem_inst__abc_19396_new_n1594_), .Y(w_mem_inst__abc_19396_new_n1594__bF_buf5));
BUFX4 BUFX4_579 ( .A(w_mem_inst__abc_19396_new_n1594_), .Y(w_mem_inst__abc_19396_new_n1594__bF_buf4));
BUFX4 BUFX4_58 ( .A(w_mem_inst__abc_19396_new_n1617_), .Y(w_mem_inst__abc_19396_new_n1617__bF_buf4));
BUFX4 BUFX4_580 ( .A(w_mem_inst__abc_19396_new_n1594_), .Y(w_mem_inst__abc_19396_new_n1594__bF_buf3));
BUFX4 BUFX4_581 ( .A(w_mem_inst__abc_19396_new_n1594_), .Y(w_mem_inst__abc_19396_new_n1594__bF_buf2));
BUFX4 BUFX4_582 ( .A(w_mem_inst__abc_19396_new_n1594_), .Y(w_mem_inst__abc_19396_new_n1594__bF_buf1));
BUFX4 BUFX4_583 ( .A(w_mem_inst__abc_19396_new_n1594_), .Y(w_mem_inst__abc_19396_new_n1594__bF_buf0));
BUFX4 BUFX4_584 ( .A(digest_update), .Y(digest_update_bF_buf8));
BUFX4 BUFX4_585 ( .A(digest_update), .Y(digest_update_bF_buf7));
BUFX4 BUFX4_586 ( .A(digest_update), .Y(digest_update_bF_buf6));
BUFX4 BUFX4_587 ( .A(digest_update), .Y(digest_update_bF_buf5));
BUFX4 BUFX4_588 ( .A(digest_update), .Y(digest_update_bF_buf4));
BUFX4 BUFX4_589 ( .A(digest_update), .Y(digest_update_bF_buf3));
BUFX4 BUFX4_59 ( .A(w_mem_inst__abc_19396_new_n1617_), .Y(w_mem_inst__abc_19396_new_n1617__bF_buf3));
BUFX4 BUFX4_590 ( .A(digest_update), .Y(digest_update_bF_buf2));
BUFX4 BUFX4_591 ( .A(digest_update), .Y(digest_update_bF_buf1));
BUFX4 BUFX4_592 ( .A(digest_update), .Y(digest_update_bF_buf0));
BUFX4 BUFX4_593 ( .A(w_mem_inst__abc_19396_new_n1606_), .Y(w_mem_inst__abc_19396_new_n1606__bF_buf4));
BUFX4 BUFX4_594 ( .A(w_mem_inst__abc_19396_new_n1606_), .Y(w_mem_inst__abc_19396_new_n1606__bF_buf3));
BUFX4 BUFX4_595 ( .A(w_mem_inst__abc_19396_new_n1606_), .Y(w_mem_inst__abc_19396_new_n1606__bF_buf2));
BUFX4 BUFX4_596 ( .A(w_mem_inst__abc_19396_new_n1606_), .Y(w_mem_inst__abc_19396_new_n1606__bF_buf1));
BUFX4 BUFX4_597 ( .A(w_mem_inst__abc_19396_new_n1606_), .Y(w_mem_inst__abc_19396_new_n1606__bF_buf0));
BUFX4 BUFX4_598 ( .A(_abc_15497_new_n2759_), .Y(_abc_15497_new_n2759__bF_buf5));
BUFX4 BUFX4_599 ( .A(_abc_15497_new_n2759_), .Y(_abc_15497_new_n2759__bF_buf4));
BUFX4 BUFX4_6 ( .A(clk), .Y(clk_hier0_bF_buf3));
BUFX4 BUFX4_60 ( .A(w_mem_inst__abc_19396_new_n1617_), .Y(w_mem_inst__abc_19396_new_n1617__bF_buf2));
BUFX4 BUFX4_600 ( .A(_abc_15497_new_n2759_), .Y(_abc_15497_new_n2759__bF_buf3));
BUFX4 BUFX4_601 ( .A(_abc_15497_new_n2759_), .Y(_abc_15497_new_n2759__bF_buf2));
BUFX4 BUFX4_602 ( .A(_abc_15497_new_n2759_), .Y(_abc_15497_new_n2759__bF_buf1));
BUFX4 BUFX4_603 ( .A(_abc_15497_new_n2759_), .Y(_abc_15497_new_n2759__bF_buf0));
BUFX4 BUFX4_604 ( .A(_abc_15497_new_n1648_), .Y(_abc_15497_new_n1648__bF_buf8));
BUFX4 BUFX4_605 ( .A(_abc_15497_new_n1648_), .Y(_abc_15497_new_n1648__bF_buf7));
BUFX4 BUFX4_606 ( .A(_abc_15497_new_n1648_), .Y(_abc_15497_new_n1648__bF_buf6));
BUFX4 BUFX4_607 ( .A(_abc_15497_new_n1648_), .Y(_abc_15497_new_n1648__bF_buf5));
BUFX4 BUFX4_608 ( .A(_abc_15497_new_n1648_), .Y(_abc_15497_new_n1648__bF_buf4));
BUFX4 BUFX4_609 ( .A(_abc_15497_new_n1648_), .Y(_abc_15497_new_n1648__bF_buf3));
BUFX4 BUFX4_61 ( .A(w_mem_inst__abc_19396_new_n1617_), .Y(w_mem_inst__abc_19396_new_n1617__bF_buf1));
BUFX4 BUFX4_610 ( .A(_abc_15497_new_n1648_), .Y(_abc_15497_new_n1648__bF_buf2));
BUFX4 BUFX4_611 ( .A(_abc_15497_new_n1648_), .Y(_abc_15497_new_n1648__bF_buf1));
BUFX4 BUFX4_612 ( .A(_abc_15497_new_n1648_), .Y(_abc_15497_new_n1648__bF_buf0));
BUFX4 BUFX4_613 ( .A(w_mem_inst__abc_19396_new_n1638_), .Y(w_mem_inst__abc_19396_new_n1638__bF_buf4));
BUFX4 BUFX4_614 ( .A(w_mem_inst__abc_19396_new_n1638_), .Y(w_mem_inst__abc_19396_new_n1638__bF_buf3));
BUFX4 BUFX4_615 ( .A(w_mem_inst__abc_19396_new_n1638_), .Y(w_mem_inst__abc_19396_new_n1638__bF_buf2));
BUFX4 BUFX4_616 ( .A(w_mem_inst__abc_19396_new_n1638_), .Y(w_mem_inst__abc_19396_new_n1638__bF_buf1));
BUFX4 BUFX4_617 ( .A(w_mem_inst__abc_19396_new_n1638_), .Y(w_mem_inst__abc_19396_new_n1638__bF_buf0));
BUFX4 BUFX4_618 ( .A(_abc_15497_new_n2756_), .Y(_abc_15497_new_n2756__bF_buf4));
BUFX4 BUFX4_619 ( .A(_abc_15497_new_n2756_), .Y(_abc_15497_new_n2756__bF_buf3));
BUFX4 BUFX4_62 ( .A(w_mem_inst__abc_19396_new_n1617_), .Y(w_mem_inst__abc_19396_new_n1617__bF_buf0));
BUFX4 BUFX4_620 ( .A(_abc_15497_new_n2756_), .Y(_abc_15497_new_n2756__bF_buf2));
BUFX4 BUFX4_621 ( .A(_abc_15497_new_n2756_), .Y(_abc_15497_new_n2756__bF_buf1));
BUFX4 BUFX4_622 ( .A(_abc_15497_new_n2756_), .Y(_abc_15497_new_n2756__bF_buf0));
BUFX4 BUFX4_623 ( .A(w_mem_inst__abc_19396_new_n1635_), .Y(w_mem_inst__abc_19396_new_n1635__bF_buf4));
BUFX4 BUFX4_624 ( .A(w_mem_inst__abc_19396_new_n1635_), .Y(w_mem_inst__abc_19396_new_n1635__bF_buf3));
BUFX4 BUFX4_625 ( .A(w_mem_inst__abc_19396_new_n1635_), .Y(w_mem_inst__abc_19396_new_n1635__bF_buf2));
BUFX4 BUFX4_626 ( .A(w_mem_inst__abc_19396_new_n1635_), .Y(w_mem_inst__abc_19396_new_n1635__bF_buf1));
BUFX4 BUFX4_627 ( .A(w_mem_inst__abc_19396_new_n1635_), .Y(w_mem_inst__abc_19396_new_n1635__bF_buf0));
BUFX4 BUFX4_628 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf6), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf60));
BUFX4 BUFX4_629 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf5), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf59));
BUFX4 BUFX4_63 ( .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf13));
BUFX4 BUFX4_630 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf4), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf58));
BUFX4 BUFX4_631 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf3), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf57));
BUFX4 BUFX4_632 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf2), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf56));
BUFX4 BUFX4_633 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf1), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf55));
BUFX4 BUFX4_634 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf0), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf54));
BUFX4 BUFX4_635 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf6), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf53));
BUFX4 BUFX4_636 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf5), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf52));
BUFX4 BUFX4_637 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf4), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf51));
BUFX4 BUFX4_638 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf3), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf50));
BUFX4 BUFX4_639 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf2), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf49));
BUFX4 BUFX4_64 ( .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf12));
BUFX4 BUFX4_640 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf1), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf48));
BUFX4 BUFX4_641 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf0), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf47));
BUFX4 BUFX4_642 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf6), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf46));
BUFX4 BUFX4_643 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf5), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf45));
BUFX4 BUFX4_644 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf4), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf44));
BUFX4 BUFX4_645 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf3), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf43));
BUFX4 BUFX4_646 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf2), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf42));
BUFX4 BUFX4_647 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf1), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf41));
BUFX4 BUFX4_648 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf0), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf40));
BUFX4 BUFX4_649 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf6), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf39));
BUFX4 BUFX4_65 ( .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf11));
BUFX4 BUFX4_650 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf5), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf38));
BUFX4 BUFX4_651 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf4), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf37));
BUFX4 BUFX4_652 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf3), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf36));
BUFX4 BUFX4_653 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf2), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf35));
BUFX4 BUFX4_654 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf1), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf34));
BUFX4 BUFX4_655 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf0), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf33));
BUFX4 BUFX4_656 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf6), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf32));
BUFX4 BUFX4_657 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf5), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf31));
BUFX4 BUFX4_658 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf4), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf30));
BUFX4 BUFX4_659 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf3), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf29));
BUFX4 BUFX4_66 ( .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf10));
BUFX4 BUFX4_660 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf2), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf28));
BUFX4 BUFX4_661 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf1), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf27));
BUFX4 BUFX4_662 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf0), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf26));
BUFX4 BUFX4_663 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf6), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf25));
BUFX4 BUFX4_664 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf5), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf24));
BUFX4 BUFX4_665 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf4), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf23));
BUFX4 BUFX4_666 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf3), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf22));
BUFX4 BUFX4_667 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf2), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf21));
BUFX4 BUFX4_668 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf1), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf20));
BUFX4 BUFX4_669 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf0), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf19));
BUFX4 BUFX4_67 ( .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf9));
BUFX4 BUFX4_670 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf6), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf18));
BUFX4 BUFX4_671 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf5), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf17));
BUFX4 BUFX4_672 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf4), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf16));
BUFX4 BUFX4_673 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf3), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf15));
BUFX4 BUFX4_674 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf2), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf14));
BUFX4 BUFX4_675 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf1), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf13));
BUFX4 BUFX4_676 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf0), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf12));
BUFX4 BUFX4_677 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf6), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf11));
BUFX4 BUFX4_678 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf5), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf10));
BUFX4 BUFX4_679 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf4), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf9));
BUFX4 BUFX4_68 ( .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf8));
BUFX4 BUFX4_680 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf3), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf8));
BUFX4 BUFX4_681 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf2), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf7));
BUFX4 BUFX4_682 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf1), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf6));
BUFX4 BUFX4_683 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf0), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf5));
BUFX4 BUFX4_684 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf6), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf4));
BUFX4 BUFX4_685 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf5), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf3));
BUFX4 BUFX4_686 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf4), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf2));
BUFX4 BUFX4_687 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf3), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf1));
BUFX4 BUFX4_688 ( .A(w_mem_inst__abc_19396_new_n2420__hier0_bF_buf2), .Y(w_mem_inst__abc_19396_new_n2420__bF_buf0));
BUFX4 BUFX4_69 ( .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf7));
BUFX4 BUFX4_7 ( .A(clk), .Y(clk_hier0_bF_buf2));
BUFX4 BUFX4_70 ( .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf6));
BUFX4 BUFX4_71 ( .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf5));
BUFX4 BUFX4_72 ( .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf4));
BUFX4 BUFX4_73 ( .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf3));
BUFX4 BUFX4_74 ( .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf2));
BUFX4 BUFX4_75 ( .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf1));
BUFX4 BUFX4_76 ( .A(round_ctr_inc), .Y(round_ctr_inc_bF_buf0));
BUFX4 BUFX4_77 ( .A(w_mem_inst__abc_19396_new_n1611_), .Y(w_mem_inst__abc_19396_new_n1611__bF_buf4));
BUFX4 BUFX4_78 ( .A(w_mem_inst__abc_19396_new_n1611_), .Y(w_mem_inst__abc_19396_new_n1611__bF_buf3));
BUFX4 BUFX4_79 ( .A(w_mem_inst__abc_19396_new_n1611_), .Y(w_mem_inst__abc_19396_new_n1611__bF_buf2));
BUFX4 BUFX4_8 ( .A(clk), .Y(clk_hier0_bF_buf1));
BUFX4 BUFX4_80 ( .A(w_mem_inst__abc_19396_new_n1611_), .Y(w_mem_inst__abc_19396_new_n1611__bF_buf1));
BUFX4 BUFX4_81 ( .A(w_mem_inst__abc_19396_new_n1611_), .Y(w_mem_inst__abc_19396_new_n1611__bF_buf0));
BUFX4 BUFX4_82 ( .A(w_mem_inst__abc_19396_new_n1587_), .Y(w_mem_inst__abc_19396_new_n1587__bF_buf4));
BUFX4 BUFX4_83 ( .A(w_mem_inst__abc_19396_new_n1587_), .Y(w_mem_inst__abc_19396_new_n1587__bF_buf3));
BUFX4 BUFX4_84 ( .A(w_mem_inst__abc_19396_new_n1587_), .Y(w_mem_inst__abc_19396_new_n1587__bF_buf2));
BUFX4 BUFX4_85 ( .A(w_mem_inst__abc_19396_new_n1587_), .Y(w_mem_inst__abc_19396_new_n1587__bF_buf1));
BUFX4 BUFX4_86 ( .A(w_mem_inst__abc_19396_new_n1587_), .Y(w_mem_inst__abc_19396_new_n1587__bF_buf0));
BUFX4 BUFX4_87 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf88));
BUFX4 BUFX4_88 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf87));
BUFX4 BUFX4_89 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf86));
BUFX4 BUFX4_9 ( .A(clk), .Y(clk_hier0_bF_buf0));
BUFX4 BUFX4_90 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf85));
BUFX4 BUFX4_91 ( .A(clk_hier0_bF_buf4), .Y(clk_bF_buf84));
BUFX4 BUFX4_92 ( .A(clk_hier0_bF_buf3), .Y(clk_bF_buf83));
BUFX4 BUFX4_93 ( .A(clk_hier0_bF_buf2), .Y(clk_bF_buf82));
BUFX4 BUFX4_94 ( .A(clk_hier0_bF_buf1), .Y(clk_bF_buf81));
BUFX4 BUFX4_95 ( .A(clk_hier0_bF_buf0), .Y(clk_bF_buf80));
BUFX4 BUFX4_96 ( .A(clk_hier0_bF_buf8), .Y(clk_bF_buf79));
BUFX4 BUFX4_97 ( .A(clk_hier0_bF_buf7), .Y(clk_bF_buf78));
BUFX4 BUFX4_98 ( .A(clk_hier0_bF_buf6), .Y(clk_bF_buf77));
BUFX4 BUFX4_99 ( .A(clk_hier0_bF_buf5), .Y(clk_bF_buf76));
DFFSR DFFSR_1 ( .CLK(clk_bF_buf88), .D(_0a_reg_31_0__0_), .Q(a_reg_0_), .R(reset_n_bF_buf88), .S(1'h1));
DFFSR DFFSR_10 ( .CLK(clk_bF_buf79), .D(_0a_reg_31_0__9_), .Q(a_reg_9_), .R(reset_n_bF_buf79), .S(1'h1));
DFFSR DFFSR_100 ( .CLK(clk_bF_buf78), .D(_0d_reg_31_0__3_), .Q(d_reg_3_), .R(reset_n_bF_buf78), .S(1'h1));
DFFSR DFFSR_101 ( .CLK(clk_bF_buf77), .D(_0d_reg_31_0__4_), .Q(d_reg_4_), .R(reset_n_bF_buf77), .S(1'h1));
DFFSR DFFSR_102 ( .CLK(clk_bF_buf76), .D(_0d_reg_31_0__5_), .Q(d_reg_5_), .R(reset_n_bF_buf76), .S(1'h1));
DFFSR DFFSR_103 ( .CLK(clk_bF_buf75), .D(_0d_reg_31_0__6_), .Q(d_reg_6_), .R(reset_n_bF_buf75), .S(1'h1));
DFFSR DFFSR_104 ( .CLK(clk_bF_buf74), .D(_0d_reg_31_0__7_), .Q(d_reg_7_), .R(reset_n_bF_buf74), .S(1'h1));
DFFSR DFFSR_105 ( .CLK(clk_bF_buf73), .D(_0d_reg_31_0__8_), .Q(d_reg_8_), .R(reset_n_bF_buf73), .S(1'h1));
DFFSR DFFSR_106 ( .CLK(clk_bF_buf72), .D(_0d_reg_31_0__9_), .Q(d_reg_9_), .R(reset_n_bF_buf72), .S(1'h1));
DFFSR DFFSR_107 ( .CLK(clk_bF_buf71), .D(_0d_reg_31_0__10_), .Q(d_reg_10_), .R(reset_n_bF_buf71), .S(1'h1));
DFFSR DFFSR_108 ( .CLK(clk_bF_buf70), .D(_0d_reg_31_0__11_), .Q(d_reg_11_), .R(reset_n_bF_buf70), .S(1'h1));
DFFSR DFFSR_109 ( .CLK(clk_bF_buf69), .D(_0d_reg_31_0__12_), .Q(d_reg_12_), .R(reset_n_bF_buf69), .S(1'h1));
DFFSR DFFSR_11 ( .CLK(clk_bF_buf78), .D(_0a_reg_31_0__10_), .Q(a_reg_10_), .R(reset_n_bF_buf78), .S(1'h1));
DFFSR DFFSR_110 ( .CLK(clk_bF_buf68), .D(_0d_reg_31_0__13_), .Q(d_reg_13_), .R(reset_n_bF_buf68), .S(1'h1));
DFFSR DFFSR_111 ( .CLK(clk_bF_buf67), .D(_0d_reg_31_0__14_), .Q(d_reg_14_), .R(reset_n_bF_buf67), .S(1'h1));
DFFSR DFFSR_112 ( .CLK(clk_bF_buf66), .D(_0d_reg_31_0__15_), .Q(d_reg_15_), .R(reset_n_bF_buf66), .S(1'h1));
DFFSR DFFSR_113 ( .CLK(clk_bF_buf65), .D(_0d_reg_31_0__16_), .Q(d_reg_16_), .R(reset_n_bF_buf65), .S(1'h1));
DFFSR DFFSR_114 ( .CLK(clk_bF_buf64), .D(_0d_reg_31_0__17_), .Q(d_reg_17_), .R(reset_n_bF_buf64), .S(1'h1));
DFFSR DFFSR_115 ( .CLK(clk_bF_buf63), .D(_0d_reg_31_0__18_), .Q(d_reg_18_), .R(reset_n_bF_buf63), .S(1'h1));
DFFSR DFFSR_116 ( .CLK(clk_bF_buf62), .D(_0d_reg_31_0__19_), .Q(d_reg_19_), .R(reset_n_bF_buf62), .S(1'h1));
DFFSR DFFSR_117 ( .CLK(clk_bF_buf61), .D(_0d_reg_31_0__20_), .Q(d_reg_20_), .R(reset_n_bF_buf61), .S(1'h1));
DFFSR DFFSR_118 ( .CLK(clk_bF_buf60), .D(_0d_reg_31_0__21_), .Q(d_reg_21_), .R(reset_n_bF_buf60), .S(1'h1));
DFFSR DFFSR_119 ( .CLK(clk_bF_buf59), .D(_0d_reg_31_0__22_), .Q(d_reg_22_), .R(reset_n_bF_buf59), .S(1'h1));
DFFSR DFFSR_12 ( .CLK(clk_bF_buf77), .D(_0a_reg_31_0__11_), .Q(a_reg_11_), .R(reset_n_bF_buf77), .S(1'h1));
DFFSR DFFSR_120 ( .CLK(clk_bF_buf58), .D(_0d_reg_31_0__23_), .Q(d_reg_23_), .R(reset_n_bF_buf58), .S(1'h1));
DFFSR DFFSR_121 ( .CLK(clk_bF_buf57), .D(_0d_reg_31_0__24_), .Q(d_reg_24_), .R(reset_n_bF_buf57), .S(1'h1));
DFFSR DFFSR_122 ( .CLK(clk_bF_buf56), .D(_0d_reg_31_0__25_), .Q(d_reg_25_), .R(reset_n_bF_buf56), .S(1'h1));
DFFSR DFFSR_123 ( .CLK(clk_bF_buf55), .D(_0d_reg_31_0__26_), .Q(d_reg_26_), .R(reset_n_bF_buf55), .S(1'h1));
DFFSR DFFSR_124 ( .CLK(clk_bF_buf54), .D(_0d_reg_31_0__27_), .Q(d_reg_27_), .R(reset_n_bF_buf54), .S(1'h1));
DFFSR DFFSR_125 ( .CLK(clk_bF_buf53), .D(_0d_reg_31_0__28_), .Q(d_reg_28_), .R(reset_n_bF_buf53), .S(1'h1));
DFFSR DFFSR_126 ( .CLK(clk_bF_buf52), .D(_0d_reg_31_0__29_), .Q(d_reg_29_), .R(reset_n_bF_buf52), .S(1'h1));
DFFSR DFFSR_127 ( .CLK(clk_bF_buf51), .D(_0d_reg_31_0__30_), .Q(d_reg_30_), .R(reset_n_bF_buf51), .S(1'h1));
DFFSR DFFSR_128 ( .CLK(clk_bF_buf50), .D(_0d_reg_31_0__31_), .Q(d_reg_31_), .R(reset_n_bF_buf50), .S(1'h1));
DFFSR DFFSR_129 ( .CLK(clk_bF_buf49), .D(_0e_reg_31_0__0_), .Q(e_reg_0_), .R(reset_n_bF_buf49), .S(1'h1));
DFFSR DFFSR_13 ( .CLK(clk_bF_buf76), .D(_0a_reg_31_0__12_), .Q(a_reg_12_), .R(reset_n_bF_buf76), .S(1'h1));
DFFSR DFFSR_130 ( .CLK(clk_bF_buf48), .D(_0e_reg_31_0__1_), .Q(e_reg_1_), .R(reset_n_bF_buf48), .S(1'h1));
DFFSR DFFSR_131 ( .CLK(clk_bF_buf47), .D(_0e_reg_31_0__2_), .Q(e_reg_2_), .R(reset_n_bF_buf47), .S(1'h1));
DFFSR DFFSR_132 ( .CLK(clk_bF_buf46), .D(_0e_reg_31_0__3_), .Q(e_reg_3_), .R(reset_n_bF_buf46), .S(1'h1));
DFFSR DFFSR_133 ( .CLK(clk_bF_buf45), .D(_0e_reg_31_0__4_), .Q(e_reg_4_), .R(reset_n_bF_buf45), .S(1'h1));
DFFSR DFFSR_134 ( .CLK(clk_bF_buf44), .D(_0e_reg_31_0__5_), .Q(e_reg_5_), .R(reset_n_bF_buf44), .S(1'h1));
DFFSR DFFSR_135 ( .CLK(clk_bF_buf43), .D(_0e_reg_31_0__6_), .Q(e_reg_6_), .R(reset_n_bF_buf43), .S(1'h1));
DFFSR DFFSR_136 ( .CLK(clk_bF_buf42), .D(_0e_reg_31_0__7_), .Q(e_reg_7_), .R(reset_n_bF_buf42), .S(1'h1));
DFFSR DFFSR_137 ( .CLK(clk_bF_buf41), .D(_0e_reg_31_0__8_), .Q(e_reg_8_), .R(reset_n_bF_buf41), .S(1'h1));
DFFSR DFFSR_138 ( .CLK(clk_bF_buf40), .D(_0e_reg_31_0__9_), .Q(e_reg_9_), .R(reset_n_bF_buf40), .S(1'h1));
DFFSR DFFSR_139 ( .CLK(clk_bF_buf39), .D(_0e_reg_31_0__10_), .Q(e_reg_10_), .R(reset_n_bF_buf39), .S(1'h1));
DFFSR DFFSR_14 ( .CLK(clk_bF_buf75), .D(_0a_reg_31_0__13_), .Q(a_reg_13_), .R(reset_n_bF_buf75), .S(1'h1));
DFFSR DFFSR_140 ( .CLK(clk_bF_buf38), .D(_0e_reg_31_0__11_), .Q(e_reg_11_), .R(reset_n_bF_buf38), .S(1'h1));
DFFSR DFFSR_141 ( .CLK(clk_bF_buf37), .D(_0e_reg_31_0__12_), .Q(e_reg_12_), .R(reset_n_bF_buf37), .S(1'h1));
DFFSR DFFSR_142 ( .CLK(clk_bF_buf36), .D(_0e_reg_31_0__13_), .Q(e_reg_13_), .R(reset_n_bF_buf36), .S(1'h1));
DFFSR DFFSR_143 ( .CLK(clk_bF_buf35), .D(_0e_reg_31_0__14_), .Q(e_reg_14_), .R(reset_n_bF_buf35), .S(1'h1));
DFFSR DFFSR_144 ( .CLK(clk_bF_buf34), .D(_0e_reg_31_0__15_), .Q(e_reg_15_), .R(reset_n_bF_buf34), .S(1'h1));
DFFSR DFFSR_145 ( .CLK(clk_bF_buf33), .D(_0e_reg_31_0__16_), .Q(e_reg_16_), .R(reset_n_bF_buf33), .S(1'h1));
DFFSR DFFSR_146 ( .CLK(clk_bF_buf32), .D(_0e_reg_31_0__17_), .Q(e_reg_17_), .R(reset_n_bF_buf32), .S(1'h1));
DFFSR DFFSR_147 ( .CLK(clk_bF_buf31), .D(_0e_reg_31_0__18_), .Q(e_reg_18_), .R(reset_n_bF_buf31), .S(1'h1));
DFFSR DFFSR_148 ( .CLK(clk_bF_buf30), .D(_0e_reg_31_0__19_), .Q(e_reg_19_), .R(reset_n_bF_buf30), .S(1'h1));
DFFSR DFFSR_149 ( .CLK(clk_bF_buf29), .D(_0e_reg_31_0__20_), .Q(e_reg_20_), .R(reset_n_bF_buf29), .S(1'h1));
DFFSR DFFSR_15 ( .CLK(clk_bF_buf74), .D(_0a_reg_31_0__14_), .Q(a_reg_14_), .R(reset_n_bF_buf74), .S(1'h1));
DFFSR DFFSR_150 ( .CLK(clk_bF_buf28), .D(_0e_reg_31_0__21_), .Q(e_reg_21_), .R(reset_n_bF_buf28), .S(1'h1));
DFFSR DFFSR_151 ( .CLK(clk_bF_buf27), .D(_0e_reg_31_0__22_), .Q(e_reg_22_), .R(reset_n_bF_buf27), .S(1'h1));
DFFSR DFFSR_152 ( .CLK(clk_bF_buf26), .D(_0e_reg_31_0__23_), .Q(e_reg_23_), .R(reset_n_bF_buf26), .S(1'h1));
DFFSR DFFSR_153 ( .CLK(clk_bF_buf25), .D(_0e_reg_31_0__24_), .Q(e_reg_24_), .R(reset_n_bF_buf25), .S(1'h1));
DFFSR DFFSR_154 ( .CLK(clk_bF_buf24), .D(_0e_reg_31_0__25_), .Q(e_reg_25_), .R(reset_n_bF_buf24), .S(1'h1));
DFFSR DFFSR_155 ( .CLK(clk_bF_buf23), .D(_0e_reg_31_0__26_), .Q(e_reg_26_), .R(reset_n_bF_buf23), .S(1'h1));
DFFSR DFFSR_156 ( .CLK(clk_bF_buf22), .D(_0e_reg_31_0__27_), .Q(e_reg_27_), .R(reset_n_bF_buf22), .S(1'h1));
DFFSR DFFSR_157 ( .CLK(clk_bF_buf21), .D(_0e_reg_31_0__28_), .Q(e_reg_28_), .R(reset_n_bF_buf21), .S(1'h1));
DFFSR DFFSR_158 ( .CLK(clk_bF_buf20), .D(_0e_reg_31_0__29_), .Q(e_reg_29_), .R(reset_n_bF_buf20), .S(1'h1));
DFFSR DFFSR_159 ( .CLK(clk_bF_buf19), .D(_0e_reg_31_0__30_), .Q(e_reg_30_), .R(reset_n_bF_buf19), .S(1'h1));
DFFSR DFFSR_16 ( .CLK(clk_bF_buf73), .D(_0a_reg_31_0__15_), .Q(a_reg_15_), .R(reset_n_bF_buf73), .S(1'h1));
DFFSR DFFSR_160 ( .CLK(clk_bF_buf18), .D(_0e_reg_31_0__31_), .Q(e_reg_31_), .R(reset_n_bF_buf18), .S(1'h1));
DFFSR DFFSR_161 ( .CLK(clk_bF_buf17), .D(_0H0_reg_31_0__0_), .Q(_auto_iopadmap_cc_368_execute_22625_128_), .R(reset_n_bF_buf17), .S(1'h1));
DFFSR DFFSR_162 ( .CLK(clk_bF_buf16), .D(_0H0_reg_31_0__1_), .Q(_auto_iopadmap_cc_368_execute_22625_129_), .R(reset_n_bF_buf16), .S(1'h1));
DFFSR DFFSR_163 ( .CLK(clk_bF_buf15), .D(_0H0_reg_31_0__2_), .Q(_auto_iopadmap_cc_368_execute_22625_130_), .R(reset_n_bF_buf15), .S(1'h1));
DFFSR DFFSR_164 ( .CLK(clk_bF_buf14), .D(_0H0_reg_31_0__3_), .Q(_auto_iopadmap_cc_368_execute_22625_131_), .R(reset_n_bF_buf14), .S(1'h1));
DFFSR DFFSR_165 ( .CLK(clk_bF_buf13), .D(_0H0_reg_31_0__4_), .Q(_auto_iopadmap_cc_368_execute_22625_132_), .R(reset_n_bF_buf13), .S(1'h1));
DFFSR DFFSR_166 ( .CLK(clk_bF_buf12), .D(_0H0_reg_31_0__5_), .Q(_auto_iopadmap_cc_368_execute_22625_133_), .R(reset_n_bF_buf12), .S(1'h1));
DFFSR DFFSR_167 ( .CLK(clk_bF_buf11), .D(_0H0_reg_31_0__6_), .Q(_auto_iopadmap_cc_368_execute_22625_134_), .R(reset_n_bF_buf11), .S(1'h1));
DFFSR DFFSR_168 ( .CLK(clk_bF_buf10), .D(_0H0_reg_31_0__7_), .Q(_auto_iopadmap_cc_368_execute_22625_135_), .R(reset_n_bF_buf10), .S(1'h1));
DFFSR DFFSR_169 ( .CLK(clk_bF_buf9), .D(_0H0_reg_31_0__8_), .Q(_auto_iopadmap_cc_368_execute_22625_136_), .R(reset_n_bF_buf9), .S(1'h1));
DFFSR DFFSR_17 ( .CLK(clk_bF_buf72), .D(_0a_reg_31_0__16_), .Q(a_reg_16_), .R(reset_n_bF_buf72), .S(1'h1));
DFFSR DFFSR_170 ( .CLK(clk_bF_buf8), .D(_0H0_reg_31_0__9_), .Q(_auto_iopadmap_cc_368_execute_22625_137_), .R(reset_n_bF_buf8), .S(1'h1));
DFFSR DFFSR_171 ( .CLK(clk_bF_buf7), .D(_0H0_reg_31_0__10_), .Q(_auto_iopadmap_cc_368_execute_22625_138_), .R(reset_n_bF_buf7), .S(1'h1));
DFFSR DFFSR_172 ( .CLK(clk_bF_buf6), .D(_0H0_reg_31_0__11_), .Q(_auto_iopadmap_cc_368_execute_22625_139_), .R(reset_n_bF_buf6), .S(1'h1));
DFFSR DFFSR_173 ( .CLK(clk_bF_buf5), .D(_0H0_reg_31_0__12_), .Q(_auto_iopadmap_cc_368_execute_22625_140_), .R(reset_n_bF_buf5), .S(1'h1));
DFFSR DFFSR_174 ( .CLK(clk_bF_buf4), .D(_0H0_reg_31_0__13_), .Q(_auto_iopadmap_cc_368_execute_22625_141_), .R(reset_n_bF_buf4), .S(1'h1));
DFFSR DFFSR_175 ( .CLK(clk_bF_buf3), .D(_0H0_reg_31_0__14_), .Q(_auto_iopadmap_cc_368_execute_22625_142_), .R(reset_n_bF_buf3), .S(1'h1));
DFFSR DFFSR_176 ( .CLK(clk_bF_buf2), .D(_0H0_reg_31_0__15_), .Q(_auto_iopadmap_cc_368_execute_22625_143_), .R(reset_n_bF_buf2), .S(1'h1));
DFFSR DFFSR_177 ( .CLK(clk_bF_buf1), .D(_0H0_reg_31_0__16_), .Q(_auto_iopadmap_cc_368_execute_22625_144_), .R(reset_n_bF_buf1), .S(1'h1));
DFFSR DFFSR_178 ( .CLK(clk_bF_buf0), .D(_0H0_reg_31_0__17_), .Q(_auto_iopadmap_cc_368_execute_22625_145_), .R(reset_n_bF_buf0), .S(1'h1));
DFFSR DFFSR_179 ( .CLK(clk_bF_buf88), .D(_0H0_reg_31_0__18_), .Q(_auto_iopadmap_cc_368_execute_22625_146_), .R(reset_n_bF_buf88), .S(1'h1));
DFFSR DFFSR_18 ( .CLK(clk_bF_buf71), .D(_0a_reg_31_0__17_), .Q(a_reg_17_), .R(reset_n_bF_buf71), .S(1'h1));
DFFSR DFFSR_180 ( .CLK(clk_bF_buf87), .D(_0H0_reg_31_0__19_), .Q(_auto_iopadmap_cc_368_execute_22625_147_), .R(reset_n_bF_buf87), .S(1'h1));
DFFSR DFFSR_181 ( .CLK(clk_bF_buf86), .D(_0H0_reg_31_0__20_), .Q(_auto_iopadmap_cc_368_execute_22625_148_), .R(reset_n_bF_buf86), .S(1'h1));
DFFSR DFFSR_182 ( .CLK(clk_bF_buf85), .D(_0H0_reg_31_0__21_), .Q(_auto_iopadmap_cc_368_execute_22625_149_), .R(reset_n_bF_buf85), .S(1'h1));
DFFSR DFFSR_183 ( .CLK(clk_bF_buf84), .D(_0H0_reg_31_0__22_), .Q(_auto_iopadmap_cc_368_execute_22625_150_), .R(reset_n_bF_buf84), .S(1'h1));
DFFSR DFFSR_184 ( .CLK(clk_bF_buf83), .D(_0H0_reg_31_0__23_), .Q(_auto_iopadmap_cc_368_execute_22625_151_), .R(reset_n_bF_buf83), .S(1'h1));
DFFSR DFFSR_185 ( .CLK(clk_bF_buf82), .D(_0H0_reg_31_0__24_), .Q(_auto_iopadmap_cc_368_execute_22625_152_), .R(reset_n_bF_buf82), .S(1'h1));
DFFSR DFFSR_186 ( .CLK(clk_bF_buf81), .D(_0H0_reg_31_0__25_), .Q(_auto_iopadmap_cc_368_execute_22625_153_), .R(reset_n_bF_buf81), .S(1'h1));
DFFSR DFFSR_187 ( .CLK(clk_bF_buf80), .D(_0H0_reg_31_0__26_), .Q(_auto_iopadmap_cc_368_execute_22625_154_), .R(reset_n_bF_buf80), .S(1'h1));
DFFSR DFFSR_188 ( .CLK(clk_bF_buf79), .D(_0H0_reg_31_0__27_), .Q(_auto_iopadmap_cc_368_execute_22625_155_), .R(reset_n_bF_buf79), .S(1'h1));
DFFSR DFFSR_189 ( .CLK(clk_bF_buf78), .D(_0H0_reg_31_0__28_), .Q(_auto_iopadmap_cc_368_execute_22625_156_), .R(reset_n_bF_buf78), .S(1'h1));
DFFSR DFFSR_19 ( .CLK(clk_bF_buf70), .D(_0a_reg_31_0__18_), .Q(a_reg_18_), .R(reset_n_bF_buf70), .S(1'h1));
DFFSR DFFSR_190 ( .CLK(clk_bF_buf77), .D(_0H0_reg_31_0__29_), .Q(_auto_iopadmap_cc_368_execute_22625_157_), .R(reset_n_bF_buf77), .S(1'h1));
DFFSR DFFSR_191 ( .CLK(clk_bF_buf76), .D(_0H0_reg_31_0__30_), .Q(_auto_iopadmap_cc_368_execute_22625_158_), .R(reset_n_bF_buf76), .S(1'h1));
DFFSR DFFSR_192 ( .CLK(clk_bF_buf75), .D(_0H0_reg_31_0__31_), .Q(_auto_iopadmap_cc_368_execute_22625_159_), .R(reset_n_bF_buf75), .S(1'h1));
DFFSR DFFSR_193 ( .CLK(clk_bF_buf74), .D(_0H1_reg_31_0__0_), .Q(_auto_iopadmap_cc_368_execute_22625_96_), .R(reset_n_bF_buf74), .S(1'h1));
DFFSR DFFSR_194 ( .CLK(clk_bF_buf73), .D(_0H1_reg_31_0__1_), .Q(_auto_iopadmap_cc_368_execute_22625_97_), .R(reset_n_bF_buf73), .S(1'h1));
DFFSR DFFSR_195 ( .CLK(clk_bF_buf72), .D(_0H1_reg_31_0__2_), .Q(_auto_iopadmap_cc_368_execute_22625_98_), .R(reset_n_bF_buf72), .S(1'h1));
DFFSR DFFSR_196 ( .CLK(clk_bF_buf71), .D(_0H1_reg_31_0__3_), .Q(_auto_iopadmap_cc_368_execute_22625_99_), .R(reset_n_bF_buf71), .S(1'h1));
DFFSR DFFSR_197 ( .CLK(clk_bF_buf70), .D(_0H1_reg_31_0__4_), .Q(_auto_iopadmap_cc_368_execute_22625_100_), .R(reset_n_bF_buf70), .S(1'h1));
DFFSR DFFSR_198 ( .CLK(clk_bF_buf69), .D(_0H1_reg_31_0__5_), .Q(_auto_iopadmap_cc_368_execute_22625_101_), .R(reset_n_bF_buf69), .S(1'h1));
DFFSR DFFSR_199 ( .CLK(clk_bF_buf68), .D(_0H1_reg_31_0__6_), .Q(_auto_iopadmap_cc_368_execute_22625_102_), .R(reset_n_bF_buf68), .S(1'h1));
DFFSR DFFSR_2 ( .CLK(clk_bF_buf87), .D(_0a_reg_31_0__1_), .Q(a_reg_1_), .R(reset_n_bF_buf87), .S(1'h1));
DFFSR DFFSR_20 ( .CLK(clk_bF_buf69), .D(_0a_reg_31_0__19_), .Q(a_reg_19_), .R(reset_n_bF_buf69), .S(1'h1));
DFFSR DFFSR_200 ( .CLK(clk_bF_buf67), .D(_0H1_reg_31_0__7_), .Q(_auto_iopadmap_cc_368_execute_22625_103_), .R(reset_n_bF_buf67), .S(1'h1));
DFFSR DFFSR_201 ( .CLK(clk_bF_buf66), .D(_0H1_reg_31_0__8_), .Q(_auto_iopadmap_cc_368_execute_22625_104_), .R(reset_n_bF_buf66), .S(1'h1));
DFFSR DFFSR_202 ( .CLK(clk_bF_buf65), .D(_0H1_reg_31_0__9_), .Q(_auto_iopadmap_cc_368_execute_22625_105_), .R(reset_n_bF_buf65), .S(1'h1));
DFFSR DFFSR_203 ( .CLK(clk_bF_buf64), .D(_0H1_reg_31_0__10_), .Q(_auto_iopadmap_cc_368_execute_22625_106_), .R(reset_n_bF_buf64), .S(1'h1));
DFFSR DFFSR_204 ( .CLK(clk_bF_buf63), .D(_0H1_reg_31_0__11_), .Q(_auto_iopadmap_cc_368_execute_22625_107_), .R(reset_n_bF_buf63), .S(1'h1));
DFFSR DFFSR_205 ( .CLK(clk_bF_buf62), .D(_0H1_reg_31_0__12_), .Q(_auto_iopadmap_cc_368_execute_22625_108_), .R(reset_n_bF_buf62), .S(1'h1));
DFFSR DFFSR_206 ( .CLK(clk_bF_buf61), .D(_0H1_reg_31_0__13_), .Q(_auto_iopadmap_cc_368_execute_22625_109_), .R(reset_n_bF_buf61), .S(1'h1));
DFFSR DFFSR_207 ( .CLK(clk_bF_buf60), .D(_0H1_reg_31_0__14_), .Q(_auto_iopadmap_cc_368_execute_22625_110_), .R(reset_n_bF_buf60), .S(1'h1));
DFFSR DFFSR_208 ( .CLK(clk_bF_buf59), .D(_0H1_reg_31_0__15_), .Q(_auto_iopadmap_cc_368_execute_22625_111_), .R(reset_n_bF_buf59), .S(1'h1));
DFFSR DFFSR_209 ( .CLK(clk_bF_buf58), .D(_0H1_reg_31_0__16_), .Q(_auto_iopadmap_cc_368_execute_22625_112_), .R(reset_n_bF_buf58), .S(1'h1));
DFFSR DFFSR_21 ( .CLK(clk_bF_buf68), .D(_0a_reg_31_0__20_), .Q(a_reg_20_), .R(reset_n_bF_buf68), .S(1'h1));
DFFSR DFFSR_210 ( .CLK(clk_bF_buf57), .D(_0H1_reg_31_0__17_), .Q(_auto_iopadmap_cc_368_execute_22625_113_), .R(reset_n_bF_buf57), .S(1'h1));
DFFSR DFFSR_211 ( .CLK(clk_bF_buf56), .D(_0H1_reg_31_0__18_), .Q(_auto_iopadmap_cc_368_execute_22625_114_), .R(reset_n_bF_buf56), .S(1'h1));
DFFSR DFFSR_212 ( .CLK(clk_bF_buf55), .D(_0H1_reg_31_0__19_), .Q(_auto_iopadmap_cc_368_execute_22625_115_), .R(reset_n_bF_buf55), .S(1'h1));
DFFSR DFFSR_213 ( .CLK(clk_bF_buf54), .D(_0H1_reg_31_0__20_), .Q(_auto_iopadmap_cc_368_execute_22625_116_), .R(reset_n_bF_buf54), .S(1'h1));
DFFSR DFFSR_214 ( .CLK(clk_bF_buf53), .D(_0H1_reg_31_0__21_), .Q(_auto_iopadmap_cc_368_execute_22625_117_), .R(reset_n_bF_buf53), .S(1'h1));
DFFSR DFFSR_215 ( .CLK(clk_bF_buf52), .D(_0H1_reg_31_0__22_), .Q(_auto_iopadmap_cc_368_execute_22625_118_), .R(reset_n_bF_buf52), .S(1'h1));
DFFSR DFFSR_216 ( .CLK(clk_bF_buf51), .D(_0H1_reg_31_0__23_), .Q(_auto_iopadmap_cc_368_execute_22625_119_), .R(reset_n_bF_buf51), .S(1'h1));
DFFSR DFFSR_217 ( .CLK(clk_bF_buf50), .D(_0H1_reg_31_0__24_), .Q(_auto_iopadmap_cc_368_execute_22625_120_), .R(reset_n_bF_buf50), .S(1'h1));
DFFSR DFFSR_218 ( .CLK(clk_bF_buf49), .D(_0H1_reg_31_0__25_), .Q(_auto_iopadmap_cc_368_execute_22625_121_), .R(reset_n_bF_buf49), .S(1'h1));
DFFSR DFFSR_219 ( .CLK(clk_bF_buf48), .D(_0H1_reg_31_0__26_), .Q(_auto_iopadmap_cc_368_execute_22625_122_), .R(reset_n_bF_buf48), .S(1'h1));
DFFSR DFFSR_22 ( .CLK(clk_bF_buf67), .D(_0a_reg_31_0__21_), .Q(a_reg_21_), .R(reset_n_bF_buf67), .S(1'h1));
DFFSR DFFSR_220 ( .CLK(clk_bF_buf47), .D(_0H1_reg_31_0__27_), .Q(_auto_iopadmap_cc_368_execute_22625_123_), .R(reset_n_bF_buf47), .S(1'h1));
DFFSR DFFSR_221 ( .CLK(clk_bF_buf46), .D(_0H1_reg_31_0__28_), .Q(_auto_iopadmap_cc_368_execute_22625_124_), .R(reset_n_bF_buf46), .S(1'h1));
DFFSR DFFSR_222 ( .CLK(clk_bF_buf45), .D(_0H1_reg_31_0__29_), .Q(_auto_iopadmap_cc_368_execute_22625_125_), .R(reset_n_bF_buf45), .S(1'h1));
DFFSR DFFSR_223 ( .CLK(clk_bF_buf44), .D(_0H1_reg_31_0__30_), .Q(_auto_iopadmap_cc_368_execute_22625_126_), .R(reset_n_bF_buf44), .S(1'h1));
DFFSR DFFSR_224 ( .CLK(clk_bF_buf43), .D(_0H1_reg_31_0__31_), .Q(_auto_iopadmap_cc_368_execute_22625_127_), .R(reset_n_bF_buf43), .S(1'h1));
DFFSR DFFSR_225 ( .CLK(clk_bF_buf42), .D(_0H2_reg_31_0__0_), .Q(_auto_iopadmap_cc_368_execute_22625_64_), .R(reset_n_bF_buf42), .S(1'h1));
DFFSR DFFSR_226 ( .CLK(clk_bF_buf41), .D(_0H2_reg_31_0__1_), .Q(_auto_iopadmap_cc_368_execute_22625_65_), .R(reset_n_bF_buf41), .S(1'h1));
DFFSR DFFSR_227 ( .CLK(clk_bF_buf40), .D(_0H2_reg_31_0__2_), .Q(_auto_iopadmap_cc_368_execute_22625_66_), .R(reset_n_bF_buf40), .S(1'h1));
DFFSR DFFSR_228 ( .CLK(clk_bF_buf39), .D(_0H2_reg_31_0__3_), .Q(_auto_iopadmap_cc_368_execute_22625_67_), .R(reset_n_bF_buf39), .S(1'h1));
DFFSR DFFSR_229 ( .CLK(clk_bF_buf38), .D(_0H2_reg_31_0__4_), .Q(_auto_iopadmap_cc_368_execute_22625_68_), .R(reset_n_bF_buf38), .S(1'h1));
DFFSR DFFSR_23 ( .CLK(clk_bF_buf66), .D(_0a_reg_31_0__22_), .Q(a_reg_22_), .R(reset_n_bF_buf66), .S(1'h1));
DFFSR DFFSR_230 ( .CLK(clk_bF_buf37), .D(_0H2_reg_31_0__5_), .Q(_auto_iopadmap_cc_368_execute_22625_69_), .R(reset_n_bF_buf37), .S(1'h1));
DFFSR DFFSR_231 ( .CLK(clk_bF_buf36), .D(_0H2_reg_31_0__6_), .Q(_auto_iopadmap_cc_368_execute_22625_70_), .R(reset_n_bF_buf36), .S(1'h1));
DFFSR DFFSR_232 ( .CLK(clk_bF_buf35), .D(_0H2_reg_31_0__7_), .Q(_auto_iopadmap_cc_368_execute_22625_71_), .R(reset_n_bF_buf35), .S(1'h1));
DFFSR DFFSR_233 ( .CLK(clk_bF_buf34), .D(_0H2_reg_31_0__8_), .Q(_auto_iopadmap_cc_368_execute_22625_72_), .R(reset_n_bF_buf34), .S(1'h1));
DFFSR DFFSR_234 ( .CLK(clk_bF_buf33), .D(_0H2_reg_31_0__9_), .Q(_auto_iopadmap_cc_368_execute_22625_73_), .R(reset_n_bF_buf33), .S(1'h1));
DFFSR DFFSR_235 ( .CLK(clk_bF_buf32), .D(_0H2_reg_31_0__10_), .Q(_auto_iopadmap_cc_368_execute_22625_74_), .R(reset_n_bF_buf32), .S(1'h1));
DFFSR DFFSR_236 ( .CLK(clk_bF_buf31), .D(_0H2_reg_31_0__11_), .Q(_auto_iopadmap_cc_368_execute_22625_75_), .R(reset_n_bF_buf31), .S(1'h1));
DFFSR DFFSR_237 ( .CLK(clk_bF_buf30), .D(_0H2_reg_31_0__12_), .Q(_auto_iopadmap_cc_368_execute_22625_76_), .R(reset_n_bF_buf30), .S(1'h1));
DFFSR DFFSR_238 ( .CLK(clk_bF_buf29), .D(_0H2_reg_31_0__13_), .Q(_auto_iopadmap_cc_368_execute_22625_77_), .R(reset_n_bF_buf29), .S(1'h1));
DFFSR DFFSR_239 ( .CLK(clk_bF_buf28), .D(_0H2_reg_31_0__14_), .Q(_auto_iopadmap_cc_368_execute_22625_78_), .R(reset_n_bF_buf28), .S(1'h1));
DFFSR DFFSR_24 ( .CLK(clk_bF_buf65), .D(_0a_reg_31_0__23_), .Q(a_reg_23_), .R(reset_n_bF_buf65), .S(1'h1));
DFFSR DFFSR_240 ( .CLK(clk_bF_buf27), .D(_0H2_reg_31_0__15_), .Q(_auto_iopadmap_cc_368_execute_22625_79_), .R(reset_n_bF_buf27), .S(1'h1));
DFFSR DFFSR_241 ( .CLK(clk_bF_buf26), .D(_0H2_reg_31_0__16_), .Q(_auto_iopadmap_cc_368_execute_22625_80_), .R(reset_n_bF_buf26), .S(1'h1));
DFFSR DFFSR_242 ( .CLK(clk_bF_buf25), .D(_0H2_reg_31_0__17_), .Q(_auto_iopadmap_cc_368_execute_22625_81_), .R(reset_n_bF_buf25), .S(1'h1));
DFFSR DFFSR_243 ( .CLK(clk_bF_buf24), .D(_0H2_reg_31_0__18_), .Q(_auto_iopadmap_cc_368_execute_22625_82_), .R(reset_n_bF_buf24), .S(1'h1));
DFFSR DFFSR_244 ( .CLK(clk_bF_buf23), .D(_0H2_reg_31_0__19_), .Q(_auto_iopadmap_cc_368_execute_22625_83_), .R(reset_n_bF_buf23), .S(1'h1));
DFFSR DFFSR_245 ( .CLK(clk_bF_buf22), .D(_0H2_reg_31_0__20_), .Q(_auto_iopadmap_cc_368_execute_22625_84_), .R(reset_n_bF_buf22), .S(1'h1));
DFFSR DFFSR_246 ( .CLK(clk_bF_buf21), .D(_0H2_reg_31_0__21_), .Q(_auto_iopadmap_cc_368_execute_22625_85_), .R(reset_n_bF_buf21), .S(1'h1));
DFFSR DFFSR_247 ( .CLK(clk_bF_buf20), .D(_0H2_reg_31_0__22_), .Q(_auto_iopadmap_cc_368_execute_22625_86_), .R(reset_n_bF_buf20), .S(1'h1));
DFFSR DFFSR_248 ( .CLK(clk_bF_buf19), .D(_0H2_reg_31_0__23_), .Q(_auto_iopadmap_cc_368_execute_22625_87_), .R(reset_n_bF_buf19), .S(1'h1));
DFFSR DFFSR_249 ( .CLK(clk_bF_buf18), .D(_0H2_reg_31_0__24_), .Q(_auto_iopadmap_cc_368_execute_22625_88_), .R(reset_n_bF_buf18), .S(1'h1));
DFFSR DFFSR_25 ( .CLK(clk_bF_buf64), .D(_0a_reg_31_0__24_), .Q(a_reg_24_), .R(reset_n_bF_buf64), .S(1'h1));
DFFSR DFFSR_250 ( .CLK(clk_bF_buf17), .D(_0H2_reg_31_0__25_), .Q(_auto_iopadmap_cc_368_execute_22625_89_), .R(reset_n_bF_buf17), .S(1'h1));
DFFSR DFFSR_251 ( .CLK(clk_bF_buf16), .D(_0H2_reg_31_0__26_), .Q(_auto_iopadmap_cc_368_execute_22625_90_), .R(reset_n_bF_buf16), .S(1'h1));
DFFSR DFFSR_252 ( .CLK(clk_bF_buf15), .D(_0H2_reg_31_0__27_), .Q(_auto_iopadmap_cc_368_execute_22625_91_), .R(reset_n_bF_buf15), .S(1'h1));
DFFSR DFFSR_253 ( .CLK(clk_bF_buf14), .D(_0H2_reg_31_0__28_), .Q(_auto_iopadmap_cc_368_execute_22625_92_), .R(reset_n_bF_buf14), .S(1'h1));
DFFSR DFFSR_254 ( .CLK(clk_bF_buf13), .D(_0H2_reg_31_0__29_), .Q(_auto_iopadmap_cc_368_execute_22625_93_), .R(reset_n_bF_buf13), .S(1'h1));
DFFSR DFFSR_255 ( .CLK(clk_bF_buf12), .D(_0H2_reg_31_0__30_), .Q(_auto_iopadmap_cc_368_execute_22625_94_), .R(reset_n_bF_buf12), .S(1'h1));
DFFSR DFFSR_256 ( .CLK(clk_bF_buf11), .D(_0H2_reg_31_0__31_), .Q(_auto_iopadmap_cc_368_execute_22625_95_), .R(reset_n_bF_buf11), .S(1'h1));
DFFSR DFFSR_257 ( .CLK(clk_bF_buf10), .D(_0H3_reg_31_0__0_), .Q(_auto_iopadmap_cc_368_execute_22625_32_), .R(reset_n_bF_buf10), .S(1'h1));
DFFSR DFFSR_258 ( .CLK(clk_bF_buf9), .D(_0H3_reg_31_0__1_), .Q(_auto_iopadmap_cc_368_execute_22625_33_), .R(reset_n_bF_buf9), .S(1'h1));
DFFSR DFFSR_259 ( .CLK(clk_bF_buf8), .D(_0H3_reg_31_0__2_), .Q(_auto_iopadmap_cc_368_execute_22625_34_), .R(reset_n_bF_buf8), .S(1'h1));
DFFSR DFFSR_26 ( .CLK(clk_bF_buf63), .D(_0a_reg_31_0__25_), .Q(a_reg_25_), .R(reset_n_bF_buf63), .S(1'h1));
DFFSR DFFSR_260 ( .CLK(clk_bF_buf7), .D(_0H3_reg_31_0__3_), .Q(_auto_iopadmap_cc_368_execute_22625_35_), .R(reset_n_bF_buf7), .S(1'h1));
DFFSR DFFSR_261 ( .CLK(clk_bF_buf6), .D(_0H3_reg_31_0__4_), .Q(_auto_iopadmap_cc_368_execute_22625_36_), .R(reset_n_bF_buf6), .S(1'h1));
DFFSR DFFSR_262 ( .CLK(clk_bF_buf5), .D(_0H3_reg_31_0__5_), .Q(_auto_iopadmap_cc_368_execute_22625_37_), .R(reset_n_bF_buf5), .S(1'h1));
DFFSR DFFSR_263 ( .CLK(clk_bF_buf4), .D(_0H3_reg_31_0__6_), .Q(_auto_iopadmap_cc_368_execute_22625_38_), .R(reset_n_bF_buf4), .S(1'h1));
DFFSR DFFSR_264 ( .CLK(clk_bF_buf3), .D(_0H3_reg_31_0__7_), .Q(_auto_iopadmap_cc_368_execute_22625_39_), .R(reset_n_bF_buf3), .S(1'h1));
DFFSR DFFSR_265 ( .CLK(clk_bF_buf2), .D(_0H3_reg_31_0__8_), .Q(_auto_iopadmap_cc_368_execute_22625_40_), .R(reset_n_bF_buf2), .S(1'h1));
DFFSR DFFSR_266 ( .CLK(clk_bF_buf1), .D(_0H3_reg_31_0__9_), .Q(_auto_iopadmap_cc_368_execute_22625_41_), .R(reset_n_bF_buf1), .S(1'h1));
DFFSR DFFSR_267 ( .CLK(clk_bF_buf0), .D(_0H3_reg_31_0__10_), .Q(_auto_iopadmap_cc_368_execute_22625_42_), .R(reset_n_bF_buf0), .S(1'h1));
DFFSR DFFSR_268 ( .CLK(clk_bF_buf88), .D(_0H3_reg_31_0__11_), .Q(_auto_iopadmap_cc_368_execute_22625_43_), .R(reset_n_bF_buf88), .S(1'h1));
DFFSR DFFSR_269 ( .CLK(clk_bF_buf87), .D(_0H3_reg_31_0__12_), .Q(_auto_iopadmap_cc_368_execute_22625_44_), .R(reset_n_bF_buf87), .S(1'h1));
DFFSR DFFSR_27 ( .CLK(clk_bF_buf62), .D(_0a_reg_31_0__26_), .Q(a_reg_26_), .R(reset_n_bF_buf62), .S(1'h1));
DFFSR DFFSR_270 ( .CLK(clk_bF_buf86), .D(_0H3_reg_31_0__13_), .Q(_auto_iopadmap_cc_368_execute_22625_45_), .R(reset_n_bF_buf86), .S(1'h1));
DFFSR DFFSR_271 ( .CLK(clk_bF_buf85), .D(_0H3_reg_31_0__14_), .Q(_auto_iopadmap_cc_368_execute_22625_46_), .R(reset_n_bF_buf85), .S(1'h1));
DFFSR DFFSR_272 ( .CLK(clk_bF_buf84), .D(_0H3_reg_31_0__15_), .Q(_auto_iopadmap_cc_368_execute_22625_47_), .R(reset_n_bF_buf84), .S(1'h1));
DFFSR DFFSR_273 ( .CLK(clk_bF_buf83), .D(_0H3_reg_31_0__16_), .Q(_auto_iopadmap_cc_368_execute_22625_48_), .R(reset_n_bF_buf83), .S(1'h1));
DFFSR DFFSR_274 ( .CLK(clk_bF_buf82), .D(_0H3_reg_31_0__17_), .Q(_auto_iopadmap_cc_368_execute_22625_49_), .R(reset_n_bF_buf82), .S(1'h1));
DFFSR DFFSR_275 ( .CLK(clk_bF_buf81), .D(_0H3_reg_31_0__18_), .Q(_auto_iopadmap_cc_368_execute_22625_50_), .R(reset_n_bF_buf81), .S(1'h1));
DFFSR DFFSR_276 ( .CLK(clk_bF_buf80), .D(_0H3_reg_31_0__19_), .Q(_auto_iopadmap_cc_368_execute_22625_51_), .R(reset_n_bF_buf80), .S(1'h1));
DFFSR DFFSR_277 ( .CLK(clk_bF_buf79), .D(_0H3_reg_31_0__20_), .Q(_auto_iopadmap_cc_368_execute_22625_52_), .R(reset_n_bF_buf79), .S(1'h1));
DFFSR DFFSR_278 ( .CLK(clk_bF_buf78), .D(_0H3_reg_31_0__21_), .Q(_auto_iopadmap_cc_368_execute_22625_53_), .R(reset_n_bF_buf78), .S(1'h1));
DFFSR DFFSR_279 ( .CLK(clk_bF_buf77), .D(_0H3_reg_31_0__22_), .Q(_auto_iopadmap_cc_368_execute_22625_54_), .R(reset_n_bF_buf77), .S(1'h1));
DFFSR DFFSR_28 ( .CLK(clk_bF_buf61), .D(_0a_reg_31_0__27_), .Q(a_reg_27_), .R(reset_n_bF_buf61), .S(1'h1));
DFFSR DFFSR_280 ( .CLK(clk_bF_buf76), .D(_0H3_reg_31_0__23_), .Q(_auto_iopadmap_cc_368_execute_22625_55_), .R(reset_n_bF_buf76), .S(1'h1));
DFFSR DFFSR_281 ( .CLK(clk_bF_buf75), .D(_0H3_reg_31_0__24_), .Q(_auto_iopadmap_cc_368_execute_22625_56_), .R(reset_n_bF_buf75), .S(1'h1));
DFFSR DFFSR_282 ( .CLK(clk_bF_buf74), .D(_0H3_reg_31_0__25_), .Q(_auto_iopadmap_cc_368_execute_22625_57_), .R(reset_n_bF_buf74), .S(1'h1));
DFFSR DFFSR_283 ( .CLK(clk_bF_buf73), .D(_0H3_reg_31_0__26_), .Q(_auto_iopadmap_cc_368_execute_22625_58_), .R(reset_n_bF_buf73), .S(1'h1));
DFFSR DFFSR_284 ( .CLK(clk_bF_buf72), .D(_0H3_reg_31_0__27_), .Q(_auto_iopadmap_cc_368_execute_22625_59_), .R(reset_n_bF_buf72), .S(1'h1));
DFFSR DFFSR_285 ( .CLK(clk_bF_buf71), .D(_0H3_reg_31_0__28_), .Q(_auto_iopadmap_cc_368_execute_22625_60_), .R(reset_n_bF_buf71), .S(1'h1));
DFFSR DFFSR_286 ( .CLK(clk_bF_buf70), .D(_0H3_reg_31_0__29_), .Q(_auto_iopadmap_cc_368_execute_22625_61_), .R(reset_n_bF_buf70), .S(1'h1));
DFFSR DFFSR_287 ( .CLK(clk_bF_buf69), .D(_0H3_reg_31_0__30_), .Q(_auto_iopadmap_cc_368_execute_22625_62_), .R(reset_n_bF_buf69), .S(1'h1));
DFFSR DFFSR_288 ( .CLK(clk_bF_buf68), .D(_0H3_reg_31_0__31_), .Q(_auto_iopadmap_cc_368_execute_22625_63_), .R(reset_n_bF_buf68), .S(1'h1));
DFFSR DFFSR_289 ( .CLK(clk_bF_buf67), .D(_0H4_reg_31_0__0_), .Q(_auto_iopadmap_cc_368_execute_22625_0_), .R(reset_n_bF_buf67), .S(1'h1));
DFFSR DFFSR_29 ( .CLK(clk_bF_buf60), .D(_0a_reg_31_0__28_), .Q(a_reg_28_), .R(reset_n_bF_buf60), .S(1'h1));
DFFSR DFFSR_290 ( .CLK(clk_bF_buf66), .D(_0H4_reg_31_0__1_), .Q(_auto_iopadmap_cc_368_execute_22625_1_), .R(reset_n_bF_buf66), .S(1'h1));
DFFSR DFFSR_291 ( .CLK(clk_bF_buf65), .D(_0H4_reg_31_0__2_), .Q(_auto_iopadmap_cc_368_execute_22625_2_), .R(reset_n_bF_buf65), .S(1'h1));
DFFSR DFFSR_292 ( .CLK(clk_bF_buf64), .D(_0H4_reg_31_0__3_), .Q(_auto_iopadmap_cc_368_execute_22625_3_), .R(reset_n_bF_buf64), .S(1'h1));
DFFSR DFFSR_293 ( .CLK(clk_bF_buf63), .D(_0H4_reg_31_0__4_), .Q(_auto_iopadmap_cc_368_execute_22625_4_), .R(reset_n_bF_buf63), .S(1'h1));
DFFSR DFFSR_294 ( .CLK(clk_bF_buf62), .D(_0H4_reg_31_0__5_), .Q(_auto_iopadmap_cc_368_execute_22625_5_), .R(reset_n_bF_buf62), .S(1'h1));
DFFSR DFFSR_295 ( .CLK(clk_bF_buf61), .D(_0H4_reg_31_0__6_), .Q(_auto_iopadmap_cc_368_execute_22625_6_), .R(reset_n_bF_buf61), .S(1'h1));
DFFSR DFFSR_296 ( .CLK(clk_bF_buf60), .D(_0H4_reg_31_0__7_), .Q(_auto_iopadmap_cc_368_execute_22625_7_), .R(reset_n_bF_buf60), .S(1'h1));
DFFSR DFFSR_297 ( .CLK(clk_bF_buf59), .D(_0H4_reg_31_0__8_), .Q(_auto_iopadmap_cc_368_execute_22625_8_), .R(reset_n_bF_buf59), .S(1'h1));
DFFSR DFFSR_298 ( .CLK(clk_bF_buf58), .D(_0H4_reg_31_0__9_), .Q(_auto_iopadmap_cc_368_execute_22625_9_), .R(reset_n_bF_buf58), .S(1'h1));
DFFSR DFFSR_299 ( .CLK(clk_bF_buf57), .D(_0H4_reg_31_0__10_), .Q(_auto_iopadmap_cc_368_execute_22625_10_), .R(reset_n_bF_buf57), .S(1'h1));
DFFSR DFFSR_3 ( .CLK(clk_bF_buf86), .D(_0a_reg_31_0__2_), .Q(a_reg_2_), .R(reset_n_bF_buf86), .S(1'h1));
DFFSR DFFSR_30 ( .CLK(clk_bF_buf59), .D(_0a_reg_31_0__29_), .Q(a_reg_29_), .R(reset_n_bF_buf59), .S(1'h1));
DFFSR DFFSR_300 ( .CLK(clk_bF_buf56), .D(_0H4_reg_31_0__11_), .Q(_auto_iopadmap_cc_368_execute_22625_11_), .R(reset_n_bF_buf56), .S(1'h1));
DFFSR DFFSR_301 ( .CLK(clk_bF_buf55), .D(_0H4_reg_31_0__12_), .Q(_auto_iopadmap_cc_368_execute_22625_12_), .R(reset_n_bF_buf55), .S(1'h1));
DFFSR DFFSR_302 ( .CLK(clk_bF_buf54), .D(_0H4_reg_31_0__13_), .Q(_auto_iopadmap_cc_368_execute_22625_13_), .R(reset_n_bF_buf54), .S(1'h1));
DFFSR DFFSR_303 ( .CLK(clk_bF_buf53), .D(_0H4_reg_31_0__14_), .Q(_auto_iopadmap_cc_368_execute_22625_14_), .R(reset_n_bF_buf53), .S(1'h1));
DFFSR DFFSR_304 ( .CLK(clk_bF_buf52), .D(_0H4_reg_31_0__15_), .Q(_auto_iopadmap_cc_368_execute_22625_15_), .R(reset_n_bF_buf52), .S(1'h1));
DFFSR DFFSR_305 ( .CLK(clk_bF_buf51), .D(_0H4_reg_31_0__16_), .Q(_auto_iopadmap_cc_368_execute_22625_16_), .R(reset_n_bF_buf51), .S(1'h1));
DFFSR DFFSR_306 ( .CLK(clk_bF_buf50), .D(_0H4_reg_31_0__17_), .Q(_auto_iopadmap_cc_368_execute_22625_17_), .R(reset_n_bF_buf50), .S(1'h1));
DFFSR DFFSR_307 ( .CLK(clk_bF_buf49), .D(_0H4_reg_31_0__18_), .Q(_auto_iopadmap_cc_368_execute_22625_18_), .R(reset_n_bF_buf49), .S(1'h1));
DFFSR DFFSR_308 ( .CLK(clk_bF_buf48), .D(_0H4_reg_31_0__19_), .Q(_auto_iopadmap_cc_368_execute_22625_19_), .R(reset_n_bF_buf48), .S(1'h1));
DFFSR DFFSR_309 ( .CLK(clk_bF_buf47), .D(_0H4_reg_31_0__20_), .Q(_auto_iopadmap_cc_368_execute_22625_20_), .R(reset_n_bF_buf47), .S(1'h1));
DFFSR DFFSR_31 ( .CLK(clk_bF_buf58), .D(_0a_reg_31_0__30_), .Q(a_reg_30_), .R(reset_n_bF_buf58), .S(1'h1));
DFFSR DFFSR_310 ( .CLK(clk_bF_buf46), .D(_0H4_reg_31_0__21_), .Q(_auto_iopadmap_cc_368_execute_22625_21_), .R(reset_n_bF_buf46), .S(1'h1));
DFFSR DFFSR_311 ( .CLK(clk_bF_buf45), .D(_0H4_reg_31_0__22_), .Q(_auto_iopadmap_cc_368_execute_22625_22_), .R(reset_n_bF_buf45), .S(1'h1));
DFFSR DFFSR_312 ( .CLK(clk_bF_buf44), .D(_0H4_reg_31_0__23_), .Q(_auto_iopadmap_cc_368_execute_22625_23_), .R(reset_n_bF_buf44), .S(1'h1));
DFFSR DFFSR_313 ( .CLK(clk_bF_buf43), .D(_0H4_reg_31_0__24_), .Q(_auto_iopadmap_cc_368_execute_22625_24_), .R(reset_n_bF_buf43), .S(1'h1));
DFFSR DFFSR_314 ( .CLK(clk_bF_buf42), .D(_0H4_reg_31_0__25_), .Q(_auto_iopadmap_cc_368_execute_22625_25_), .R(reset_n_bF_buf42), .S(1'h1));
DFFSR DFFSR_315 ( .CLK(clk_bF_buf41), .D(_0H4_reg_31_0__26_), .Q(_auto_iopadmap_cc_368_execute_22625_26_), .R(reset_n_bF_buf41), .S(1'h1));
DFFSR DFFSR_316 ( .CLK(clk_bF_buf40), .D(_0H4_reg_31_0__27_), .Q(_auto_iopadmap_cc_368_execute_22625_27_), .R(reset_n_bF_buf40), .S(1'h1));
DFFSR DFFSR_317 ( .CLK(clk_bF_buf39), .D(_0H4_reg_31_0__28_), .Q(_auto_iopadmap_cc_368_execute_22625_28_), .R(reset_n_bF_buf39), .S(1'h1));
DFFSR DFFSR_318 ( .CLK(clk_bF_buf38), .D(_0H4_reg_31_0__29_), .Q(_auto_iopadmap_cc_368_execute_22625_29_), .R(reset_n_bF_buf38), .S(1'h1));
DFFSR DFFSR_319 ( .CLK(clk_bF_buf37), .D(_0H4_reg_31_0__30_), .Q(_auto_iopadmap_cc_368_execute_22625_30_), .R(reset_n_bF_buf37), .S(1'h1));
DFFSR DFFSR_32 ( .CLK(clk_bF_buf57), .D(_0a_reg_31_0__31_), .Q(a_reg_31_), .R(reset_n_bF_buf57), .S(1'h1));
DFFSR DFFSR_320 ( .CLK(clk_bF_buf36), .D(_0H4_reg_31_0__31_), .Q(_auto_iopadmap_cc_368_execute_22625_31_), .R(reset_n_bF_buf36), .S(1'h1));
DFFSR DFFSR_321 ( .CLK(clk_bF_buf35), .D(_0round_ctr_reg_6_0__0_), .Q(round_ctr_reg_0_), .R(reset_n_bF_buf35), .S(1'h1));
DFFSR DFFSR_322 ( .CLK(clk_bF_buf34), .D(_0round_ctr_reg_6_0__1_), .Q(round_ctr_reg_1_), .R(reset_n_bF_buf34), .S(1'h1));
DFFSR DFFSR_323 ( .CLK(clk_bF_buf33), .D(_0round_ctr_reg_6_0__2_), .Q(round_ctr_reg_2_), .R(reset_n_bF_buf33), .S(1'h1));
DFFSR DFFSR_324 ( .CLK(clk_bF_buf32), .D(_0round_ctr_reg_6_0__3_), .Q(round_ctr_reg_3_), .R(reset_n_bF_buf32), .S(1'h1));
DFFSR DFFSR_325 ( .CLK(clk_bF_buf31), .D(_0round_ctr_reg_6_0__4_), .Q(round_ctr_reg_4_), .R(reset_n_bF_buf31), .S(1'h1));
DFFSR DFFSR_326 ( .CLK(clk_bF_buf30), .D(_0round_ctr_reg_6_0__5_), .Q(round_ctr_reg_5_), .R(reset_n_bF_buf30), .S(1'h1));
DFFSR DFFSR_327 ( .CLK(clk_bF_buf29), .D(_0round_ctr_reg_6_0__6_), .Q(round_ctr_reg_6_), .R(reset_n_bF_buf29), .S(1'h1));
DFFSR DFFSR_328 ( .CLK(clk_bF_buf28), .D(_0digest_valid_reg_0_0_), .Q(_auto_iopadmap_cc_368_execute_22786), .R(reset_n_bF_buf28), .S(1'h1));
DFFSR DFFSR_329 ( .CLK(clk_bF_buf27), .D(_abc_15497_abc_9717_auto_fsm_map_cc_170_map_fsm_844_0_), .Q(_auto_iopadmap_cc_368_execute_22788), .R(1'h1), .S(reset_n_bF_buf27));
DFFSR DFFSR_33 ( .CLK(clk_bF_buf56), .D(_0b_reg_31_0__0_), .Q(b_reg_0_), .R(reset_n_bF_buf56), .S(1'h1));
DFFSR DFFSR_330 ( .CLK(clk_bF_buf26), .D(_abc_15497_abc_9717_auto_fsm_map_cc_118_implement_pattern_cache_863), .Q(digest_update), .R(reset_n_bF_buf26), .S(1'h1));
DFFSR DFFSR_331 ( .CLK(clk_bF_buf25), .D(_abc_15497_abc_9717_auto_fsm_map_cc_170_map_fsm_844_2_), .Q(round_ctr_inc), .R(reset_n_bF_buf25), .S(1'h1));
DFFSR DFFSR_332 ( .CLK(clk_bF_buf24), .D(w_mem_inst__0w_ctr_reg_6_0__0_), .Q(w_mem_inst_w_ctr_reg_0_), .R(reset_n_bF_buf24), .S(1'h1));
DFFSR DFFSR_333 ( .CLK(clk_bF_buf23), .D(w_mem_inst__0w_ctr_reg_6_0__1_), .Q(w_mem_inst_w_ctr_reg_1_), .R(reset_n_bF_buf23), .S(1'h1));
DFFSR DFFSR_334 ( .CLK(clk_bF_buf22), .D(w_mem_inst__0w_ctr_reg_6_0__2_), .Q(w_mem_inst_w_ctr_reg_2_), .R(reset_n_bF_buf22), .S(1'h1));
DFFSR DFFSR_335 ( .CLK(clk_bF_buf21), .D(w_mem_inst__0w_ctr_reg_6_0__3_), .Q(w_mem_inst_w_ctr_reg_3_), .R(reset_n_bF_buf21), .S(1'h1));
DFFSR DFFSR_336 ( .CLK(clk_bF_buf20), .D(w_mem_inst__0w_ctr_reg_6_0__4_), .Q(w_mem_inst_w_ctr_reg_4_), .R(reset_n_bF_buf20), .S(1'h1));
DFFSR DFFSR_337 ( .CLK(clk_bF_buf19), .D(w_mem_inst__0w_ctr_reg_6_0__5_), .Q(w_mem_inst_w_ctr_reg_5_), .R(reset_n_bF_buf19), .S(1'h1));
DFFSR DFFSR_338 ( .CLK(clk_bF_buf18), .D(w_mem_inst__0w_ctr_reg_6_0__6_), .Q(w_mem_inst_w_ctr_reg_6_), .R(reset_n_bF_buf18), .S(1'h1));
DFFSR DFFSR_339 ( .CLK(clk_bF_buf17), .D(w_mem_inst__0w_mem_0__31_0__0_), .Q(w_mem_inst_w_mem_0__0_), .R(reset_n_bF_buf17), .S(1'h1));
DFFSR DFFSR_34 ( .CLK(clk_bF_buf55), .D(_0b_reg_31_0__1_), .Q(b_reg_1_), .R(reset_n_bF_buf55), .S(1'h1));
DFFSR DFFSR_340 ( .CLK(clk_bF_buf16), .D(w_mem_inst__0w_mem_0__31_0__1_), .Q(w_mem_inst_w_mem_0__1_), .R(reset_n_bF_buf16), .S(1'h1));
DFFSR DFFSR_341 ( .CLK(clk_bF_buf15), .D(w_mem_inst__0w_mem_0__31_0__2_), .Q(w_mem_inst_w_mem_0__2_), .R(reset_n_bF_buf15), .S(1'h1));
DFFSR DFFSR_342 ( .CLK(clk_bF_buf14), .D(w_mem_inst__0w_mem_0__31_0__3_), .Q(w_mem_inst_w_mem_0__3_), .R(reset_n_bF_buf14), .S(1'h1));
DFFSR DFFSR_343 ( .CLK(clk_bF_buf13), .D(w_mem_inst__0w_mem_0__31_0__4_), .Q(w_mem_inst_w_mem_0__4_), .R(reset_n_bF_buf13), .S(1'h1));
DFFSR DFFSR_344 ( .CLK(clk_bF_buf12), .D(w_mem_inst__0w_mem_0__31_0__5_), .Q(w_mem_inst_w_mem_0__5_), .R(reset_n_bF_buf12), .S(1'h1));
DFFSR DFFSR_345 ( .CLK(clk_bF_buf11), .D(w_mem_inst__0w_mem_0__31_0__6_), .Q(w_mem_inst_w_mem_0__6_), .R(reset_n_bF_buf11), .S(1'h1));
DFFSR DFFSR_346 ( .CLK(clk_bF_buf10), .D(w_mem_inst__0w_mem_0__31_0__7_), .Q(w_mem_inst_w_mem_0__7_), .R(reset_n_bF_buf10), .S(1'h1));
DFFSR DFFSR_347 ( .CLK(clk_bF_buf9), .D(w_mem_inst__0w_mem_0__31_0__8_), .Q(w_mem_inst_w_mem_0__8_), .R(reset_n_bF_buf9), .S(1'h1));
DFFSR DFFSR_348 ( .CLK(clk_bF_buf8), .D(w_mem_inst__0w_mem_0__31_0__9_), .Q(w_mem_inst_w_mem_0__9_), .R(reset_n_bF_buf8), .S(1'h1));
DFFSR DFFSR_349 ( .CLK(clk_bF_buf7), .D(w_mem_inst__0w_mem_0__31_0__10_), .Q(w_mem_inst_w_mem_0__10_), .R(reset_n_bF_buf7), .S(1'h1));
DFFSR DFFSR_35 ( .CLK(clk_bF_buf54), .D(_0b_reg_31_0__2_), .Q(b_reg_2_), .R(reset_n_bF_buf54), .S(1'h1));
DFFSR DFFSR_350 ( .CLK(clk_bF_buf6), .D(w_mem_inst__0w_mem_0__31_0__11_), .Q(w_mem_inst_w_mem_0__11_), .R(reset_n_bF_buf6), .S(1'h1));
DFFSR DFFSR_351 ( .CLK(clk_bF_buf5), .D(w_mem_inst__0w_mem_0__31_0__12_), .Q(w_mem_inst_w_mem_0__12_), .R(reset_n_bF_buf5), .S(1'h1));
DFFSR DFFSR_352 ( .CLK(clk_bF_buf4), .D(w_mem_inst__0w_mem_0__31_0__13_), .Q(w_mem_inst_w_mem_0__13_), .R(reset_n_bF_buf4), .S(1'h1));
DFFSR DFFSR_353 ( .CLK(clk_bF_buf3), .D(w_mem_inst__0w_mem_0__31_0__14_), .Q(w_mem_inst_w_mem_0__14_), .R(reset_n_bF_buf3), .S(1'h1));
DFFSR DFFSR_354 ( .CLK(clk_bF_buf2), .D(w_mem_inst__0w_mem_0__31_0__15_), .Q(w_mem_inst_w_mem_0__15_), .R(reset_n_bF_buf2), .S(1'h1));
DFFSR DFFSR_355 ( .CLK(clk_bF_buf1), .D(w_mem_inst__0w_mem_0__31_0__16_), .Q(w_mem_inst_w_mem_0__16_), .R(reset_n_bF_buf1), .S(1'h1));
DFFSR DFFSR_356 ( .CLK(clk_bF_buf0), .D(w_mem_inst__0w_mem_0__31_0__17_), .Q(w_mem_inst_w_mem_0__17_), .R(reset_n_bF_buf0), .S(1'h1));
DFFSR DFFSR_357 ( .CLK(clk_bF_buf88), .D(w_mem_inst__0w_mem_0__31_0__18_), .Q(w_mem_inst_w_mem_0__18_), .R(reset_n_bF_buf88), .S(1'h1));
DFFSR DFFSR_358 ( .CLK(clk_bF_buf87), .D(w_mem_inst__0w_mem_0__31_0__19_), .Q(w_mem_inst_w_mem_0__19_), .R(reset_n_bF_buf87), .S(1'h1));
DFFSR DFFSR_359 ( .CLK(clk_bF_buf86), .D(w_mem_inst__0w_mem_0__31_0__20_), .Q(w_mem_inst_w_mem_0__20_), .R(reset_n_bF_buf86), .S(1'h1));
DFFSR DFFSR_36 ( .CLK(clk_bF_buf53), .D(_0b_reg_31_0__3_), .Q(b_reg_3_), .R(reset_n_bF_buf53), .S(1'h1));
DFFSR DFFSR_360 ( .CLK(clk_bF_buf85), .D(w_mem_inst__0w_mem_0__31_0__21_), .Q(w_mem_inst_w_mem_0__21_), .R(reset_n_bF_buf85), .S(1'h1));
DFFSR DFFSR_361 ( .CLK(clk_bF_buf84), .D(w_mem_inst__0w_mem_0__31_0__22_), .Q(w_mem_inst_w_mem_0__22_), .R(reset_n_bF_buf84), .S(1'h1));
DFFSR DFFSR_362 ( .CLK(clk_bF_buf83), .D(w_mem_inst__0w_mem_0__31_0__23_), .Q(w_mem_inst_w_mem_0__23_), .R(reset_n_bF_buf83), .S(1'h1));
DFFSR DFFSR_363 ( .CLK(clk_bF_buf82), .D(w_mem_inst__0w_mem_0__31_0__24_), .Q(w_mem_inst_w_mem_0__24_), .R(reset_n_bF_buf82), .S(1'h1));
DFFSR DFFSR_364 ( .CLK(clk_bF_buf81), .D(w_mem_inst__0w_mem_0__31_0__25_), .Q(w_mem_inst_w_mem_0__25_), .R(reset_n_bF_buf81), .S(1'h1));
DFFSR DFFSR_365 ( .CLK(clk_bF_buf80), .D(w_mem_inst__0w_mem_0__31_0__26_), .Q(w_mem_inst_w_mem_0__26_), .R(reset_n_bF_buf80), .S(1'h1));
DFFSR DFFSR_366 ( .CLK(clk_bF_buf79), .D(w_mem_inst__0w_mem_0__31_0__27_), .Q(w_mem_inst_w_mem_0__27_), .R(reset_n_bF_buf79), .S(1'h1));
DFFSR DFFSR_367 ( .CLK(clk_bF_buf78), .D(w_mem_inst__0w_mem_0__31_0__28_), .Q(w_mem_inst_w_mem_0__28_), .R(reset_n_bF_buf78), .S(1'h1));
DFFSR DFFSR_368 ( .CLK(clk_bF_buf77), .D(w_mem_inst__0w_mem_0__31_0__29_), .Q(w_mem_inst_w_mem_0__29_), .R(reset_n_bF_buf77), .S(1'h1));
DFFSR DFFSR_369 ( .CLK(clk_bF_buf76), .D(w_mem_inst__0w_mem_0__31_0__30_), .Q(w_mem_inst_w_mem_0__30_), .R(reset_n_bF_buf76), .S(1'h1));
DFFSR DFFSR_37 ( .CLK(clk_bF_buf52), .D(_0b_reg_31_0__4_), .Q(b_reg_4_), .R(reset_n_bF_buf52), .S(1'h1));
DFFSR DFFSR_370 ( .CLK(clk_bF_buf75), .D(w_mem_inst__0w_mem_0__31_0__31_), .Q(w_mem_inst_w_mem_0__31_), .R(reset_n_bF_buf75), .S(1'h1));
DFFSR DFFSR_371 ( .CLK(clk_bF_buf74), .D(w_mem_inst__0w_mem_1__31_0__0_), .Q(w_mem_inst_w_mem_1__0_), .R(reset_n_bF_buf74), .S(1'h1));
DFFSR DFFSR_372 ( .CLK(clk_bF_buf73), .D(w_mem_inst__0w_mem_1__31_0__1_), .Q(w_mem_inst_w_mem_1__1_), .R(reset_n_bF_buf73), .S(1'h1));
DFFSR DFFSR_373 ( .CLK(clk_bF_buf72), .D(w_mem_inst__0w_mem_1__31_0__2_), .Q(w_mem_inst_w_mem_1__2_), .R(reset_n_bF_buf72), .S(1'h1));
DFFSR DFFSR_374 ( .CLK(clk_bF_buf71), .D(w_mem_inst__0w_mem_1__31_0__3_), .Q(w_mem_inst_w_mem_1__3_), .R(reset_n_bF_buf71), .S(1'h1));
DFFSR DFFSR_375 ( .CLK(clk_bF_buf70), .D(w_mem_inst__0w_mem_1__31_0__4_), .Q(w_mem_inst_w_mem_1__4_), .R(reset_n_bF_buf70), .S(1'h1));
DFFSR DFFSR_376 ( .CLK(clk_bF_buf69), .D(w_mem_inst__0w_mem_1__31_0__5_), .Q(w_mem_inst_w_mem_1__5_), .R(reset_n_bF_buf69), .S(1'h1));
DFFSR DFFSR_377 ( .CLK(clk_bF_buf68), .D(w_mem_inst__0w_mem_1__31_0__6_), .Q(w_mem_inst_w_mem_1__6_), .R(reset_n_bF_buf68), .S(1'h1));
DFFSR DFFSR_378 ( .CLK(clk_bF_buf67), .D(w_mem_inst__0w_mem_1__31_0__7_), .Q(w_mem_inst_w_mem_1__7_), .R(reset_n_bF_buf67), .S(1'h1));
DFFSR DFFSR_379 ( .CLK(clk_bF_buf66), .D(w_mem_inst__0w_mem_1__31_0__8_), .Q(w_mem_inst_w_mem_1__8_), .R(reset_n_bF_buf66), .S(1'h1));
DFFSR DFFSR_38 ( .CLK(clk_bF_buf51), .D(_0b_reg_31_0__5_), .Q(b_reg_5_), .R(reset_n_bF_buf51), .S(1'h1));
DFFSR DFFSR_380 ( .CLK(clk_bF_buf65), .D(w_mem_inst__0w_mem_1__31_0__9_), .Q(w_mem_inst_w_mem_1__9_), .R(reset_n_bF_buf65), .S(1'h1));
DFFSR DFFSR_381 ( .CLK(clk_bF_buf64), .D(w_mem_inst__0w_mem_1__31_0__10_), .Q(w_mem_inst_w_mem_1__10_), .R(reset_n_bF_buf64), .S(1'h1));
DFFSR DFFSR_382 ( .CLK(clk_bF_buf63), .D(w_mem_inst__0w_mem_1__31_0__11_), .Q(w_mem_inst_w_mem_1__11_), .R(reset_n_bF_buf63), .S(1'h1));
DFFSR DFFSR_383 ( .CLK(clk_bF_buf62), .D(w_mem_inst__0w_mem_1__31_0__12_), .Q(w_mem_inst_w_mem_1__12_), .R(reset_n_bF_buf62), .S(1'h1));
DFFSR DFFSR_384 ( .CLK(clk_bF_buf61), .D(w_mem_inst__0w_mem_1__31_0__13_), .Q(w_mem_inst_w_mem_1__13_), .R(reset_n_bF_buf61), .S(1'h1));
DFFSR DFFSR_385 ( .CLK(clk_bF_buf60), .D(w_mem_inst__0w_mem_1__31_0__14_), .Q(w_mem_inst_w_mem_1__14_), .R(reset_n_bF_buf60), .S(1'h1));
DFFSR DFFSR_386 ( .CLK(clk_bF_buf59), .D(w_mem_inst__0w_mem_1__31_0__15_), .Q(w_mem_inst_w_mem_1__15_), .R(reset_n_bF_buf59), .S(1'h1));
DFFSR DFFSR_387 ( .CLK(clk_bF_buf58), .D(w_mem_inst__0w_mem_1__31_0__16_), .Q(w_mem_inst_w_mem_1__16_), .R(reset_n_bF_buf58), .S(1'h1));
DFFSR DFFSR_388 ( .CLK(clk_bF_buf57), .D(w_mem_inst__0w_mem_1__31_0__17_), .Q(w_mem_inst_w_mem_1__17_), .R(reset_n_bF_buf57), .S(1'h1));
DFFSR DFFSR_389 ( .CLK(clk_bF_buf56), .D(w_mem_inst__0w_mem_1__31_0__18_), .Q(w_mem_inst_w_mem_1__18_), .R(reset_n_bF_buf56), .S(1'h1));
DFFSR DFFSR_39 ( .CLK(clk_bF_buf50), .D(_0b_reg_31_0__6_), .Q(b_reg_6_), .R(reset_n_bF_buf50), .S(1'h1));
DFFSR DFFSR_390 ( .CLK(clk_bF_buf55), .D(w_mem_inst__0w_mem_1__31_0__19_), .Q(w_mem_inst_w_mem_1__19_), .R(reset_n_bF_buf55), .S(1'h1));
DFFSR DFFSR_391 ( .CLK(clk_bF_buf54), .D(w_mem_inst__0w_mem_1__31_0__20_), .Q(w_mem_inst_w_mem_1__20_), .R(reset_n_bF_buf54), .S(1'h1));
DFFSR DFFSR_392 ( .CLK(clk_bF_buf53), .D(w_mem_inst__0w_mem_1__31_0__21_), .Q(w_mem_inst_w_mem_1__21_), .R(reset_n_bF_buf53), .S(1'h1));
DFFSR DFFSR_393 ( .CLK(clk_bF_buf52), .D(w_mem_inst__0w_mem_1__31_0__22_), .Q(w_mem_inst_w_mem_1__22_), .R(reset_n_bF_buf52), .S(1'h1));
DFFSR DFFSR_394 ( .CLK(clk_bF_buf51), .D(w_mem_inst__0w_mem_1__31_0__23_), .Q(w_mem_inst_w_mem_1__23_), .R(reset_n_bF_buf51), .S(1'h1));
DFFSR DFFSR_395 ( .CLK(clk_bF_buf50), .D(w_mem_inst__0w_mem_1__31_0__24_), .Q(w_mem_inst_w_mem_1__24_), .R(reset_n_bF_buf50), .S(1'h1));
DFFSR DFFSR_396 ( .CLK(clk_bF_buf49), .D(w_mem_inst__0w_mem_1__31_0__25_), .Q(w_mem_inst_w_mem_1__25_), .R(reset_n_bF_buf49), .S(1'h1));
DFFSR DFFSR_397 ( .CLK(clk_bF_buf48), .D(w_mem_inst__0w_mem_1__31_0__26_), .Q(w_mem_inst_w_mem_1__26_), .R(reset_n_bF_buf48), .S(1'h1));
DFFSR DFFSR_398 ( .CLK(clk_bF_buf47), .D(w_mem_inst__0w_mem_1__31_0__27_), .Q(w_mem_inst_w_mem_1__27_), .R(reset_n_bF_buf47), .S(1'h1));
DFFSR DFFSR_399 ( .CLK(clk_bF_buf46), .D(w_mem_inst__0w_mem_1__31_0__28_), .Q(w_mem_inst_w_mem_1__28_), .R(reset_n_bF_buf46), .S(1'h1));
DFFSR DFFSR_4 ( .CLK(clk_bF_buf85), .D(_0a_reg_31_0__3_), .Q(a_reg_3_), .R(reset_n_bF_buf85), .S(1'h1));
DFFSR DFFSR_40 ( .CLK(clk_bF_buf49), .D(_0b_reg_31_0__7_), .Q(b_reg_7_), .R(reset_n_bF_buf49), .S(1'h1));
DFFSR DFFSR_400 ( .CLK(clk_bF_buf45), .D(w_mem_inst__0w_mem_1__31_0__29_), .Q(w_mem_inst_w_mem_1__29_), .R(reset_n_bF_buf45), .S(1'h1));
DFFSR DFFSR_401 ( .CLK(clk_bF_buf44), .D(w_mem_inst__0w_mem_1__31_0__30_), .Q(w_mem_inst_w_mem_1__30_), .R(reset_n_bF_buf44), .S(1'h1));
DFFSR DFFSR_402 ( .CLK(clk_bF_buf43), .D(w_mem_inst__0w_mem_1__31_0__31_), .Q(w_mem_inst_w_mem_1__31_), .R(reset_n_bF_buf43), .S(1'h1));
DFFSR DFFSR_403 ( .CLK(clk_bF_buf42), .D(w_mem_inst__0w_mem_2__31_0__0_), .Q(w_mem_inst_w_mem_2__0_), .R(reset_n_bF_buf42), .S(1'h1));
DFFSR DFFSR_404 ( .CLK(clk_bF_buf41), .D(w_mem_inst__0w_mem_2__31_0__1_), .Q(w_mem_inst_w_mem_2__1_), .R(reset_n_bF_buf41), .S(1'h1));
DFFSR DFFSR_405 ( .CLK(clk_bF_buf40), .D(w_mem_inst__0w_mem_2__31_0__2_), .Q(w_mem_inst_w_mem_2__2_), .R(reset_n_bF_buf40), .S(1'h1));
DFFSR DFFSR_406 ( .CLK(clk_bF_buf39), .D(w_mem_inst__0w_mem_2__31_0__3_), .Q(w_mem_inst_w_mem_2__3_), .R(reset_n_bF_buf39), .S(1'h1));
DFFSR DFFSR_407 ( .CLK(clk_bF_buf38), .D(w_mem_inst__0w_mem_2__31_0__4_), .Q(w_mem_inst_w_mem_2__4_), .R(reset_n_bF_buf38), .S(1'h1));
DFFSR DFFSR_408 ( .CLK(clk_bF_buf37), .D(w_mem_inst__0w_mem_2__31_0__5_), .Q(w_mem_inst_w_mem_2__5_), .R(reset_n_bF_buf37), .S(1'h1));
DFFSR DFFSR_409 ( .CLK(clk_bF_buf36), .D(w_mem_inst__0w_mem_2__31_0__6_), .Q(w_mem_inst_w_mem_2__6_), .R(reset_n_bF_buf36), .S(1'h1));
DFFSR DFFSR_41 ( .CLK(clk_bF_buf48), .D(_0b_reg_31_0__8_), .Q(b_reg_8_), .R(reset_n_bF_buf48), .S(1'h1));
DFFSR DFFSR_410 ( .CLK(clk_bF_buf35), .D(w_mem_inst__0w_mem_2__31_0__7_), .Q(w_mem_inst_w_mem_2__7_), .R(reset_n_bF_buf35), .S(1'h1));
DFFSR DFFSR_411 ( .CLK(clk_bF_buf34), .D(w_mem_inst__0w_mem_2__31_0__8_), .Q(w_mem_inst_w_mem_2__8_), .R(reset_n_bF_buf34), .S(1'h1));
DFFSR DFFSR_412 ( .CLK(clk_bF_buf33), .D(w_mem_inst__0w_mem_2__31_0__9_), .Q(w_mem_inst_w_mem_2__9_), .R(reset_n_bF_buf33), .S(1'h1));
DFFSR DFFSR_413 ( .CLK(clk_bF_buf32), .D(w_mem_inst__0w_mem_2__31_0__10_), .Q(w_mem_inst_w_mem_2__10_), .R(reset_n_bF_buf32), .S(1'h1));
DFFSR DFFSR_414 ( .CLK(clk_bF_buf31), .D(w_mem_inst__0w_mem_2__31_0__11_), .Q(w_mem_inst_w_mem_2__11_), .R(reset_n_bF_buf31), .S(1'h1));
DFFSR DFFSR_415 ( .CLK(clk_bF_buf30), .D(w_mem_inst__0w_mem_2__31_0__12_), .Q(w_mem_inst_w_mem_2__12_), .R(reset_n_bF_buf30), .S(1'h1));
DFFSR DFFSR_416 ( .CLK(clk_bF_buf29), .D(w_mem_inst__0w_mem_2__31_0__13_), .Q(w_mem_inst_w_mem_2__13_), .R(reset_n_bF_buf29), .S(1'h1));
DFFSR DFFSR_417 ( .CLK(clk_bF_buf28), .D(w_mem_inst__0w_mem_2__31_0__14_), .Q(w_mem_inst_w_mem_2__14_), .R(reset_n_bF_buf28), .S(1'h1));
DFFSR DFFSR_418 ( .CLK(clk_bF_buf27), .D(w_mem_inst__0w_mem_2__31_0__15_), .Q(w_mem_inst_w_mem_2__15_), .R(reset_n_bF_buf27), .S(1'h1));
DFFSR DFFSR_419 ( .CLK(clk_bF_buf26), .D(w_mem_inst__0w_mem_2__31_0__16_), .Q(w_mem_inst_w_mem_2__16_), .R(reset_n_bF_buf26), .S(1'h1));
DFFSR DFFSR_42 ( .CLK(clk_bF_buf47), .D(_0b_reg_31_0__9_), .Q(b_reg_9_), .R(reset_n_bF_buf47), .S(1'h1));
DFFSR DFFSR_420 ( .CLK(clk_bF_buf25), .D(w_mem_inst__0w_mem_2__31_0__17_), .Q(w_mem_inst_w_mem_2__17_), .R(reset_n_bF_buf25), .S(1'h1));
DFFSR DFFSR_421 ( .CLK(clk_bF_buf24), .D(w_mem_inst__0w_mem_2__31_0__18_), .Q(w_mem_inst_w_mem_2__18_), .R(reset_n_bF_buf24), .S(1'h1));
DFFSR DFFSR_422 ( .CLK(clk_bF_buf23), .D(w_mem_inst__0w_mem_2__31_0__19_), .Q(w_mem_inst_w_mem_2__19_), .R(reset_n_bF_buf23), .S(1'h1));
DFFSR DFFSR_423 ( .CLK(clk_bF_buf22), .D(w_mem_inst__0w_mem_2__31_0__20_), .Q(w_mem_inst_w_mem_2__20_), .R(reset_n_bF_buf22), .S(1'h1));
DFFSR DFFSR_424 ( .CLK(clk_bF_buf21), .D(w_mem_inst__0w_mem_2__31_0__21_), .Q(w_mem_inst_w_mem_2__21_), .R(reset_n_bF_buf21), .S(1'h1));
DFFSR DFFSR_425 ( .CLK(clk_bF_buf20), .D(w_mem_inst__0w_mem_2__31_0__22_), .Q(w_mem_inst_w_mem_2__22_), .R(reset_n_bF_buf20), .S(1'h1));
DFFSR DFFSR_426 ( .CLK(clk_bF_buf19), .D(w_mem_inst__0w_mem_2__31_0__23_), .Q(w_mem_inst_w_mem_2__23_), .R(reset_n_bF_buf19), .S(1'h1));
DFFSR DFFSR_427 ( .CLK(clk_bF_buf18), .D(w_mem_inst__0w_mem_2__31_0__24_), .Q(w_mem_inst_w_mem_2__24_), .R(reset_n_bF_buf18), .S(1'h1));
DFFSR DFFSR_428 ( .CLK(clk_bF_buf17), .D(w_mem_inst__0w_mem_2__31_0__25_), .Q(w_mem_inst_w_mem_2__25_), .R(reset_n_bF_buf17), .S(1'h1));
DFFSR DFFSR_429 ( .CLK(clk_bF_buf16), .D(w_mem_inst__0w_mem_2__31_0__26_), .Q(w_mem_inst_w_mem_2__26_), .R(reset_n_bF_buf16), .S(1'h1));
DFFSR DFFSR_43 ( .CLK(clk_bF_buf46), .D(_0b_reg_31_0__10_), .Q(b_reg_10_), .R(reset_n_bF_buf46), .S(1'h1));
DFFSR DFFSR_430 ( .CLK(clk_bF_buf15), .D(w_mem_inst__0w_mem_2__31_0__27_), .Q(w_mem_inst_w_mem_2__27_), .R(reset_n_bF_buf15), .S(1'h1));
DFFSR DFFSR_431 ( .CLK(clk_bF_buf14), .D(w_mem_inst__0w_mem_2__31_0__28_), .Q(w_mem_inst_w_mem_2__28_), .R(reset_n_bF_buf14), .S(1'h1));
DFFSR DFFSR_432 ( .CLK(clk_bF_buf13), .D(w_mem_inst__0w_mem_2__31_0__29_), .Q(w_mem_inst_w_mem_2__29_), .R(reset_n_bF_buf13), .S(1'h1));
DFFSR DFFSR_433 ( .CLK(clk_bF_buf12), .D(w_mem_inst__0w_mem_2__31_0__30_), .Q(w_mem_inst_w_mem_2__30_), .R(reset_n_bF_buf12), .S(1'h1));
DFFSR DFFSR_434 ( .CLK(clk_bF_buf11), .D(w_mem_inst__0w_mem_2__31_0__31_), .Q(w_mem_inst_w_mem_2__31_), .R(reset_n_bF_buf11), .S(1'h1));
DFFSR DFFSR_435 ( .CLK(clk_bF_buf10), .D(w_mem_inst__0w_mem_3__31_0__0_), .Q(w_mem_inst_w_mem_3__0_), .R(reset_n_bF_buf10), .S(1'h1));
DFFSR DFFSR_436 ( .CLK(clk_bF_buf9), .D(w_mem_inst__0w_mem_3__31_0__1_), .Q(w_mem_inst_w_mem_3__1_), .R(reset_n_bF_buf9), .S(1'h1));
DFFSR DFFSR_437 ( .CLK(clk_bF_buf8), .D(w_mem_inst__0w_mem_3__31_0__2_), .Q(w_mem_inst_w_mem_3__2_), .R(reset_n_bF_buf8), .S(1'h1));
DFFSR DFFSR_438 ( .CLK(clk_bF_buf7), .D(w_mem_inst__0w_mem_3__31_0__3_), .Q(w_mem_inst_w_mem_3__3_), .R(reset_n_bF_buf7), .S(1'h1));
DFFSR DFFSR_439 ( .CLK(clk_bF_buf6), .D(w_mem_inst__0w_mem_3__31_0__4_), .Q(w_mem_inst_w_mem_3__4_), .R(reset_n_bF_buf6), .S(1'h1));
DFFSR DFFSR_44 ( .CLK(clk_bF_buf45), .D(_0b_reg_31_0__11_), .Q(b_reg_11_), .R(reset_n_bF_buf45), .S(1'h1));
DFFSR DFFSR_440 ( .CLK(clk_bF_buf5), .D(w_mem_inst__0w_mem_3__31_0__5_), .Q(w_mem_inst_w_mem_3__5_), .R(reset_n_bF_buf5), .S(1'h1));
DFFSR DFFSR_441 ( .CLK(clk_bF_buf4), .D(w_mem_inst__0w_mem_3__31_0__6_), .Q(w_mem_inst_w_mem_3__6_), .R(reset_n_bF_buf4), .S(1'h1));
DFFSR DFFSR_442 ( .CLK(clk_bF_buf3), .D(w_mem_inst__0w_mem_3__31_0__7_), .Q(w_mem_inst_w_mem_3__7_), .R(reset_n_bF_buf3), .S(1'h1));
DFFSR DFFSR_443 ( .CLK(clk_bF_buf2), .D(w_mem_inst__0w_mem_3__31_0__8_), .Q(w_mem_inst_w_mem_3__8_), .R(reset_n_bF_buf2), .S(1'h1));
DFFSR DFFSR_444 ( .CLK(clk_bF_buf1), .D(w_mem_inst__0w_mem_3__31_0__9_), .Q(w_mem_inst_w_mem_3__9_), .R(reset_n_bF_buf1), .S(1'h1));
DFFSR DFFSR_445 ( .CLK(clk_bF_buf0), .D(w_mem_inst__0w_mem_3__31_0__10_), .Q(w_mem_inst_w_mem_3__10_), .R(reset_n_bF_buf0), .S(1'h1));
DFFSR DFFSR_446 ( .CLK(clk_bF_buf88), .D(w_mem_inst__0w_mem_3__31_0__11_), .Q(w_mem_inst_w_mem_3__11_), .R(reset_n_bF_buf88), .S(1'h1));
DFFSR DFFSR_447 ( .CLK(clk_bF_buf87), .D(w_mem_inst__0w_mem_3__31_0__12_), .Q(w_mem_inst_w_mem_3__12_), .R(reset_n_bF_buf87), .S(1'h1));
DFFSR DFFSR_448 ( .CLK(clk_bF_buf86), .D(w_mem_inst__0w_mem_3__31_0__13_), .Q(w_mem_inst_w_mem_3__13_), .R(reset_n_bF_buf86), .S(1'h1));
DFFSR DFFSR_449 ( .CLK(clk_bF_buf85), .D(w_mem_inst__0w_mem_3__31_0__14_), .Q(w_mem_inst_w_mem_3__14_), .R(reset_n_bF_buf85), .S(1'h1));
DFFSR DFFSR_45 ( .CLK(clk_bF_buf44), .D(_0b_reg_31_0__12_), .Q(b_reg_12_), .R(reset_n_bF_buf44), .S(1'h1));
DFFSR DFFSR_450 ( .CLK(clk_bF_buf84), .D(w_mem_inst__0w_mem_3__31_0__15_), .Q(w_mem_inst_w_mem_3__15_), .R(reset_n_bF_buf84), .S(1'h1));
DFFSR DFFSR_451 ( .CLK(clk_bF_buf83), .D(w_mem_inst__0w_mem_3__31_0__16_), .Q(w_mem_inst_w_mem_3__16_), .R(reset_n_bF_buf83), .S(1'h1));
DFFSR DFFSR_452 ( .CLK(clk_bF_buf82), .D(w_mem_inst__0w_mem_3__31_0__17_), .Q(w_mem_inst_w_mem_3__17_), .R(reset_n_bF_buf82), .S(1'h1));
DFFSR DFFSR_453 ( .CLK(clk_bF_buf81), .D(w_mem_inst__0w_mem_3__31_0__18_), .Q(w_mem_inst_w_mem_3__18_), .R(reset_n_bF_buf81), .S(1'h1));
DFFSR DFFSR_454 ( .CLK(clk_bF_buf80), .D(w_mem_inst__0w_mem_3__31_0__19_), .Q(w_mem_inst_w_mem_3__19_), .R(reset_n_bF_buf80), .S(1'h1));
DFFSR DFFSR_455 ( .CLK(clk_bF_buf79), .D(w_mem_inst__0w_mem_3__31_0__20_), .Q(w_mem_inst_w_mem_3__20_), .R(reset_n_bF_buf79), .S(1'h1));
DFFSR DFFSR_456 ( .CLK(clk_bF_buf78), .D(w_mem_inst__0w_mem_3__31_0__21_), .Q(w_mem_inst_w_mem_3__21_), .R(reset_n_bF_buf78), .S(1'h1));
DFFSR DFFSR_457 ( .CLK(clk_bF_buf77), .D(w_mem_inst__0w_mem_3__31_0__22_), .Q(w_mem_inst_w_mem_3__22_), .R(reset_n_bF_buf77), .S(1'h1));
DFFSR DFFSR_458 ( .CLK(clk_bF_buf76), .D(w_mem_inst__0w_mem_3__31_0__23_), .Q(w_mem_inst_w_mem_3__23_), .R(reset_n_bF_buf76), .S(1'h1));
DFFSR DFFSR_459 ( .CLK(clk_bF_buf75), .D(w_mem_inst__0w_mem_3__31_0__24_), .Q(w_mem_inst_w_mem_3__24_), .R(reset_n_bF_buf75), .S(1'h1));
DFFSR DFFSR_46 ( .CLK(clk_bF_buf43), .D(_0b_reg_31_0__13_), .Q(b_reg_13_), .R(reset_n_bF_buf43), .S(1'h1));
DFFSR DFFSR_460 ( .CLK(clk_bF_buf74), .D(w_mem_inst__0w_mem_3__31_0__25_), .Q(w_mem_inst_w_mem_3__25_), .R(reset_n_bF_buf74), .S(1'h1));
DFFSR DFFSR_461 ( .CLK(clk_bF_buf73), .D(w_mem_inst__0w_mem_3__31_0__26_), .Q(w_mem_inst_w_mem_3__26_), .R(reset_n_bF_buf73), .S(1'h1));
DFFSR DFFSR_462 ( .CLK(clk_bF_buf72), .D(w_mem_inst__0w_mem_3__31_0__27_), .Q(w_mem_inst_w_mem_3__27_), .R(reset_n_bF_buf72), .S(1'h1));
DFFSR DFFSR_463 ( .CLK(clk_bF_buf71), .D(w_mem_inst__0w_mem_3__31_0__28_), .Q(w_mem_inst_w_mem_3__28_), .R(reset_n_bF_buf71), .S(1'h1));
DFFSR DFFSR_464 ( .CLK(clk_bF_buf70), .D(w_mem_inst__0w_mem_3__31_0__29_), .Q(w_mem_inst_w_mem_3__29_), .R(reset_n_bF_buf70), .S(1'h1));
DFFSR DFFSR_465 ( .CLK(clk_bF_buf69), .D(w_mem_inst__0w_mem_3__31_0__30_), .Q(w_mem_inst_w_mem_3__30_), .R(reset_n_bF_buf69), .S(1'h1));
DFFSR DFFSR_466 ( .CLK(clk_bF_buf68), .D(w_mem_inst__0w_mem_3__31_0__31_), .Q(w_mem_inst_w_mem_3__31_), .R(reset_n_bF_buf68), .S(1'h1));
DFFSR DFFSR_467 ( .CLK(clk_bF_buf67), .D(w_mem_inst__0w_mem_4__31_0__0_), .Q(w_mem_inst_w_mem_4__0_), .R(reset_n_bF_buf67), .S(1'h1));
DFFSR DFFSR_468 ( .CLK(clk_bF_buf66), .D(w_mem_inst__0w_mem_4__31_0__1_), .Q(w_mem_inst_w_mem_4__1_), .R(reset_n_bF_buf66), .S(1'h1));
DFFSR DFFSR_469 ( .CLK(clk_bF_buf65), .D(w_mem_inst__0w_mem_4__31_0__2_), .Q(w_mem_inst_w_mem_4__2_), .R(reset_n_bF_buf65), .S(1'h1));
DFFSR DFFSR_47 ( .CLK(clk_bF_buf42), .D(_0b_reg_31_0__14_), .Q(b_reg_14_), .R(reset_n_bF_buf42), .S(1'h1));
DFFSR DFFSR_470 ( .CLK(clk_bF_buf64), .D(w_mem_inst__0w_mem_4__31_0__3_), .Q(w_mem_inst_w_mem_4__3_), .R(reset_n_bF_buf64), .S(1'h1));
DFFSR DFFSR_471 ( .CLK(clk_bF_buf63), .D(w_mem_inst__0w_mem_4__31_0__4_), .Q(w_mem_inst_w_mem_4__4_), .R(reset_n_bF_buf63), .S(1'h1));
DFFSR DFFSR_472 ( .CLK(clk_bF_buf62), .D(w_mem_inst__0w_mem_4__31_0__5_), .Q(w_mem_inst_w_mem_4__5_), .R(reset_n_bF_buf62), .S(1'h1));
DFFSR DFFSR_473 ( .CLK(clk_bF_buf61), .D(w_mem_inst__0w_mem_4__31_0__6_), .Q(w_mem_inst_w_mem_4__6_), .R(reset_n_bF_buf61), .S(1'h1));
DFFSR DFFSR_474 ( .CLK(clk_bF_buf60), .D(w_mem_inst__0w_mem_4__31_0__7_), .Q(w_mem_inst_w_mem_4__7_), .R(reset_n_bF_buf60), .S(1'h1));
DFFSR DFFSR_475 ( .CLK(clk_bF_buf59), .D(w_mem_inst__0w_mem_4__31_0__8_), .Q(w_mem_inst_w_mem_4__8_), .R(reset_n_bF_buf59), .S(1'h1));
DFFSR DFFSR_476 ( .CLK(clk_bF_buf58), .D(w_mem_inst__0w_mem_4__31_0__9_), .Q(w_mem_inst_w_mem_4__9_), .R(reset_n_bF_buf58), .S(1'h1));
DFFSR DFFSR_477 ( .CLK(clk_bF_buf57), .D(w_mem_inst__0w_mem_4__31_0__10_), .Q(w_mem_inst_w_mem_4__10_), .R(reset_n_bF_buf57), .S(1'h1));
DFFSR DFFSR_478 ( .CLK(clk_bF_buf56), .D(w_mem_inst__0w_mem_4__31_0__11_), .Q(w_mem_inst_w_mem_4__11_), .R(reset_n_bF_buf56), .S(1'h1));
DFFSR DFFSR_479 ( .CLK(clk_bF_buf55), .D(w_mem_inst__0w_mem_4__31_0__12_), .Q(w_mem_inst_w_mem_4__12_), .R(reset_n_bF_buf55), .S(1'h1));
DFFSR DFFSR_48 ( .CLK(clk_bF_buf41), .D(_0b_reg_31_0__15_), .Q(b_reg_15_), .R(reset_n_bF_buf41), .S(1'h1));
DFFSR DFFSR_480 ( .CLK(clk_bF_buf54), .D(w_mem_inst__0w_mem_4__31_0__13_), .Q(w_mem_inst_w_mem_4__13_), .R(reset_n_bF_buf54), .S(1'h1));
DFFSR DFFSR_481 ( .CLK(clk_bF_buf53), .D(w_mem_inst__0w_mem_4__31_0__14_), .Q(w_mem_inst_w_mem_4__14_), .R(reset_n_bF_buf53), .S(1'h1));
DFFSR DFFSR_482 ( .CLK(clk_bF_buf52), .D(w_mem_inst__0w_mem_4__31_0__15_), .Q(w_mem_inst_w_mem_4__15_), .R(reset_n_bF_buf52), .S(1'h1));
DFFSR DFFSR_483 ( .CLK(clk_bF_buf51), .D(w_mem_inst__0w_mem_4__31_0__16_), .Q(w_mem_inst_w_mem_4__16_), .R(reset_n_bF_buf51), .S(1'h1));
DFFSR DFFSR_484 ( .CLK(clk_bF_buf50), .D(w_mem_inst__0w_mem_4__31_0__17_), .Q(w_mem_inst_w_mem_4__17_), .R(reset_n_bF_buf50), .S(1'h1));
DFFSR DFFSR_485 ( .CLK(clk_bF_buf49), .D(w_mem_inst__0w_mem_4__31_0__18_), .Q(w_mem_inst_w_mem_4__18_), .R(reset_n_bF_buf49), .S(1'h1));
DFFSR DFFSR_486 ( .CLK(clk_bF_buf48), .D(w_mem_inst__0w_mem_4__31_0__19_), .Q(w_mem_inst_w_mem_4__19_), .R(reset_n_bF_buf48), .S(1'h1));
DFFSR DFFSR_487 ( .CLK(clk_bF_buf47), .D(w_mem_inst__0w_mem_4__31_0__20_), .Q(w_mem_inst_w_mem_4__20_), .R(reset_n_bF_buf47), .S(1'h1));
DFFSR DFFSR_488 ( .CLK(clk_bF_buf46), .D(w_mem_inst__0w_mem_4__31_0__21_), .Q(w_mem_inst_w_mem_4__21_), .R(reset_n_bF_buf46), .S(1'h1));
DFFSR DFFSR_489 ( .CLK(clk_bF_buf45), .D(w_mem_inst__0w_mem_4__31_0__22_), .Q(w_mem_inst_w_mem_4__22_), .R(reset_n_bF_buf45), .S(1'h1));
DFFSR DFFSR_49 ( .CLK(clk_bF_buf40), .D(_0b_reg_31_0__16_), .Q(b_reg_16_), .R(reset_n_bF_buf40), .S(1'h1));
DFFSR DFFSR_490 ( .CLK(clk_bF_buf44), .D(w_mem_inst__0w_mem_4__31_0__23_), .Q(w_mem_inst_w_mem_4__23_), .R(reset_n_bF_buf44), .S(1'h1));
DFFSR DFFSR_491 ( .CLK(clk_bF_buf43), .D(w_mem_inst__0w_mem_4__31_0__24_), .Q(w_mem_inst_w_mem_4__24_), .R(reset_n_bF_buf43), .S(1'h1));
DFFSR DFFSR_492 ( .CLK(clk_bF_buf42), .D(w_mem_inst__0w_mem_4__31_0__25_), .Q(w_mem_inst_w_mem_4__25_), .R(reset_n_bF_buf42), .S(1'h1));
DFFSR DFFSR_493 ( .CLK(clk_bF_buf41), .D(w_mem_inst__0w_mem_4__31_0__26_), .Q(w_mem_inst_w_mem_4__26_), .R(reset_n_bF_buf41), .S(1'h1));
DFFSR DFFSR_494 ( .CLK(clk_bF_buf40), .D(w_mem_inst__0w_mem_4__31_0__27_), .Q(w_mem_inst_w_mem_4__27_), .R(reset_n_bF_buf40), .S(1'h1));
DFFSR DFFSR_495 ( .CLK(clk_bF_buf39), .D(w_mem_inst__0w_mem_4__31_0__28_), .Q(w_mem_inst_w_mem_4__28_), .R(reset_n_bF_buf39), .S(1'h1));
DFFSR DFFSR_496 ( .CLK(clk_bF_buf38), .D(w_mem_inst__0w_mem_4__31_0__29_), .Q(w_mem_inst_w_mem_4__29_), .R(reset_n_bF_buf38), .S(1'h1));
DFFSR DFFSR_497 ( .CLK(clk_bF_buf37), .D(w_mem_inst__0w_mem_4__31_0__30_), .Q(w_mem_inst_w_mem_4__30_), .R(reset_n_bF_buf37), .S(1'h1));
DFFSR DFFSR_498 ( .CLK(clk_bF_buf36), .D(w_mem_inst__0w_mem_4__31_0__31_), .Q(w_mem_inst_w_mem_4__31_), .R(reset_n_bF_buf36), .S(1'h1));
DFFSR DFFSR_499 ( .CLK(clk_bF_buf35), .D(w_mem_inst__0w_mem_5__31_0__0_), .Q(w_mem_inst_w_mem_5__0_), .R(reset_n_bF_buf35), .S(1'h1));
DFFSR DFFSR_5 ( .CLK(clk_bF_buf84), .D(_0a_reg_31_0__4_), .Q(a_reg_4_), .R(reset_n_bF_buf84), .S(1'h1));
DFFSR DFFSR_50 ( .CLK(clk_bF_buf39), .D(_0b_reg_31_0__17_), .Q(b_reg_17_), .R(reset_n_bF_buf39), .S(1'h1));
DFFSR DFFSR_500 ( .CLK(clk_bF_buf34), .D(w_mem_inst__0w_mem_5__31_0__1_), .Q(w_mem_inst_w_mem_5__1_), .R(reset_n_bF_buf34), .S(1'h1));
DFFSR DFFSR_501 ( .CLK(clk_bF_buf33), .D(w_mem_inst__0w_mem_5__31_0__2_), .Q(w_mem_inst_w_mem_5__2_), .R(reset_n_bF_buf33), .S(1'h1));
DFFSR DFFSR_502 ( .CLK(clk_bF_buf32), .D(w_mem_inst__0w_mem_5__31_0__3_), .Q(w_mem_inst_w_mem_5__3_), .R(reset_n_bF_buf32), .S(1'h1));
DFFSR DFFSR_503 ( .CLK(clk_bF_buf31), .D(w_mem_inst__0w_mem_5__31_0__4_), .Q(w_mem_inst_w_mem_5__4_), .R(reset_n_bF_buf31), .S(1'h1));
DFFSR DFFSR_504 ( .CLK(clk_bF_buf30), .D(w_mem_inst__0w_mem_5__31_0__5_), .Q(w_mem_inst_w_mem_5__5_), .R(reset_n_bF_buf30), .S(1'h1));
DFFSR DFFSR_505 ( .CLK(clk_bF_buf29), .D(w_mem_inst__0w_mem_5__31_0__6_), .Q(w_mem_inst_w_mem_5__6_), .R(reset_n_bF_buf29), .S(1'h1));
DFFSR DFFSR_506 ( .CLK(clk_bF_buf28), .D(w_mem_inst__0w_mem_5__31_0__7_), .Q(w_mem_inst_w_mem_5__7_), .R(reset_n_bF_buf28), .S(1'h1));
DFFSR DFFSR_507 ( .CLK(clk_bF_buf27), .D(w_mem_inst__0w_mem_5__31_0__8_), .Q(w_mem_inst_w_mem_5__8_), .R(reset_n_bF_buf27), .S(1'h1));
DFFSR DFFSR_508 ( .CLK(clk_bF_buf26), .D(w_mem_inst__0w_mem_5__31_0__9_), .Q(w_mem_inst_w_mem_5__9_), .R(reset_n_bF_buf26), .S(1'h1));
DFFSR DFFSR_509 ( .CLK(clk_bF_buf25), .D(w_mem_inst__0w_mem_5__31_0__10_), .Q(w_mem_inst_w_mem_5__10_), .R(reset_n_bF_buf25), .S(1'h1));
DFFSR DFFSR_51 ( .CLK(clk_bF_buf38), .D(_0b_reg_31_0__18_), .Q(b_reg_18_), .R(reset_n_bF_buf38), .S(1'h1));
DFFSR DFFSR_510 ( .CLK(clk_bF_buf24), .D(w_mem_inst__0w_mem_5__31_0__11_), .Q(w_mem_inst_w_mem_5__11_), .R(reset_n_bF_buf24), .S(1'h1));
DFFSR DFFSR_511 ( .CLK(clk_bF_buf23), .D(w_mem_inst__0w_mem_5__31_0__12_), .Q(w_mem_inst_w_mem_5__12_), .R(reset_n_bF_buf23), .S(1'h1));
DFFSR DFFSR_512 ( .CLK(clk_bF_buf22), .D(w_mem_inst__0w_mem_5__31_0__13_), .Q(w_mem_inst_w_mem_5__13_), .R(reset_n_bF_buf22), .S(1'h1));
DFFSR DFFSR_513 ( .CLK(clk_bF_buf21), .D(w_mem_inst__0w_mem_5__31_0__14_), .Q(w_mem_inst_w_mem_5__14_), .R(reset_n_bF_buf21), .S(1'h1));
DFFSR DFFSR_514 ( .CLK(clk_bF_buf20), .D(w_mem_inst__0w_mem_5__31_0__15_), .Q(w_mem_inst_w_mem_5__15_), .R(reset_n_bF_buf20), .S(1'h1));
DFFSR DFFSR_515 ( .CLK(clk_bF_buf19), .D(w_mem_inst__0w_mem_5__31_0__16_), .Q(w_mem_inst_w_mem_5__16_), .R(reset_n_bF_buf19), .S(1'h1));
DFFSR DFFSR_516 ( .CLK(clk_bF_buf18), .D(w_mem_inst__0w_mem_5__31_0__17_), .Q(w_mem_inst_w_mem_5__17_), .R(reset_n_bF_buf18), .S(1'h1));
DFFSR DFFSR_517 ( .CLK(clk_bF_buf17), .D(w_mem_inst__0w_mem_5__31_0__18_), .Q(w_mem_inst_w_mem_5__18_), .R(reset_n_bF_buf17), .S(1'h1));
DFFSR DFFSR_518 ( .CLK(clk_bF_buf16), .D(w_mem_inst__0w_mem_5__31_0__19_), .Q(w_mem_inst_w_mem_5__19_), .R(reset_n_bF_buf16), .S(1'h1));
DFFSR DFFSR_519 ( .CLK(clk_bF_buf15), .D(w_mem_inst__0w_mem_5__31_0__20_), .Q(w_mem_inst_w_mem_5__20_), .R(reset_n_bF_buf15), .S(1'h1));
DFFSR DFFSR_52 ( .CLK(clk_bF_buf37), .D(_0b_reg_31_0__19_), .Q(b_reg_19_), .R(reset_n_bF_buf37), .S(1'h1));
DFFSR DFFSR_520 ( .CLK(clk_bF_buf14), .D(w_mem_inst__0w_mem_5__31_0__21_), .Q(w_mem_inst_w_mem_5__21_), .R(reset_n_bF_buf14), .S(1'h1));
DFFSR DFFSR_521 ( .CLK(clk_bF_buf13), .D(w_mem_inst__0w_mem_5__31_0__22_), .Q(w_mem_inst_w_mem_5__22_), .R(reset_n_bF_buf13), .S(1'h1));
DFFSR DFFSR_522 ( .CLK(clk_bF_buf12), .D(w_mem_inst__0w_mem_5__31_0__23_), .Q(w_mem_inst_w_mem_5__23_), .R(reset_n_bF_buf12), .S(1'h1));
DFFSR DFFSR_523 ( .CLK(clk_bF_buf11), .D(w_mem_inst__0w_mem_5__31_0__24_), .Q(w_mem_inst_w_mem_5__24_), .R(reset_n_bF_buf11), .S(1'h1));
DFFSR DFFSR_524 ( .CLK(clk_bF_buf10), .D(w_mem_inst__0w_mem_5__31_0__25_), .Q(w_mem_inst_w_mem_5__25_), .R(reset_n_bF_buf10), .S(1'h1));
DFFSR DFFSR_525 ( .CLK(clk_bF_buf9), .D(w_mem_inst__0w_mem_5__31_0__26_), .Q(w_mem_inst_w_mem_5__26_), .R(reset_n_bF_buf9), .S(1'h1));
DFFSR DFFSR_526 ( .CLK(clk_bF_buf8), .D(w_mem_inst__0w_mem_5__31_0__27_), .Q(w_mem_inst_w_mem_5__27_), .R(reset_n_bF_buf8), .S(1'h1));
DFFSR DFFSR_527 ( .CLK(clk_bF_buf7), .D(w_mem_inst__0w_mem_5__31_0__28_), .Q(w_mem_inst_w_mem_5__28_), .R(reset_n_bF_buf7), .S(1'h1));
DFFSR DFFSR_528 ( .CLK(clk_bF_buf6), .D(w_mem_inst__0w_mem_5__31_0__29_), .Q(w_mem_inst_w_mem_5__29_), .R(reset_n_bF_buf6), .S(1'h1));
DFFSR DFFSR_529 ( .CLK(clk_bF_buf5), .D(w_mem_inst__0w_mem_5__31_0__30_), .Q(w_mem_inst_w_mem_5__30_), .R(reset_n_bF_buf5), .S(1'h1));
DFFSR DFFSR_53 ( .CLK(clk_bF_buf36), .D(_0b_reg_31_0__20_), .Q(b_reg_20_), .R(reset_n_bF_buf36), .S(1'h1));
DFFSR DFFSR_530 ( .CLK(clk_bF_buf4), .D(w_mem_inst__0w_mem_5__31_0__31_), .Q(w_mem_inst_w_mem_5__31_), .R(reset_n_bF_buf4), .S(1'h1));
DFFSR DFFSR_531 ( .CLK(clk_bF_buf3), .D(w_mem_inst__0w_mem_6__31_0__0_), .Q(w_mem_inst_w_mem_6__0_), .R(reset_n_bF_buf3), .S(1'h1));
DFFSR DFFSR_532 ( .CLK(clk_bF_buf2), .D(w_mem_inst__0w_mem_6__31_0__1_), .Q(w_mem_inst_w_mem_6__1_), .R(reset_n_bF_buf2), .S(1'h1));
DFFSR DFFSR_533 ( .CLK(clk_bF_buf1), .D(w_mem_inst__0w_mem_6__31_0__2_), .Q(w_mem_inst_w_mem_6__2_), .R(reset_n_bF_buf1), .S(1'h1));
DFFSR DFFSR_534 ( .CLK(clk_bF_buf0), .D(w_mem_inst__0w_mem_6__31_0__3_), .Q(w_mem_inst_w_mem_6__3_), .R(reset_n_bF_buf0), .S(1'h1));
DFFSR DFFSR_535 ( .CLK(clk_bF_buf88), .D(w_mem_inst__0w_mem_6__31_0__4_), .Q(w_mem_inst_w_mem_6__4_), .R(reset_n_bF_buf88), .S(1'h1));
DFFSR DFFSR_536 ( .CLK(clk_bF_buf87), .D(w_mem_inst__0w_mem_6__31_0__5_), .Q(w_mem_inst_w_mem_6__5_), .R(reset_n_bF_buf87), .S(1'h1));
DFFSR DFFSR_537 ( .CLK(clk_bF_buf86), .D(w_mem_inst__0w_mem_6__31_0__6_), .Q(w_mem_inst_w_mem_6__6_), .R(reset_n_bF_buf86), .S(1'h1));
DFFSR DFFSR_538 ( .CLK(clk_bF_buf85), .D(w_mem_inst__0w_mem_6__31_0__7_), .Q(w_mem_inst_w_mem_6__7_), .R(reset_n_bF_buf85), .S(1'h1));
DFFSR DFFSR_539 ( .CLK(clk_bF_buf84), .D(w_mem_inst__0w_mem_6__31_0__8_), .Q(w_mem_inst_w_mem_6__8_), .R(reset_n_bF_buf84), .S(1'h1));
DFFSR DFFSR_54 ( .CLK(clk_bF_buf35), .D(_0b_reg_31_0__21_), .Q(b_reg_21_), .R(reset_n_bF_buf35), .S(1'h1));
DFFSR DFFSR_540 ( .CLK(clk_bF_buf83), .D(w_mem_inst__0w_mem_6__31_0__9_), .Q(w_mem_inst_w_mem_6__9_), .R(reset_n_bF_buf83), .S(1'h1));
DFFSR DFFSR_541 ( .CLK(clk_bF_buf82), .D(w_mem_inst__0w_mem_6__31_0__10_), .Q(w_mem_inst_w_mem_6__10_), .R(reset_n_bF_buf82), .S(1'h1));
DFFSR DFFSR_542 ( .CLK(clk_bF_buf81), .D(w_mem_inst__0w_mem_6__31_0__11_), .Q(w_mem_inst_w_mem_6__11_), .R(reset_n_bF_buf81), .S(1'h1));
DFFSR DFFSR_543 ( .CLK(clk_bF_buf80), .D(w_mem_inst__0w_mem_6__31_0__12_), .Q(w_mem_inst_w_mem_6__12_), .R(reset_n_bF_buf80), .S(1'h1));
DFFSR DFFSR_544 ( .CLK(clk_bF_buf79), .D(w_mem_inst__0w_mem_6__31_0__13_), .Q(w_mem_inst_w_mem_6__13_), .R(reset_n_bF_buf79), .S(1'h1));
DFFSR DFFSR_545 ( .CLK(clk_bF_buf78), .D(w_mem_inst__0w_mem_6__31_0__14_), .Q(w_mem_inst_w_mem_6__14_), .R(reset_n_bF_buf78), .S(1'h1));
DFFSR DFFSR_546 ( .CLK(clk_bF_buf77), .D(w_mem_inst__0w_mem_6__31_0__15_), .Q(w_mem_inst_w_mem_6__15_), .R(reset_n_bF_buf77), .S(1'h1));
DFFSR DFFSR_547 ( .CLK(clk_bF_buf76), .D(w_mem_inst__0w_mem_6__31_0__16_), .Q(w_mem_inst_w_mem_6__16_), .R(reset_n_bF_buf76), .S(1'h1));
DFFSR DFFSR_548 ( .CLK(clk_bF_buf75), .D(w_mem_inst__0w_mem_6__31_0__17_), .Q(w_mem_inst_w_mem_6__17_), .R(reset_n_bF_buf75), .S(1'h1));
DFFSR DFFSR_549 ( .CLK(clk_bF_buf74), .D(w_mem_inst__0w_mem_6__31_0__18_), .Q(w_mem_inst_w_mem_6__18_), .R(reset_n_bF_buf74), .S(1'h1));
DFFSR DFFSR_55 ( .CLK(clk_bF_buf34), .D(_0b_reg_31_0__22_), .Q(b_reg_22_), .R(reset_n_bF_buf34), .S(1'h1));
DFFSR DFFSR_550 ( .CLK(clk_bF_buf73), .D(w_mem_inst__0w_mem_6__31_0__19_), .Q(w_mem_inst_w_mem_6__19_), .R(reset_n_bF_buf73), .S(1'h1));
DFFSR DFFSR_551 ( .CLK(clk_bF_buf72), .D(w_mem_inst__0w_mem_6__31_0__20_), .Q(w_mem_inst_w_mem_6__20_), .R(reset_n_bF_buf72), .S(1'h1));
DFFSR DFFSR_552 ( .CLK(clk_bF_buf71), .D(w_mem_inst__0w_mem_6__31_0__21_), .Q(w_mem_inst_w_mem_6__21_), .R(reset_n_bF_buf71), .S(1'h1));
DFFSR DFFSR_553 ( .CLK(clk_bF_buf70), .D(w_mem_inst__0w_mem_6__31_0__22_), .Q(w_mem_inst_w_mem_6__22_), .R(reset_n_bF_buf70), .S(1'h1));
DFFSR DFFSR_554 ( .CLK(clk_bF_buf69), .D(w_mem_inst__0w_mem_6__31_0__23_), .Q(w_mem_inst_w_mem_6__23_), .R(reset_n_bF_buf69), .S(1'h1));
DFFSR DFFSR_555 ( .CLK(clk_bF_buf68), .D(w_mem_inst__0w_mem_6__31_0__24_), .Q(w_mem_inst_w_mem_6__24_), .R(reset_n_bF_buf68), .S(1'h1));
DFFSR DFFSR_556 ( .CLK(clk_bF_buf67), .D(w_mem_inst__0w_mem_6__31_0__25_), .Q(w_mem_inst_w_mem_6__25_), .R(reset_n_bF_buf67), .S(1'h1));
DFFSR DFFSR_557 ( .CLK(clk_bF_buf66), .D(w_mem_inst__0w_mem_6__31_0__26_), .Q(w_mem_inst_w_mem_6__26_), .R(reset_n_bF_buf66), .S(1'h1));
DFFSR DFFSR_558 ( .CLK(clk_bF_buf65), .D(w_mem_inst__0w_mem_6__31_0__27_), .Q(w_mem_inst_w_mem_6__27_), .R(reset_n_bF_buf65), .S(1'h1));
DFFSR DFFSR_559 ( .CLK(clk_bF_buf64), .D(w_mem_inst__0w_mem_6__31_0__28_), .Q(w_mem_inst_w_mem_6__28_), .R(reset_n_bF_buf64), .S(1'h1));
DFFSR DFFSR_56 ( .CLK(clk_bF_buf33), .D(_0b_reg_31_0__23_), .Q(b_reg_23_), .R(reset_n_bF_buf33), .S(1'h1));
DFFSR DFFSR_560 ( .CLK(clk_bF_buf63), .D(w_mem_inst__0w_mem_6__31_0__29_), .Q(w_mem_inst_w_mem_6__29_), .R(reset_n_bF_buf63), .S(1'h1));
DFFSR DFFSR_561 ( .CLK(clk_bF_buf62), .D(w_mem_inst__0w_mem_6__31_0__30_), .Q(w_mem_inst_w_mem_6__30_), .R(reset_n_bF_buf62), .S(1'h1));
DFFSR DFFSR_562 ( .CLK(clk_bF_buf61), .D(w_mem_inst__0w_mem_6__31_0__31_), .Q(w_mem_inst_w_mem_6__31_), .R(reset_n_bF_buf61), .S(1'h1));
DFFSR DFFSR_563 ( .CLK(clk_bF_buf60), .D(w_mem_inst__0w_mem_7__31_0__0_), .Q(w_mem_inst_w_mem_7__0_), .R(reset_n_bF_buf60), .S(1'h1));
DFFSR DFFSR_564 ( .CLK(clk_bF_buf59), .D(w_mem_inst__0w_mem_7__31_0__1_), .Q(w_mem_inst_w_mem_7__1_), .R(reset_n_bF_buf59), .S(1'h1));
DFFSR DFFSR_565 ( .CLK(clk_bF_buf58), .D(w_mem_inst__0w_mem_7__31_0__2_), .Q(w_mem_inst_w_mem_7__2_), .R(reset_n_bF_buf58), .S(1'h1));
DFFSR DFFSR_566 ( .CLK(clk_bF_buf57), .D(w_mem_inst__0w_mem_7__31_0__3_), .Q(w_mem_inst_w_mem_7__3_), .R(reset_n_bF_buf57), .S(1'h1));
DFFSR DFFSR_567 ( .CLK(clk_bF_buf56), .D(w_mem_inst__0w_mem_7__31_0__4_), .Q(w_mem_inst_w_mem_7__4_), .R(reset_n_bF_buf56), .S(1'h1));
DFFSR DFFSR_568 ( .CLK(clk_bF_buf55), .D(w_mem_inst__0w_mem_7__31_0__5_), .Q(w_mem_inst_w_mem_7__5_), .R(reset_n_bF_buf55), .S(1'h1));
DFFSR DFFSR_569 ( .CLK(clk_bF_buf54), .D(w_mem_inst__0w_mem_7__31_0__6_), .Q(w_mem_inst_w_mem_7__6_), .R(reset_n_bF_buf54), .S(1'h1));
DFFSR DFFSR_57 ( .CLK(clk_bF_buf32), .D(_0b_reg_31_0__24_), .Q(b_reg_24_), .R(reset_n_bF_buf32), .S(1'h1));
DFFSR DFFSR_570 ( .CLK(clk_bF_buf53), .D(w_mem_inst__0w_mem_7__31_0__7_), .Q(w_mem_inst_w_mem_7__7_), .R(reset_n_bF_buf53), .S(1'h1));
DFFSR DFFSR_571 ( .CLK(clk_bF_buf52), .D(w_mem_inst__0w_mem_7__31_0__8_), .Q(w_mem_inst_w_mem_7__8_), .R(reset_n_bF_buf52), .S(1'h1));
DFFSR DFFSR_572 ( .CLK(clk_bF_buf51), .D(w_mem_inst__0w_mem_7__31_0__9_), .Q(w_mem_inst_w_mem_7__9_), .R(reset_n_bF_buf51), .S(1'h1));
DFFSR DFFSR_573 ( .CLK(clk_bF_buf50), .D(w_mem_inst__0w_mem_7__31_0__10_), .Q(w_mem_inst_w_mem_7__10_), .R(reset_n_bF_buf50), .S(1'h1));
DFFSR DFFSR_574 ( .CLK(clk_bF_buf49), .D(w_mem_inst__0w_mem_7__31_0__11_), .Q(w_mem_inst_w_mem_7__11_), .R(reset_n_bF_buf49), .S(1'h1));
DFFSR DFFSR_575 ( .CLK(clk_bF_buf48), .D(w_mem_inst__0w_mem_7__31_0__12_), .Q(w_mem_inst_w_mem_7__12_), .R(reset_n_bF_buf48), .S(1'h1));
DFFSR DFFSR_576 ( .CLK(clk_bF_buf47), .D(w_mem_inst__0w_mem_7__31_0__13_), .Q(w_mem_inst_w_mem_7__13_), .R(reset_n_bF_buf47), .S(1'h1));
DFFSR DFFSR_577 ( .CLK(clk_bF_buf46), .D(w_mem_inst__0w_mem_7__31_0__14_), .Q(w_mem_inst_w_mem_7__14_), .R(reset_n_bF_buf46), .S(1'h1));
DFFSR DFFSR_578 ( .CLK(clk_bF_buf45), .D(w_mem_inst__0w_mem_7__31_0__15_), .Q(w_mem_inst_w_mem_7__15_), .R(reset_n_bF_buf45), .S(1'h1));
DFFSR DFFSR_579 ( .CLK(clk_bF_buf44), .D(w_mem_inst__0w_mem_7__31_0__16_), .Q(w_mem_inst_w_mem_7__16_), .R(reset_n_bF_buf44), .S(1'h1));
DFFSR DFFSR_58 ( .CLK(clk_bF_buf31), .D(_0b_reg_31_0__25_), .Q(b_reg_25_), .R(reset_n_bF_buf31), .S(1'h1));
DFFSR DFFSR_580 ( .CLK(clk_bF_buf43), .D(w_mem_inst__0w_mem_7__31_0__17_), .Q(w_mem_inst_w_mem_7__17_), .R(reset_n_bF_buf43), .S(1'h1));
DFFSR DFFSR_581 ( .CLK(clk_bF_buf42), .D(w_mem_inst__0w_mem_7__31_0__18_), .Q(w_mem_inst_w_mem_7__18_), .R(reset_n_bF_buf42), .S(1'h1));
DFFSR DFFSR_582 ( .CLK(clk_bF_buf41), .D(w_mem_inst__0w_mem_7__31_0__19_), .Q(w_mem_inst_w_mem_7__19_), .R(reset_n_bF_buf41), .S(1'h1));
DFFSR DFFSR_583 ( .CLK(clk_bF_buf40), .D(w_mem_inst__0w_mem_7__31_0__20_), .Q(w_mem_inst_w_mem_7__20_), .R(reset_n_bF_buf40), .S(1'h1));
DFFSR DFFSR_584 ( .CLK(clk_bF_buf39), .D(w_mem_inst__0w_mem_7__31_0__21_), .Q(w_mem_inst_w_mem_7__21_), .R(reset_n_bF_buf39), .S(1'h1));
DFFSR DFFSR_585 ( .CLK(clk_bF_buf38), .D(w_mem_inst__0w_mem_7__31_0__22_), .Q(w_mem_inst_w_mem_7__22_), .R(reset_n_bF_buf38), .S(1'h1));
DFFSR DFFSR_586 ( .CLK(clk_bF_buf37), .D(w_mem_inst__0w_mem_7__31_0__23_), .Q(w_mem_inst_w_mem_7__23_), .R(reset_n_bF_buf37), .S(1'h1));
DFFSR DFFSR_587 ( .CLK(clk_bF_buf36), .D(w_mem_inst__0w_mem_7__31_0__24_), .Q(w_mem_inst_w_mem_7__24_), .R(reset_n_bF_buf36), .S(1'h1));
DFFSR DFFSR_588 ( .CLK(clk_bF_buf35), .D(w_mem_inst__0w_mem_7__31_0__25_), .Q(w_mem_inst_w_mem_7__25_), .R(reset_n_bF_buf35), .S(1'h1));
DFFSR DFFSR_589 ( .CLK(clk_bF_buf34), .D(w_mem_inst__0w_mem_7__31_0__26_), .Q(w_mem_inst_w_mem_7__26_), .R(reset_n_bF_buf34), .S(1'h1));
DFFSR DFFSR_59 ( .CLK(clk_bF_buf30), .D(_0b_reg_31_0__26_), .Q(b_reg_26_), .R(reset_n_bF_buf30), .S(1'h1));
DFFSR DFFSR_590 ( .CLK(clk_bF_buf33), .D(w_mem_inst__0w_mem_7__31_0__27_), .Q(w_mem_inst_w_mem_7__27_), .R(reset_n_bF_buf33), .S(1'h1));
DFFSR DFFSR_591 ( .CLK(clk_bF_buf32), .D(w_mem_inst__0w_mem_7__31_0__28_), .Q(w_mem_inst_w_mem_7__28_), .R(reset_n_bF_buf32), .S(1'h1));
DFFSR DFFSR_592 ( .CLK(clk_bF_buf31), .D(w_mem_inst__0w_mem_7__31_0__29_), .Q(w_mem_inst_w_mem_7__29_), .R(reset_n_bF_buf31), .S(1'h1));
DFFSR DFFSR_593 ( .CLK(clk_bF_buf30), .D(w_mem_inst__0w_mem_7__31_0__30_), .Q(w_mem_inst_w_mem_7__30_), .R(reset_n_bF_buf30), .S(1'h1));
DFFSR DFFSR_594 ( .CLK(clk_bF_buf29), .D(w_mem_inst__0w_mem_7__31_0__31_), .Q(w_mem_inst_w_mem_7__31_), .R(reset_n_bF_buf29), .S(1'h1));
DFFSR DFFSR_595 ( .CLK(clk_bF_buf28), .D(w_mem_inst__0w_mem_8__31_0__0_), .Q(w_mem_inst_w_mem_8__0_), .R(reset_n_bF_buf28), .S(1'h1));
DFFSR DFFSR_596 ( .CLK(clk_bF_buf27), .D(w_mem_inst__0w_mem_8__31_0__1_), .Q(w_mem_inst_w_mem_8__1_), .R(reset_n_bF_buf27), .S(1'h1));
DFFSR DFFSR_597 ( .CLK(clk_bF_buf26), .D(w_mem_inst__0w_mem_8__31_0__2_), .Q(w_mem_inst_w_mem_8__2_), .R(reset_n_bF_buf26), .S(1'h1));
DFFSR DFFSR_598 ( .CLK(clk_bF_buf25), .D(w_mem_inst__0w_mem_8__31_0__3_), .Q(w_mem_inst_w_mem_8__3_), .R(reset_n_bF_buf25), .S(1'h1));
DFFSR DFFSR_599 ( .CLK(clk_bF_buf24), .D(w_mem_inst__0w_mem_8__31_0__4_), .Q(w_mem_inst_w_mem_8__4_), .R(reset_n_bF_buf24), .S(1'h1));
DFFSR DFFSR_6 ( .CLK(clk_bF_buf83), .D(_0a_reg_31_0__5_), .Q(a_reg_5_), .R(reset_n_bF_buf83), .S(1'h1));
DFFSR DFFSR_60 ( .CLK(clk_bF_buf29), .D(_0b_reg_31_0__27_), .Q(b_reg_27_), .R(reset_n_bF_buf29), .S(1'h1));
DFFSR DFFSR_600 ( .CLK(clk_bF_buf23), .D(w_mem_inst__0w_mem_8__31_0__5_), .Q(w_mem_inst_w_mem_8__5_), .R(reset_n_bF_buf23), .S(1'h1));
DFFSR DFFSR_601 ( .CLK(clk_bF_buf22), .D(w_mem_inst__0w_mem_8__31_0__6_), .Q(w_mem_inst_w_mem_8__6_), .R(reset_n_bF_buf22), .S(1'h1));
DFFSR DFFSR_602 ( .CLK(clk_bF_buf21), .D(w_mem_inst__0w_mem_8__31_0__7_), .Q(w_mem_inst_w_mem_8__7_), .R(reset_n_bF_buf21), .S(1'h1));
DFFSR DFFSR_603 ( .CLK(clk_bF_buf20), .D(w_mem_inst__0w_mem_8__31_0__8_), .Q(w_mem_inst_w_mem_8__8_), .R(reset_n_bF_buf20), .S(1'h1));
DFFSR DFFSR_604 ( .CLK(clk_bF_buf19), .D(w_mem_inst__0w_mem_8__31_0__9_), .Q(w_mem_inst_w_mem_8__9_), .R(reset_n_bF_buf19), .S(1'h1));
DFFSR DFFSR_605 ( .CLK(clk_bF_buf18), .D(w_mem_inst__0w_mem_8__31_0__10_), .Q(w_mem_inst_w_mem_8__10_), .R(reset_n_bF_buf18), .S(1'h1));
DFFSR DFFSR_606 ( .CLK(clk_bF_buf17), .D(w_mem_inst__0w_mem_8__31_0__11_), .Q(w_mem_inst_w_mem_8__11_), .R(reset_n_bF_buf17), .S(1'h1));
DFFSR DFFSR_607 ( .CLK(clk_bF_buf16), .D(w_mem_inst__0w_mem_8__31_0__12_), .Q(w_mem_inst_w_mem_8__12_), .R(reset_n_bF_buf16), .S(1'h1));
DFFSR DFFSR_608 ( .CLK(clk_bF_buf15), .D(w_mem_inst__0w_mem_8__31_0__13_), .Q(w_mem_inst_w_mem_8__13_), .R(reset_n_bF_buf15), .S(1'h1));
DFFSR DFFSR_609 ( .CLK(clk_bF_buf14), .D(w_mem_inst__0w_mem_8__31_0__14_), .Q(w_mem_inst_w_mem_8__14_), .R(reset_n_bF_buf14), .S(1'h1));
DFFSR DFFSR_61 ( .CLK(clk_bF_buf28), .D(_0b_reg_31_0__28_), .Q(b_reg_28_), .R(reset_n_bF_buf28), .S(1'h1));
DFFSR DFFSR_610 ( .CLK(clk_bF_buf13), .D(w_mem_inst__0w_mem_8__31_0__15_), .Q(w_mem_inst_w_mem_8__15_), .R(reset_n_bF_buf13), .S(1'h1));
DFFSR DFFSR_611 ( .CLK(clk_bF_buf12), .D(w_mem_inst__0w_mem_8__31_0__16_), .Q(w_mem_inst_w_mem_8__16_), .R(reset_n_bF_buf12), .S(1'h1));
DFFSR DFFSR_612 ( .CLK(clk_bF_buf11), .D(w_mem_inst__0w_mem_8__31_0__17_), .Q(w_mem_inst_w_mem_8__17_), .R(reset_n_bF_buf11), .S(1'h1));
DFFSR DFFSR_613 ( .CLK(clk_bF_buf10), .D(w_mem_inst__0w_mem_8__31_0__18_), .Q(w_mem_inst_w_mem_8__18_), .R(reset_n_bF_buf10), .S(1'h1));
DFFSR DFFSR_614 ( .CLK(clk_bF_buf9), .D(w_mem_inst__0w_mem_8__31_0__19_), .Q(w_mem_inst_w_mem_8__19_), .R(reset_n_bF_buf9), .S(1'h1));
DFFSR DFFSR_615 ( .CLK(clk_bF_buf8), .D(w_mem_inst__0w_mem_8__31_0__20_), .Q(w_mem_inst_w_mem_8__20_), .R(reset_n_bF_buf8), .S(1'h1));
DFFSR DFFSR_616 ( .CLK(clk_bF_buf7), .D(w_mem_inst__0w_mem_8__31_0__21_), .Q(w_mem_inst_w_mem_8__21_), .R(reset_n_bF_buf7), .S(1'h1));
DFFSR DFFSR_617 ( .CLK(clk_bF_buf6), .D(w_mem_inst__0w_mem_8__31_0__22_), .Q(w_mem_inst_w_mem_8__22_), .R(reset_n_bF_buf6), .S(1'h1));
DFFSR DFFSR_618 ( .CLK(clk_bF_buf5), .D(w_mem_inst__0w_mem_8__31_0__23_), .Q(w_mem_inst_w_mem_8__23_), .R(reset_n_bF_buf5), .S(1'h1));
DFFSR DFFSR_619 ( .CLK(clk_bF_buf4), .D(w_mem_inst__0w_mem_8__31_0__24_), .Q(w_mem_inst_w_mem_8__24_), .R(reset_n_bF_buf4), .S(1'h1));
DFFSR DFFSR_62 ( .CLK(clk_bF_buf27), .D(_0b_reg_31_0__29_), .Q(b_reg_29_), .R(reset_n_bF_buf27), .S(1'h1));
DFFSR DFFSR_620 ( .CLK(clk_bF_buf3), .D(w_mem_inst__0w_mem_8__31_0__25_), .Q(w_mem_inst_w_mem_8__25_), .R(reset_n_bF_buf3), .S(1'h1));
DFFSR DFFSR_621 ( .CLK(clk_bF_buf2), .D(w_mem_inst__0w_mem_8__31_0__26_), .Q(w_mem_inst_w_mem_8__26_), .R(reset_n_bF_buf2), .S(1'h1));
DFFSR DFFSR_622 ( .CLK(clk_bF_buf1), .D(w_mem_inst__0w_mem_8__31_0__27_), .Q(w_mem_inst_w_mem_8__27_), .R(reset_n_bF_buf1), .S(1'h1));
DFFSR DFFSR_623 ( .CLK(clk_bF_buf0), .D(w_mem_inst__0w_mem_8__31_0__28_), .Q(w_mem_inst_w_mem_8__28_), .R(reset_n_bF_buf0), .S(1'h1));
DFFSR DFFSR_624 ( .CLK(clk_bF_buf88), .D(w_mem_inst__0w_mem_8__31_0__29_), .Q(w_mem_inst_w_mem_8__29_), .R(reset_n_bF_buf88), .S(1'h1));
DFFSR DFFSR_625 ( .CLK(clk_bF_buf87), .D(w_mem_inst__0w_mem_8__31_0__30_), .Q(w_mem_inst_w_mem_8__30_), .R(reset_n_bF_buf87), .S(1'h1));
DFFSR DFFSR_626 ( .CLK(clk_bF_buf86), .D(w_mem_inst__0w_mem_8__31_0__31_), .Q(w_mem_inst_w_mem_8__31_), .R(reset_n_bF_buf86), .S(1'h1));
DFFSR DFFSR_627 ( .CLK(clk_bF_buf85), .D(w_mem_inst__0w_mem_9__31_0__0_), .Q(w_mem_inst_w_mem_9__0_), .R(reset_n_bF_buf85), .S(1'h1));
DFFSR DFFSR_628 ( .CLK(clk_bF_buf84), .D(w_mem_inst__0w_mem_9__31_0__1_), .Q(w_mem_inst_w_mem_9__1_), .R(reset_n_bF_buf84), .S(1'h1));
DFFSR DFFSR_629 ( .CLK(clk_bF_buf83), .D(w_mem_inst__0w_mem_9__31_0__2_), .Q(w_mem_inst_w_mem_9__2_), .R(reset_n_bF_buf83), .S(1'h1));
DFFSR DFFSR_63 ( .CLK(clk_bF_buf26), .D(_0b_reg_31_0__30_), .Q(b_reg_30_), .R(reset_n_bF_buf26), .S(1'h1));
DFFSR DFFSR_630 ( .CLK(clk_bF_buf82), .D(w_mem_inst__0w_mem_9__31_0__3_), .Q(w_mem_inst_w_mem_9__3_), .R(reset_n_bF_buf82), .S(1'h1));
DFFSR DFFSR_631 ( .CLK(clk_bF_buf81), .D(w_mem_inst__0w_mem_9__31_0__4_), .Q(w_mem_inst_w_mem_9__4_), .R(reset_n_bF_buf81), .S(1'h1));
DFFSR DFFSR_632 ( .CLK(clk_bF_buf80), .D(w_mem_inst__0w_mem_9__31_0__5_), .Q(w_mem_inst_w_mem_9__5_), .R(reset_n_bF_buf80), .S(1'h1));
DFFSR DFFSR_633 ( .CLK(clk_bF_buf79), .D(w_mem_inst__0w_mem_9__31_0__6_), .Q(w_mem_inst_w_mem_9__6_), .R(reset_n_bF_buf79), .S(1'h1));
DFFSR DFFSR_634 ( .CLK(clk_bF_buf78), .D(w_mem_inst__0w_mem_9__31_0__7_), .Q(w_mem_inst_w_mem_9__7_), .R(reset_n_bF_buf78), .S(1'h1));
DFFSR DFFSR_635 ( .CLK(clk_bF_buf77), .D(w_mem_inst__0w_mem_9__31_0__8_), .Q(w_mem_inst_w_mem_9__8_), .R(reset_n_bF_buf77), .S(1'h1));
DFFSR DFFSR_636 ( .CLK(clk_bF_buf76), .D(w_mem_inst__0w_mem_9__31_0__9_), .Q(w_mem_inst_w_mem_9__9_), .R(reset_n_bF_buf76), .S(1'h1));
DFFSR DFFSR_637 ( .CLK(clk_bF_buf75), .D(w_mem_inst__0w_mem_9__31_0__10_), .Q(w_mem_inst_w_mem_9__10_), .R(reset_n_bF_buf75), .S(1'h1));
DFFSR DFFSR_638 ( .CLK(clk_bF_buf74), .D(w_mem_inst__0w_mem_9__31_0__11_), .Q(w_mem_inst_w_mem_9__11_), .R(reset_n_bF_buf74), .S(1'h1));
DFFSR DFFSR_639 ( .CLK(clk_bF_buf73), .D(w_mem_inst__0w_mem_9__31_0__12_), .Q(w_mem_inst_w_mem_9__12_), .R(reset_n_bF_buf73), .S(1'h1));
DFFSR DFFSR_64 ( .CLK(clk_bF_buf25), .D(_0b_reg_31_0__31_), .Q(b_reg_31_), .R(reset_n_bF_buf25), .S(1'h1));
DFFSR DFFSR_640 ( .CLK(clk_bF_buf72), .D(w_mem_inst__0w_mem_9__31_0__13_), .Q(w_mem_inst_w_mem_9__13_), .R(reset_n_bF_buf72), .S(1'h1));
DFFSR DFFSR_641 ( .CLK(clk_bF_buf71), .D(w_mem_inst__0w_mem_9__31_0__14_), .Q(w_mem_inst_w_mem_9__14_), .R(reset_n_bF_buf71), .S(1'h1));
DFFSR DFFSR_642 ( .CLK(clk_bF_buf70), .D(w_mem_inst__0w_mem_9__31_0__15_), .Q(w_mem_inst_w_mem_9__15_), .R(reset_n_bF_buf70), .S(1'h1));
DFFSR DFFSR_643 ( .CLK(clk_bF_buf69), .D(w_mem_inst__0w_mem_9__31_0__16_), .Q(w_mem_inst_w_mem_9__16_), .R(reset_n_bF_buf69), .S(1'h1));
DFFSR DFFSR_644 ( .CLK(clk_bF_buf68), .D(w_mem_inst__0w_mem_9__31_0__17_), .Q(w_mem_inst_w_mem_9__17_), .R(reset_n_bF_buf68), .S(1'h1));
DFFSR DFFSR_645 ( .CLK(clk_bF_buf67), .D(w_mem_inst__0w_mem_9__31_0__18_), .Q(w_mem_inst_w_mem_9__18_), .R(reset_n_bF_buf67), .S(1'h1));
DFFSR DFFSR_646 ( .CLK(clk_bF_buf66), .D(w_mem_inst__0w_mem_9__31_0__19_), .Q(w_mem_inst_w_mem_9__19_), .R(reset_n_bF_buf66), .S(1'h1));
DFFSR DFFSR_647 ( .CLK(clk_bF_buf65), .D(w_mem_inst__0w_mem_9__31_0__20_), .Q(w_mem_inst_w_mem_9__20_), .R(reset_n_bF_buf65), .S(1'h1));
DFFSR DFFSR_648 ( .CLK(clk_bF_buf64), .D(w_mem_inst__0w_mem_9__31_0__21_), .Q(w_mem_inst_w_mem_9__21_), .R(reset_n_bF_buf64), .S(1'h1));
DFFSR DFFSR_649 ( .CLK(clk_bF_buf63), .D(w_mem_inst__0w_mem_9__31_0__22_), .Q(w_mem_inst_w_mem_9__22_), .R(reset_n_bF_buf63), .S(1'h1));
DFFSR DFFSR_65 ( .CLK(clk_bF_buf24), .D(_0c_reg_31_0__0_), .Q(c_reg_0_), .R(reset_n_bF_buf24), .S(1'h1));
DFFSR DFFSR_650 ( .CLK(clk_bF_buf62), .D(w_mem_inst__0w_mem_9__31_0__23_), .Q(w_mem_inst_w_mem_9__23_), .R(reset_n_bF_buf62), .S(1'h1));
DFFSR DFFSR_651 ( .CLK(clk_bF_buf61), .D(w_mem_inst__0w_mem_9__31_0__24_), .Q(w_mem_inst_w_mem_9__24_), .R(reset_n_bF_buf61), .S(1'h1));
DFFSR DFFSR_652 ( .CLK(clk_bF_buf60), .D(w_mem_inst__0w_mem_9__31_0__25_), .Q(w_mem_inst_w_mem_9__25_), .R(reset_n_bF_buf60), .S(1'h1));
DFFSR DFFSR_653 ( .CLK(clk_bF_buf59), .D(w_mem_inst__0w_mem_9__31_0__26_), .Q(w_mem_inst_w_mem_9__26_), .R(reset_n_bF_buf59), .S(1'h1));
DFFSR DFFSR_654 ( .CLK(clk_bF_buf58), .D(w_mem_inst__0w_mem_9__31_0__27_), .Q(w_mem_inst_w_mem_9__27_), .R(reset_n_bF_buf58), .S(1'h1));
DFFSR DFFSR_655 ( .CLK(clk_bF_buf57), .D(w_mem_inst__0w_mem_9__31_0__28_), .Q(w_mem_inst_w_mem_9__28_), .R(reset_n_bF_buf57), .S(1'h1));
DFFSR DFFSR_656 ( .CLK(clk_bF_buf56), .D(w_mem_inst__0w_mem_9__31_0__29_), .Q(w_mem_inst_w_mem_9__29_), .R(reset_n_bF_buf56), .S(1'h1));
DFFSR DFFSR_657 ( .CLK(clk_bF_buf55), .D(w_mem_inst__0w_mem_9__31_0__30_), .Q(w_mem_inst_w_mem_9__30_), .R(reset_n_bF_buf55), .S(1'h1));
DFFSR DFFSR_658 ( .CLK(clk_bF_buf54), .D(w_mem_inst__0w_mem_9__31_0__31_), .Q(w_mem_inst_w_mem_9__31_), .R(reset_n_bF_buf54), .S(1'h1));
DFFSR DFFSR_659 ( .CLK(clk_bF_buf53), .D(w_mem_inst__0w_mem_10__31_0__0_), .Q(w_mem_inst_w_mem_10__0_), .R(reset_n_bF_buf53), .S(1'h1));
DFFSR DFFSR_66 ( .CLK(clk_bF_buf23), .D(_0c_reg_31_0__1_), .Q(c_reg_1_), .R(reset_n_bF_buf23), .S(1'h1));
DFFSR DFFSR_660 ( .CLK(clk_bF_buf52), .D(w_mem_inst__0w_mem_10__31_0__1_), .Q(w_mem_inst_w_mem_10__1_), .R(reset_n_bF_buf52), .S(1'h1));
DFFSR DFFSR_661 ( .CLK(clk_bF_buf51), .D(w_mem_inst__0w_mem_10__31_0__2_), .Q(w_mem_inst_w_mem_10__2_), .R(reset_n_bF_buf51), .S(1'h1));
DFFSR DFFSR_662 ( .CLK(clk_bF_buf50), .D(w_mem_inst__0w_mem_10__31_0__3_), .Q(w_mem_inst_w_mem_10__3_), .R(reset_n_bF_buf50), .S(1'h1));
DFFSR DFFSR_663 ( .CLK(clk_bF_buf49), .D(w_mem_inst__0w_mem_10__31_0__4_), .Q(w_mem_inst_w_mem_10__4_), .R(reset_n_bF_buf49), .S(1'h1));
DFFSR DFFSR_664 ( .CLK(clk_bF_buf48), .D(w_mem_inst__0w_mem_10__31_0__5_), .Q(w_mem_inst_w_mem_10__5_), .R(reset_n_bF_buf48), .S(1'h1));
DFFSR DFFSR_665 ( .CLK(clk_bF_buf47), .D(w_mem_inst__0w_mem_10__31_0__6_), .Q(w_mem_inst_w_mem_10__6_), .R(reset_n_bF_buf47), .S(1'h1));
DFFSR DFFSR_666 ( .CLK(clk_bF_buf46), .D(w_mem_inst__0w_mem_10__31_0__7_), .Q(w_mem_inst_w_mem_10__7_), .R(reset_n_bF_buf46), .S(1'h1));
DFFSR DFFSR_667 ( .CLK(clk_bF_buf45), .D(w_mem_inst__0w_mem_10__31_0__8_), .Q(w_mem_inst_w_mem_10__8_), .R(reset_n_bF_buf45), .S(1'h1));
DFFSR DFFSR_668 ( .CLK(clk_bF_buf44), .D(w_mem_inst__0w_mem_10__31_0__9_), .Q(w_mem_inst_w_mem_10__9_), .R(reset_n_bF_buf44), .S(1'h1));
DFFSR DFFSR_669 ( .CLK(clk_bF_buf43), .D(w_mem_inst__0w_mem_10__31_0__10_), .Q(w_mem_inst_w_mem_10__10_), .R(reset_n_bF_buf43), .S(1'h1));
DFFSR DFFSR_67 ( .CLK(clk_bF_buf22), .D(_0c_reg_31_0__2_), .Q(c_reg_2_), .R(reset_n_bF_buf22), .S(1'h1));
DFFSR DFFSR_670 ( .CLK(clk_bF_buf42), .D(w_mem_inst__0w_mem_10__31_0__11_), .Q(w_mem_inst_w_mem_10__11_), .R(reset_n_bF_buf42), .S(1'h1));
DFFSR DFFSR_671 ( .CLK(clk_bF_buf41), .D(w_mem_inst__0w_mem_10__31_0__12_), .Q(w_mem_inst_w_mem_10__12_), .R(reset_n_bF_buf41), .S(1'h1));
DFFSR DFFSR_672 ( .CLK(clk_bF_buf40), .D(w_mem_inst__0w_mem_10__31_0__13_), .Q(w_mem_inst_w_mem_10__13_), .R(reset_n_bF_buf40), .S(1'h1));
DFFSR DFFSR_673 ( .CLK(clk_bF_buf39), .D(w_mem_inst__0w_mem_10__31_0__14_), .Q(w_mem_inst_w_mem_10__14_), .R(reset_n_bF_buf39), .S(1'h1));
DFFSR DFFSR_674 ( .CLK(clk_bF_buf38), .D(w_mem_inst__0w_mem_10__31_0__15_), .Q(w_mem_inst_w_mem_10__15_), .R(reset_n_bF_buf38), .S(1'h1));
DFFSR DFFSR_675 ( .CLK(clk_bF_buf37), .D(w_mem_inst__0w_mem_10__31_0__16_), .Q(w_mem_inst_w_mem_10__16_), .R(reset_n_bF_buf37), .S(1'h1));
DFFSR DFFSR_676 ( .CLK(clk_bF_buf36), .D(w_mem_inst__0w_mem_10__31_0__17_), .Q(w_mem_inst_w_mem_10__17_), .R(reset_n_bF_buf36), .S(1'h1));
DFFSR DFFSR_677 ( .CLK(clk_bF_buf35), .D(w_mem_inst__0w_mem_10__31_0__18_), .Q(w_mem_inst_w_mem_10__18_), .R(reset_n_bF_buf35), .S(1'h1));
DFFSR DFFSR_678 ( .CLK(clk_bF_buf34), .D(w_mem_inst__0w_mem_10__31_0__19_), .Q(w_mem_inst_w_mem_10__19_), .R(reset_n_bF_buf34), .S(1'h1));
DFFSR DFFSR_679 ( .CLK(clk_bF_buf33), .D(w_mem_inst__0w_mem_10__31_0__20_), .Q(w_mem_inst_w_mem_10__20_), .R(reset_n_bF_buf33), .S(1'h1));
DFFSR DFFSR_68 ( .CLK(clk_bF_buf21), .D(_0c_reg_31_0__3_), .Q(c_reg_3_), .R(reset_n_bF_buf21), .S(1'h1));
DFFSR DFFSR_680 ( .CLK(clk_bF_buf32), .D(w_mem_inst__0w_mem_10__31_0__21_), .Q(w_mem_inst_w_mem_10__21_), .R(reset_n_bF_buf32), .S(1'h1));
DFFSR DFFSR_681 ( .CLK(clk_bF_buf31), .D(w_mem_inst__0w_mem_10__31_0__22_), .Q(w_mem_inst_w_mem_10__22_), .R(reset_n_bF_buf31), .S(1'h1));
DFFSR DFFSR_682 ( .CLK(clk_bF_buf30), .D(w_mem_inst__0w_mem_10__31_0__23_), .Q(w_mem_inst_w_mem_10__23_), .R(reset_n_bF_buf30), .S(1'h1));
DFFSR DFFSR_683 ( .CLK(clk_bF_buf29), .D(w_mem_inst__0w_mem_10__31_0__24_), .Q(w_mem_inst_w_mem_10__24_), .R(reset_n_bF_buf29), .S(1'h1));
DFFSR DFFSR_684 ( .CLK(clk_bF_buf28), .D(w_mem_inst__0w_mem_10__31_0__25_), .Q(w_mem_inst_w_mem_10__25_), .R(reset_n_bF_buf28), .S(1'h1));
DFFSR DFFSR_685 ( .CLK(clk_bF_buf27), .D(w_mem_inst__0w_mem_10__31_0__26_), .Q(w_mem_inst_w_mem_10__26_), .R(reset_n_bF_buf27), .S(1'h1));
DFFSR DFFSR_686 ( .CLK(clk_bF_buf26), .D(w_mem_inst__0w_mem_10__31_0__27_), .Q(w_mem_inst_w_mem_10__27_), .R(reset_n_bF_buf26), .S(1'h1));
DFFSR DFFSR_687 ( .CLK(clk_bF_buf25), .D(w_mem_inst__0w_mem_10__31_0__28_), .Q(w_mem_inst_w_mem_10__28_), .R(reset_n_bF_buf25), .S(1'h1));
DFFSR DFFSR_688 ( .CLK(clk_bF_buf24), .D(w_mem_inst__0w_mem_10__31_0__29_), .Q(w_mem_inst_w_mem_10__29_), .R(reset_n_bF_buf24), .S(1'h1));
DFFSR DFFSR_689 ( .CLK(clk_bF_buf23), .D(w_mem_inst__0w_mem_10__31_0__30_), .Q(w_mem_inst_w_mem_10__30_), .R(reset_n_bF_buf23), .S(1'h1));
DFFSR DFFSR_69 ( .CLK(clk_bF_buf20), .D(_0c_reg_31_0__4_), .Q(c_reg_4_), .R(reset_n_bF_buf20), .S(1'h1));
DFFSR DFFSR_690 ( .CLK(clk_bF_buf22), .D(w_mem_inst__0w_mem_10__31_0__31_), .Q(w_mem_inst_w_mem_10__31_), .R(reset_n_bF_buf22), .S(1'h1));
DFFSR DFFSR_691 ( .CLK(clk_bF_buf21), .D(w_mem_inst__0w_mem_11__31_0__0_), .Q(w_mem_inst_w_mem_11__0_), .R(reset_n_bF_buf21), .S(1'h1));
DFFSR DFFSR_692 ( .CLK(clk_bF_buf20), .D(w_mem_inst__0w_mem_11__31_0__1_), .Q(w_mem_inst_w_mem_11__1_), .R(reset_n_bF_buf20), .S(1'h1));
DFFSR DFFSR_693 ( .CLK(clk_bF_buf19), .D(w_mem_inst__0w_mem_11__31_0__2_), .Q(w_mem_inst_w_mem_11__2_), .R(reset_n_bF_buf19), .S(1'h1));
DFFSR DFFSR_694 ( .CLK(clk_bF_buf18), .D(w_mem_inst__0w_mem_11__31_0__3_), .Q(w_mem_inst_w_mem_11__3_), .R(reset_n_bF_buf18), .S(1'h1));
DFFSR DFFSR_695 ( .CLK(clk_bF_buf17), .D(w_mem_inst__0w_mem_11__31_0__4_), .Q(w_mem_inst_w_mem_11__4_), .R(reset_n_bF_buf17), .S(1'h1));
DFFSR DFFSR_696 ( .CLK(clk_bF_buf16), .D(w_mem_inst__0w_mem_11__31_0__5_), .Q(w_mem_inst_w_mem_11__5_), .R(reset_n_bF_buf16), .S(1'h1));
DFFSR DFFSR_697 ( .CLK(clk_bF_buf15), .D(w_mem_inst__0w_mem_11__31_0__6_), .Q(w_mem_inst_w_mem_11__6_), .R(reset_n_bF_buf15), .S(1'h1));
DFFSR DFFSR_698 ( .CLK(clk_bF_buf14), .D(w_mem_inst__0w_mem_11__31_0__7_), .Q(w_mem_inst_w_mem_11__7_), .R(reset_n_bF_buf14), .S(1'h1));
DFFSR DFFSR_699 ( .CLK(clk_bF_buf13), .D(w_mem_inst__0w_mem_11__31_0__8_), .Q(w_mem_inst_w_mem_11__8_), .R(reset_n_bF_buf13), .S(1'h1));
DFFSR DFFSR_7 ( .CLK(clk_bF_buf82), .D(_0a_reg_31_0__6_), .Q(a_reg_6_), .R(reset_n_bF_buf82), .S(1'h1));
DFFSR DFFSR_70 ( .CLK(clk_bF_buf19), .D(_0c_reg_31_0__5_), .Q(c_reg_5_), .R(reset_n_bF_buf19), .S(1'h1));
DFFSR DFFSR_700 ( .CLK(clk_bF_buf12), .D(w_mem_inst__0w_mem_11__31_0__9_), .Q(w_mem_inst_w_mem_11__9_), .R(reset_n_bF_buf12), .S(1'h1));
DFFSR DFFSR_701 ( .CLK(clk_bF_buf11), .D(w_mem_inst__0w_mem_11__31_0__10_), .Q(w_mem_inst_w_mem_11__10_), .R(reset_n_bF_buf11), .S(1'h1));
DFFSR DFFSR_702 ( .CLK(clk_bF_buf10), .D(w_mem_inst__0w_mem_11__31_0__11_), .Q(w_mem_inst_w_mem_11__11_), .R(reset_n_bF_buf10), .S(1'h1));
DFFSR DFFSR_703 ( .CLK(clk_bF_buf9), .D(w_mem_inst__0w_mem_11__31_0__12_), .Q(w_mem_inst_w_mem_11__12_), .R(reset_n_bF_buf9), .S(1'h1));
DFFSR DFFSR_704 ( .CLK(clk_bF_buf8), .D(w_mem_inst__0w_mem_11__31_0__13_), .Q(w_mem_inst_w_mem_11__13_), .R(reset_n_bF_buf8), .S(1'h1));
DFFSR DFFSR_705 ( .CLK(clk_bF_buf7), .D(w_mem_inst__0w_mem_11__31_0__14_), .Q(w_mem_inst_w_mem_11__14_), .R(reset_n_bF_buf7), .S(1'h1));
DFFSR DFFSR_706 ( .CLK(clk_bF_buf6), .D(w_mem_inst__0w_mem_11__31_0__15_), .Q(w_mem_inst_w_mem_11__15_), .R(reset_n_bF_buf6), .S(1'h1));
DFFSR DFFSR_707 ( .CLK(clk_bF_buf5), .D(w_mem_inst__0w_mem_11__31_0__16_), .Q(w_mem_inst_w_mem_11__16_), .R(reset_n_bF_buf5), .S(1'h1));
DFFSR DFFSR_708 ( .CLK(clk_bF_buf4), .D(w_mem_inst__0w_mem_11__31_0__17_), .Q(w_mem_inst_w_mem_11__17_), .R(reset_n_bF_buf4), .S(1'h1));
DFFSR DFFSR_709 ( .CLK(clk_bF_buf3), .D(w_mem_inst__0w_mem_11__31_0__18_), .Q(w_mem_inst_w_mem_11__18_), .R(reset_n_bF_buf3), .S(1'h1));
DFFSR DFFSR_71 ( .CLK(clk_bF_buf18), .D(_0c_reg_31_0__6_), .Q(c_reg_6_), .R(reset_n_bF_buf18), .S(1'h1));
DFFSR DFFSR_710 ( .CLK(clk_bF_buf2), .D(w_mem_inst__0w_mem_11__31_0__19_), .Q(w_mem_inst_w_mem_11__19_), .R(reset_n_bF_buf2), .S(1'h1));
DFFSR DFFSR_711 ( .CLK(clk_bF_buf1), .D(w_mem_inst__0w_mem_11__31_0__20_), .Q(w_mem_inst_w_mem_11__20_), .R(reset_n_bF_buf1), .S(1'h1));
DFFSR DFFSR_712 ( .CLK(clk_bF_buf0), .D(w_mem_inst__0w_mem_11__31_0__21_), .Q(w_mem_inst_w_mem_11__21_), .R(reset_n_bF_buf0), .S(1'h1));
DFFSR DFFSR_713 ( .CLK(clk_bF_buf88), .D(w_mem_inst__0w_mem_11__31_0__22_), .Q(w_mem_inst_w_mem_11__22_), .R(reset_n_bF_buf88), .S(1'h1));
DFFSR DFFSR_714 ( .CLK(clk_bF_buf87), .D(w_mem_inst__0w_mem_11__31_0__23_), .Q(w_mem_inst_w_mem_11__23_), .R(reset_n_bF_buf87), .S(1'h1));
DFFSR DFFSR_715 ( .CLK(clk_bF_buf86), .D(w_mem_inst__0w_mem_11__31_0__24_), .Q(w_mem_inst_w_mem_11__24_), .R(reset_n_bF_buf86), .S(1'h1));
DFFSR DFFSR_716 ( .CLK(clk_bF_buf85), .D(w_mem_inst__0w_mem_11__31_0__25_), .Q(w_mem_inst_w_mem_11__25_), .R(reset_n_bF_buf85), .S(1'h1));
DFFSR DFFSR_717 ( .CLK(clk_bF_buf84), .D(w_mem_inst__0w_mem_11__31_0__26_), .Q(w_mem_inst_w_mem_11__26_), .R(reset_n_bF_buf84), .S(1'h1));
DFFSR DFFSR_718 ( .CLK(clk_bF_buf83), .D(w_mem_inst__0w_mem_11__31_0__27_), .Q(w_mem_inst_w_mem_11__27_), .R(reset_n_bF_buf83), .S(1'h1));
DFFSR DFFSR_719 ( .CLK(clk_bF_buf82), .D(w_mem_inst__0w_mem_11__31_0__28_), .Q(w_mem_inst_w_mem_11__28_), .R(reset_n_bF_buf82), .S(1'h1));
DFFSR DFFSR_72 ( .CLK(clk_bF_buf17), .D(_0c_reg_31_0__7_), .Q(c_reg_7_), .R(reset_n_bF_buf17), .S(1'h1));
DFFSR DFFSR_720 ( .CLK(clk_bF_buf81), .D(w_mem_inst__0w_mem_11__31_0__29_), .Q(w_mem_inst_w_mem_11__29_), .R(reset_n_bF_buf81), .S(1'h1));
DFFSR DFFSR_721 ( .CLK(clk_bF_buf80), .D(w_mem_inst__0w_mem_11__31_0__30_), .Q(w_mem_inst_w_mem_11__30_), .R(reset_n_bF_buf80), .S(1'h1));
DFFSR DFFSR_722 ( .CLK(clk_bF_buf79), .D(w_mem_inst__0w_mem_11__31_0__31_), .Q(w_mem_inst_w_mem_11__31_), .R(reset_n_bF_buf79), .S(1'h1));
DFFSR DFFSR_723 ( .CLK(clk_bF_buf78), .D(w_mem_inst__0w_mem_12__31_0__0_), .Q(w_mem_inst_w_mem_12__0_), .R(reset_n_bF_buf78), .S(1'h1));
DFFSR DFFSR_724 ( .CLK(clk_bF_buf77), .D(w_mem_inst__0w_mem_12__31_0__1_), .Q(w_mem_inst_w_mem_12__1_), .R(reset_n_bF_buf77), .S(1'h1));
DFFSR DFFSR_725 ( .CLK(clk_bF_buf76), .D(w_mem_inst__0w_mem_12__31_0__2_), .Q(w_mem_inst_w_mem_12__2_), .R(reset_n_bF_buf76), .S(1'h1));
DFFSR DFFSR_726 ( .CLK(clk_bF_buf75), .D(w_mem_inst__0w_mem_12__31_0__3_), .Q(w_mem_inst_w_mem_12__3_), .R(reset_n_bF_buf75), .S(1'h1));
DFFSR DFFSR_727 ( .CLK(clk_bF_buf74), .D(w_mem_inst__0w_mem_12__31_0__4_), .Q(w_mem_inst_w_mem_12__4_), .R(reset_n_bF_buf74), .S(1'h1));
DFFSR DFFSR_728 ( .CLK(clk_bF_buf73), .D(w_mem_inst__0w_mem_12__31_0__5_), .Q(w_mem_inst_w_mem_12__5_), .R(reset_n_bF_buf73), .S(1'h1));
DFFSR DFFSR_729 ( .CLK(clk_bF_buf72), .D(w_mem_inst__0w_mem_12__31_0__6_), .Q(w_mem_inst_w_mem_12__6_), .R(reset_n_bF_buf72), .S(1'h1));
DFFSR DFFSR_73 ( .CLK(clk_bF_buf16), .D(_0c_reg_31_0__8_), .Q(c_reg_8_), .R(reset_n_bF_buf16), .S(1'h1));
DFFSR DFFSR_730 ( .CLK(clk_bF_buf71), .D(w_mem_inst__0w_mem_12__31_0__7_), .Q(w_mem_inst_w_mem_12__7_), .R(reset_n_bF_buf71), .S(1'h1));
DFFSR DFFSR_731 ( .CLK(clk_bF_buf70), .D(w_mem_inst__0w_mem_12__31_0__8_), .Q(w_mem_inst_w_mem_12__8_), .R(reset_n_bF_buf70), .S(1'h1));
DFFSR DFFSR_732 ( .CLK(clk_bF_buf69), .D(w_mem_inst__0w_mem_12__31_0__9_), .Q(w_mem_inst_w_mem_12__9_), .R(reset_n_bF_buf69), .S(1'h1));
DFFSR DFFSR_733 ( .CLK(clk_bF_buf68), .D(w_mem_inst__0w_mem_12__31_0__10_), .Q(w_mem_inst_w_mem_12__10_), .R(reset_n_bF_buf68), .S(1'h1));
DFFSR DFFSR_734 ( .CLK(clk_bF_buf67), .D(w_mem_inst__0w_mem_12__31_0__11_), .Q(w_mem_inst_w_mem_12__11_), .R(reset_n_bF_buf67), .S(1'h1));
DFFSR DFFSR_735 ( .CLK(clk_bF_buf66), .D(w_mem_inst__0w_mem_12__31_0__12_), .Q(w_mem_inst_w_mem_12__12_), .R(reset_n_bF_buf66), .S(1'h1));
DFFSR DFFSR_736 ( .CLK(clk_bF_buf65), .D(w_mem_inst__0w_mem_12__31_0__13_), .Q(w_mem_inst_w_mem_12__13_), .R(reset_n_bF_buf65), .S(1'h1));
DFFSR DFFSR_737 ( .CLK(clk_bF_buf64), .D(w_mem_inst__0w_mem_12__31_0__14_), .Q(w_mem_inst_w_mem_12__14_), .R(reset_n_bF_buf64), .S(1'h1));
DFFSR DFFSR_738 ( .CLK(clk_bF_buf63), .D(w_mem_inst__0w_mem_12__31_0__15_), .Q(w_mem_inst_w_mem_12__15_), .R(reset_n_bF_buf63), .S(1'h1));
DFFSR DFFSR_739 ( .CLK(clk_bF_buf62), .D(w_mem_inst__0w_mem_12__31_0__16_), .Q(w_mem_inst_w_mem_12__16_), .R(reset_n_bF_buf62), .S(1'h1));
DFFSR DFFSR_74 ( .CLK(clk_bF_buf15), .D(_0c_reg_31_0__9_), .Q(c_reg_9_), .R(reset_n_bF_buf15), .S(1'h1));
DFFSR DFFSR_740 ( .CLK(clk_bF_buf61), .D(w_mem_inst__0w_mem_12__31_0__17_), .Q(w_mem_inst_w_mem_12__17_), .R(reset_n_bF_buf61), .S(1'h1));
DFFSR DFFSR_741 ( .CLK(clk_bF_buf60), .D(w_mem_inst__0w_mem_12__31_0__18_), .Q(w_mem_inst_w_mem_12__18_), .R(reset_n_bF_buf60), .S(1'h1));
DFFSR DFFSR_742 ( .CLK(clk_bF_buf59), .D(w_mem_inst__0w_mem_12__31_0__19_), .Q(w_mem_inst_w_mem_12__19_), .R(reset_n_bF_buf59), .S(1'h1));
DFFSR DFFSR_743 ( .CLK(clk_bF_buf58), .D(w_mem_inst__0w_mem_12__31_0__20_), .Q(w_mem_inst_w_mem_12__20_), .R(reset_n_bF_buf58), .S(1'h1));
DFFSR DFFSR_744 ( .CLK(clk_bF_buf57), .D(w_mem_inst__0w_mem_12__31_0__21_), .Q(w_mem_inst_w_mem_12__21_), .R(reset_n_bF_buf57), .S(1'h1));
DFFSR DFFSR_745 ( .CLK(clk_bF_buf56), .D(w_mem_inst__0w_mem_12__31_0__22_), .Q(w_mem_inst_w_mem_12__22_), .R(reset_n_bF_buf56), .S(1'h1));
DFFSR DFFSR_746 ( .CLK(clk_bF_buf55), .D(w_mem_inst__0w_mem_12__31_0__23_), .Q(w_mem_inst_w_mem_12__23_), .R(reset_n_bF_buf55), .S(1'h1));
DFFSR DFFSR_747 ( .CLK(clk_bF_buf54), .D(w_mem_inst__0w_mem_12__31_0__24_), .Q(w_mem_inst_w_mem_12__24_), .R(reset_n_bF_buf54), .S(1'h1));
DFFSR DFFSR_748 ( .CLK(clk_bF_buf53), .D(w_mem_inst__0w_mem_12__31_0__25_), .Q(w_mem_inst_w_mem_12__25_), .R(reset_n_bF_buf53), .S(1'h1));
DFFSR DFFSR_749 ( .CLK(clk_bF_buf52), .D(w_mem_inst__0w_mem_12__31_0__26_), .Q(w_mem_inst_w_mem_12__26_), .R(reset_n_bF_buf52), .S(1'h1));
DFFSR DFFSR_75 ( .CLK(clk_bF_buf14), .D(_0c_reg_31_0__10_), .Q(c_reg_10_), .R(reset_n_bF_buf14), .S(1'h1));
DFFSR DFFSR_750 ( .CLK(clk_bF_buf51), .D(w_mem_inst__0w_mem_12__31_0__27_), .Q(w_mem_inst_w_mem_12__27_), .R(reset_n_bF_buf51), .S(1'h1));
DFFSR DFFSR_751 ( .CLK(clk_bF_buf50), .D(w_mem_inst__0w_mem_12__31_0__28_), .Q(w_mem_inst_w_mem_12__28_), .R(reset_n_bF_buf50), .S(1'h1));
DFFSR DFFSR_752 ( .CLK(clk_bF_buf49), .D(w_mem_inst__0w_mem_12__31_0__29_), .Q(w_mem_inst_w_mem_12__29_), .R(reset_n_bF_buf49), .S(1'h1));
DFFSR DFFSR_753 ( .CLK(clk_bF_buf48), .D(w_mem_inst__0w_mem_12__31_0__30_), .Q(w_mem_inst_w_mem_12__30_), .R(reset_n_bF_buf48), .S(1'h1));
DFFSR DFFSR_754 ( .CLK(clk_bF_buf47), .D(w_mem_inst__0w_mem_12__31_0__31_), .Q(w_mem_inst_w_mem_12__31_), .R(reset_n_bF_buf47), .S(1'h1));
DFFSR DFFSR_755 ( .CLK(clk_bF_buf46), .D(w_mem_inst__0w_mem_13__31_0__0_), .Q(w_mem_inst_w_mem_13__0_), .R(reset_n_bF_buf46), .S(1'h1));
DFFSR DFFSR_756 ( .CLK(clk_bF_buf45), .D(w_mem_inst__0w_mem_13__31_0__1_), .Q(w_mem_inst_w_mem_13__1_), .R(reset_n_bF_buf45), .S(1'h1));
DFFSR DFFSR_757 ( .CLK(clk_bF_buf44), .D(w_mem_inst__0w_mem_13__31_0__2_), .Q(w_mem_inst_w_mem_13__2_), .R(reset_n_bF_buf44), .S(1'h1));
DFFSR DFFSR_758 ( .CLK(clk_bF_buf43), .D(w_mem_inst__0w_mem_13__31_0__3_), .Q(w_mem_inst_w_mem_13__3_), .R(reset_n_bF_buf43), .S(1'h1));
DFFSR DFFSR_759 ( .CLK(clk_bF_buf42), .D(w_mem_inst__0w_mem_13__31_0__4_), .Q(w_mem_inst_w_mem_13__4_), .R(reset_n_bF_buf42), .S(1'h1));
DFFSR DFFSR_76 ( .CLK(clk_bF_buf13), .D(_0c_reg_31_0__11_), .Q(c_reg_11_), .R(reset_n_bF_buf13), .S(1'h1));
DFFSR DFFSR_760 ( .CLK(clk_bF_buf41), .D(w_mem_inst__0w_mem_13__31_0__5_), .Q(w_mem_inst_w_mem_13__5_), .R(reset_n_bF_buf41), .S(1'h1));
DFFSR DFFSR_761 ( .CLK(clk_bF_buf40), .D(w_mem_inst__0w_mem_13__31_0__6_), .Q(w_mem_inst_w_mem_13__6_), .R(reset_n_bF_buf40), .S(1'h1));
DFFSR DFFSR_762 ( .CLK(clk_bF_buf39), .D(w_mem_inst__0w_mem_13__31_0__7_), .Q(w_mem_inst_w_mem_13__7_), .R(reset_n_bF_buf39), .S(1'h1));
DFFSR DFFSR_763 ( .CLK(clk_bF_buf38), .D(w_mem_inst__0w_mem_13__31_0__8_), .Q(w_mem_inst_w_mem_13__8_), .R(reset_n_bF_buf38), .S(1'h1));
DFFSR DFFSR_764 ( .CLK(clk_bF_buf37), .D(w_mem_inst__0w_mem_13__31_0__9_), .Q(w_mem_inst_w_mem_13__9_), .R(reset_n_bF_buf37), .S(1'h1));
DFFSR DFFSR_765 ( .CLK(clk_bF_buf36), .D(w_mem_inst__0w_mem_13__31_0__10_), .Q(w_mem_inst_w_mem_13__10_), .R(reset_n_bF_buf36), .S(1'h1));
DFFSR DFFSR_766 ( .CLK(clk_bF_buf35), .D(w_mem_inst__0w_mem_13__31_0__11_), .Q(w_mem_inst_w_mem_13__11_), .R(reset_n_bF_buf35), .S(1'h1));
DFFSR DFFSR_767 ( .CLK(clk_bF_buf34), .D(w_mem_inst__0w_mem_13__31_0__12_), .Q(w_mem_inst_w_mem_13__12_), .R(reset_n_bF_buf34), .S(1'h1));
DFFSR DFFSR_768 ( .CLK(clk_bF_buf33), .D(w_mem_inst__0w_mem_13__31_0__13_), .Q(w_mem_inst_w_mem_13__13_), .R(reset_n_bF_buf33), .S(1'h1));
DFFSR DFFSR_769 ( .CLK(clk_bF_buf32), .D(w_mem_inst__0w_mem_13__31_0__14_), .Q(w_mem_inst_w_mem_13__14_), .R(reset_n_bF_buf32), .S(1'h1));
DFFSR DFFSR_77 ( .CLK(clk_bF_buf12), .D(_0c_reg_31_0__12_), .Q(c_reg_12_), .R(reset_n_bF_buf12), .S(1'h1));
DFFSR DFFSR_770 ( .CLK(clk_bF_buf31), .D(w_mem_inst__0w_mem_13__31_0__15_), .Q(w_mem_inst_w_mem_13__15_), .R(reset_n_bF_buf31), .S(1'h1));
DFFSR DFFSR_771 ( .CLK(clk_bF_buf30), .D(w_mem_inst__0w_mem_13__31_0__16_), .Q(w_mem_inst_w_mem_13__16_), .R(reset_n_bF_buf30), .S(1'h1));
DFFSR DFFSR_772 ( .CLK(clk_bF_buf29), .D(w_mem_inst__0w_mem_13__31_0__17_), .Q(w_mem_inst_w_mem_13__17_), .R(reset_n_bF_buf29), .S(1'h1));
DFFSR DFFSR_773 ( .CLK(clk_bF_buf28), .D(w_mem_inst__0w_mem_13__31_0__18_), .Q(w_mem_inst_w_mem_13__18_), .R(reset_n_bF_buf28), .S(1'h1));
DFFSR DFFSR_774 ( .CLK(clk_bF_buf27), .D(w_mem_inst__0w_mem_13__31_0__19_), .Q(w_mem_inst_w_mem_13__19_), .R(reset_n_bF_buf27), .S(1'h1));
DFFSR DFFSR_775 ( .CLK(clk_bF_buf26), .D(w_mem_inst__0w_mem_13__31_0__20_), .Q(w_mem_inst_w_mem_13__20_), .R(reset_n_bF_buf26), .S(1'h1));
DFFSR DFFSR_776 ( .CLK(clk_bF_buf25), .D(w_mem_inst__0w_mem_13__31_0__21_), .Q(w_mem_inst_w_mem_13__21_), .R(reset_n_bF_buf25), .S(1'h1));
DFFSR DFFSR_777 ( .CLK(clk_bF_buf24), .D(w_mem_inst__0w_mem_13__31_0__22_), .Q(w_mem_inst_w_mem_13__22_), .R(reset_n_bF_buf24), .S(1'h1));
DFFSR DFFSR_778 ( .CLK(clk_bF_buf23), .D(w_mem_inst__0w_mem_13__31_0__23_), .Q(w_mem_inst_w_mem_13__23_), .R(reset_n_bF_buf23), .S(1'h1));
DFFSR DFFSR_779 ( .CLK(clk_bF_buf22), .D(w_mem_inst__0w_mem_13__31_0__24_), .Q(w_mem_inst_w_mem_13__24_), .R(reset_n_bF_buf22), .S(1'h1));
DFFSR DFFSR_78 ( .CLK(clk_bF_buf11), .D(_0c_reg_31_0__13_), .Q(c_reg_13_), .R(reset_n_bF_buf11), .S(1'h1));
DFFSR DFFSR_780 ( .CLK(clk_bF_buf21), .D(w_mem_inst__0w_mem_13__31_0__25_), .Q(w_mem_inst_w_mem_13__25_), .R(reset_n_bF_buf21), .S(1'h1));
DFFSR DFFSR_781 ( .CLK(clk_bF_buf20), .D(w_mem_inst__0w_mem_13__31_0__26_), .Q(w_mem_inst_w_mem_13__26_), .R(reset_n_bF_buf20), .S(1'h1));
DFFSR DFFSR_782 ( .CLK(clk_bF_buf19), .D(w_mem_inst__0w_mem_13__31_0__27_), .Q(w_mem_inst_w_mem_13__27_), .R(reset_n_bF_buf19), .S(1'h1));
DFFSR DFFSR_783 ( .CLK(clk_bF_buf18), .D(w_mem_inst__0w_mem_13__31_0__28_), .Q(w_mem_inst_w_mem_13__28_), .R(reset_n_bF_buf18), .S(1'h1));
DFFSR DFFSR_784 ( .CLK(clk_bF_buf17), .D(w_mem_inst__0w_mem_13__31_0__29_), .Q(w_mem_inst_w_mem_13__29_), .R(reset_n_bF_buf17), .S(1'h1));
DFFSR DFFSR_785 ( .CLK(clk_bF_buf16), .D(w_mem_inst__0w_mem_13__31_0__30_), .Q(w_mem_inst_w_mem_13__30_), .R(reset_n_bF_buf16), .S(1'h1));
DFFSR DFFSR_786 ( .CLK(clk_bF_buf15), .D(w_mem_inst__0w_mem_13__31_0__31_), .Q(w_mem_inst_w_mem_13__31_), .R(reset_n_bF_buf15), .S(1'h1));
DFFSR DFFSR_787 ( .CLK(clk_bF_buf14), .D(w_mem_inst__0w_mem_14__31_0__0_), .Q(w_mem_inst_w_mem_14__0_), .R(reset_n_bF_buf14), .S(1'h1));
DFFSR DFFSR_788 ( .CLK(clk_bF_buf13), .D(w_mem_inst__0w_mem_14__31_0__1_), .Q(w_mem_inst_w_mem_14__1_), .R(reset_n_bF_buf13), .S(1'h1));
DFFSR DFFSR_789 ( .CLK(clk_bF_buf12), .D(w_mem_inst__0w_mem_14__31_0__2_), .Q(w_mem_inst_w_mem_14__2_), .R(reset_n_bF_buf12), .S(1'h1));
DFFSR DFFSR_79 ( .CLK(clk_bF_buf10), .D(_0c_reg_31_0__14_), .Q(c_reg_14_), .R(reset_n_bF_buf10), .S(1'h1));
DFFSR DFFSR_790 ( .CLK(clk_bF_buf11), .D(w_mem_inst__0w_mem_14__31_0__3_), .Q(w_mem_inst_w_mem_14__3_), .R(reset_n_bF_buf11), .S(1'h1));
DFFSR DFFSR_791 ( .CLK(clk_bF_buf10), .D(w_mem_inst__0w_mem_14__31_0__4_), .Q(w_mem_inst_w_mem_14__4_), .R(reset_n_bF_buf10), .S(1'h1));
DFFSR DFFSR_792 ( .CLK(clk_bF_buf9), .D(w_mem_inst__0w_mem_14__31_0__5_), .Q(w_mem_inst_w_mem_14__5_), .R(reset_n_bF_buf9), .S(1'h1));
DFFSR DFFSR_793 ( .CLK(clk_bF_buf8), .D(w_mem_inst__0w_mem_14__31_0__6_), .Q(w_mem_inst_w_mem_14__6_), .R(reset_n_bF_buf8), .S(1'h1));
DFFSR DFFSR_794 ( .CLK(clk_bF_buf7), .D(w_mem_inst__0w_mem_14__31_0__7_), .Q(w_mem_inst_w_mem_14__7_), .R(reset_n_bF_buf7), .S(1'h1));
DFFSR DFFSR_795 ( .CLK(clk_bF_buf6), .D(w_mem_inst__0w_mem_14__31_0__8_), .Q(w_mem_inst_w_mem_14__8_), .R(reset_n_bF_buf6), .S(1'h1));
DFFSR DFFSR_796 ( .CLK(clk_bF_buf5), .D(w_mem_inst__0w_mem_14__31_0__9_), .Q(w_mem_inst_w_mem_14__9_), .R(reset_n_bF_buf5), .S(1'h1));
DFFSR DFFSR_797 ( .CLK(clk_bF_buf4), .D(w_mem_inst__0w_mem_14__31_0__10_), .Q(w_mem_inst_w_mem_14__10_), .R(reset_n_bF_buf4), .S(1'h1));
DFFSR DFFSR_798 ( .CLK(clk_bF_buf3), .D(w_mem_inst__0w_mem_14__31_0__11_), .Q(w_mem_inst_w_mem_14__11_), .R(reset_n_bF_buf3), .S(1'h1));
DFFSR DFFSR_799 ( .CLK(clk_bF_buf2), .D(w_mem_inst__0w_mem_14__31_0__12_), .Q(w_mem_inst_w_mem_14__12_), .R(reset_n_bF_buf2), .S(1'h1));
DFFSR DFFSR_8 ( .CLK(clk_bF_buf81), .D(_0a_reg_31_0__7_), .Q(a_reg_7_), .R(reset_n_bF_buf81), .S(1'h1));
DFFSR DFFSR_80 ( .CLK(clk_bF_buf9), .D(_0c_reg_31_0__15_), .Q(c_reg_15_), .R(reset_n_bF_buf9), .S(1'h1));
DFFSR DFFSR_800 ( .CLK(clk_bF_buf1), .D(w_mem_inst__0w_mem_14__31_0__13_), .Q(w_mem_inst_w_mem_14__13_), .R(reset_n_bF_buf1), .S(1'h1));
DFFSR DFFSR_801 ( .CLK(clk_bF_buf0), .D(w_mem_inst__0w_mem_14__31_0__14_), .Q(w_mem_inst_w_mem_14__14_), .R(reset_n_bF_buf0), .S(1'h1));
DFFSR DFFSR_802 ( .CLK(clk_bF_buf88), .D(w_mem_inst__0w_mem_14__31_0__15_), .Q(w_mem_inst_w_mem_14__15_), .R(reset_n_bF_buf88), .S(1'h1));
DFFSR DFFSR_803 ( .CLK(clk_bF_buf87), .D(w_mem_inst__0w_mem_14__31_0__16_), .Q(w_mem_inst_w_mem_14__16_), .R(reset_n_bF_buf87), .S(1'h1));
DFFSR DFFSR_804 ( .CLK(clk_bF_buf86), .D(w_mem_inst__0w_mem_14__31_0__17_), .Q(w_mem_inst_w_mem_14__17_), .R(reset_n_bF_buf86), .S(1'h1));
DFFSR DFFSR_805 ( .CLK(clk_bF_buf85), .D(w_mem_inst__0w_mem_14__31_0__18_), .Q(w_mem_inst_w_mem_14__18_), .R(reset_n_bF_buf85), .S(1'h1));
DFFSR DFFSR_806 ( .CLK(clk_bF_buf84), .D(w_mem_inst__0w_mem_14__31_0__19_), .Q(w_mem_inst_w_mem_14__19_), .R(reset_n_bF_buf84), .S(1'h1));
DFFSR DFFSR_807 ( .CLK(clk_bF_buf83), .D(w_mem_inst__0w_mem_14__31_0__20_), .Q(w_mem_inst_w_mem_14__20_), .R(reset_n_bF_buf83), .S(1'h1));
DFFSR DFFSR_808 ( .CLK(clk_bF_buf82), .D(w_mem_inst__0w_mem_14__31_0__21_), .Q(w_mem_inst_w_mem_14__21_), .R(reset_n_bF_buf82), .S(1'h1));
DFFSR DFFSR_809 ( .CLK(clk_bF_buf81), .D(w_mem_inst__0w_mem_14__31_0__22_), .Q(w_mem_inst_w_mem_14__22_), .R(reset_n_bF_buf81), .S(1'h1));
DFFSR DFFSR_81 ( .CLK(clk_bF_buf8), .D(_0c_reg_31_0__16_), .Q(c_reg_16_), .R(reset_n_bF_buf8), .S(1'h1));
DFFSR DFFSR_810 ( .CLK(clk_bF_buf80), .D(w_mem_inst__0w_mem_14__31_0__23_), .Q(w_mem_inst_w_mem_14__23_), .R(reset_n_bF_buf80), .S(1'h1));
DFFSR DFFSR_811 ( .CLK(clk_bF_buf79), .D(w_mem_inst__0w_mem_14__31_0__24_), .Q(w_mem_inst_w_mem_14__24_), .R(reset_n_bF_buf79), .S(1'h1));
DFFSR DFFSR_812 ( .CLK(clk_bF_buf78), .D(w_mem_inst__0w_mem_14__31_0__25_), .Q(w_mem_inst_w_mem_14__25_), .R(reset_n_bF_buf78), .S(1'h1));
DFFSR DFFSR_813 ( .CLK(clk_bF_buf77), .D(w_mem_inst__0w_mem_14__31_0__26_), .Q(w_mem_inst_w_mem_14__26_), .R(reset_n_bF_buf77), .S(1'h1));
DFFSR DFFSR_814 ( .CLK(clk_bF_buf76), .D(w_mem_inst__0w_mem_14__31_0__27_), .Q(w_mem_inst_w_mem_14__27_), .R(reset_n_bF_buf76), .S(1'h1));
DFFSR DFFSR_815 ( .CLK(clk_bF_buf75), .D(w_mem_inst__0w_mem_14__31_0__28_), .Q(w_mem_inst_w_mem_14__28_), .R(reset_n_bF_buf75), .S(1'h1));
DFFSR DFFSR_816 ( .CLK(clk_bF_buf74), .D(w_mem_inst__0w_mem_14__31_0__29_), .Q(w_mem_inst_w_mem_14__29_), .R(reset_n_bF_buf74), .S(1'h1));
DFFSR DFFSR_817 ( .CLK(clk_bF_buf73), .D(w_mem_inst__0w_mem_14__31_0__30_), .Q(w_mem_inst_w_mem_14__30_), .R(reset_n_bF_buf73), .S(1'h1));
DFFSR DFFSR_818 ( .CLK(clk_bF_buf72), .D(w_mem_inst__0w_mem_14__31_0__31_), .Q(w_mem_inst_w_mem_14__31_), .R(reset_n_bF_buf72), .S(1'h1));
DFFSR DFFSR_819 ( .CLK(clk_bF_buf71), .D(w_mem_inst__0w_mem_15__31_0__0_), .Q(w_mem_inst_w_mem_15__0_), .R(reset_n_bF_buf71), .S(1'h1));
DFFSR DFFSR_82 ( .CLK(clk_bF_buf7), .D(_0c_reg_31_0__17_), .Q(c_reg_17_), .R(reset_n_bF_buf7), .S(1'h1));
DFFSR DFFSR_820 ( .CLK(clk_bF_buf70), .D(w_mem_inst__0w_mem_15__31_0__1_), .Q(w_mem_inst_w_mem_15__1_), .R(reset_n_bF_buf70), .S(1'h1));
DFFSR DFFSR_821 ( .CLK(clk_bF_buf69), .D(w_mem_inst__0w_mem_15__31_0__2_), .Q(w_mem_inst_w_mem_15__2_), .R(reset_n_bF_buf69), .S(1'h1));
DFFSR DFFSR_822 ( .CLK(clk_bF_buf68), .D(w_mem_inst__0w_mem_15__31_0__3_), .Q(w_mem_inst_w_mem_15__3_), .R(reset_n_bF_buf68), .S(1'h1));
DFFSR DFFSR_823 ( .CLK(clk_bF_buf67), .D(w_mem_inst__0w_mem_15__31_0__4_), .Q(w_mem_inst_w_mem_15__4_), .R(reset_n_bF_buf67), .S(1'h1));
DFFSR DFFSR_824 ( .CLK(clk_bF_buf66), .D(w_mem_inst__0w_mem_15__31_0__5_), .Q(w_mem_inst_w_mem_15__5_), .R(reset_n_bF_buf66), .S(1'h1));
DFFSR DFFSR_825 ( .CLK(clk_bF_buf65), .D(w_mem_inst__0w_mem_15__31_0__6_), .Q(w_mem_inst_w_mem_15__6_), .R(reset_n_bF_buf65), .S(1'h1));
DFFSR DFFSR_826 ( .CLK(clk_bF_buf64), .D(w_mem_inst__0w_mem_15__31_0__7_), .Q(w_mem_inst_w_mem_15__7_), .R(reset_n_bF_buf64), .S(1'h1));
DFFSR DFFSR_827 ( .CLK(clk_bF_buf63), .D(w_mem_inst__0w_mem_15__31_0__8_), .Q(w_mem_inst_w_mem_15__8_), .R(reset_n_bF_buf63), .S(1'h1));
DFFSR DFFSR_828 ( .CLK(clk_bF_buf62), .D(w_mem_inst__0w_mem_15__31_0__9_), .Q(w_mem_inst_w_mem_15__9_), .R(reset_n_bF_buf62), .S(1'h1));
DFFSR DFFSR_829 ( .CLK(clk_bF_buf61), .D(w_mem_inst__0w_mem_15__31_0__10_), .Q(w_mem_inst_w_mem_15__10_), .R(reset_n_bF_buf61), .S(1'h1));
DFFSR DFFSR_83 ( .CLK(clk_bF_buf6), .D(_0c_reg_31_0__18_), .Q(c_reg_18_), .R(reset_n_bF_buf6), .S(1'h1));
DFFSR DFFSR_830 ( .CLK(clk_bF_buf60), .D(w_mem_inst__0w_mem_15__31_0__11_), .Q(w_mem_inst_w_mem_15__11_), .R(reset_n_bF_buf60), .S(1'h1));
DFFSR DFFSR_831 ( .CLK(clk_bF_buf59), .D(w_mem_inst__0w_mem_15__31_0__12_), .Q(w_mem_inst_w_mem_15__12_), .R(reset_n_bF_buf59), .S(1'h1));
DFFSR DFFSR_832 ( .CLK(clk_bF_buf58), .D(w_mem_inst__0w_mem_15__31_0__13_), .Q(w_mem_inst_w_mem_15__13_), .R(reset_n_bF_buf58), .S(1'h1));
DFFSR DFFSR_833 ( .CLK(clk_bF_buf57), .D(w_mem_inst__0w_mem_15__31_0__14_), .Q(w_mem_inst_w_mem_15__14_), .R(reset_n_bF_buf57), .S(1'h1));
DFFSR DFFSR_834 ( .CLK(clk_bF_buf56), .D(w_mem_inst__0w_mem_15__31_0__15_), .Q(w_mem_inst_w_mem_15__15_), .R(reset_n_bF_buf56), .S(1'h1));
DFFSR DFFSR_835 ( .CLK(clk_bF_buf55), .D(w_mem_inst__0w_mem_15__31_0__16_), .Q(w_mem_inst_w_mem_15__16_), .R(reset_n_bF_buf55), .S(1'h1));
DFFSR DFFSR_836 ( .CLK(clk_bF_buf54), .D(w_mem_inst__0w_mem_15__31_0__17_), .Q(w_mem_inst_w_mem_15__17_), .R(reset_n_bF_buf54), .S(1'h1));
DFFSR DFFSR_837 ( .CLK(clk_bF_buf53), .D(w_mem_inst__0w_mem_15__31_0__18_), .Q(w_mem_inst_w_mem_15__18_), .R(reset_n_bF_buf53), .S(1'h1));
DFFSR DFFSR_838 ( .CLK(clk_bF_buf52), .D(w_mem_inst__0w_mem_15__31_0__19_), .Q(w_mem_inst_w_mem_15__19_), .R(reset_n_bF_buf52), .S(1'h1));
DFFSR DFFSR_839 ( .CLK(clk_bF_buf51), .D(w_mem_inst__0w_mem_15__31_0__20_), .Q(w_mem_inst_w_mem_15__20_), .R(reset_n_bF_buf51), .S(1'h1));
DFFSR DFFSR_84 ( .CLK(clk_bF_buf5), .D(_0c_reg_31_0__19_), .Q(c_reg_19_), .R(reset_n_bF_buf5), .S(1'h1));
DFFSR DFFSR_840 ( .CLK(clk_bF_buf50), .D(w_mem_inst__0w_mem_15__31_0__21_), .Q(w_mem_inst_w_mem_15__21_), .R(reset_n_bF_buf50), .S(1'h1));
DFFSR DFFSR_841 ( .CLK(clk_bF_buf49), .D(w_mem_inst__0w_mem_15__31_0__22_), .Q(w_mem_inst_w_mem_15__22_), .R(reset_n_bF_buf49), .S(1'h1));
DFFSR DFFSR_842 ( .CLK(clk_bF_buf48), .D(w_mem_inst__0w_mem_15__31_0__23_), .Q(w_mem_inst_w_mem_15__23_), .R(reset_n_bF_buf48), .S(1'h1));
DFFSR DFFSR_843 ( .CLK(clk_bF_buf47), .D(w_mem_inst__0w_mem_15__31_0__24_), .Q(w_mem_inst_w_mem_15__24_), .R(reset_n_bF_buf47), .S(1'h1));
DFFSR DFFSR_844 ( .CLK(clk_bF_buf46), .D(w_mem_inst__0w_mem_15__31_0__25_), .Q(w_mem_inst_w_mem_15__25_), .R(reset_n_bF_buf46), .S(1'h1));
DFFSR DFFSR_845 ( .CLK(clk_bF_buf45), .D(w_mem_inst__0w_mem_15__31_0__26_), .Q(w_mem_inst_w_mem_15__26_), .R(reset_n_bF_buf45), .S(1'h1));
DFFSR DFFSR_846 ( .CLK(clk_bF_buf44), .D(w_mem_inst__0w_mem_15__31_0__27_), .Q(w_mem_inst_w_mem_15__27_), .R(reset_n_bF_buf44), .S(1'h1));
DFFSR DFFSR_847 ( .CLK(clk_bF_buf43), .D(w_mem_inst__0w_mem_15__31_0__28_), .Q(w_mem_inst_w_mem_15__28_), .R(reset_n_bF_buf43), .S(1'h1));
DFFSR DFFSR_848 ( .CLK(clk_bF_buf42), .D(w_mem_inst__0w_mem_15__31_0__29_), .Q(w_mem_inst_w_mem_15__29_), .R(reset_n_bF_buf42), .S(1'h1));
DFFSR DFFSR_849 ( .CLK(clk_bF_buf41), .D(w_mem_inst__0w_mem_15__31_0__30_), .Q(w_mem_inst_w_mem_15__30_), .R(reset_n_bF_buf41), .S(1'h1));
DFFSR DFFSR_85 ( .CLK(clk_bF_buf4), .D(_0c_reg_31_0__20_), .Q(c_reg_20_), .R(reset_n_bF_buf4), .S(1'h1));
DFFSR DFFSR_850 ( .CLK(clk_bF_buf40), .D(w_mem_inst__0w_mem_15__31_0__31_), .Q(w_mem_inst_w_mem_15__31_), .R(reset_n_bF_buf40), .S(1'h1));
DFFSR DFFSR_86 ( .CLK(clk_bF_buf3), .D(_0c_reg_31_0__21_), .Q(c_reg_21_), .R(reset_n_bF_buf3), .S(1'h1));
DFFSR DFFSR_87 ( .CLK(clk_bF_buf2), .D(_0c_reg_31_0__22_), .Q(c_reg_22_), .R(reset_n_bF_buf2), .S(1'h1));
DFFSR DFFSR_88 ( .CLK(clk_bF_buf1), .D(_0c_reg_31_0__23_), .Q(c_reg_23_), .R(reset_n_bF_buf1), .S(1'h1));
DFFSR DFFSR_89 ( .CLK(clk_bF_buf0), .D(_0c_reg_31_0__24_), .Q(c_reg_24_), .R(reset_n_bF_buf0), .S(1'h1));
DFFSR DFFSR_9 ( .CLK(clk_bF_buf80), .D(_0a_reg_31_0__8_), .Q(a_reg_8_), .R(reset_n_bF_buf80), .S(1'h1));
DFFSR DFFSR_90 ( .CLK(clk_bF_buf88), .D(_0c_reg_31_0__25_), .Q(c_reg_25_), .R(reset_n_bF_buf88), .S(1'h1));
DFFSR DFFSR_91 ( .CLK(clk_bF_buf87), .D(_0c_reg_31_0__26_), .Q(c_reg_26_), .R(reset_n_bF_buf87), .S(1'h1));
DFFSR DFFSR_92 ( .CLK(clk_bF_buf86), .D(_0c_reg_31_0__27_), .Q(c_reg_27_), .R(reset_n_bF_buf86), .S(1'h1));
DFFSR DFFSR_93 ( .CLK(clk_bF_buf85), .D(_0c_reg_31_0__28_), .Q(c_reg_28_), .R(reset_n_bF_buf85), .S(1'h1));
DFFSR DFFSR_94 ( .CLK(clk_bF_buf84), .D(_0c_reg_31_0__29_), .Q(c_reg_29_), .R(reset_n_bF_buf84), .S(1'h1));
DFFSR DFFSR_95 ( .CLK(clk_bF_buf83), .D(_0c_reg_31_0__30_), .Q(c_reg_30_), .R(reset_n_bF_buf83), .S(1'h1));
DFFSR DFFSR_96 ( .CLK(clk_bF_buf82), .D(_0c_reg_31_0__31_), .Q(c_reg_31_), .R(reset_n_bF_buf82), .S(1'h1));
DFFSR DFFSR_97 ( .CLK(clk_bF_buf81), .D(_0d_reg_31_0__0_), .Q(d_reg_0_), .R(reset_n_bF_buf81), .S(1'h1));
DFFSR DFFSR_98 ( .CLK(clk_bF_buf80), .D(_0d_reg_31_0__1_), .Q(d_reg_1_), .R(reset_n_bF_buf80), .S(1'h1));
DFFSR DFFSR_99 ( .CLK(clk_bF_buf79), .D(_0d_reg_31_0__2_), .Q(d_reg_2_), .R(reset_n_bF_buf79), .S(1'h1));
INVX1 INVX1_1 ( .A(_auto_iopadmap_cc_368_execute_22625_78_), .Y(_abc_15497_new_n703_));
INVX1 INVX1_10 ( .A(_auto_iopadmap_cc_368_execute_22625_74_), .Y(_abc_15497_new_n728_));
INVX1 INVX1_100 ( .A(_auto_iopadmap_cc_368_execute_22625_19_), .Y(_abc_15497_new_n1142_));
INVX1 INVX1_1000 ( .A(\block[204] ), .Y(w_mem_inst__abc_19396_new_n3476_));
INVX1 INVX1_1001 ( .A(w_mem_inst_w_mem_9__13_), .Y(w_mem_inst__abc_19396_new_n3480_));
INVX1 INVX1_1002 ( .A(\block[205] ), .Y(w_mem_inst__abc_19396_new_n3481_));
INVX1 INVX1_1003 ( .A(w_mem_inst_w_mem_9__14_), .Y(w_mem_inst__abc_19396_new_n3485_));
INVX1 INVX1_1004 ( .A(\block[206] ), .Y(w_mem_inst__abc_19396_new_n3486_));
INVX1 INVX1_1005 ( .A(w_mem_inst_w_mem_9__15_), .Y(w_mem_inst__abc_19396_new_n3490_));
INVX1 INVX1_1006 ( .A(\block[207] ), .Y(w_mem_inst__abc_19396_new_n3491_));
INVX1 INVX1_1007 ( .A(w_mem_inst_w_mem_9__16_), .Y(w_mem_inst__abc_19396_new_n3495_));
INVX1 INVX1_1008 ( .A(\block[208] ), .Y(w_mem_inst__abc_19396_new_n3496_));
INVX1 INVX1_1009 ( .A(w_mem_inst_w_mem_9__17_), .Y(w_mem_inst__abc_19396_new_n3500_));
INVX1 INVX1_101 ( .A(_abc_15497_new_n1131_), .Y(_abc_15497_new_n1143_));
INVX1 INVX1_1010 ( .A(\block[209] ), .Y(w_mem_inst__abc_19396_new_n3501_));
INVX1 INVX1_1011 ( .A(w_mem_inst_w_mem_9__18_), .Y(w_mem_inst__abc_19396_new_n3505_));
INVX1 INVX1_1012 ( .A(\block[210] ), .Y(w_mem_inst__abc_19396_new_n3506_));
INVX1 INVX1_1013 ( .A(w_mem_inst_w_mem_9__19_), .Y(w_mem_inst__abc_19396_new_n3510_));
INVX1 INVX1_1014 ( .A(\block[211] ), .Y(w_mem_inst__abc_19396_new_n3511_));
INVX1 INVX1_1015 ( .A(w_mem_inst_w_mem_9__20_), .Y(w_mem_inst__abc_19396_new_n3515_));
INVX1 INVX1_1016 ( .A(\block[212] ), .Y(w_mem_inst__abc_19396_new_n3516_));
INVX1 INVX1_1017 ( .A(w_mem_inst_w_mem_9__21_), .Y(w_mem_inst__abc_19396_new_n3520_));
INVX1 INVX1_1018 ( .A(\block[213] ), .Y(w_mem_inst__abc_19396_new_n3521_));
INVX1 INVX1_1019 ( .A(w_mem_inst_w_mem_9__22_), .Y(w_mem_inst__abc_19396_new_n3525_));
INVX1 INVX1_102 ( .A(_abc_15497_new_n1154_), .Y(_abc_15497_new_n1155_));
INVX1 INVX1_1020 ( .A(\block[214] ), .Y(w_mem_inst__abc_19396_new_n3526_));
INVX1 INVX1_1021 ( .A(w_mem_inst_w_mem_9__23_), .Y(w_mem_inst__abc_19396_new_n3530_));
INVX1 INVX1_1022 ( .A(\block[215] ), .Y(w_mem_inst__abc_19396_new_n3531_));
INVX1 INVX1_1023 ( .A(w_mem_inst_w_mem_9__24_), .Y(w_mem_inst__abc_19396_new_n3535_));
INVX1 INVX1_1024 ( .A(\block[216] ), .Y(w_mem_inst__abc_19396_new_n3536_));
INVX1 INVX1_1025 ( .A(w_mem_inst_w_mem_9__25_), .Y(w_mem_inst__abc_19396_new_n3540_));
INVX1 INVX1_1026 ( .A(\block[217] ), .Y(w_mem_inst__abc_19396_new_n3541_));
INVX1 INVX1_1027 ( .A(w_mem_inst_w_mem_9__26_), .Y(w_mem_inst__abc_19396_new_n3545_));
INVX1 INVX1_1028 ( .A(\block[218] ), .Y(w_mem_inst__abc_19396_new_n3546_));
INVX1 INVX1_1029 ( .A(w_mem_inst_w_mem_9__27_), .Y(w_mem_inst__abc_19396_new_n3550_));
INVX1 INVX1_103 ( .A(_abc_15497_new_n1158_), .Y(_abc_15497_new_n1159_));
INVX1 INVX1_1030 ( .A(\block[219] ), .Y(w_mem_inst__abc_19396_new_n3551_));
INVX1 INVX1_1031 ( .A(w_mem_inst_w_mem_9__28_), .Y(w_mem_inst__abc_19396_new_n3555_));
INVX1 INVX1_1032 ( .A(\block[220] ), .Y(w_mem_inst__abc_19396_new_n3556_));
INVX1 INVX1_1033 ( .A(w_mem_inst_w_mem_9__29_), .Y(w_mem_inst__abc_19396_new_n3560_));
INVX1 INVX1_1034 ( .A(\block[221] ), .Y(w_mem_inst__abc_19396_new_n3561_));
INVX1 INVX1_1035 ( .A(w_mem_inst_w_mem_9__30_), .Y(w_mem_inst__abc_19396_new_n3565_));
INVX1 INVX1_1036 ( .A(\block[222] ), .Y(w_mem_inst__abc_19396_new_n3566_));
INVX1 INVX1_1037 ( .A(w_mem_inst_w_mem_9__31_), .Y(w_mem_inst__abc_19396_new_n3570_));
INVX1 INVX1_1038 ( .A(\block[223] ), .Y(w_mem_inst__abc_19396_new_n3571_));
INVX1 INVX1_1039 ( .A(\block[224] ), .Y(w_mem_inst__abc_19396_new_n3575_));
INVX1 INVX1_104 ( .A(_auto_iopadmap_cc_368_execute_22625_20_), .Y(_abc_15497_new_n1163_));
INVX1 INVX1_1040 ( .A(\block[225] ), .Y(w_mem_inst__abc_19396_new_n3579_));
INVX1 INVX1_1041 ( .A(\block[226] ), .Y(w_mem_inst__abc_19396_new_n3583_));
INVX1 INVX1_1042 ( .A(\block[227] ), .Y(w_mem_inst__abc_19396_new_n3587_));
INVX1 INVX1_1043 ( .A(\block[228] ), .Y(w_mem_inst__abc_19396_new_n3591_));
INVX1 INVX1_1044 ( .A(\block[229] ), .Y(w_mem_inst__abc_19396_new_n3595_));
INVX1 INVX1_1045 ( .A(\block[230] ), .Y(w_mem_inst__abc_19396_new_n3599_));
INVX1 INVX1_1046 ( .A(\block[231] ), .Y(w_mem_inst__abc_19396_new_n3603_));
INVX1 INVX1_1047 ( .A(\block[232] ), .Y(w_mem_inst__abc_19396_new_n3607_));
INVX1 INVX1_1048 ( .A(\block[233] ), .Y(w_mem_inst__abc_19396_new_n3611_));
INVX1 INVX1_1049 ( .A(\block[234] ), .Y(w_mem_inst__abc_19396_new_n3615_));
INVX1 INVX1_105 ( .A(_abc_15497_new_n1179_), .Y(_abc_15497_new_n1180_));
INVX1 INVX1_1050 ( .A(\block[235] ), .Y(w_mem_inst__abc_19396_new_n3619_));
INVX1 INVX1_1051 ( .A(\block[236] ), .Y(w_mem_inst__abc_19396_new_n3623_));
INVX1 INVX1_1052 ( .A(\block[237] ), .Y(w_mem_inst__abc_19396_new_n3627_));
INVX1 INVX1_1053 ( .A(\block[238] ), .Y(w_mem_inst__abc_19396_new_n3631_));
INVX1 INVX1_1054 ( .A(\block[239] ), .Y(w_mem_inst__abc_19396_new_n3635_));
INVX1 INVX1_1055 ( .A(\block[240] ), .Y(w_mem_inst__abc_19396_new_n3639_));
INVX1 INVX1_1056 ( .A(\block[241] ), .Y(w_mem_inst__abc_19396_new_n3643_));
INVX1 INVX1_1057 ( .A(\block[242] ), .Y(w_mem_inst__abc_19396_new_n3647_));
INVX1 INVX1_1058 ( .A(\block[243] ), .Y(w_mem_inst__abc_19396_new_n3651_));
INVX1 INVX1_1059 ( .A(\block[244] ), .Y(w_mem_inst__abc_19396_new_n3655_));
INVX1 INVX1_106 ( .A(_abc_15497_new_n1185_), .Y(_abc_15497_new_n1186_));
INVX1 INVX1_1060 ( .A(\block[245] ), .Y(w_mem_inst__abc_19396_new_n3659_));
INVX1 INVX1_1061 ( .A(\block[246] ), .Y(w_mem_inst__abc_19396_new_n3663_));
INVX1 INVX1_1062 ( .A(\block[247] ), .Y(w_mem_inst__abc_19396_new_n3667_));
INVX1 INVX1_1063 ( .A(\block[248] ), .Y(w_mem_inst__abc_19396_new_n3671_));
INVX1 INVX1_1064 ( .A(\block[249] ), .Y(w_mem_inst__abc_19396_new_n3675_));
INVX1 INVX1_1065 ( .A(\block[250] ), .Y(w_mem_inst__abc_19396_new_n3679_));
INVX1 INVX1_1066 ( .A(\block[251] ), .Y(w_mem_inst__abc_19396_new_n3683_));
INVX1 INVX1_1067 ( .A(\block[252] ), .Y(w_mem_inst__abc_19396_new_n3687_));
INVX1 INVX1_1068 ( .A(\block[253] ), .Y(w_mem_inst__abc_19396_new_n3691_));
INVX1 INVX1_1069 ( .A(\block[254] ), .Y(w_mem_inst__abc_19396_new_n3695_));
INVX1 INVX1_107 ( .A(_abc_15497_new_n1187_), .Y(_abc_15497_new_n1188_));
INVX1 INVX1_1070 ( .A(\block[255] ), .Y(w_mem_inst__abc_19396_new_n3699_));
INVX1 INVX1_1071 ( .A(w_mem_inst_w_mem_4__0_), .Y(w_mem_inst__abc_19396_new_n3703_));
INVX1 INVX1_1072 ( .A(\block[352] ), .Y(w_mem_inst__abc_19396_new_n3704_));
INVX1 INVX1_1073 ( .A(w_mem_inst_w_mem_4__1_), .Y(w_mem_inst__abc_19396_new_n3708_));
INVX1 INVX1_1074 ( .A(\block[353] ), .Y(w_mem_inst__abc_19396_new_n3709_));
INVX1 INVX1_1075 ( .A(w_mem_inst_w_mem_4__2_), .Y(w_mem_inst__abc_19396_new_n3713_));
INVX1 INVX1_1076 ( .A(\block[354] ), .Y(w_mem_inst__abc_19396_new_n3714_));
INVX1 INVX1_1077 ( .A(w_mem_inst_w_mem_4__3_), .Y(w_mem_inst__abc_19396_new_n3718_));
INVX1 INVX1_1078 ( .A(\block[355] ), .Y(w_mem_inst__abc_19396_new_n3719_));
INVX1 INVX1_1079 ( .A(w_mem_inst_w_mem_4__4_), .Y(w_mem_inst__abc_19396_new_n3723_));
INVX1 INVX1_108 ( .A(_abc_15497_new_n1195_), .Y(_abc_15497_new_n1196_));
INVX1 INVX1_1080 ( .A(\block[356] ), .Y(w_mem_inst__abc_19396_new_n3724_));
INVX1 INVX1_1081 ( .A(w_mem_inst_w_mem_4__5_), .Y(w_mem_inst__abc_19396_new_n3728_));
INVX1 INVX1_1082 ( .A(\block[357] ), .Y(w_mem_inst__abc_19396_new_n3729_));
INVX1 INVX1_1083 ( .A(w_mem_inst_w_mem_4__6_), .Y(w_mem_inst__abc_19396_new_n3733_));
INVX1 INVX1_1084 ( .A(\block[358] ), .Y(w_mem_inst__abc_19396_new_n3734_));
INVX1 INVX1_1085 ( .A(w_mem_inst_w_mem_4__7_), .Y(w_mem_inst__abc_19396_new_n3738_));
INVX1 INVX1_1086 ( .A(\block[359] ), .Y(w_mem_inst__abc_19396_new_n3739_));
INVX1 INVX1_1087 ( .A(w_mem_inst_w_mem_4__8_), .Y(w_mem_inst__abc_19396_new_n3743_));
INVX1 INVX1_1088 ( .A(\block[360] ), .Y(w_mem_inst__abc_19396_new_n3744_));
INVX1 INVX1_1089 ( .A(w_mem_inst_w_mem_4__9_), .Y(w_mem_inst__abc_19396_new_n3748_));
INVX1 INVX1_109 ( .A(_abc_15497_new_n1202_), .Y(_abc_15497_new_n1203_));
INVX1 INVX1_1090 ( .A(\block[361] ), .Y(w_mem_inst__abc_19396_new_n3749_));
INVX1 INVX1_1091 ( .A(w_mem_inst_w_mem_4__10_), .Y(w_mem_inst__abc_19396_new_n3753_));
INVX1 INVX1_1092 ( .A(\block[362] ), .Y(w_mem_inst__abc_19396_new_n3754_));
INVX1 INVX1_1093 ( .A(w_mem_inst_w_mem_4__11_), .Y(w_mem_inst__abc_19396_new_n3758_));
INVX1 INVX1_1094 ( .A(\block[363] ), .Y(w_mem_inst__abc_19396_new_n3759_));
INVX1 INVX1_1095 ( .A(w_mem_inst_w_mem_4__12_), .Y(w_mem_inst__abc_19396_new_n3763_));
INVX1 INVX1_1096 ( .A(\block[364] ), .Y(w_mem_inst__abc_19396_new_n3764_));
INVX1 INVX1_1097 ( .A(w_mem_inst_w_mem_4__13_), .Y(w_mem_inst__abc_19396_new_n3768_));
INVX1 INVX1_1098 ( .A(\block[365] ), .Y(w_mem_inst__abc_19396_new_n3769_));
INVX1 INVX1_1099 ( .A(w_mem_inst_w_mem_4__14_), .Y(w_mem_inst__abc_19396_new_n3773_));
INVX1 INVX1_11 ( .A(_abc_15497_new_n732_), .Y(_abc_15497_new_n733_));
INVX1 INVX1_110 ( .A(_abc_15497_new_n1208_), .Y(_abc_15497_new_n1209_));
INVX1 INVX1_1100 ( .A(\block[366] ), .Y(w_mem_inst__abc_19396_new_n3774_));
INVX1 INVX1_1101 ( .A(w_mem_inst_w_mem_4__15_), .Y(w_mem_inst__abc_19396_new_n3778_));
INVX1 INVX1_1102 ( .A(\block[367] ), .Y(w_mem_inst__abc_19396_new_n3779_));
INVX1 INVX1_1103 ( .A(w_mem_inst_w_mem_4__16_), .Y(w_mem_inst__abc_19396_new_n3783_));
INVX1 INVX1_1104 ( .A(\block[368] ), .Y(w_mem_inst__abc_19396_new_n3784_));
INVX1 INVX1_1105 ( .A(w_mem_inst_w_mem_4__17_), .Y(w_mem_inst__abc_19396_new_n3788_));
INVX1 INVX1_1106 ( .A(\block[369] ), .Y(w_mem_inst__abc_19396_new_n3789_));
INVX1 INVX1_1107 ( .A(w_mem_inst_w_mem_4__18_), .Y(w_mem_inst__abc_19396_new_n3793_));
INVX1 INVX1_1108 ( .A(\block[370] ), .Y(w_mem_inst__abc_19396_new_n3794_));
INVX1 INVX1_1109 ( .A(w_mem_inst_w_mem_4__19_), .Y(w_mem_inst__abc_19396_new_n3798_));
INVX1 INVX1_111 ( .A(_abc_15497_new_n1210_), .Y(_abc_15497_new_n1211_));
INVX1 INVX1_1110 ( .A(\block[371] ), .Y(w_mem_inst__abc_19396_new_n3799_));
INVX1 INVX1_1111 ( .A(w_mem_inst_w_mem_4__20_), .Y(w_mem_inst__abc_19396_new_n3803_));
INVX1 INVX1_1112 ( .A(\block[372] ), .Y(w_mem_inst__abc_19396_new_n3804_));
INVX1 INVX1_1113 ( .A(w_mem_inst_w_mem_4__21_), .Y(w_mem_inst__abc_19396_new_n3808_));
INVX1 INVX1_1114 ( .A(\block[373] ), .Y(w_mem_inst__abc_19396_new_n3809_));
INVX1 INVX1_1115 ( .A(w_mem_inst_w_mem_4__22_), .Y(w_mem_inst__abc_19396_new_n3813_));
INVX1 INVX1_1116 ( .A(\block[374] ), .Y(w_mem_inst__abc_19396_new_n3814_));
INVX1 INVX1_1117 ( .A(w_mem_inst_w_mem_4__23_), .Y(w_mem_inst__abc_19396_new_n3818_));
INVX1 INVX1_1118 ( .A(\block[375] ), .Y(w_mem_inst__abc_19396_new_n3819_));
INVX1 INVX1_1119 ( .A(w_mem_inst_w_mem_4__24_), .Y(w_mem_inst__abc_19396_new_n3823_));
INVX1 INVX1_112 ( .A(e_reg_24_), .Y(_abc_15497_new_n1213_));
INVX1 INVX1_1120 ( .A(\block[376] ), .Y(w_mem_inst__abc_19396_new_n3824_));
INVX1 INVX1_1121 ( .A(w_mem_inst_w_mem_4__25_), .Y(w_mem_inst__abc_19396_new_n3828_));
INVX1 INVX1_1122 ( .A(\block[377] ), .Y(w_mem_inst__abc_19396_new_n3829_));
INVX1 INVX1_1123 ( .A(w_mem_inst_w_mem_4__26_), .Y(w_mem_inst__abc_19396_new_n3833_));
INVX1 INVX1_1124 ( .A(\block[378] ), .Y(w_mem_inst__abc_19396_new_n3834_));
INVX1 INVX1_1125 ( .A(w_mem_inst_w_mem_4__27_), .Y(w_mem_inst__abc_19396_new_n3838_));
INVX1 INVX1_1126 ( .A(\block[379] ), .Y(w_mem_inst__abc_19396_new_n3839_));
INVX1 INVX1_1127 ( .A(w_mem_inst_w_mem_4__28_), .Y(w_mem_inst__abc_19396_new_n3843_));
INVX1 INVX1_1128 ( .A(\block[380] ), .Y(w_mem_inst__abc_19396_new_n3844_));
INVX1 INVX1_1129 ( .A(w_mem_inst_w_mem_4__29_), .Y(w_mem_inst__abc_19396_new_n3848_));
INVX1 INVX1_113 ( .A(_auto_iopadmap_cc_368_execute_22625_24_), .Y(_abc_15497_new_n1214_));
INVX1 INVX1_1130 ( .A(\block[381] ), .Y(w_mem_inst__abc_19396_new_n3849_));
INVX1 INVX1_1131 ( .A(w_mem_inst_w_mem_4__30_), .Y(w_mem_inst__abc_19396_new_n3853_));
INVX1 INVX1_1132 ( .A(\block[382] ), .Y(w_mem_inst__abc_19396_new_n3854_));
INVX1 INVX1_1133 ( .A(w_mem_inst_w_mem_4__31_), .Y(w_mem_inst__abc_19396_new_n3858_));
INVX1 INVX1_1134 ( .A(\block[383] ), .Y(w_mem_inst__abc_19396_new_n3859_));
INVX1 INVX1_1135 ( .A(w_mem_inst_w_mem_6__0_), .Y(w_mem_inst__abc_19396_new_n3863_));
INVX1 INVX1_1136 ( .A(\block[288] ), .Y(w_mem_inst__abc_19396_new_n3864_));
INVX1 INVX1_1137 ( .A(w_mem_inst_w_mem_6__1_), .Y(w_mem_inst__abc_19396_new_n3868_));
INVX1 INVX1_1138 ( .A(\block[289] ), .Y(w_mem_inst__abc_19396_new_n3869_));
INVX1 INVX1_1139 ( .A(w_mem_inst_w_mem_6__2_), .Y(w_mem_inst__abc_19396_new_n3873_));
INVX1 INVX1_114 ( .A(_abc_15497_new_n1216_), .Y(_abc_15497_new_n1218_));
INVX1 INVX1_1140 ( .A(\block[290] ), .Y(w_mem_inst__abc_19396_new_n3874_));
INVX1 INVX1_1141 ( .A(w_mem_inst_w_mem_6__3_), .Y(w_mem_inst__abc_19396_new_n3878_));
INVX1 INVX1_1142 ( .A(\block[291] ), .Y(w_mem_inst__abc_19396_new_n3879_));
INVX1 INVX1_1143 ( .A(w_mem_inst_w_mem_6__4_), .Y(w_mem_inst__abc_19396_new_n3883_));
INVX1 INVX1_1144 ( .A(\block[292] ), .Y(w_mem_inst__abc_19396_new_n3884_));
INVX1 INVX1_1145 ( .A(w_mem_inst_w_mem_6__5_), .Y(w_mem_inst__abc_19396_new_n3888_));
INVX1 INVX1_1146 ( .A(\block[293] ), .Y(w_mem_inst__abc_19396_new_n3889_));
INVX1 INVX1_1147 ( .A(w_mem_inst_w_mem_6__6_), .Y(w_mem_inst__abc_19396_new_n3893_));
INVX1 INVX1_1148 ( .A(\block[294] ), .Y(w_mem_inst__abc_19396_new_n3894_));
INVX1 INVX1_1149 ( .A(w_mem_inst_w_mem_6__7_), .Y(w_mem_inst__abc_19396_new_n3898_));
INVX1 INVX1_115 ( .A(_abc_15497_new_n1215_), .Y(_abc_15497_new_n1222_));
INVX1 INVX1_1150 ( .A(\block[295] ), .Y(w_mem_inst__abc_19396_new_n3899_));
INVX1 INVX1_1151 ( .A(w_mem_inst_w_mem_6__8_), .Y(w_mem_inst__abc_19396_new_n3903_));
INVX1 INVX1_1152 ( .A(\block[296] ), .Y(w_mem_inst__abc_19396_new_n3904_));
INVX1 INVX1_1153 ( .A(w_mem_inst_w_mem_6__9_), .Y(w_mem_inst__abc_19396_new_n3908_));
INVX1 INVX1_1154 ( .A(\block[297] ), .Y(w_mem_inst__abc_19396_new_n3909_));
INVX1 INVX1_1155 ( .A(w_mem_inst_w_mem_6__10_), .Y(w_mem_inst__abc_19396_new_n3913_));
INVX1 INVX1_1156 ( .A(\block[298] ), .Y(w_mem_inst__abc_19396_new_n3914_));
INVX1 INVX1_1157 ( .A(w_mem_inst_w_mem_6__11_), .Y(w_mem_inst__abc_19396_new_n3918_));
INVX1 INVX1_1158 ( .A(\block[299] ), .Y(w_mem_inst__abc_19396_new_n3919_));
INVX1 INVX1_1159 ( .A(w_mem_inst_w_mem_6__12_), .Y(w_mem_inst__abc_19396_new_n3923_));
INVX1 INVX1_116 ( .A(_abc_15497_new_n1225_), .Y(_abc_15497_new_n1226_));
INVX1 INVX1_1160 ( .A(\block[300] ), .Y(w_mem_inst__abc_19396_new_n3924_));
INVX1 INVX1_1161 ( .A(w_mem_inst_w_mem_6__13_), .Y(w_mem_inst__abc_19396_new_n3928_));
INVX1 INVX1_1162 ( .A(\block[301] ), .Y(w_mem_inst__abc_19396_new_n3929_));
INVX1 INVX1_1163 ( .A(w_mem_inst_w_mem_6__14_), .Y(w_mem_inst__abc_19396_new_n3933_));
INVX1 INVX1_1164 ( .A(\block[302] ), .Y(w_mem_inst__abc_19396_new_n3934_));
INVX1 INVX1_1165 ( .A(w_mem_inst_w_mem_6__15_), .Y(w_mem_inst__abc_19396_new_n3938_));
INVX1 INVX1_1166 ( .A(\block[303] ), .Y(w_mem_inst__abc_19396_new_n3939_));
INVX1 INVX1_1167 ( .A(w_mem_inst_w_mem_6__16_), .Y(w_mem_inst__abc_19396_new_n3943_));
INVX1 INVX1_1168 ( .A(\block[304] ), .Y(w_mem_inst__abc_19396_new_n3944_));
INVX1 INVX1_1169 ( .A(w_mem_inst_w_mem_6__17_), .Y(w_mem_inst__abc_19396_new_n3948_));
INVX1 INVX1_117 ( .A(_abc_15497_new_n1227_), .Y(_abc_15497_new_n1232_));
INVX1 INVX1_1170 ( .A(\block[305] ), .Y(w_mem_inst__abc_19396_new_n3949_));
INVX1 INVX1_1171 ( .A(w_mem_inst_w_mem_6__18_), .Y(w_mem_inst__abc_19396_new_n3953_));
INVX1 INVX1_1172 ( .A(\block[306] ), .Y(w_mem_inst__abc_19396_new_n3954_));
INVX1 INVX1_1173 ( .A(w_mem_inst_w_mem_6__19_), .Y(w_mem_inst__abc_19396_new_n3958_));
INVX1 INVX1_1174 ( .A(\block[307] ), .Y(w_mem_inst__abc_19396_new_n3959_));
INVX1 INVX1_1175 ( .A(w_mem_inst_w_mem_6__20_), .Y(w_mem_inst__abc_19396_new_n3963_));
INVX1 INVX1_1176 ( .A(\block[308] ), .Y(w_mem_inst__abc_19396_new_n3964_));
INVX1 INVX1_1177 ( .A(w_mem_inst_w_mem_6__21_), .Y(w_mem_inst__abc_19396_new_n3968_));
INVX1 INVX1_1178 ( .A(\block[309] ), .Y(w_mem_inst__abc_19396_new_n3969_));
INVX1 INVX1_1179 ( .A(w_mem_inst_w_mem_6__22_), .Y(w_mem_inst__abc_19396_new_n3973_));
INVX1 INVX1_118 ( .A(_abc_15497_new_n1233_), .Y(_abc_15497_new_n1234_));
INVX1 INVX1_1180 ( .A(\block[310] ), .Y(w_mem_inst__abc_19396_new_n3974_));
INVX1 INVX1_1181 ( .A(w_mem_inst_w_mem_6__23_), .Y(w_mem_inst__abc_19396_new_n3978_));
INVX1 INVX1_1182 ( .A(\block[311] ), .Y(w_mem_inst__abc_19396_new_n3979_));
INVX1 INVX1_1183 ( .A(w_mem_inst_w_mem_6__24_), .Y(w_mem_inst__abc_19396_new_n3983_));
INVX1 INVX1_1184 ( .A(\block[312] ), .Y(w_mem_inst__abc_19396_new_n3984_));
INVX1 INVX1_1185 ( .A(w_mem_inst_w_mem_6__25_), .Y(w_mem_inst__abc_19396_new_n3988_));
INVX1 INVX1_1186 ( .A(\block[313] ), .Y(w_mem_inst__abc_19396_new_n3989_));
INVX1 INVX1_1187 ( .A(w_mem_inst_w_mem_6__26_), .Y(w_mem_inst__abc_19396_new_n3993_));
INVX1 INVX1_1188 ( .A(\block[314] ), .Y(w_mem_inst__abc_19396_new_n3994_));
INVX1 INVX1_1189 ( .A(w_mem_inst_w_mem_6__27_), .Y(w_mem_inst__abc_19396_new_n3998_));
INVX1 INVX1_119 ( .A(_abc_15497_new_n1235_), .Y(_abc_15497_new_n1236_));
INVX1 INVX1_1190 ( .A(\block[315] ), .Y(w_mem_inst__abc_19396_new_n3999_));
INVX1 INVX1_1191 ( .A(w_mem_inst_w_mem_6__28_), .Y(w_mem_inst__abc_19396_new_n4003_));
INVX1 INVX1_1192 ( .A(\block[316] ), .Y(w_mem_inst__abc_19396_new_n4004_));
INVX1 INVX1_1193 ( .A(w_mem_inst_w_mem_6__29_), .Y(w_mem_inst__abc_19396_new_n4008_));
INVX1 INVX1_1194 ( .A(\block[317] ), .Y(w_mem_inst__abc_19396_new_n4009_));
INVX1 INVX1_1195 ( .A(w_mem_inst_w_mem_6__30_), .Y(w_mem_inst__abc_19396_new_n4013_));
INVX1 INVX1_1196 ( .A(\block[318] ), .Y(w_mem_inst__abc_19396_new_n4014_));
INVX1 INVX1_1197 ( .A(w_mem_inst_w_mem_6__31_), .Y(w_mem_inst__abc_19396_new_n4018_));
INVX1 INVX1_1198 ( .A(\block[319] ), .Y(w_mem_inst__abc_19396_new_n4019_));
INVX1 INVX1_1199 ( .A(\block[320] ), .Y(w_mem_inst__abc_19396_new_n4023_));
INVX1 INVX1_12 ( .A(_abc_15497_new_n736_), .Y(_abc_15497_new_n737_));
INVX1 INVX1_120 ( .A(_abc_15497_new_n1237_), .Y(_abc_15497_new_n1243_));
INVX1 INVX1_1200 ( .A(\block[321] ), .Y(w_mem_inst__abc_19396_new_n4027_));
INVX1 INVX1_1201 ( .A(\block[322] ), .Y(w_mem_inst__abc_19396_new_n4031_));
INVX1 INVX1_1202 ( .A(\block[323] ), .Y(w_mem_inst__abc_19396_new_n4035_));
INVX1 INVX1_1203 ( .A(\block[324] ), .Y(w_mem_inst__abc_19396_new_n4039_));
INVX1 INVX1_1204 ( .A(\block[325] ), .Y(w_mem_inst__abc_19396_new_n4043_));
INVX1 INVX1_1205 ( .A(\block[326] ), .Y(w_mem_inst__abc_19396_new_n4047_));
INVX1 INVX1_1206 ( .A(\block[327] ), .Y(w_mem_inst__abc_19396_new_n4051_));
INVX1 INVX1_1207 ( .A(\block[328] ), .Y(w_mem_inst__abc_19396_new_n4055_));
INVX1 INVX1_1208 ( .A(\block[329] ), .Y(w_mem_inst__abc_19396_new_n4059_));
INVX1 INVX1_1209 ( .A(\block[330] ), .Y(w_mem_inst__abc_19396_new_n4063_));
INVX1 INVX1_121 ( .A(_abc_15497_new_n1241_), .Y(_abc_15497_new_n1244_));
INVX1 INVX1_1210 ( .A(\block[331] ), .Y(w_mem_inst__abc_19396_new_n4067_));
INVX1 INVX1_1211 ( .A(\block[332] ), .Y(w_mem_inst__abc_19396_new_n4071_));
INVX1 INVX1_1212 ( .A(\block[333] ), .Y(w_mem_inst__abc_19396_new_n4075_));
INVX1 INVX1_1213 ( .A(\block[334] ), .Y(w_mem_inst__abc_19396_new_n4079_));
INVX1 INVX1_1214 ( .A(\block[335] ), .Y(w_mem_inst__abc_19396_new_n4083_));
INVX1 INVX1_1215 ( .A(\block[336] ), .Y(w_mem_inst__abc_19396_new_n4087_));
INVX1 INVX1_1216 ( .A(\block[337] ), .Y(w_mem_inst__abc_19396_new_n4091_));
INVX1 INVX1_1217 ( .A(\block[338] ), .Y(w_mem_inst__abc_19396_new_n4095_));
INVX1 INVX1_1218 ( .A(\block[339] ), .Y(w_mem_inst__abc_19396_new_n4099_));
INVX1 INVX1_1219 ( .A(\block[340] ), .Y(w_mem_inst__abc_19396_new_n4103_));
INVX1 INVX1_122 ( .A(_abc_15497_new_n1252_), .Y(_abc_15497_new_n1253_));
INVX1 INVX1_1220 ( .A(\block[341] ), .Y(w_mem_inst__abc_19396_new_n4107_));
INVX1 INVX1_1221 ( .A(\block[342] ), .Y(w_mem_inst__abc_19396_new_n4111_));
INVX1 INVX1_1222 ( .A(\block[343] ), .Y(w_mem_inst__abc_19396_new_n4115_));
INVX1 INVX1_1223 ( .A(\block[344] ), .Y(w_mem_inst__abc_19396_new_n4119_));
INVX1 INVX1_1224 ( .A(\block[345] ), .Y(w_mem_inst__abc_19396_new_n4123_));
INVX1 INVX1_1225 ( .A(\block[346] ), .Y(w_mem_inst__abc_19396_new_n4127_));
INVX1 INVX1_1226 ( .A(\block[347] ), .Y(w_mem_inst__abc_19396_new_n4131_));
INVX1 INVX1_1227 ( .A(\block[348] ), .Y(w_mem_inst__abc_19396_new_n4135_));
INVX1 INVX1_1228 ( .A(\block[349] ), .Y(w_mem_inst__abc_19396_new_n4139_));
INVX1 INVX1_1229 ( .A(\block[350] ), .Y(w_mem_inst__abc_19396_new_n4143_));
INVX1 INVX1_123 ( .A(_auto_iopadmap_cc_368_execute_22625_28_), .Y(_abc_15497_new_n1258_));
INVX1 INVX1_1230 ( .A(\block[351] ), .Y(w_mem_inst__abc_19396_new_n4147_));
INVX1 INVX1_1231 ( .A(w_mem_inst_w_mem_1__0_), .Y(w_mem_inst__abc_19396_new_n4151_));
INVX1 INVX1_1232 ( .A(\block[448] ), .Y(w_mem_inst__abc_19396_new_n4152_));
INVX1 INVX1_1233 ( .A(w_mem_inst_w_mem_1__1_), .Y(w_mem_inst__abc_19396_new_n4156_));
INVX1 INVX1_1234 ( .A(\block[449] ), .Y(w_mem_inst__abc_19396_new_n4157_));
INVX1 INVX1_1235 ( .A(w_mem_inst_w_mem_1__2_), .Y(w_mem_inst__abc_19396_new_n4161_));
INVX1 INVX1_1236 ( .A(\block[450] ), .Y(w_mem_inst__abc_19396_new_n4162_));
INVX1 INVX1_1237 ( .A(w_mem_inst_w_mem_1__3_), .Y(w_mem_inst__abc_19396_new_n4166_));
INVX1 INVX1_1238 ( .A(\block[451] ), .Y(w_mem_inst__abc_19396_new_n4167_));
INVX1 INVX1_1239 ( .A(w_mem_inst_w_mem_1__4_), .Y(w_mem_inst__abc_19396_new_n4171_));
INVX1 INVX1_124 ( .A(_auto_iopadmap_cc_368_execute_22625_29_), .Y(_abc_15497_new_n1274_));
INVX1 INVX1_1240 ( .A(\block[452] ), .Y(w_mem_inst__abc_19396_new_n4172_));
INVX1 INVX1_1241 ( .A(w_mem_inst_w_mem_1__5_), .Y(w_mem_inst__abc_19396_new_n4176_));
INVX1 INVX1_1242 ( .A(\block[453] ), .Y(w_mem_inst__abc_19396_new_n4177_));
INVX1 INVX1_1243 ( .A(w_mem_inst_w_mem_1__6_), .Y(w_mem_inst__abc_19396_new_n4181_));
INVX1 INVX1_1244 ( .A(\block[454] ), .Y(w_mem_inst__abc_19396_new_n4182_));
INVX1 INVX1_1245 ( .A(w_mem_inst_w_mem_1__7_), .Y(w_mem_inst__abc_19396_new_n4186_));
INVX1 INVX1_1246 ( .A(\block[455] ), .Y(w_mem_inst__abc_19396_new_n4187_));
INVX1 INVX1_1247 ( .A(w_mem_inst_w_mem_1__8_), .Y(w_mem_inst__abc_19396_new_n4191_));
INVX1 INVX1_1248 ( .A(\block[456] ), .Y(w_mem_inst__abc_19396_new_n4192_));
INVX1 INVX1_1249 ( .A(w_mem_inst_w_mem_1__9_), .Y(w_mem_inst__abc_19396_new_n4196_));
INVX1 INVX1_125 ( .A(_abc_15497_new_n1280_), .Y(_abc_15497_new_n1281_));
INVX1 INVX1_1250 ( .A(\block[457] ), .Y(w_mem_inst__abc_19396_new_n4197_));
INVX1 INVX1_1251 ( .A(w_mem_inst_w_mem_1__10_), .Y(w_mem_inst__abc_19396_new_n4201_));
INVX1 INVX1_1252 ( .A(\block[458] ), .Y(w_mem_inst__abc_19396_new_n4202_));
INVX1 INVX1_1253 ( .A(w_mem_inst_w_mem_1__11_), .Y(w_mem_inst__abc_19396_new_n4206_));
INVX1 INVX1_1254 ( .A(\block[459] ), .Y(w_mem_inst__abc_19396_new_n4207_));
INVX1 INVX1_1255 ( .A(w_mem_inst_w_mem_1__12_), .Y(w_mem_inst__abc_19396_new_n4211_));
INVX1 INVX1_1256 ( .A(\block[460] ), .Y(w_mem_inst__abc_19396_new_n4212_));
INVX1 INVX1_1257 ( .A(w_mem_inst_w_mem_1__13_), .Y(w_mem_inst__abc_19396_new_n4216_));
INVX1 INVX1_1258 ( .A(\block[461] ), .Y(w_mem_inst__abc_19396_new_n4217_));
INVX1 INVX1_1259 ( .A(w_mem_inst_w_mem_1__14_), .Y(w_mem_inst__abc_19396_new_n4221_));
INVX1 INVX1_126 ( .A(_abc_15497_new_n1275_), .Y(_abc_15497_new_n1282_));
INVX1 INVX1_1260 ( .A(\block[462] ), .Y(w_mem_inst__abc_19396_new_n4222_));
INVX1 INVX1_1261 ( .A(w_mem_inst_w_mem_1__15_), .Y(w_mem_inst__abc_19396_new_n4226_));
INVX1 INVX1_1262 ( .A(\block[463] ), .Y(w_mem_inst__abc_19396_new_n4227_));
INVX1 INVX1_1263 ( .A(w_mem_inst_w_mem_1__16_), .Y(w_mem_inst__abc_19396_new_n4231_));
INVX1 INVX1_1264 ( .A(\block[464] ), .Y(w_mem_inst__abc_19396_new_n4232_));
INVX1 INVX1_1265 ( .A(w_mem_inst_w_mem_1__17_), .Y(w_mem_inst__abc_19396_new_n4236_));
INVX1 INVX1_1266 ( .A(\block[465] ), .Y(w_mem_inst__abc_19396_new_n4237_));
INVX1 INVX1_1267 ( .A(w_mem_inst_w_mem_1__18_), .Y(w_mem_inst__abc_19396_new_n4241_));
INVX1 INVX1_1268 ( .A(\block[466] ), .Y(w_mem_inst__abc_19396_new_n4242_));
INVX1 INVX1_1269 ( .A(w_mem_inst_w_mem_1__19_), .Y(w_mem_inst__abc_19396_new_n4246_));
INVX1 INVX1_127 ( .A(_auto_iopadmap_cc_368_execute_22625_32_), .Y(_abc_15497_new_n1298_));
INVX1 INVX1_1270 ( .A(\block[467] ), .Y(w_mem_inst__abc_19396_new_n4247_));
INVX1 INVX1_1271 ( .A(w_mem_inst_w_mem_1__20_), .Y(w_mem_inst__abc_19396_new_n4251_));
INVX1 INVX1_1272 ( .A(\block[468] ), .Y(w_mem_inst__abc_19396_new_n4252_));
INVX1 INVX1_1273 ( .A(w_mem_inst_w_mem_1__21_), .Y(w_mem_inst__abc_19396_new_n4256_));
INVX1 INVX1_1274 ( .A(\block[469] ), .Y(w_mem_inst__abc_19396_new_n4257_));
INVX1 INVX1_1275 ( .A(w_mem_inst_w_mem_1__22_), .Y(w_mem_inst__abc_19396_new_n4261_));
INVX1 INVX1_1276 ( .A(\block[470] ), .Y(w_mem_inst__abc_19396_new_n4262_));
INVX1 INVX1_1277 ( .A(w_mem_inst_w_mem_1__23_), .Y(w_mem_inst__abc_19396_new_n4266_));
INVX1 INVX1_1278 ( .A(\block[471] ), .Y(w_mem_inst__abc_19396_new_n4267_));
INVX1 INVX1_1279 ( .A(w_mem_inst_w_mem_1__24_), .Y(w_mem_inst__abc_19396_new_n4271_));
INVX1 INVX1_128 ( .A(_auto_iopadmap_cc_368_execute_22625_33_), .Y(_abc_15497_new_n1307_));
INVX1 INVX1_1280 ( .A(\block[472] ), .Y(w_mem_inst__abc_19396_new_n4272_));
INVX1 INVX1_1281 ( .A(w_mem_inst_w_mem_1__25_), .Y(w_mem_inst__abc_19396_new_n4276_));
INVX1 INVX1_1282 ( .A(\block[473] ), .Y(w_mem_inst__abc_19396_new_n4277_));
INVX1 INVX1_1283 ( .A(w_mem_inst_w_mem_1__26_), .Y(w_mem_inst__abc_19396_new_n4281_));
INVX1 INVX1_1284 ( .A(\block[474] ), .Y(w_mem_inst__abc_19396_new_n4282_));
INVX1 INVX1_1285 ( .A(w_mem_inst_w_mem_1__27_), .Y(w_mem_inst__abc_19396_new_n4286_));
INVX1 INVX1_1286 ( .A(\block[475] ), .Y(w_mem_inst__abc_19396_new_n4287_));
INVX1 INVX1_1287 ( .A(w_mem_inst_w_mem_1__28_), .Y(w_mem_inst__abc_19396_new_n4291_));
INVX1 INVX1_1288 ( .A(\block[476] ), .Y(w_mem_inst__abc_19396_new_n4292_));
INVX1 INVX1_1289 ( .A(w_mem_inst_w_mem_1__29_), .Y(w_mem_inst__abc_19396_new_n4296_));
INVX1 INVX1_129 ( .A(_auto_iopadmap_cc_368_execute_22625_35_), .Y(_abc_15497_new_n1317_));
INVX1 INVX1_1290 ( .A(\block[477] ), .Y(w_mem_inst__abc_19396_new_n4297_));
INVX1 INVX1_1291 ( .A(w_mem_inst_w_mem_1__30_), .Y(w_mem_inst__abc_19396_new_n4301_));
INVX1 INVX1_1292 ( .A(\block[478] ), .Y(w_mem_inst__abc_19396_new_n4302_));
INVX1 INVX1_1293 ( .A(w_mem_inst_w_mem_1__31_), .Y(w_mem_inst__abc_19396_new_n4306_));
INVX1 INVX1_1294 ( .A(\block[479] ), .Y(w_mem_inst__abc_19396_new_n4307_));
INVX1 INVX1_1295 ( .A(w_mem_inst_w_mem_3__0_), .Y(w_mem_inst__abc_19396_new_n4311_));
INVX1 INVX1_1296 ( .A(\block[384] ), .Y(w_mem_inst__abc_19396_new_n4312_));
INVX1 INVX1_1297 ( .A(w_mem_inst_w_mem_3__1_), .Y(w_mem_inst__abc_19396_new_n4316_));
INVX1 INVX1_1298 ( .A(\block[385] ), .Y(w_mem_inst__abc_19396_new_n4317_));
INVX1 INVX1_1299 ( .A(w_mem_inst_w_mem_3__2_), .Y(w_mem_inst__abc_19396_new_n4321_));
INVX1 INVX1_13 ( .A(c_reg_9_), .Y(_abc_15497_new_n738_));
INVX1 INVX1_130 ( .A(_abc_15497_new_n1321_), .Y(_abc_15497_new_n1327_));
INVX1 INVX1_1300 ( .A(\block[386] ), .Y(w_mem_inst__abc_19396_new_n4322_));
INVX1 INVX1_1301 ( .A(w_mem_inst_w_mem_3__3_), .Y(w_mem_inst__abc_19396_new_n4326_));
INVX1 INVX1_1302 ( .A(\block[387] ), .Y(w_mem_inst__abc_19396_new_n4327_));
INVX1 INVX1_1303 ( .A(w_mem_inst_w_mem_3__4_), .Y(w_mem_inst__abc_19396_new_n4331_));
INVX1 INVX1_1304 ( .A(\block[388] ), .Y(w_mem_inst__abc_19396_new_n4332_));
INVX1 INVX1_1305 ( .A(w_mem_inst_w_mem_3__5_), .Y(w_mem_inst__abc_19396_new_n4336_));
INVX1 INVX1_1306 ( .A(\block[389] ), .Y(w_mem_inst__abc_19396_new_n4337_));
INVX1 INVX1_1307 ( .A(w_mem_inst_w_mem_3__6_), .Y(w_mem_inst__abc_19396_new_n4341_));
INVX1 INVX1_1308 ( .A(\block[390] ), .Y(w_mem_inst__abc_19396_new_n4342_));
INVX1 INVX1_1309 ( .A(w_mem_inst_w_mem_3__7_), .Y(w_mem_inst__abc_19396_new_n4346_));
INVX1 INVX1_131 ( .A(_auto_iopadmap_cc_368_execute_22625_36_), .Y(_abc_15497_new_n1332_));
INVX1 INVX1_1310 ( .A(\block[391] ), .Y(w_mem_inst__abc_19396_new_n4347_));
INVX1 INVX1_1311 ( .A(w_mem_inst_w_mem_3__8_), .Y(w_mem_inst__abc_19396_new_n4351_));
INVX1 INVX1_1312 ( .A(\block[392] ), .Y(w_mem_inst__abc_19396_new_n4352_));
INVX1 INVX1_1313 ( .A(w_mem_inst_w_mem_3__9_), .Y(w_mem_inst__abc_19396_new_n4356_));
INVX1 INVX1_1314 ( .A(\block[393] ), .Y(w_mem_inst__abc_19396_new_n4357_));
INVX1 INVX1_1315 ( .A(w_mem_inst_w_mem_3__10_), .Y(w_mem_inst__abc_19396_new_n4361_));
INVX1 INVX1_1316 ( .A(\block[394] ), .Y(w_mem_inst__abc_19396_new_n4362_));
INVX1 INVX1_1317 ( .A(w_mem_inst_w_mem_3__11_), .Y(w_mem_inst__abc_19396_new_n4366_));
INVX1 INVX1_1318 ( .A(\block[395] ), .Y(w_mem_inst__abc_19396_new_n4367_));
INVX1 INVX1_1319 ( .A(w_mem_inst_w_mem_3__12_), .Y(w_mem_inst__abc_19396_new_n4371_));
INVX1 INVX1_132 ( .A(_auto_iopadmap_cc_368_execute_22625_37_), .Y(_abc_15497_new_n1342_));
INVX1 INVX1_1320 ( .A(\block[396] ), .Y(w_mem_inst__abc_19396_new_n4372_));
INVX1 INVX1_1321 ( .A(w_mem_inst_w_mem_3__13_), .Y(w_mem_inst__abc_19396_new_n4376_));
INVX1 INVX1_1322 ( .A(\block[397] ), .Y(w_mem_inst__abc_19396_new_n4377_));
INVX1 INVX1_1323 ( .A(w_mem_inst_w_mem_3__14_), .Y(w_mem_inst__abc_19396_new_n4381_));
INVX1 INVX1_1324 ( .A(\block[398] ), .Y(w_mem_inst__abc_19396_new_n4382_));
INVX1 INVX1_1325 ( .A(w_mem_inst_w_mem_3__15_), .Y(w_mem_inst__abc_19396_new_n4386_));
INVX1 INVX1_1326 ( .A(\block[399] ), .Y(w_mem_inst__abc_19396_new_n4387_));
INVX1 INVX1_1327 ( .A(w_mem_inst_w_mem_3__16_), .Y(w_mem_inst__abc_19396_new_n4391_));
INVX1 INVX1_1328 ( .A(\block[400] ), .Y(w_mem_inst__abc_19396_new_n4392_));
INVX1 INVX1_1329 ( .A(w_mem_inst_w_mem_3__17_), .Y(w_mem_inst__abc_19396_new_n4396_));
INVX1 INVX1_133 ( .A(_auto_iopadmap_cc_368_execute_22625_39_), .Y(_abc_15497_new_n1351_));
INVX1 INVX1_1330 ( .A(\block[401] ), .Y(w_mem_inst__abc_19396_new_n4397_));
INVX1 INVX1_1331 ( .A(w_mem_inst_w_mem_3__18_), .Y(w_mem_inst__abc_19396_new_n4401_));
INVX1 INVX1_1332 ( .A(\block[402] ), .Y(w_mem_inst__abc_19396_new_n4402_));
INVX1 INVX1_1333 ( .A(w_mem_inst_w_mem_3__19_), .Y(w_mem_inst__abc_19396_new_n4406_));
INVX1 INVX1_1334 ( .A(\block[403] ), .Y(w_mem_inst__abc_19396_new_n4407_));
INVX1 INVX1_1335 ( .A(w_mem_inst_w_mem_3__20_), .Y(w_mem_inst__abc_19396_new_n4411_));
INVX1 INVX1_1336 ( .A(\block[404] ), .Y(w_mem_inst__abc_19396_new_n4412_));
INVX1 INVX1_1337 ( .A(w_mem_inst_w_mem_3__21_), .Y(w_mem_inst__abc_19396_new_n4416_));
INVX1 INVX1_1338 ( .A(\block[405] ), .Y(w_mem_inst__abc_19396_new_n4417_));
INVX1 INVX1_1339 ( .A(w_mem_inst_w_mem_3__22_), .Y(w_mem_inst__abc_19396_new_n4421_));
INVX1 INVX1_134 ( .A(_auto_iopadmap_cc_368_execute_22625_38_), .Y(_abc_15497_new_n1356_));
INVX1 INVX1_1340 ( .A(\block[406] ), .Y(w_mem_inst__abc_19396_new_n4422_));
INVX1 INVX1_1341 ( .A(w_mem_inst_w_mem_3__23_), .Y(w_mem_inst__abc_19396_new_n4426_));
INVX1 INVX1_1342 ( .A(\block[407] ), .Y(w_mem_inst__abc_19396_new_n4427_));
INVX1 INVX1_1343 ( .A(w_mem_inst_w_mem_3__24_), .Y(w_mem_inst__abc_19396_new_n4431_));
INVX1 INVX1_1344 ( .A(\block[408] ), .Y(w_mem_inst__abc_19396_new_n4432_));
INVX1 INVX1_1345 ( .A(w_mem_inst_w_mem_3__25_), .Y(w_mem_inst__abc_19396_new_n4436_));
INVX1 INVX1_1346 ( .A(\block[409] ), .Y(w_mem_inst__abc_19396_new_n4437_));
INVX1 INVX1_1347 ( .A(w_mem_inst_w_mem_3__26_), .Y(w_mem_inst__abc_19396_new_n4441_));
INVX1 INVX1_1348 ( .A(\block[410] ), .Y(w_mem_inst__abc_19396_new_n4442_));
INVX1 INVX1_1349 ( .A(w_mem_inst_w_mem_3__27_), .Y(w_mem_inst__abc_19396_new_n4446_));
INVX1 INVX1_135 ( .A(_auto_iopadmap_cc_368_execute_22625_41_), .Y(_abc_15497_new_n1371_));
INVX1 INVX1_1350 ( .A(\block[411] ), .Y(w_mem_inst__abc_19396_new_n4447_));
INVX1 INVX1_1351 ( .A(w_mem_inst_w_mem_3__28_), .Y(w_mem_inst__abc_19396_new_n4451_));
INVX1 INVX1_1352 ( .A(\block[412] ), .Y(w_mem_inst__abc_19396_new_n4452_));
INVX1 INVX1_1353 ( .A(w_mem_inst_w_mem_3__29_), .Y(w_mem_inst__abc_19396_new_n4456_));
INVX1 INVX1_1354 ( .A(\block[413] ), .Y(w_mem_inst__abc_19396_new_n4457_));
INVX1 INVX1_1355 ( .A(w_mem_inst_w_mem_3__30_), .Y(w_mem_inst__abc_19396_new_n4461_));
INVX1 INVX1_1356 ( .A(\block[414] ), .Y(w_mem_inst__abc_19396_new_n4462_));
INVX1 INVX1_1357 ( .A(w_mem_inst_w_mem_3__31_), .Y(w_mem_inst__abc_19396_new_n4466_));
INVX1 INVX1_1358 ( .A(\block[415] ), .Y(w_mem_inst__abc_19396_new_n4467_));
INVX1 INVX1_1359 ( .A(w_mem_inst_w_mem_2__0_), .Y(w_mem_inst__abc_19396_new_n4471_));
INVX1 INVX1_136 ( .A(_abc_15497_new_n1376_), .Y(_abc_15497_new_n1377_));
INVX1 INVX1_1360 ( .A(\block[416] ), .Y(w_mem_inst__abc_19396_new_n4472_));
INVX1 INVX1_1361 ( .A(w_mem_inst_w_mem_2__1_), .Y(w_mem_inst__abc_19396_new_n4476_));
INVX1 INVX1_1362 ( .A(\block[417] ), .Y(w_mem_inst__abc_19396_new_n4477_));
INVX1 INVX1_1363 ( .A(w_mem_inst_w_mem_2__2_), .Y(w_mem_inst__abc_19396_new_n4481_));
INVX1 INVX1_1364 ( .A(\block[418] ), .Y(w_mem_inst__abc_19396_new_n4482_));
INVX1 INVX1_1365 ( .A(w_mem_inst_w_mem_2__3_), .Y(w_mem_inst__abc_19396_new_n4486_));
INVX1 INVX1_1366 ( .A(\block[419] ), .Y(w_mem_inst__abc_19396_new_n4487_));
INVX1 INVX1_1367 ( .A(w_mem_inst_w_mem_2__4_), .Y(w_mem_inst__abc_19396_new_n4491_));
INVX1 INVX1_1368 ( .A(\block[420] ), .Y(w_mem_inst__abc_19396_new_n4492_));
INVX1 INVX1_1369 ( .A(w_mem_inst_w_mem_2__5_), .Y(w_mem_inst__abc_19396_new_n4496_));
INVX1 INVX1_137 ( .A(_abc_15497_new_n1382_), .Y(_abc_15497_new_n1383_));
INVX1 INVX1_1370 ( .A(\block[421] ), .Y(w_mem_inst__abc_19396_new_n4497_));
INVX1 INVX1_1371 ( .A(w_mem_inst_w_mem_2__6_), .Y(w_mem_inst__abc_19396_new_n4501_));
INVX1 INVX1_1372 ( .A(\block[422] ), .Y(w_mem_inst__abc_19396_new_n4502_));
INVX1 INVX1_1373 ( .A(w_mem_inst_w_mem_2__7_), .Y(w_mem_inst__abc_19396_new_n4506_));
INVX1 INVX1_1374 ( .A(\block[423] ), .Y(w_mem_inst__abc_19396_new_n4507_));
INVX1 INVX1_1375 ( .A(w_mem_inst_w_mem_2__8_), .Y(w_mem_inst__abc_19396_new_n4511_));
INVX1 INVX1_1376 ( .A(\block[424] ), .Y(w_mem_inst__abc_19396_new_n4512_));
INVX1 INVX1_1377 ( .A(w_mem_inst_w_mem_2__9_), .Y(w_mem_inst__abc_19396_new_n4516_));
INVX1 INVX1_1378 ( .A(\block[425] ), .Y(w_mem_inst__abc_19396_new_n4517_));
INVX1 INVX1_1379 ( .A(w_mem_inst_w_mem_2__10_), .Y(w_mem_inst__abc_19396_new_n4521_));
INVX1 INVX1_138 ( .A(_abc_15497_new_n1387_), .Y(_abc_15497_new_n1388_));
INVX1 INVX1_1380 ( .A(\block[426] ), .Y(w_mem_inst__abc_19396_new_n4522_));
INVX1 INVX1_1381 ( .A(w_mem_inst_w_mem_2__11_), .Y(w_mem_inst__abc_19396_new_n4526_));
INVX1 INVX1_1382 ( .A(\block[427] ), .Y(w_mem_inst__abc_19396_new_n4527_));
INVX1 INVX1_1383 ( .A(w_mem_inst_w_mem_2__12_), .Y(w_mem_inst__abc_19396_new_n4531_));
INVX1 INVX1_1384 ( .A(\block[428] ), .Y(w_mem_inst__abc_19396_new_n4532_));
INVX1 INVX1_1385 ( .A(w_mem_inst_w_mem_2__13_), .Y(w_mem_inst__abc_19396_new_n4536_));
INVX1 INVX1_1386 ( .A(\block[429] ), .Y(w_mem_inst__abc_19396_new_n4537_));
INVX1 INVX1_1387 ( .A(w_mem_inst_w_mem_2__14_), .Y(w_mem_inst__abc_19396_new_n4541_));
INVX1 INVX1_1388 ( .A(\block[430] ), .Y(w_mem_inst__abc_19396_new_n4542_));
INVX1 INVX1_1389 ( .A(w_mem_inst_w_mem_2__15_), .Y(w_mem_inst__abc_19396_new_n4546_));
INVX1 INVX1_139 ( .A(_auto_iopadmap_cc_368_execute_22625_43_), .Y(_abc_15497_new_n1395_));
INVX1 INVX1_1390 ( .A(\block[431] ), .Y(w_mem_inst__abc_19396_new_n4547_));
INVX1 INVX1_1391 ( .A(w_mem_inst_w_mem_2__16_), .Y(w_mem_inst__abc_19396_new_n4551_));
INVX1 INVX1_1392 ( .A(\block[432] ), .Y(w_mem_inst__abc_19396_new_n4552_));
INVX1 INVX1_1393 ( .A(w_mem_inst_w_mem_2__17_), .Y(w_mem_inst__abc_19396_new_n4556_));
INVX1 INVX1_1394 ( .A(\block[433] ), .Y(w_mem_inst__abc_19396_new_n4557_));
INVX1 INVX1_1395 ( .A(w_mem_inst_w_mem_2__18_), .Y(w_mem_inst__abc_19396_new_n4561_));
INVX1 INVX1_1396 ( .A(\block[434] ), .Y(w_mem_inst__abc_19396_new_n4562_));
INVX1 INVX1_1397 ( .A(w_mem_inst_w_mem_2__19_), .Y(w_mem_inst__abc_19396_new_n4566_));
INVX1 INVX1_1398 ( .A(\block[435] ), .Y(w_mem_inst__abc_19396_new_n4567_));
INVX1 INVX1_1399 ( .A(w_mem_inst_w_mem_2__20_), .Y(w_mem_inst__abc_19396_new_n4571_));
INVX1 INVX1_14 ( .A(_auto_iopadmap_cc_368_execute_22625_73_), .Y(_abc_15497_new_n739_));
INVX1 INVX1_140 ( .A(_abc_15497_new_n1400_), .Y(_abc_15497_new_n1401_));
INVX1 INVX1_1400 ( .A(\block[436] ), .Y(w_mem_inst__abc_19396_new_n4572_));
INVX1 INVX1_1401 ( .A(w_mem_inst_w_mem_2__21_), .Y(w_mem_inst__abc_19396_new_n4576_));
INVX1 INVX1_1402 ( .A(\block[437] ), .Y(w_mem_inst__abc_19396_new_n4577_));
INVX1 INVX1_1403 ( .A(w_mem_inst_w_mem_2__22_), .Y(w_mem_inst__abc_19396_new_n4581_));
INVX1 INVX1_1404 ( .A(\block[438] ), .Y(w_mem_inst__abc_19396_new_n4582_));
INVX1 INVX1_1405 ( .A(w_mem_inst_w_mem_2__23_), .Y(w_mem_inst__abc_19396_new_n4586_));
INVX1 INVX1_1406 ( .A(\block[439] ), .Y(w_mem_inst__abc_19396_new_n4587_));
INVX1 INVX1_1407 ( .A(w_mem_inst_w_mem_2__24_), .Y(w_mem_inst__abc_19396_new_n4591_));
INVX1 INVX1_1408 ( .A(\block[440] ), .Y(w_mem_inst__abc_19396_new_n4592_));
INVX1 INVX1_1409 ( .A(w_mem_inst_w_mem_2__25_), .Y(w_mem_inst__abc_19396_new_n4596_));
INVX1 INVX1_141 ( .A(_abc_15497_new_n1406_), .Y(_abc_15497_new_n1407_));
INVX1 INVX1_1410 ( .A(\block[441] ), .Y(w_mem_inst__abc_19396_new_n4597_));
INVX1 INVX1_1411 ( .A(w_mem_inst_w_mem_2__26_), .Y(w_mem_inst__abc_19396_new_n4601_));
INVX1 INVX1_1412 ( .A(\block[442] ), .Y(w_mem_inst__abc_19396_new_n4602_));
INVX1 INVX1_1413 ( .A(w_mem_inst_w_mem_2__27_), .Y(w_mem_inst__abc_19396_new_n4606_));
INVX1 INVX1_1414 ( .A(\block[443] ), .Y(w_mem_inst__abc_19396_new_n4607_));
INVX1 INVX1_1415 ( .A(w_mem_inst_w_mem_2__28_), .Y(w_mem_inst__abc_19396_new_n4611_));
INVX1 INVX1_1416 ( .A(\block[444] ), .Y(w_mem_inst__abc_19396_new_n4612_));
INVX1 INVX1_1417 ( .A(w_mem_inst_w_mem_2__29_), .Y(w_mem_inst__abc_19396_new_n4616_));
INVX1 INVX1_1418 ( .A(\block[445] ), .Y(w_mem_inst__abc_19396_new_n4617_));
INVX1 INVX1_1419 ( .A(w_mem_inst_w_mem_2__30_), .Y(w_mem_inst__abc_19396_new_n4621_));
INVX1 INVX1_142 ( .A(_abc_15497_new_n1409_), .Y(_abc_15497_new_n1410_));
INVX1 INVX1_1420 ( .A(\block[446] ), .Y(w_mem_inst__abc_19396_new_n4622_));
INVX1 INVX1_1421 ( .A(w_mem_inst_w_mem_2__31_), .Y(w_mem_inst__abc_19396_new_n4626_));
INVX1 INVX1_1422 ( .A(\block[447] ), .Y(w_mem_inst__abc_19396_new_n4627_));
INVX1 INVX1_1423 ( .A(w_mem_inst_w_mem_0__0_), .Y(w_mem_inst__abc_19396_new_n4631_));
INVX1 INVX1_1424 ( .A(\block[480] ), .Y(w_mem_inst__abc_19396_new_n4632_));
INVX1 INVX1_1425 ( .A(w_mem_inst_w_mem_0__1_), .Y(w_mem_inst__abc_19396_new_n4636_));
INVX1 INVX1_1426 ( .A(\block[481] ), .Y(w_mem_inst__abc_19396_new_n4637_));
INVX1 INVX1_1427 ( .A(w_mem_inst_w_mem_0__2_), .Y(w_mem_inst__abc_19396_new_n4641_));
INVX1 INVX1_1428 ( .A(\block[482] ), .Y(w_mem_inst__abc_19396_new_n4642_));
INVX1 INVX1_1429 ( .A(w_mem_inst_w_mem_0__3_), .Y(w_mem_inst__abc_19396_new_n4646_));
INVX1 INVX1_143 ( .A(_auto_iopadmap_cc_368_execute_22625_44_), .Y(_abc_15497_new_n1413_));
INVX1 INVX1_1430 ( .A(\block[483] ), .Y(w_mem_inst__abc_19396_new_n4647_));
INVX1 INVX1_1431 ( .A(w_mem_inst_w_mem_0__4_), .Y(w_mem_inst__abc_19396_new_n4651_));
INVX1 INVX1_1432 ( .A(\block[484] ), .Y(w_mem_inst__abc_19396_new_n4652_));
INVX1 INVX1_1433 ( .A(w_mem_inst_w_mem_0__5_), .Y(w_mem_inst__abc_19396_new_n4656_));
INVX1 INVX1_1434 ( .A(\block[485] ), .Y(w_mem_inst__abc_19396_new_n4657_));
INVX1 INVX1_1435 ( .A(w_mem_inst_w_mem_0__6_), .Y(w_mem_inst__abc_19396_new_n4661_));
INVX1 INVX1_1436 ( .A(\block[486] ), .Y(w_mem_inst__abc_19396_new_n4662_));
INVX1 INVX1_1437 ( .A(w_mem_inst_w_mem_0__7_), .Y(w_mem_inst__abc_19396_new_n4666_));
INVX1 INVX1_1438 ( .A(\block[487] ), .Y(w_mem_inst__abc_19396_new_n4667_));
INVX1 INVX1_1439 ( .A(w_mem_inst_w_mem_0__8_), .Y(w_mem_inst__abc_19396_new_n4671_));
INVX1 INVX1_144 ( .A(_auto_iopadmap_cc_368_execute_22625_45_), .Y(_abc_15497_new_n1422_));
INVX1 INVX1_1440 ( .A(\block[488] ), .Y(w_mem_inst__abc_19396_new_n4672_));
INVX1 INVX1_1441 ( .A(w_mem_inst_w_mem_0__9_), .Y(w_mem_inst__abc_19396_new_n4676_));
INVX1 INVX1_1442 ( .A(\block[489] ), .Y(w_mem_inst__abc_19396_new_n4677_));
INVX1 INVX1_1443 ( .A(w_mem_inst_w_mem_0__10_), .Y(w_mem_inst__abc_19396_new_n4681_));
INVX1 INVX1_1444 ( .A(\block[490] ), .Y(w_mem_inst__abc_19396_new_n4682_));
INVX1 INVX1_1445 ( .A(w_mem_inst_w_mem_0__11_), .Y(w_mem_inst__abc_19396_new_n4686_));
INVX1 INVX1_1446 ( .A(\block[491] ), .Y(w_mem_inst__abc_19396_new_n4687_));
INVX1 INVX1_1447 ( .A(w_mem_inst_w_mem_0__12_), .Y(w_mem_inst__abc_19396_new_n4691_));
INVX1 INVX1_1448 ( .A(\block[492] ), .Y(w_mem_inst__abc_19396_new_n4692_));
INVX1 INVX1_1449 ( .A(w_mem_inst_w_mem_0__13_), .Y(w_mem_inst__abc_19396_new_n4696_));
INVX1 INVX1_145 ( .A(_abc_15497_new_n1418_), .Y(_abc_15497_new_n1423_));
INVX1 INVX1_1450 ( .A(\block[493] ), .Y(w_mem_inst__abc_19396_new_n4697_));
INVX1 INVX1_1451 ( .A(w_mem_inst_w_mem_0__14_), .Y(w_mem_inst__abc_19396_new_n4701_));
INVX1 INVX1_1452 ( .A(\block[494] ), .Y(w_mem_inst__abc_19396_new_n4702_));
INVX1 INVX1_1453 ( .A(w_mem_inst_w_mem_0__15_), .Y(w_mem_inst__abc_19396_new_n4706_));
INVX1 INVX1_1454 ( .A(\block[495] ), .Y(w_mem_inst__abc_19396_new_n4707_));
INVX1 INVX1_1455 ( .A(w_mem_inst_w_mem_0__16_), .Y(w_mem_inst__abc_19396_new_n4711_));
INVX1 INVX1_1456 ( .A(\block[496] ), .Y(w_mem_inst__abc_19396_new_n4712_));
INVX1 INVX1_1457 ( .A(w_mem_inst_w_mem_0__17_), .Y(w_mem_inst__abc_19396_new_n4716_));
INVX1 INVX1_1458 ( .A(\block[497] ), .Y(w_mem_inst__abc_19396_new_n4717_));
INVX1 INVX1_1459 ( .A(w_mem_inst_w_mem_0__18_), .Y(w_mem_inst__abc_19396_new_n4721_));
INVX1 INVX1_146 ( .A(_abc_15497_new_n1432_), .Y(_abc_15497_new_n1433_));
INVX1 INVX1_1460 ( .A(\block[498] ), .Y(w_mem_inst__abc_19396_new_n4722_));
INVX1 INVX1_1461 ( .A(w_mem_inst_w_mem_0__19_), .Y(w_mem_inst__abc_19396_new_n4726_));
INVX1 INVX1_1462 ( .A(\block[499] ), .Y(w_mem_inst__abc_19396_new_n4727_));
INVX1 INVX1_1463 ( .A(w_mem_inst_w_mem_0__20_), .Y(w_mem_inst__abc_19396_new_n4731_));
INVX1 INVX1_1464 ( .A(\block[500] ), .Y(w_mem_inst__abc_19396_new_n4732_));
INVX1 INVX1_1465 ( .A(w_mem_inst_w_mem_0__21_), .Y(w_mem_inst__abc_19396_new_n4736_));
INVX1 INVX1_1466 ( .A(\block[501] ), .Y(w_mem_inst__abc_19396_new_n4737_));
INVX1 INVX1_1467 ( .A(w_mem_inst_w_mem_0__22_), .Y(w_mem_inst__abc_19396_new_n4741_));
INVX1 INVX1_1468 ( .A(\block[502] ), .Y(w_mem_inst__abc_19396_new_n4742_));
INVX1 INVX1_1469 ( .A(w_mem_inst_w_mem_0__23_), .Y(w_mem_inst__abc_19396_new_n4746_));
INVX1 INVX1_147 ( .A(_abc_15497_new_n1436_), .Y(_abc_15497_new_n1437_));
INVX1 INVX1_1470 ( .A(\block[503] ), .Y(w_mem_inst__abc_19396_new_n4747_));
INVX1 INVX1_1471 ( .A(w_mem_inst_w_mem_0__24_), .Y(w_mem_inst__abc_19396_new_n4751_));
INVX1 INVX1_1472 ( .A(\block[504] ), .Y(w_mem_inst__abc_19396_new_n4752_));
INVX1 INVX1_1473 ( .A(w_mem_inst_w_mem_0__25_), .Y(w_mem_inst__abc_19396_new_n4756_));
INVX1 INVX1_1474 ( .A(\block[505] ), .Y(w_mem_inst__abc_19396_new_n4757_));
INVX1 INVX1_1475 ( .A(w_mem_inst_w_mem_0__26_), .Y(w_mem_inst__abc_19396_new_n4761_));
INVX1 INVX1_1476 ( .A(\block[506] ), .Y(w_mem_inst__abc_19396_new_n4762_));
INVX1 INVX1_1477 ( .A(w_mem_inst_w_mem_0__27_), .Y(w_mem_inst__abc_19396_new_n4766_));
INVX1 INVX1_1478 ( .A(\block[507] ), .Y(w_mem_inst__abc_19396_new_n4767_));
INVX1 INVX1_1479 ( .A(w_mem_inst_w_mem_0__28_), .Y(w_mem_inst__abc_19396_new_n4771_));
INVX1 INVX1_148 ( .A(_abc_15497_new_n1438_), .Y(_abc_15497_new_n1439_));
INVX1 INVX1_1480 ( .A(\block[508] ), .Y(w_mem_inst__abc_19396_new_n4772_));
INVX1 INVX1_1481 ( .A(w_mem_inst_w_mem_0__29_), .Y(w_mem_inst__abc_19396_new_n4776_));
INVX1 INVX1_1482 ( .A(\block[509] ), .Y(w_mem_inst__abc_19396_new_n4777_));
INVX1 INVX1_1483 ( .A(w_mem_inst_w_mem_0__30_), .Y(w_mem_inst__abc_19396_new_n4781_));
INVX1 INVX1_1484 ( .A(\block[510] ), .Y(w_mem_inst__abc_19396_new_n4782_));
INVX1 INVX1_1485 ( .A(w_mem_inst_w_mem_0__31_), .Y(w_mem_inst__abc_19396_new_n4786_));
INVX1 INVX1_1486 ( .A(\block[511] ), .Y(w_mem_inst__abc_19396_new_n4787_));
INVX1 INVX1_1487 ( .A(w_mem_inst_w_ctr_reg_4_), .Y(w_mem_inst__abc_19396_new_n4804_));
INVX1 INVX1_149 ( .A(_auto_iopadmap_cc_368_execute_22625_47_), .Y(_abc_15497_new_n1444_));
INVX1 INVX1_15 ( .A(c_reg_8_), .Y(_abc_15497_new_n741_));
INVX1 INVX1_150 ( .A(_auto_iopadmap_cc_368_execute_22625_48_), .Y(_abc_15497_new_n1452_));
INVX1 INVX1_151 ( .A(_abc_15497_new_n1469_), .Y(_abc_15497_new_n1470_));
INVX1 INVX1_152 ( .A(_auto_iopadmap_cc_368_execute_22625_50_), .Y(_abc_15497_new_n1477_));
INVX1 INVX1_153 ( .A(_abc_15497_new_n1478_), .Y(_abc_15497_new_n1479_));
INVX1 INVX1_154 ( .A(_abc_15497_new_n1480_), .Y(_abc_15497_new_n1481_));
INVX1 INVX1_155 ( .A(_abc_15497_new_n1482_), .Y(_abc_15497_new_n1483_));
INVX1 INVX1_156 ( .A(d_reg_18_), .Y(_abc_15497_new_n1485_));
INVX1 INVX1_157 ( .A(_abc_15497_new_n1487_), .Y(_abc_15497_new_n1489_));
INVX1 INVX1_158 ( .A(_auto_iopadmap_cc_368_execute_22625_51_), .Y(_abc_15497_new_n1492_));
INVX1 INVX1_159 ( .A(_abc_15497_new_n1497_), .Y(_abc_15497_new_n1498_));
INVX1 INVX1_16 ( .A(_auto_iopadmap_cc_368_execute_22625_72_), .Y(_abc_15497_new_n742_));
INVX1 INVX1_160 ( .A(_abc_15497_new_n1502_), .Y(_abc_15497_new_n1503_));
INVX1 INVX1_161 ( .A(_abc_15497_new_n1507_), .Y(_abc_15497_new_n1508_));
INVX1 INVX1_162 ( .A(_auto_iopadmap_cc_368_execute_22625_52_), .Y(_abc_15497_new_n1510_));
INVX1 INVX1_163 ( .A(_abc_15497_new_n1513_), .Y(_abc_15497_new_n1515_));
INVX1 INVX1_164 ( .A(_abc_15497_new_n1512_), .Y(_abc_15497_new_n1519_));
INVX1 INVX1_165 ( .A(_abc_15497_new_n1521_), .Y(_abc_15497_new_n1522_));
INVX1 INVX1_166 ( .A(_auto_iopadmap_cc_368_execute_22625_55_), .Y(_abc_15497_new_n1540_));
INVX1 INVX1_167 ( .A(_abc_15497_new_n1506_), .Y(_abc_15497_new_n1551_));
INVX1 INVX1_168 ( .A(_abc_15497_new_n1504_), .Y(_abc_15497_new_n1557_));
INVX1 INVX1_169 ( .A(_abc_15497_new_n1559_), .Y(_abc_15497_new_n1560_));
INVX1 INVX1_17 ( .A(c_reg_6_), .Y(_abc_15497_new_n748_));
INVX1 INVX1_170 ( .A(_abc_15497_new_n1564_), .Y(_abc_15497_new_n1566_));
INVX1 INVX1_171 ( .A(_auto_iopadmap_cc_368_execute_22625_57_), .Y(_abc_15497_new_n1569_));
INVX1 INVX1_172 ( .A(_abc_15497_new_n1574_), .Y(_abc_15497_new_n1575_));
INVX1 INVX1_173 ( .A(_abc_15497_new_n1582_), .Y(_abc_15497_new_n1583_));
INVX1 INVX1_174 ( .A(_auto_iopadmap_cc_368_execute_22625_59_), .Y(_abc_15497_new_n1593_));
INVX1 INVX1_175 ( .A(_abc_15497_new_n1598_), .Y(_abc_15497_new_n1599_));
INVX1 INVX1_176 ( .A(_abc_15497_new_n1604_), .Y(_abc_15497_new_n1606_));
INVX1 INVX1_177 ( .A(_abc_15497_new_n1608_), .Y(_abc_15497_new_n1609_));
INVX1 INVX1_178 ( .A(_auto_iopadmap_cc_368_execute_22625_61_), .Y(_abc_15497_new_n1621_));
INVX1 INVX1_179 ( .A(d_reg_29_), .Y(_abc_15497_new_n1622_));
INVX1 INVX1_18 ( .A(_auto_iopadmap_cc_368_execute_22625_70_), .Y(_abc_15497_new_n749_));
INVX1 INVX1_180 ( .A(_auto_iopadmap_cc_368_execute_22625_62_), .Y(_abc_15497_new_n1628_));
INVX1 INVX1_181 ( .A(_abc_15497_new_n1629_), .Y(_abc_15497_new_n1630_));
INVX1 INVX1_182 ( .A(_abc_15497_new_n1623_), .Y(_abc_15497_new_n1631_));
INVX1 INVX1_183 ( .A(_auto_iopadmap_cc_368_execute_22625_63_), .Y(_abc_15497_new_n1637_));
INVX1 INVX1_184 ( .A(e_reg_11_), .Y(_abc_15497_new_n1684_));
INVX1 INVX1_185 ( .A(e_reg_28_), .Y(_abc_15497_new_n1736_));
INVX1 INVX1_186 ( .A(_auto_iopadmap_cc_368_execute_22625_96_), .Y(_abc_15497_new_n1751_));
INVX1 INVX1_187 ( .A(_auto_iopadmap_cc_368_execute_22625_97_), .Y(_abc_15497_new_n1756_));
INVX1 INVX1_188 ( .A(_auto_iopadmap_cc_368_execute_22625_98_), .Y(_abc_15497_new_n1762_));
INVX1 INVX1_189 ( .A(b_reg_1_), .Y(_abc_15497_new_n1763_));
INVX1 INVX1_19 ( .A(_abc_15497_new_n753_), .Y(_abc_15497_new_n754_));
INVX1 INVX1_190 ( .A(_abc_15497_new_n1767_), .Y(_abc_15497_new_n1768_));
INVX1 INVX1_191 ( .A(b_reg_2_), .Y(_abc_15497_new_n1771_));
INVX1 INVX1_192 ( .A(_auto_iopadmap_cc_368_execute_22625_100_), .Y(_abc_15497_new_n1779_));
INVX1 INVX1_193 ( .A(_abc_15497_new_n1773_), .Y(_abc_15497_new_n1781_));
INVX1 INVX1_194 ( .A(b_reg_4_), .Y(_abc_15497_new_n1788_));
INVX1 INVX1_195 ( .A(b_reg_5_), .Y(_abc_15497_new_n1792_));
INVX1 INVX1_196 ( .A(_auto_iopadmap_cc_368_execute_22625_102_), .Y(_abc_15497_new_n1799_));
INVX1 INVX1_197 ( .A(b_reg_6_), .Y(_abc_15497_new_n1802_));
INVX1 INVX1_198 ( .A(_abc_15497_new_n1809_), .Y(_abc_15497_new_n1810_));
INVX1 INVX1_199 ( .A(_abc_15497_new_n1812_), .Y(_abc_15497_new_n1813_));
INVX1 INVX1_2 ( .A(c_reg_13_), .Y(_abc_15497_new_n708_));
INVX1 INVX1_20 ( .A(_abc_15497_new_n757_), .Y(_abc_15497_new_n758_));
INVX1 INVX1_200 ( .A(_auto_iopadmap_cc_368_execute_22625_104_), .Y(_abc_15497_new_n1819_));
INVX1 INVX1_201 ( .A(b_reg_8_), .Y(_abc_15497_new_n1820_));
INVX1 INVX1_202 ( .A(b_reg_10_), .Y(_abc_15497_new_n1841_));
INVX1 INVX1_203 ( .A(_abc_15497_new_n1850_), .Y(_abc_15497_new_n1851_));
INVX1 INVX1_204 ( .A(_auto_iopadmap_cc_368_execute_22625_108_), .Y(_abc_15497_new_n1856_));
INVX1 INVX1_205 ( .A(b_reg_12_), .Y(_abc_15497_new_n1858_));
INVX1 INVX1_206 ( .A(_abc_15497_new_n1859_), .Y(_abc_15497_new_n1868_));
INVX1 INVX1_207 ( .A(_auto_iopadmap_cc_368_execute_22625_110_), .Y(_abc_15497_new_n1874_));
INVX1 INVX1_208 ( .A(b_reg_14_), .Y(_abc_15497_new_n1876_));
INVX1 INVX1_209 ( .A(_abc_15497_new_n1878_), .Y(_abc_15497_new_n1879_));
INVX1 INVX1_21 ( .A(c_reg_5_), .Y(_abc_15497_new_n759_));
INVX1 INVX1_210 ( .A(_auto_iopadmap_cc_368_execute_22625_109_), .Y(_abc_15497_new_n1880_));
INVX1 INVX1_211 ( .A(b_reg_13_), .Y(_abc_15497_new_n1881_));
INVX1 INVX1_212 ( .A(_abc_15497_new_n1877_), .Y(_abc_15497_new_n1890_));
INVX1 INVX1_213 ( .A(_abc_15497_new_n1893_), .Y(_abc_15497_new_n1894_));
INVX1 INVX1_214 ( .A(_auto_iopadmap_cc_368_execute_22625_112_), .Y(_abc_15497_new_n1907_));
INVX1 INVX1_215 ( .A(b_reg_17_), .Y(_abc_15497_new_n1918_));
INVX1 INVX1_216 ( .A(_abc_15497_new_n1920_), .Y(_abc_15497_new_n1924_));
INVX1 INVX1_217 ( .A(_abc_15497_new_n1930_), .Y(_abc_15497_new_n1931_));
INVX1 INVX1_218 ( .A(_abc_15497_new_n1940_), .Y(_abc_15497_new_n1941_));
INVX1 INVX1_219 ( .A(_abc_15497_new_n1942_), .Y(_abc_15497_new_n1943_));
INVX1 INVX1_22 ( .A(_auto_iopadmap_cc_368_execute_22625_69_), .Y(_abc_15497_new_n760_));
INVX1 INVX1_220 ( .A(_auto_iopadmap_cc_368_execute_22625_116_), .Y(_abc_15497_new_n1949_));
INVX1 INVX1_221 ( .A(b_reg_20_), .Y(_abc_15497_new_n1958_));
INVX1 INVX1_222 ( .A(_abc_15497_new_n1960_), .Y(_abc_15497_new_n1961_));
INVX1 INVX1_223 ( .A(_auto_iopadmap_cc_368_execute_22625_117_), .Y(_abc_15497_new_n1965_));
INVX1 INVX1_224 ( .A(b_reg_21_), .Y(_abc_15497_new_n1967_));
INVX1 INVX1_225 ( .A(_abc_15497_new_n1959_), .Y(_abc_15497_new_n1970_));
INVX1 INVX1_226 ( .A(_abc_15497_new_n1969_), .Y(_abc_15497_new_n1974_));
INVX1 INVX1_227 ( .A(_abc_15497_new_n1975_), .Y(_abc_15497_new_n1976_));
INVX1 INVX1_228 ( .A(_abc_15497_new_n1980_), .Y(_abc_15497_new_n1981_));
INVX1 INVX1_229 ( .A(_abc_15497_new_n1988_), .Y(_abc_15497_new_n1989_));
INVX1 INVX1_23 ( .A(_abc_15497_new_n761_), .Y(_abc_15497_new_n762_));
INVX1 INVX1_230 ( .A(_abc_15497_new_n1996_), .Y(_abc_15497_new_n1997_));
INVX1 INVX1_231 ( .A(_abc_15497_new_n2000_), .Y(_abc_15497_new_n2001_));
INVX1 INVX1_232 ( .A(_auto_iopadmap_cc_368_execute_22625_120_), .Y(_abc_15497_new_n2005_));
INVX1 INVX1_233 ( .A(b_reg_24_), .Y(_abc_15497_new_n2006_));
INVX1 INVX1_234 ( .A(_abc_15497_new_n2008_), .Y(_abc_15497_new_n2009_));
INVX1 INVX1_235 ( .A(_abc_15497_new_n2007_), .Y(_abc_15497_new_n2014_));
INVX1 INVX1_236 ( .A(_abc_15497_new_n2017_), .Y(_abc_15497_new_n2018_));
INVX1 INVX1_237 ( .A(_abc_15497_new_n2019_), .Y(_abc_15497_new_n2023_));
INVX1 INVX1_238 ( .A(_abc_15497_new_n2024_), .Y(_abc_15497_new_n2025_));
INVX1 INVX1_239 ( .A(_abc_15497_new_n2026_), .Y(_abc_15497_new_n2027_));
INVX1 INVX1_24 ( .A(_abc_15497_new_n745_), .Y(_abc_15497_new_n784_));
INVX1 INVX1_240 ( .A(_auto_iopadmap_cc_368_execute_22625_122_), .Y(_abc_15497_new_n2030_));
INVX1 INVX1_241 ( .A(_abc_15497_new_n2041_), .Y(_abc_15497_new_n2042_));
INVX1 INVX1_242 ( .A(_auto_iopadmap_cc_368_execute_22625_124_), .Y(_abc_15497_new_n2047_));
INVX1 INVX1_243 ( .A(_abc_15497_new_n2032_), .Y(_abc_15497_new_n2050_));
INVX1 INVX1_244 ( .A(b_reg_28_), .Y(_abc_15497_new_n2054_));
INVX1 INVX1_245 ( .A(_abc_15497_new_n2053_), .Y(_abc_15497_new_n2058_));
INVX1 INVX1_246 ( .A(_abc_15497_new_n2065_), .Y(_abc_15497_new_n2066_));
INVX1 INVX1_247 ( .A(_abc_15497_new_n2067_), .Y(_abc_15497_new_n2068_));
INVX1 INVX1_248 ( .A(_abc_15497_new_n2072_), .Y(_abc_15497_new_n2073_));
INVX1 INVX1_249 ( .A(_abc_15497_new_n2083_), .Y(_abc_15497_new_n2086_));
INVX1 INVX1_25 ( .A(_abc_15497_new_n786_), .Y(_abc_15497_new_n787_));
INVX1 INVX1_250 ( .A(_auto_iopadmap_cc_368_execute_22625_128_), .Y(_abc_15497_new_n2092_));
INVX1 INVX1_251 ( .A(a_reg_0_), .Y(_abc_15497_new_n2093_));
INVX1 INVX1_252 ( .A(_auto_iopadmap_cc_368_execute_22625_129_), .Y(_abc_15497_new_n2097_));
INVX1 INVX1_253 ( .A(_auto_iopadmap_cc_368_execute_22625_130_), .Y(_abc_15497_new_n2103_));
INVX1 INVX1_254 ( .A(a_reg_1_), .Y(_abc_15497_new_n2104_));
INVX1 INVX1_255 ( .A(_abc_15497_new_n2108_), .Y(_abc_15497_new_n2109_));
INVX1 INVX1_256 ( .A(a_reg_2_), .Y(_abc_15497_new_n2113_));
INVX1 INVX1_257 ( .A(a_reg_3_), .Y(_abc_15497_new_n2115_));
INVX1 INVX1_258 ( .A(_abc_15497_new_n2117_), .Y(_abc_15497_new_n2118_));
INVX1 INVX1_259 ( .A(_auto_iopadmap_cc_368_execute_22625_132_), .Y(_abc_15497_new_n2122_));
INVX1 INVX1_26 ( .A(_abc_15497_new_n788_), .Y(_abc_15497_new_n789_));
INVX1 INVX1_260 ( .A(a_reg_4_), .Y(_abc_15497_new_n2130_));
INVX1 INVX1_261 ( .A(a_reg_5_), .Y(_abc_15497_new_n2134_));
INVX1 INVX1_262 ( .A(a_reg_6_), .Y(_abc_15497_new_n2144_));
INVX1 INVX1_263 ( .A(_auto_iopadmap_cc_368_execute_22625_135_), .Y(_abc_15497_new_n2151_));
INVX1 INVX1_264 ( .A(_abc_15497_new_n2152_), .Y(_abc_15497_new_n2153_));
INVX1 INVX1_265 ( .A(a_reg_7_), .Y(_abc_15497_new_n2159_));
INVX1 INVX1_266 ( .A(_abc_15497_new_n2162_), .Y(_abc_15497_new_n2163_));
INVX1 INVX1_267 ( .A(_auto_iopadmap_cc_368_execute_22625_136_), .Y(_abc_15497_new_n2165_));
INVX1 INVX1_268 ( .A(a_reg_8_), .Y(_abc_15497_new_n2166_));
INVX1 INVX1_269 ( .A(_abc_15497_new_n2168_), .Y(_abc_15497_new_n2170_));
INVX1 INVX1_27 ( .A(_abc_15497_new_n794_), .Y(_abc_15497_new_n795_));
INVX1 INVX1_270 ( .A(_abc_15497_new_n2167_), .Y(_abc_15497_new_n2174_));
INVX1 INVX1_271 ( .A(_auto_iopadmap_cc_368_execute_22625_138_), .Y(_abc_15497_new_n2180_));
INVX1 INVX1_272 ( .A(a_reg_10_), .Y(_abc_15497_new_n2182_));
INVX1 INVX1_273 ( .A(_abc_15497_new_n2184_), .Y(_abc_15497_new_n2185_));
INVX1 INVX1_274 ( .A(_auto_iopadmap_cc_368_execute_22625_137_), .Y(_abc_15497_new_n2186_));
INVX1 INVX1_275 ( .A(a_reg_9_), .Y(_abc_15497_new_n2187_));
INVX1 INVX1_276 ( .A(_abc_15497_new_n2189_), .Y(_abc_15497_new_n2190_));
INVX1 INVX1_277 ( .A(_abc_15497_new_n2191_), .Y(_abc_15497_new_n2192_));
INVX1 INVX1_278 ( .A(_auto_iopadmap_cc_368_execute_22625_139_), .Y(_abc_15497_new_n2197_));
INVX1 INVX1_279 ( .A(_abc_15497_new_n2183_), .Y(_abc_15497_new_n2198_));
INVX1 INVX1_28 ( .A(_abc_15497_new_n796_), .Y(_abc_15497_new_n797_));
INVX1 INVX1_280 ( .A(_abc_15497_new_n2205_), .Y(_abc_15497_new_n2206_));
INVX1 INVX1_281 ( .A(a_reg_11_), .Y(_abc_15497_new_n2207_));
INVX1 INVX1_282 ( .A(_abc_15497_new_n2210_), .Y(_abc_15497_new_n2211_));
INVX1 INVX1_283 ( .A(_auto_iopadmap_cc_368_execute_22625_143_), .Y(_abc_15497_new_n2241_));
INVX1 INVX1_284 ( .A(a_reg_15_), .Y(_abc_15497_new_n2244_));
INVX1 INVX1_285 ( .A(_auto_iopadmap_cc_368_execute_22625_144_), .Y(_abc_15497_new_n2257_));
INVX1 INVX1_286 ( .A(_abc_15497_new_n2255_), .Y(_abc_15497_new_n2262_));
INVX1 INVX1_287 ( .A(_abc_15497_new_n2260_), .Y(_abc_15497_new_n2263_));
INVX1 INVX1_288 ( .A(_auto_iopadmap_cc_368_execute_22625_145_), .Y(_abc_15497_new_n2267_));
INVX1 INVX1_289 ( .A(a_reg_17_), .Y(_abc_15497_new_n2270_));
INVX1 INVX1_29 ( .A(c_reg_22_), .Y(_abc_15497_new_n798_));
INVX1 INVX1_290 ( .A(_abc_15497_new_n2272_), .Y(_abc_15497_new_n2273_));
INVX1 INVX1_291 ( .A(_abc_15497_new_n2278_), .Y(_abc_15497_new_n2279_));
INVX1 INVX1_292 ( .A(_auto_iopadmap_cc_368_execute_22625_146_), .Y(_abc_15497_new_n2283_));
INVX1 INVX1_293 ( .A(a_reg_18_), .Y(_abc_15497_new_n2284_));
INVX1 INVX1_294 ( .A(_abc_15497_new_n2290_), .Y(_abc_15497_new_n2291_));
INVX1 INVX1_295 ( .A(_auto_iopadmap_cc_368_execute_22625_147_), .Y(_abc_15497_new_n2293_));
INVX1 INVX1_296 ( .A(a_reg_19_), .Y(_abc_15497_new_n2296_));
INVX1 INVX1_297 ( .A(_abc_15497_new_n2298_), .Y(_abc_15497_new_n2299_));
INVX1 INVX1_298 ( .A(_auto_iopadmap_cc_368_execute_22625_148_), .Y(_abc_15497_new_n2303_));
INVX1 INVX1_299 ( .A(a_reg_20_), .Y(_abc_15497_new_n2310_));
INVX1 INVX1_3 ( .A(_auto_iopadmap_cc_368_execute_22625_77_), .Y(_abc_15497_new_n709_));
INVX1 INVX1_30 ( .A(_auto_iopadmap_cc_368_execute_22625_86_), .Y(_abc_15497_new_n799_));
INVX1 INVX1_300 ( .A(_abc_15497_new_n2312_), .Y(_abc_15497_new_n2313_));
INVX1 INVX1_301 ( .A(_auto_iopadmap_cc_368_execute_22625_149_), .Y(_abc_15497_new_n2317_));
INVX1 INVX1_302 ( .A(_abc_15497_new_n2311_), .Y(_abc_15497_new_n2319_));
INVX1 INVX1_303 ( .A(a_reg_21_), .Y(_abc_15497_new_n2321_));
INVX1 INVX1_304 ( .A(_abc_15497_new_n2322_), .Y(_abc_15497_new_n2328_));
INVX1 INVX1_305 ( .A(_auto_iopadmap_cc_368_execute_22625_150_), .Y(_abc_15497_new_n2331_));
INVX1 INVX1_306 ( .A(a_reg_22_), .Y(_abc_15497_new_n2332_));
INVX1 INVX1_307 ( .A(_auto_iopadmap_cc_368_execute_22625_151_), .Y(_abc_15497_new_n2341_));
INVX1 INVX1_308 ( .A(_abc_15497_new_n2307_), .Y(_abc_15497_new_n2345_));
INVX1 INVX1_309 ( .A(_abc_15497_new_n2334_), .Y(_abc_15497_new_n2347_));
INVX1 INVX1_31 ( .A(_abc_15497_new_n802_), .Y(_abc_15497_new_n803_));
INVX1 INVX1_310 ( .A(a_reg_23_), .Y(_abc_15497_new_n2349_));
INVX1 INVX1_311 ( .A(_abc_15497_new_n2305_), .Y(_abc_15497_new_n2355_));
INVX1 INVX1_312 ( .A(_auto_iopadmap_cc_368_execute_22625_152_), .Y(_abc_15497_new_n2359_));
INVX1 INVX1_313 ( .A(_abc_15497_new_n2362_), .Y(_abc_15497_new_n2363_));
INVX1 INVX1_314 ( .A(_abc_15497_new_n2361_), .Y(_abc_15497_new_n2368_));
INVX1 INVX1_315 ( .A(_auto_iopadmap_cc_368_execute_22625_153_), .Y(_abc_15497_new_n2371_));
INVX1 INVX1_316 ( .A(a_reg_25_), .Y(_abc_15497_new_n2372_));
INVX1 INVX1_317 ( .A(_abc_15497_new_n2374_), .Y(_abc_15497_new_n2378_));
INVX1 INVX1_318 ( .A(_abc_15497_new_n2379_), .Y(_abc_15497_new_n2380_));
INVX1 INVX1_319 ( .A(_auto_iopadmap_cc_368_execute_22625_154_), .Y(_abc_15497_new_n2384_));
INVX1 INVX1_32 ( .A(_abc_15497_new_n804_), .Y(_abc_15497_new_n805_));
INVX1 INVX1_320 ( .A(a_reg_26_), .Y(_abc_15497_new_n2385_));
INVX1 INVX1_321 ( .A(_auto_iopadmap_cc_368_execute_22625_155_), .Y(_abc_15497_new_n2393_));
INVX1 INVX1_322 ( .A(a_reg_27_), .Y(_abc_15497_new_n2395_));
INVX1 INVX1_323 ( .A(_auto_iopadmap_cc_368_execute_22625_156_), .Y(_abc_15497_new_n2401_));
INVX1 INVX1_324 ( .A(_abc_15497_new_n2381_), .Y(_abc_15497_new_n2404_));
INVX1 INVX1_325 ( .A(_abc_15497_new_n2405_), .Y(_abc_15497_new_n2406_));
INVX1 INVX1_326 ( .A(a_reg_28_), .Y(_abc_15497_new_n2414_));
INVX1 INVX1_327 ( .A(_auto_iopadmap_cc_368_execute_22625_157_), .Y(_abc_15497_new_n2417_));
INVX1 INVX1_328 ( .A(a_reg_29_), .Y(_abc_15497_new_n2418_));
INVX1 INVX1_329 ( .A(_auto_iopadmap_cc_368_execute_22625_158_), .Y(_abc_15497_new_n2425_));
INVX1 INVX1_33 ( .A(_abc_15497_new_n809_), .Y(_abc_15497_new_n813_));
INVX1 INVX1_330 ( .A(a_reg_30_), .Y(_abc_15497_new_n2426_));
INVX1 INVX1_331 ( .A(_auto_iopadmap_cc_368_execute_22625_159_), .Y(_abc_15497_new_n2438_));
INVX1 INVX1_332 ( .A(d_reg_30_), .Y(_abc_15497_new_n2630_));
INVX1 INVX1_333 ( .A(_abc_15497_new_n883__bF_buf13), .Y(_abc_15497_new_n2634_));
INVX1 INVX1_334 ( .A(w_0_), .Y(_abc_15497_new_n2762_));
INVX1 INVX1_335 ( .A(_abc_15497_new_n2764_), .Y(_abc_15497_new_n2765_));
INVX1 INVX1_336 ( .A(_abc_15497_new_n2771_), .Y(_abc_15497_new_n2772_));
INVX1 INVX1_337 ( .A(w_1_), .Y(_abc_15497_new_n2792_));
INVX1 INVX1_338 ( .A(_abc_15497_new_n2794_), .Y(_abc_15497_new_n2795_));
INVX1 INVX1_339 ( .A(_abc_15497_new_n2793_), .Y(_abc_15497_new_n2797_));
INVX1 INVX1_34 ( .A(_abc_15497_new_n815_), .Y(_abc_15497_new_n816_));
INVX1 INVX1_340 ( .A(_abc_15497_new_n2791_), .Y(_abc_15497_new_n2800_));
INVX1 INVX1_341 ( .A(w_2_), .Y(_abc_15497_new_n2840_));
INVX1 INVX1_342 ( .A(_abc_15497_new_n2842_), .Y(_abc_15497_new_n2843_));
INVX1 INVX1_343 ( .A(_abc_15497_new_n2841_), .Y(_abc_15497_new_n2845_));
INVX1 INVX1_344 ( .A(_abc_15497_new_n2839_), .Y(_abc_15497_new_n2848_));
INVX1 INVX1_345 ( .A(_abc_15497_new_n2799_), .Y(_abc_15497_new_n2857_));
INVX1 INVX1_346 ( .A(_abc_15497_new_n2885_), .Y(_abc_15497_new_n2886_));
INVX1 INVX1_347 ( .A(_abc_15497_new_n2847_), .Y(_abc_15497_new_n2887_));
INVX1 INVX1_348 ( .A(_abc_15497_new_n2901_), .Y(_abc_15497_new_n2902_));
INVX1 INVX1_349 ( .A(w_3_), .Y(_abc_15497_new_n2903_));
INVX1 INVX1_35 ( .A(_abc_15497_new_n817_), .Y(_abc_15497_new_n818_));
INVX1 INVX1_350 ( .A(_abc_15497_new_n2898_), .Y(_abc_15497_new_n2907_));
INVX1 INVX1_351 ( .A(_abc_15497_new_n2899_), .Y(_abc_15497_new_n2955_));
INVX1 INVX1_352 ( .A(w_4_), .Y(_abc_15497_new_n2957_));
INVX1 INVX1_353 ( .A(_abc_15497_new_n2959_), .Y(_abc_15497_new_n2960_));
INVX1 INVX1_354 ( .A(_abc_15497_new_n2958_), .Y(_abc_15497_new_n2962_));
INVX1 INVX1_355 ( .A(_abc_15497_new_n2900_), .Y(_abc_15497_new_n2965_));
INVX1 INVX1_356 ( .A(_abc_15497_new_n2969_), .Y(_abc_15497_new_n2970_));
INVX1 INVX1_357 ( .A(_abc_15497_new_n2906_), .Y(_abc_15497_new_n2974_));
INVX1 INVX1_358 ( .A(_abc_15497_new_n2949_), .Y(_abc_15497_new_n2977_));
INVX1 INVX1_359 ( .A(_abc_15497_new_n2952_), .Y(_abc_15497_new_n2978_));
INVX1 INVX1_36 ( .A(c_reg_18_), .Y(_abc_15497_new_n823_));
INVX1 INVX1_360 ( .A(w_5_), .Y(_abc_15497_new_n3018_));
INVX1 INVX1_361 ( .A(_abc_15497_new_n3020_), .Y(_abc_15497_new_n3021_));
INVX1 INVX1_362 ( .A(_abc_15497_new_n3019_), .Y(_abc_15497_new_n3023_));
INVX1 INVX1_363 ( .A(_abc_15497_new_n3017_), .Y(_abc_15497_new_n3026_));
INVX1 INVX1_364 ( .A(_abc_15497_new_n2964_), .Y(_abc_15497_new_n3036_));
INVX1 INVX1_365 ( .A(_abc_15497_new_n3061_), .Y(_abc_15497_new_n3062_));
INVX1 INVX1_366 ( .A(w_6_), .Y(_abc_15497_new_n3076_));
INVX1 INVX1_367 ( .A(_abc_15497_new_n3078_), .Y(_abc_15497_new_n3079_));
INVX1 INVX1_368 ( .A(_abc_15497_new_n3077_), .Y(_abc_15497_new_n3081_));
INVX1 INVX1_369 ( .A(_abc_15497_new_n3075_), .Y(_abc_15497_new_n3084_));
INVX1 INVX1_37 ( .A(_auto_iopadmap_cc_368_execute_22625_82_), .Y(_abc_15497_new_n824_));
INVX1 INVX1_370 ( .A(_abc_15497_new_n3025_), .Y(_abc_15497_new_n3094_));
INVX1 INVX1_371 ( .A(_abc_15497_new_n3064_), .Y(_abc_15497_new_n3104_));
INVX1 INVX1_372 ( .A(_abc_15497_new_n3063_), .Y(_abc_15497_new_n3110_));
INVX1 INVX1_373 ( .A(_abc_15497_new_n3108_), .Y(_abc_15497_new_n3111_));
INVX1 INVX1_374 ( .A(_abc_15497_new_n3122_), .Y(_abc_15497_new_n3125_));
INVX1 INVX1_375 ( .A(_abc_15497_new_n3126_), .Y(_abc_15497_new_n3127_));
INVX1 INVX1_376 ( .A(w_7_), .Y(_abc_15497_new_n3131_));
INVX1 INVX1_377 ( .A(_abc_15497_new_n3133_), .Y(_abc_15497_new_n3134_));
INVX1 INVX1_378 ( .A(_abc_15497_new_n3132_), .Y(_abc_15497_new_n3136_));
INVX1 INVX1_379 ( .A(_abc_15497_new_n3130_), .Y(_abc_15497_new_n3139_));
INVX1 INVX1_38 ( .A(c_reg_16_), .Y(_abc_15497_new_n832_));
INVX1 INVX1_380 ( .A(_abc_15497_new_n3083_), .Y(_abc_15497_new_n3153_));
INVX1 INVX1_381 ( .A(_abc_15497_new_n3167_), .Y(_abc_15497_new_n3168_));
INVX1 INVX1_382 ( .A(w_8_), .Y(_abc_15497_new_n3179_));
INVX1 INVX1_383 ( .A(_abc_15497_new_n3181_), .Y(_abc_15497_new_n3182_));
INVX1 INVX1_384 ( .A(_abc_15497_new_n3180_), .Y(_abc_15497_new_n3184_));
INVX1 INVX1_385 ( .A(_abc_15497_new_n3178_), .Y(_abc_15497_new_n3192_));
INVX1 INVX1_386 ( .A(_abc_15497_new_n3138_), .Y(_abc_15497_new_n3196_));
INVX1 INVX1_387 ( .A(_abc_15497_new_n3225_), .Y(_abc_15497_new_n3226_));
INVX1 INVX1_388 ( .A(b_reg_9_), .Y(_abc_15497_new_n3232_));
INVX1 INVX1_389 ( .A(w_9_), .Y(_abc_15497_new_n3242_));
INVX1 INVX1_39 ( .A(_auto_iopadmap_cc_368_execute_22625_80_), .Y(_abc_15497_new_n833_));
INVX1 INVX1_390 ( .A(_abc_15497_new_n3244_), .Y(_abc_15497_new_n3245_));
INVX1 INVX1_391 ( .A(_abc_15497_new_n3241_), .Y(_abc_15497_new_n3251_));
INVX1 INVX1_392 ( .A(_abc_15497_new_n3229_), .Y(_abc_15497_new_n3275_));
INVX1 INVX1_393 ( .A(_abc_15497_new_n3285_), .Y(_abc_15497_new_n3286_));
INVX1 INVX1_394 ( .A(_abc_15497_new_n3300_), .Y(_abc_15497_new_n3301_));
INVX1 INVX1_395 ( .A(w_10_), .Y(_abc_15497_new_n3302_));
INVX1 INVX1_396 ( .A(_abc_15497_new_n3304_), .Y(_abc_15497_new_n3305_));
INVX1 INVX1_397 ( .A(_abc_15497_new_n3303_), .Y(_abc_15497_new_n3307_));
INVX1 INVX1_398 ( .A(_abc_15497_new_n3293_), .Y(_abc_15497_new_n3315_));
INVX1 INVX1_399 ( .A(_abc_15497_new_n3297_), .Y(_abc_15497_new_n3316_));
INVX1 INVX1_4 ( .A(_abc_15497_new_n716_), .Y(_abc_15497_new_n717_));
INVX1 INVX1_40 ( .A(_abc_15497_new_n838_), .Y(_abc_15497_new_n839_));
INVX1 INVX1_400 ( .A(_abc_15497_new_n3259_), .Y(_abc_15497_new_n3331_));
INVX1 INVX1_401 ( .A(_abc_15497_new_n3341_), .Y(_abc_15497_new_n3342_));
INVX1 INVX1_402 ( .A(w_11_), .Y(_abc_15497_new_n3361_));
INVX1 INVX1_403 ( .A(_abc_15497_new_n3360_), .Y(_abc_15497_new_n3369_));
INVX1 INVX1_404 ( .A(_abc_15497_new_n3319_), .Y(_abc_15497_new_n3381_));
INVX1 INVX1_405 ( .A(_abc_15497_new_n3217_), .Y(_abc_15497_new_n3403_));
INVX1 INVX1_406 ( .A(_abc_15497_new_n3354_), .Y(_abc_15497_new_n3411_));
INVX1 INVX1_407 ( .A(_abc_15497_new_n3358_), .Y(_abc_15497_new_n3412_));
INVX1 INVX1_408 ( .A(_abc_15497_new_n3429_), .Y(_abc_15497_new_n3430_));
INVX1 INVX1_409 ( .A(w_12_), .Y(_abc_15497_new_n3431_));
INVX1 INVX1_41 ( .A(_abc_15497_new_n831_), .Y(_abc_15497_new_n840_));
INVX1 INVX1_410 ( .A(_abc_15497_new_n3433_), .Y(_abc_15497_new_n3434_));
INVX1 INVX1_411 ( .A(_abc_15497_new_n3426_), .Y(_abc_15497_new_n3446_));
INVX1 INVX1_412 ( .A(_abc_15497_new_n3368_), .Y(_abc_15497_new_n3454_));
INVX1 INVX1_413 ( .A(_abc_15497_new_n3490_), .Y(_abc_15497_new_n3491_));
INVX1 INVX1_414 ( .A(w_13_), .Y(_abc_15497_new_n3494_));
INVX1 INVX1_415 ( .A(_abc_15497_new_n3493_), .Y(_abc_15497_new_n3503_));
INVX1 INVX1_416 ( .A(_abc_15497_new_n3449_), .Y(_abc_15497_new_n3517_));
INVX1 INVX1_417 ( .A(_abc_15497_new_n3527_), .Y(_abc_15497_new_n3528_));
INVX1 INVX1_418 ( .A(a_reg_13_), .Y(_abc_15497_new_n3531_));
INVX1 INVX1_419 ( .A(d_reg_14_), .Y(_abc_15497_new_n3543_));
INVX1 INVX1_42 ( .A(_abc_15497_new_n842_), .Y(_abc_15497_new_n843_));
INVX1 INVX1_420 ( .A(_abc_15497_new_n3552_), .Y(_abc_15497_new_n3553_));
INVX1 INVX1_421 ( .A(_abc_15497_new_n3554_), .Y(_abc_15497_new_n3555_));
INVX1 INVX1_422 ( .A(_abc_15497_new_n3557_), .Y(_abc_15497_new_n3558_));
INVX1 INVX1_423 ( .A(w_14_), .Y(_abc_15497_new_n3559_));
INVX1 INVX1_424 ( .A(_abc_15497_new_n3508_), .Y(_abc_15497_new_n3586_));
INVX1 INVX1_425 ( .A(b_reg_15_), .Y(_abc_15497_new_n3608_));
INVX1 INVX1_426 ( .A(c_reg_15_), .Y(_abc_15497_new_n3609_));
INVX1 INVX1_427 ( .A(_abc_15497_new_n3620_), .Y(_abc_15497_new_n3621_));
INVX1 INVX1_428 ( .A(w_15_), .Y(_abc_15497_new_n3622_));
INVX1 INVX1_429 ( .A(_abc_15497_new_n3624_), .Y(_abc_15497_new_n3625_));
INVX1 INVX1_43 ( .A(_abc_15497_new_n844_), .Y(_abc_15497_new_n845_));
INVX1 INVX1_430 ( .A(_abc_15497_new_n3574_), .Y(_abc_15497_new_n3650_));
INVX1 INVX1_431 ( .A(_abc_15497_new_n3660_), .Y(_abc_15497_new_n3663_));
INVX1 INVX1_432 ( .A(_abc_15497_new_n3675_), .Y(_abc_15497_new_n3676_));
INVX1 INVX1_433 ( .A(_abc_15497_new_n3680_), .Y(_abc_15497_new_n3681_));
INVX1 INVX1_434 ( .A(w_16_), .Y(_abc_15497_new_n3692_));
INVX1 INVX1_435 ( .A(_abc_15497_new_n3690_), .Y(_abc_15497_new_n3699_));
INVX1 INVX1_436 ( .A(_abc_15497_new_n3711_), .Y(_abc_15497_new_n3712_));
INVX1 INVX1_437 ( .A(w_17_), .Y(_abc_15497_new_n3738_));
INVX1 INVX1_438 ( .A(_abc_15497_new_n3735_), .Y(_abc_15497_new_n3751_));
INVX1 INVX1_439 ( .A(_abc_15497_new_n3724_), .Y(_abc_15497_new_n3755_));
INVX1 INVX1_44 ( .A(c_reg_25_), .Y(_abc_15497_new_n849_));
INVX1 INVX1_440 ( .A(_abc_15497_new_n3722_), .Y(_abc_15497_new_n3765_));
INVX1 INVX1_441 ( .A(_abc_15497_new_n3769_), .Y(_abc_15497_new_n3770_));
INVX1 INVX1_442 ( .A(_abc_15497_new_n3779_), .Y(_abc_15497_new_n3780_));
INVX1 INVX1_443 ( .A(b_reg_18_), .Y(_abc_15497_new_n3785_));
INVX1 INVX1_444 ( .A(w_18_), .Y(_abc_15497_new_n3797_));
INVX1 INVX1_445 ( .A(_abc_15497_new_n3801_), .Y(_abc_15497_new_n3805_));
INVX1 INVX1_446 ( .A(_abc_15497_new_n3783_), .Y(_abc_15497_new_n3811_));
INVX1 INVX1_447 ( .A(_abc_15497_new_n3818_), .Y(_abc_15497_new_n3819_));
INVX1 INVX1_448 ( .A(_abc_15497_new_n3824_), .Y(_abc_15497_new_n3825_));
INVX1 INVX1_449 ( .A(_abc_15497_new_n3810_), .Y(_abc_15497_new_n3827_));
INVX1 INVX1_45 ( .A(_auto_iopadmap_cc_368_execute_22625_89_), .Y(_abc_15497_new_n850_));
INVX1 INVX1_450 ( .A(_abc_15497_new_n3806_), .Y(_abc_15497_new_n3828_));
INVX1 INVX1_451 ( .A(b_reg_19_), .Y(_abc_15497_new_n3833_));
INVX1 INVX1_452 ( .A(w_19_), .Y(_abc_15497_new_n3841_));
INVX1 INVX1_453 ( .A(_abc_15497_new_n3881_), .Y(_abc_15497_new_n3882_));
INVX1 INVX1_454 ( .A(_abc_15497_new_n3800_), .Y(_abc_15497_new_n3889_));
INVX1 INVX1_455 ( .A(_abc_15497_new_n3845_), .Y(_abc_15497_new_n3890_));
INVX1 INVX1_456 ( .A(_abc_15497_new_n3891_), .Y(_abc_15497_new_n3892_));
INVX1 INVX1_457 ( .A(w_20_), .Y(_abc_15497_new_n3904_));
INVX1 INVX1_458 ( .A(_abc_15497_new_n3902_), .Y(_abc_15497_new_n3911_));
INVX1 INVX1_459 ( .A(_abc_15497_new_n3844_), .Y(_abc_15497_new_n3939_));
INVX1 INVX1_46 ( .A(_abc_15497_new_n853_), .Y(_abc_15497_new_n854_));
INVX1 INVX1_460 ( .A(_abc_15497_new_n3908_), .Y(_abc_15497_new_n3940_));
INVX1 INVX1_461 ( .A(_abc_15497_new_n3941_), .Y(_abc_15497_new_n3942_));
INVX1 INVX1_462 ( .A(d_reg_21_), .Y(_abc_15497_new_n3948_));
INVX1 INVX1_463 ( .A(w_21_), .Y(_abc_15497_new_n3955_));
INVX1 INVX1_464 ( .A(_abc_15497_new_n3953_), .Y(_abc_15497_new_n3962_));
INVX1 INVX1_465 ( .A(_abc_15497_new_n3979_), .Y(_abc_15497_new_n3980_));
INVX1 INVX1_466 ( .A(_abc_15497_new_n3907_), .Y(_abc_15497_new_n3994_));
INVX1 INVX1_467 ( .A(_abc_15497_new_n3959_), .Y(_abc_15497_new_n3995_));
INVX1 INVX1_468 ( .A(_abc_15497_new_n3996_), .Y(_abc_15497_new_n3997_));
INVX1 INVX1_469 ( .A(b_reg_22_), .Y(_abc_15497_new_n4005_));
INVX1 INVX1_47 ( .A(c_reg_24_), .Y(_abc_15497_new_n855_));
INVX1 INVX1_470 ( .A(w_22_), .Y(_abc_15497_new_n4010_));
INVX1 INVX1_471 ( .A(_abc_15497_new_n4008_), .Y(_abc_15497_new_n4017_));
INVX1 INVX1_472 ( .A(_abc_15497_new_n4034_), .Y(_abc_15497_new_n4035_));
INVX1 INVX1_473 ( .A(_abc_15497_new_n3958_), .Y(_abc_15497_new_n4046_));
INVX1 INVX1_474 ( .A(_abc_15497_new_n4014_), .Y(_abc_15497_new_n4047_));
INVX1 INVX1_475 ( .A(_abc_15497_new_n4058_), .Y(_abc_15497_new_n4059_));
INVX1 INVX1_476 ( .A(e_reg_22_), .Y(_abc_15497_new_n4060_));
INVX1 INVX1_477 ( .A(_abc_15497_new_n4061_), .Y(_abc_15497_new_n4062_));
INVX1 INVX1_478 ( .A(w_23_), .Y(_abc_15497_new_n4064_));
INVX1 INVX1_479 ( .A(_abc_15497_new_n4048_), .Y(_abc_15497_new_n4075_));
INVX1 INVX1_48 ( .A(_auto_iopadmap_cc_368_execute_22625_88_), .Y(_abc_15497_new_n856_));
INVX1 INVX1_480 ( .A(_abc_15497_new_n4089_), .Y(_abc_15497_new_n4090_));
INVX1 INVX1_481 ( .A(e_reg_23_), .Y(_abc_15497_new_n4118_));
INVX1 INVX1_482 ( .A(_abc_15497_new_n4119_), .Y(_abc_15497_new_n4120_));
INVX1 INVX1_483 ( .A(w_24_), .Y(_abc_15497_new_n4122_));
INVX1 INVX1_484 ( .A(_abc_15497_new_n4134_), .Y(_abc_15497_new_n4135_));
INVX1 INVX1_485 ( .A(_abc_15497_new_n4107_), .Y(_abc_15497_new_n4141_));
INVX1 INVX1_486 ( .A(_abc_15497_new_n4117_), .Y(_abc_15497_new_n4152_));
INVX1 INVX1_487 ( .A(_abc_15497_new_n4154_), .Y(_abc_15497_new_n4155_));
INVX1 INVX1_488 ( .A(e_reg_25_), .Y(_abc_15497_new_n4165_));
INVX1 INVX1_489 ( .A(_abc_15497_new_n4173_), .Y(_abc_15497_new_n4174_));
INVX1 INVX1_49 ( .A(_abc_15497_new_n861_), .Y(_abc_15497_new_n862_));
INVX1 INVX1_490 ( .A(w_26_), .Y(_abc_15497_new_n4207_));
INVX1 INVX1_491 ( .A(_abc_15497_new_n4220_), .Y(_abc_15497_new_n4221_));
INVX1 INVX1_492 ( .A(_abc_15497_new_n4217_), .Y(_abc_15497_new_n4234_));
INVX1 INVX1_493 ( .A(_abc_15497_new_n4204_), .Y(_abc_15497_new_n4236_));
INVX1 INVX1_494 ( .A(c_reg_27_), .Y(_abc_15497_new_n4239_));
INVX1 INVX1_495 ( .A(b_reg_27_), .Y(_abc_15497_new_n4240_));
INVX1 INVX1_496 ( .A(w_27_), .Y(_abc_15497_new_n4251_));
INVX1 INVX1_497 ( .A(_abc_15497_new_n4238_), .Y(_abc_15497_new_n4276_));
INVX1 INVX1_498 ( .A(_abc_15497_new_n4280_), .Y(_abc_15497_new_n4281_));
INVX1 INVX1_499 ( .A(_abc_15497_new_n4303_), .Y(_abc_15497_new_n4324_));
INVX1 INVX1_5 ( .A(_abc_15497_new_n713_), .Y(_abc_15497_new_n718_));
INVX1 INVX1_50 ( .A(_abc_15497_new_n879_), .Y(_abc_15497_new_n880_));
INVX1 INVX1_500 ( .A(b_reg_29_), .Y(_abc_15497_new_n4330_));
INVX1 INVX1_501 ( .A(_abc_15497_new_n4334_), .Y(_abc_15497_new_n4339_));
INVX1 INVX1_502 ( .A(_abc_15497_new_n4348_), .Y(_abc_15497_new_n4349_));
INVX1 INVX1_503 ( .A(_abc_15497_new_n4358_), .Y(_abc_15497_new_n4366_));
INVX1 INVX1_504 ( .A(b_reg_30_), .Y(_abc_15497_new_n4372_));
INVX1 INVX1_505 ( .A(_abc_15497_new_n4376_), .Y(_abc_15497_new_n4381_));
INVX1 INVX1_506 ( .A(e_reg_30_), .Y(_abc_15497_new_n4388_));
INVX1 INVX1_507 ( .A(_abc_15497_new_n4394_), .Y(_abc_15497_new_n4395_));
INVX1 INVX1_508 ( .A(_abc_15497_new_n4401_), .Y(_abc_15497_new_n4409_));
INVX1 INVX1_509 ( .A(_abc_15497_new_n4399_), .Y(_abc_15497_new_n4412_));
INVX1 INVX1_51 ( .A(_abc_15497_new_n863_), .Y(_abc_15497_new_n888_));
INVX1 INVX1_510 ( .A(_abc_15497_new_n4419_), .Y(_abc_15497_new_n4422_));
INVX1 INVX1_511 ( .A(_abc_15497_new_n4433_), .Y(_abc_15497_new_n4436_));
INVX1 INVX1_512 ( .A(round_ctr_reg_1_), .Y(_abc_15497_new_n4442_));
INVX1 INVX1_513 ( .A(_abc_15497_new_n4445_), .Y(_abc_15497_new_n4446_));
INVX1 INVX1_514 ( .A(_auto_iopadmap_cc_368_execute_22786), .Y(_abc_15497_new_n4474_));
INVX1 INVX1_515 ( .A(_abc_15497_new_n765_), .Y(_abc_15497_new_n4485_));
INVX1 INVX1_516 ( .A(_abc_15497_new_n763_), .Y(_abc_15497_new_n4499_));
INVX1 INVX1_517 ( .A(_abc_15497_new_n746_), .Y(_abc_15497_new_n4519_));
INVX1 INVX1_518 ( .A(_abc_15497_new_n4577_), .Y(_abc_15497_new_n4579_));
INVX1 INVX1_519 ( .A(_abc_15497_new_n800_), .Y(_abc_15497_new_n4583_));
INVX1 INVX1_52 ( .A(_abc_15497_new_n867_), .Y(_abc_15497_new_n889_));
INVX1 INVX1_520 ( .A(w_mem_inst_w_mem_5__0_), .Y(w_mem_inst__abc_19396_new_n1591_));
INVX1 INVX1_521 ( .A(w_mem_inst_w_ctr_reg_1_), .Y(w_mem_inst__abc_19396_new_n1592_));
INVX1 INVX1_522 ( .A(w_mem_inst_w_ctr_reg_3_), .Y(w_mem_inst__abc_19396_new_n1595_));
INVX1 INVX1_523 ( .A(w_mem_inst__abc_19396_new_n1596_), .Y(w_mem_inst__abc_19396_new_n1597_));
INVX1 INVX1_524 ( .A(w_mem_inst_w_mem_8__0_), .Y(w_mem_inst__abc_19396_new_n1600_));
INVX1 INVX1_525 ( .A(w_mem_inst_w_ctr_reg_2_), .Y(w_mem_inst__abc_19396_new_n1602_));
INVX1 INVX1_526 ( .A(w_mem_inst_w_mem_7__0_), .Y(w_mem_inst__abc_19396_new_n1609_));
INVX1 INVX1_527 ( .A(w_mem_inst__abc_19396_new_n1605_), .Y(w_mem_inst__abc_19396_new_n1610_));
INVX1 INVX1_528 ( .A(w_mem_inst_w_ctr_reg_0_), .Y(w_mem_inst__abc_19396_new_n1626_));
INVX1 INVX1_529 ( .A(w_mem_inst_w_mem_5__1_), .Y(w_mem_inst__abc_19396_new_n1646_));
INVX1 INVX1_53 ( .A(_abc_15497_new_n894_), .Y(_abc_15497_new_n895_));
INVX1 INVX1_530 ( .A(w_mem_inst_w_mem_8__1_), .Y(w_mem_inst__abc_19396_new_n1648_));
INVX1 INVX1_531 ( .A(w_mem_inst_w_mem_7__1_), .Y(w_mem_inst__abc_19396_new_n1651_));
INVX1 INVX1_532 ( .A(w_mem_inst_w_mem_5__2_), .Y(w_mem_inst__abc_19396_new_n1671_));
INVX1 INVX1_533 ( .A(w_mem_inst_w_mem_8__2_), .Y(w_mem_inst__abc_19396_new_n1673_));
INVX1 INVX1_534 ( .A(w_mem_inst_w_mem_7__2_), .Y(w_mem_inst__abc_19396_new_n1676_));
INVX1 INVX1_535 ( .A(w_mem_inst_w_mem_5__3_), .Y(w_mem_inst__abc_19396_new_n1696_));
INVX1 INVX1_536 ( .A(w_mem_inst_w_mem_8__3_), .Y(w_mem_inst__abc_19396_new_n1698_));
INVX1 INVX1_537 ( .A(w_mem_inst_w_mem_7__3_), .Y(w_mem_inst__abc_19396_new_n1701_));
INVX1 INVX1_538 ( .A(w_mem_inst_w_mem_5__4_), .Y(w_mem_inst__abc_19396_new_n1721_));
INVX1 INVX1_539 ( .A(w_mem_inst_w_mem_8__4_), .Y(w_mem_inst__abc_19396_new_n1723_));
INVX1 INVX1_54 ( .A(_auto_iopadmap_cc_368_execute_22625_93_), .Y(_abc_15497_new_n901_));
INVX1 INVX1_540 ( .A(w_mem_inst_w_mem_7__4_), .Y(w_mem_inst__abc_19396_new_n1726_));
INVX1 INVX1_541 ( .A(w_mem_inst_w_mem_5__5_), .Y(w_mem_inst__abc_19396_new_n1746_));
INVX1 INVX1_542 ( .A(w_mem_inst_w_mem_8__5_), .Y(w_mem_inst__abc_19396_new_n1748_));
INVX1 INVX1_543 ( .A(w_mem_inst_w_mem_7__5_), .Y(w_mem_inst__abc_19396_new_n1751_));
INVX1 INVX1_544 ( .A(w_mem_inst_w_mem_5__6_), .Y(w_mem_inst__abc_19396_new_n1771_));
INVX1 INVX1_545 ( .A(w_mem_inst_w_mem_8__6_), .Y(w_mem_inst__abc_19396_new_n1773_));
INVX1 INVX1_546 ( .A(w_mem_inst_w_mem_7__6_), .Y(w_mem_inst__abc_19396_new_n1776_));
INVX1 INVX1_547 ( .A(w_mem_inst_w_mem_5__7_), .Y(w_mem_inst__abc_19396_new_n1796_));
INVX1 INVX1_548 ( .A(w_mem_inst_w_mem_8__7_), .Y(w_mem_inst__abc_19396_new_n1798_));
INVX1 INVX1_549 ( .A(w_mem_inst_w_mem_7__7_), .Y(w_mem_inst__abc_19396_new_n1801_));
INVX1 INVX1_55 ( .A(c_reg_29_), .Y(_abc_15497_new_n904_));
INVX1 INVX1_550 ( .A(w_mem_inst_w_mem_5__8_), .Y(w_mem_inst__abc_19396_new_n1821_));
INVX1 INVX1_551 ( .A(w_mem_inst_w_mem_8__8_), .Y(w_mem_inst__abc_19396_new_n1823_));
INVX1 INVX1_552 ( .A(w_mem_inst_w_mem_7__8_), .Y(w_mem_inst__abc_19396_new_n1826_));
INVX1 INVX1_553 ( .A(w_mem_inst_w_mem_5__9_), .Y(w_mem_inst__abc_19396_new_n1846_));
INVX1 INVX1_554 ( .A(w_mem_inst_w_mem_8__9_), .Y(w_mem_inst__abc_19396_new_n1848_));
INVX1 INVX1_555 ( .A(w_mem_inst_w_mem_7__9_), .Y(w_mem_inst__abc_19396_new_n1851_));
INVX1 INVX1_556 ( .A(w_mem_inst_w_mem_5__10_), .Y(w_mem_inst__abc_19396_new_n1871_));
INVX1 INVX1_557 ( .A(w_mem_inst_w_mem_8__10_), .Y(w_mem_inst__abc_19396_new_n1873_));
INVX1 INVX1_558 ( .A(w_mem_inst_w_mem_7__10_), .Y(w_mem_inst__abc_19396_new_n1876_));
INVX1 INVX1_559 ( .A(w_mem_inst_w_mem_5__11_), .Y(w_mem_inst__abc_19396_new_n1896_));
INVX1 INVX1_56 ( .A(_abc_15497_new_n906_), .Y(_abc_15497_new_n907_));
INVX1 INVX1_560 ( .A(w_mem_inst_w_mem_8__11_), .Y(w_mem_inst__abc_19396_new_n1898_));
INVX1 INVX1_561 ( .A(w_mem_inst_w_mem_7__11_), .Y(w_mem_inst__abc_19396_new_n1901_));
INVX1 INVX1_562 ( .A(w_mem_inst_w_mem_5__12_), .Y(w_mem_inst__abc_19396_new_n1921_));
INVX1 INVX1_563 ( .A(w_mem_inst_w_mem_8__12_), .Y(w_mem_inst__abc_19396_new_n1923_));
INVX1 INVX1_564 ( .A(w_mem_inst_w_mem_7__12_), .Y(w_mem_inst__abc_19396_new_n1926_));
INVX1 INVX1_565 ( .A(w_mem_inst_w_mem_5__13_), .Y(w_mem_inst__abc_19396_new_n1946_));
INVX1 INVX1_566 ( .A(w_mem_inst_w_mem_8__13_), .Y(w_mem_inst__abc_19396_new_n1948_));
INVX1 INVX1_567 ( .A(w_mem_inst_w_mem_7__13_), .Y(w_mem_inst__abc_19396_new_n1951_));
INVX1 INVX1_568 ( .A(w_mem_inst_w_mem_5__14_), .Y(w_mem_inst__abc_19396_new_n1971_));
INVX1 INVX1_569 ( .A(w_mem_inst_w_mem_8__14_), .Y(w_mem_inst__abc_19396_new_n1973_));
INVX1 INVX1_57 ( .A(_abc_15497_new_n905_), .Y(_abc_15497_new_n915_));
INVX1 INVX1_570 ( .A(w_mem_inst_w_mem_7__14_), .Y(w_mem_inst__abc_19396_new_n1976_));
INVX1 INVX1_571 ( .A(w_mem_inst_w_mem_5__15_), .Y(w_mem_inst__abc_19396_new_n1996_));
INVX1 INVX1_572 ( .A(w_mem_inst_w_mem_8__15_), .Y(w_mem_inst__abc_19396_new_n1998_));
INVX1 INVX1_573 ( .A(w_mem_inst_w_mem_7__15_), .Y(w_mem_inst__abc_19396_new_n2001_));
INVX1 INVX1_574 ( .A(w_mem_inst_w_mem_5__16_), .Y(w_mem_inst__abc_19396_new_n2021_));
INVX1 INVX1_575 ( .A(w_mem_inst_w_mem_8__16_), .Y(w_mem_inst__abc_19396_new_n2023_));
INVX1 INVX1_576 ( .A(w_mem_inst_w_mem_7__16_), .Y(w_mem_inst__abc_19396_new_n2026_));
INVX1 INVX1_577 ( .A(w_mem_inst_w_mem_5__17_), .Y(w_mem_inst__abc_19396_new_n2046_));
INVX1 INVX1_578 ( .A(w_mem_inst_w_mem_8__17_), .Y(w_mem_inst__abc_19396_new_n2048_));
INVX1 INVX1_579 ( .A(w_mem_inst_w_mem_7__17_), .Y(w_mem_inst__abc_19396_new_n2051_));
INVX1 INVX1_58 ( .A(_abc_15497_new_n916_), .Y(_abc_15497_new_n917_));
INVX1 INVX1_580 ( .A(w_mem_inst_w_mem_5__18_), .Y(w_mem_inst__abc_19396_new_n2071_));
INVX1 INVX1_581 ( .A(w_mem_inst_w_mem_8__18_), .Y(w_mem_inst__abc_19396_new_n2073_));
INVX1 INVX1_582 ( .A(w_mem_inst_w_mem_7__18_), .Y(w_mem_inst__abc_19396_new_n2076_));
INVX1 INVX1_583 ( .A(w_mem_inst_w_mem_5__19_), .Y(w_mem_inst__abc_19396_new_n2096_));
INVX1 INVX1_584 ( .A(w_mem_inst_w_mem_8__19_), .Y(w_mem_inst__abc_19396_new_n2098_));
INVX1 INVX1_585 ( .A(w_mem_inst_w_mem_7__19_), .Y(w_mem_inst__abc_19396_new_n2101_));
INVX1 INVX1_586 ( .A(w_mem_inst_w_mem_5__20_), .Y(w_mem_inst__abc_19396_new_n2121_));
INVX1 INVX1_587 ( .A(w_mem_inst_w_mem_8__20_), .Y(w_mem_inst__abc_19396_new_n2123_));
INVX1 INVX1_588 ( .A(w_mem_inst_w_mem_7__20_), .Y(w_mem_inst__abc_19396_new_n2126_));
INVX1 INVX1_589 ( .A(w_mem_inst_w_mem_5__21_), .Y(w_mem_inst__abc_19396_new_n2146_));
INVX1 INVX1_59 ( .A(_abc_15497_new_n925_), .Y(_abc_15497_new_n926_));
INVX1 INVX1_590 ( .A(w_mem_inst_w_mem_8__21_), .Y(w_mem_inst__abc_19396_new_n2148_));
INVX1 INVX1_591 ( .A(w_mem_inst_w_mem_7__21_), .Y(w_mem_inst__abc_19396_new_n2151_));
INVX1 INVX1_592 ( .A(w_mem_inst_w_mem_5__22_), .Y(w_mem_inst__abc_19396_new_n2171_));
INVX1 INVX1_593 ( .A(w_mem_inst_w_mem_8__22_), .Y(w_mem_inst__abc_19396_new_n2173_));
INVX1 INVX1_594 ( .A(w_mem_inst_w_mem_7__22_), .Y(w_mem_inst__abc_19396_new_n2176_));
INVX1 INVX1_595 ( .A(w_mem_inst_w_mem_5__23_), .Y(w_mem_inst__abc_19396_new_n2196_));
INVX1 INVX1_596 ( .A(w_mem_inst_w_mem_8__23_), .Y(w_mem_inst__abc_19396_new_n2198_));
INVX1 INVX1_597 ( .A(w_mem_inst_w_mem_7__23_), .Y(w_mem_inst__abc_19396_new_n2201_));
INVX1 INVX1_598 ( .A(w_mem_inst_w_mem_5__24_), .Y(w_mem_inst__abc_19396_new_n2221_));
INVX1 INVX1_599 ( .A(w_mem_inst_w_mem_8__24_), .Y(w_mem_inst__abc_19396_new_n2223_));
INVX1 INVX1_6 ( .A(_abc_15497_new_n720_), .Y(_abc_15497_new_n721_));
INVX1 INVX1_60 ( .A(_abc_15497_new_n929_), .Y(_abc_15497_new_n931_));
INVX1 INVX1_600 ( .A(w_mem_inst_w_mem_7__24_), .Y(w_mem_inst__abc_19396_new_n2226_));
INVX1 INVX1_601 ( .A(w_mem_inst_w_mem_5__25_), .Y(w_mem_inst__abc_19396_new_n2246_));
INVX1 INVX1_602 ( .A(w_mem_inst_w_mem_8__25_), .Y(w_mem_inst__abc_19396_new_n2248_));
INVX1 INVX1_603 ( .A(w_mem_inst_w_mem_7__25_), .Y(w_mem_inst__abc_19396_new_n2251_));
INVX1 INVX1_604 ( .A(w_mem_inst_w_mem_5__26_), .Y(w_mem_inst__abc_19396_new_n2271_));
INVX1 INVX1_605 ( .A(w_mem_inst_w_mem_8__26_), .Y(w_mem_inst__abc_19396_new_n2273_));
INVX1 INVX1_606 ( .A(w_mem_inst_w_mem_7__26_), .Y(w_mem_inst__abc_19396_new_n2276_));
INVX1 INVX1_607 ( .A(w_mem_inst_w_mem_5__27_), .Y(w_mem_inst__abc_19396_new_n2296_));
INVX1 INVX1_608 ( .A(w_mem_inst_w_mem_8__27_), .Y(w_mem_inst__abc_19396_new_n2298_));
INVX1 INVX1_609 ( .A(w_mem_inst_w_mem_7__27_), .Y(w_mem_inst__abc_19396_new_n2301_));
INVX1 INVX1_61 ( .A(_auto_iopadmap_cc_368_execute_22625_0_), .Y(_abc_15497_new_n936_));
INVX1 INVX1_610 ( .A(w_mem_inst_w_mem_5__28_), .Y(w_mem_inst__abc_19396_new_n2321_));
INVX1 INVX1_611 ( .A(w_mem_inst_w_mem_8__28_), .Y(w_mem_inst__abc_19396_new_n2323_));
INVX1 INVX1_612 ( .A(w_mem_inst_w_mem_7__28_), .Y(w_mem_inst__abc_19396_new_n2326_));
INVX1 INVX1_613 ( .A(w_mem_inst_w_mem_5__29_), .Y(w_mem_inst__abc_19396_new_n2346_));
INVX1 INVX1_614 ( .A(w_mem_inst_w_mem_8__29_), .Y(w_mem_inst__abc_19396_new_n2348_));
INVX1 INVX1_615 ( .A(w_mem_inst_w_mem_7__29_), .Y(w_mem_inst__abc_19396_new_n2351_));
INVX1 INVX1_616 ( .A(w_mem_inst_w_mem_5__30_), .Y(w_mem_inst__abc_19396_new_n2371_));
INVX1 INVX1_617 ( .A(w_mem_inst_w_mem_8__30_), .Y(w_mem_inst__abc_19396_new_n2373_));
INVX1 INVX1_618 ( .A(w_mem_inst_w_mem_7__30_), .Y(w_mem_inst__abc_19396_new_n2376_));
INVX1 INVX1_619 ( .A(w_mem_inst_w_mem_5__31_), .Y(w_mem_inst__abc_19396_new_n2396_));
INVX1 INVX1_62 ( .A(e_reg_0_), .Y(_abc_15497_new_n937_));
INVX1 INVX1_620 ( .A(w_mem_inst_w_mem_8__31_), .Y(w_mem_inst__abc_19396_new_n2398_));
INVX1 INVX1_621 ( .A(w_mem_inst_w_mem_7__31_), .Y(w_mem_inst__abc_19396_new_n2401_));
INVX1 INVX1_622 ( .A(w_mem_inst_w_mem_13__0_), .Y(w_mem_inst__abc_19396_new_n2418_));
INVX1 INVX1_623 ( .A(round_ctr_inc_bF_buf2), .Y(w_mem_inst__abc_19396_new_n2419_));
INVX1 INVX1_624 ( .A(\block[64] ), .Y(w_mem_inst__abc_19396_new_n2423_));
INVX1 INVX1_625 ( .A(w_mem_inst_w_mem_13__1_), .Y(w_mem_inst__abc_19396_new_n2427_));
INVX1 INVX1_626 ( .A(\block[65] ), .Y(w_mem_inst__abc_19396_new_n2428_));
INVX1 INVX1_627 ( .A(w_mem_inst_w_mem_13__2_), .Y(w_mem_inst__abc_19396_new_n2432_));
INVX1 INVX1_628 ( .A(\block[66] ), .Y(w_mem_inst__abc_19396_new_n2433_));
INVX1 INVX1_629 ( .A(w_mem_inst_w_mem_13__3_), .Y(w_mem_inst__abc_19396_new_n2437_));
INVX1 INVX1_63 ( .A(_auto_iopadmap_cc_368_execute_22625_1_), .Y(_abc_15497_new_n941_));
INVX1 INVX1_630 ( .A(\block[67] ), .Y(w_mem_inst__abc_19396_new_n2438_));
INVX1 INVX1_631 ( .A(w_mem_inst_w_mem_13__4_), .Y(w_mem_inst__abc_19396_new_n2442_));
INVX1 INVX1_632 ( .A(\block[68] ), .Y(w_mem_inst__abc_19396_new_n2443_));
INVX1 INVX1_633 ( .A(w_mem_inst_w_mem_13__5_), .Y(w_mem_inst__abc_19396_new_n2447_));
INVX1 INVX1_634 ( .A(\block[69] ), .Y(w_mem_inst__abc_19396_new_n2448_));
INVX1 INVX1_635 ( .A(w_mem_inst_w_mem_13__6_), .Y(w_mem_inst__abc_19396_new_n2452_));
INVX1 INVX1_636 ( .A(\block[70] ), .Y(w_mem_inst__abc_19396_new_n2453_));
INVX1 INVX1_637 ( .A(w_mem_inst_w_mem_13__7_), .Y(w_mem_inst__abc_19396_new_n2457_));
INVX1 INVX1_638 ( .A(\block[71] ), .Y(w_mem_inst__abc_19396_new_n2458_));
INVX1 INVX1_639 ( .A(w_mem_inst_w_mem_13__8_), .Y(w_mem_inst__abc_19396_new_n2462_));
INVX1 INVX1_64 ( .A(_auto_iopadmap_cc_368_execute_22625_2_), .Y(_abc_15497_new_n946_));
INVX1 INVX1_640 ( .A(\block[72] ), .Y(w_mem_inst__abc_19396_new_n2463_));
INVX1 INVX1_641 ( .A(w_mem_inst_w_mem_13__9_), .Y(w_mem_inst__abc_19396_new_n2467_));
INVX1 INVX1_642 ( .A(\block[73] ), .Y(w_mem_inst__abc_19396_new_n2468_));
INVX1 INVX1_643 ( .A(w_mem_inst_w_mem_13__10_), .Y(w_mem_inst__abc_19396_new_n2472_));
INVX1 INVX1_644 ( .A(\block[74] ), .Y(w_mem_inst__abc_19396_new_n2473_));
INVX1 INVX1_645 ( .A(w_mem_inst_w_mem_13__11_), .Y(w_mem_inst__abc_19396_new_n2477_));
INVX1 INVX1_646 ( .A(\block[75] ), .Y(w_mem_inst__abc_19396_new_n2478_));
INVX1 INVX1_647 ( .A(w_mem_inst_w_mem_13__12_), .Y(w_mem_inst__abc_19396_new_n2482_));
INVX1 INVX1_648 ( .A(\block[76] ), .Y(w_mem_inst__abc_19396_new_n2483_));
INVX1 INVX1_649 ( .A(w_mem_inst_w_mem_13__13_), .Y(w_mem_inst__abc_19396_new_n2487_));
INVX1 INVX1_65 ( .A(e_reg_1_), .Y(_abc_15497_new_n947_));
INVX1 INVX1_650 ( .A(\block[77] ), .Y(w_mem_inst__abc_19396_new_n2488_));
INVX1 INVX1_651 ( .A(w_mem_inst_w_mem_13__14_), .Y(w_mem_inst__abc_19396_new_n2492_));
INVX1 INVX1_652 ( .A(\block[78] ), .Y(w_mem_inst__abc_19396_new_n2493_));
INVX1 INVX1_653 ( .A(w_mem_inst_w_mem_13__15_), .Y(w_mem_inst__abc_19396_new_n2497_));
INVX1 INVX1_654 ( .A(\block[79] ), .Y(w_mem_inst__abc_19396_new_n2498_));
INVX1 INVX1_655 ( .A(w_mem_inst_w_mem_13__16_), .Y(w_mem_inst__abc_19396_new_n2502_));
INVX1 INVX1_656 ( .A(\block[80] ), .Y(w_mem_inst__abc_19396_new_n2503_));
INVX1 INVX1_657 ( .A(w_mem_inst_w_mem_13__17_), .Y(w_mem_inst__abc_19396_new_n2507_));
INVX1 INVX1_658 ( .A(\block[81] ), .Y(w_mem_inst__abc_19396_new_n2508_));
INVX1 INVX1_659 ( .A(w_mem_inst_w_mem_13__18_), .Y(w_mem_inst__abc_19396_new_n2512_));
INVX1 INVX1_66 ( .A(_abc_15497_new_n951_), .Y(_abc_15497_new_n952_));
INVX1 INVX1_660 ( .A(\block[82] ), .Y(w_mem_inst__abc_19396_new_n2513_));
INVX1 INVX1_661 ( .A(w_mem_inst_w_mem_13__19_), .Y(w_mem_inst__abc_19396_new_n2517_));
INVX1 INVX1_662 ( .A(\block[83] ), .Y(w_mem_inst__abc_19396_new_n2518_));
INVX1 INVX1_663 ( .A(w_mem_inst_w_mem_13__20_), .Y(w_mem_inst__abc_19396_new_n2522_));
INVX1 INVX1_664 ( .A(\block[84] ), .Y(w_mem_inst__abc_19396_new_n2523_));
INVX1 INVX1_665 ( .A(w_mem_inst_w_mem_13__21_), .Y(w_mem_inst__abc_19396_new_n2527_));
INVX1 INVX1_666 ( .A(\block[85] ), .Y(w_mem_inst__abc_19396_new_n2528_));
INVX1 INVX1_667 ( .A(w_mem_inst_w_mem_13__22_), .Y(w_mem_inst__abc_19396_new_n2532_));
INVX1 INVX1_668 ( .A(\block[86] ), .Y(w_mem_inst__abc_19396_new_n2533_));
INVX1 INVX1_669 ( .A(w_mem_inst_w_mem_13__23_), .Y(w_mem_inst__abc_19396_new_n2537_));
INVX1 INVX1_67 ( .A(_auto_iopadmap_cc_368_execute_22625_3_), .Y(_abc_15497_new_n955_));
INVX1 INVX1_670 ( .A(\block[87] ), .Y(w_mem_inst__abc_19396_new_n2538_));
INVX1 INVX1_671 ( .A(w_mem_inst_w_mem_13__24_), .Y(w_mem_inst__abc_19396_new_n2542_));
INVX1 INVX1_672 ( .A(\block[88] ), .Y(w_mem_inst__abc_19396_new_n2543_));
INVX1 INVX1_673 ( .A(w_mem_inst_w_mem_13__25_), .Y(w_mem_inst__abc_19396_new_n2547_));
INVX1 INVX1_674 ( .A(\block[89] ), .Y(w_mem_inst__abc_19396_new_n2548_));
INVX1 INVX1_675 ( .A(w_mem_inst_w_mem_13__26_), .Y(w_mem_inst__abc_19396_new_n2552_));
INVX1 INVX1_676 ( .A(\block[90] ), .Y(w_mem_inst__abc_19396_new_n2553_));
INVX1 INVX1_677 ( .A(w_mem_inst_w_mem_13__27_), .Y(w_mem_inst__abc_19396_new_n2557_));
INVX1 INVX1_678 ( .A(\block[91] ), .Y(w_mem_inst__abc_19396_new_n2558_));
INVX1 INVX1_679 ( .A(w_mem_inst_w_mem_13__28_), .Y(w_mem_inst__abc_19396_new_n2562_));
INVX1 INVX1_68 ( .A(e_reg_2_), .Y(_abc_15497_new_n956_));
INVX1 INVX1_680 ( .A(\block[92] ), .Y(w_mem_inst__abc_19396_new_n2563_));
INVX1 INVX1_681 ( .A(w_mem_inst_w_mem_13__29_), .Y(w_mem_inst__abc_19396_new_n2567_));
INVX1 INVX1_682 ( .A(\block[93] ), .Y(w_mem_inst__abc_19396_new_n2568_));
INVX1 INVX1_683 ( .A(w_mem_inst_w_mem_13__30_), .Y(w_mem_inst__abc_19396_new_n2572_));
INVX1 INVX1_684 ( .A(\block[94] ), .Y(w_mem_inst__abc_19396_new_n2573_));
INVX1 INVX1_685 ( .A(w_mem_inst_w_mem_13__31_), .Y(w_mem_inst__abc_19396_new_n2577_));
INVX1 INVX1_686 ( .A(\block[95] ), .Y(w_mem_inst__abc_19396_new_n2578_));
INVX1 INVX1_687 ( .A(w_mem_inst_w_mem_14__0_), .Y(w_mem_inst__abc_19396_new_n2647_));
INVX1 INVX1_688 ( .A(\block[32] ), .Y(w_mem_inst__abc_19396_new_n2648_));
INVX1 INVX1_689 ( .A(w_mem_inst_w_mem_14__1_), .Y(w_mem_inst__abc_19396_new_n2652_));
INVX1 INVX1_69 ( .A(_abc_15497_new_n958_), .Y(_abc_15497_new_n959_));
INVX1 INVX1_690 ( .A(\block[33] ), .Y(w_mem_inst__abc_19396_new_n2653_));
INVX1 INVX1_691 ( .A(w_mem_inst_w_mem_14__2_), .Y(w_mem_inst__abc_19396_new_n2657_));
INVX1 INVX1_692 ( .A(\block[34] ), .Y(w_mem_inst__abc_19396_new_n2658_));
INVX1 INVX1_693 ( .A(w_mem_inst_w_mem_14__3_), .Y(w_mem_inst__abc_19396_new_n2662_));
INVX1 INVX1_694 ( .A(\block[35] ), .Y(w_mem_inst__abc_19396_new_n2663_));
INVX1 INVX1_695 ( .A(w_mem_inst_w_mem_14__4_), .Y(w_mem_inst__abc_19396_new_n2667_));
INVX1 INVX1_696 ( .A(\block[36] ), .Y(w_mem_inst__abc_19396_new_n2668_));
INVX1 INVX1_697 ( .A(w_mem_inst_w_mem_14__5_), .Y(w_mem_inst__abc_19396_new_n2672_));
INVX1 INVX1_698 ( .A(\block[37] ), .Y(w_mem_inst__abc_19396_new_n2673_));
INVX1 INVX1_699 ( .A(w_mem_inst_w_mem_14__6_), .Y(w_mem_inst__abc_19396_new_n2677_));
INVX1 INVX1_7 ( .A(_abc_15497_new_n722_), .Y(_abc_15497_new_n723_));
INVX1 INVX1_70 ( .A(e_reg_3_), .Y(_abc_15497_new_n960_));
INVX1 INVX1_700 ( .A(\block[38] ), .Y(w_mem_inst__abc_19396_new_n2678_));
INVX1 INVX1_701 ( .A(w_mem_inst_w_mem_14__7_), .Y(w_mem_inst__abc_19396_new_n2682_));
INVX1 INVX1_702 ( .A(\block[39] ), .Y(w_mem_inst__abc_19396_new_n2683_));
INVX1 INVX1_703 ( .A(w_mem_inst_w_mem_14__8_), .Y(w_mem_inst__abc_19396_new_n2687_));
INVX1 INVX1_704 ( .A(\block[40] ), .Y(w_mem_inst__abc_19396_new_n2688_));
INVX1 INVX1_705 ( .A(w_mem_inst_w_mem_14__9_), .Y(w_mem_inst__abc_19396_new_n2692_));
INVX1 INVX1_706 ( .A(\block[41] ), .Y(w_mem_inst__abc_19396_new_n2693_));
INVX1 INVX1_707 ( .A(w_mem_inst_w_mem_14__10_), .Y(w_mem_inst__abc_19396_new_n2697_));
INVX1 INVX1_708 ( .A(\block[42] ), .Y(w_mem_inst__abc_19396_new_n2698_));
INVX1 INVX1_709 ( .A(w_mem_inst_w_mem_14__11_), .Y(w_mem_inst__abc_19396_new_n2702_));
INVX1 INVX1_71 ( .A(_abc_15497_new_n961_), .Y(_abc_15497_new_n962_));
INVX1 INVX1_710 ( .A(\block[43] ), .Y(w_mem_inst__abc_19396_new_n2703_));
INVX1 INVX1_711 ( .A(w_mem_inst_w_mem_14__12_), .Y(w_mem_inst__abc_19396_new_n2707_));
INVX1 INVX1_712 ( .A(\block[44] ), .Y(w_mem_inst__abc_19396_new_n2708_));
INVX1 INVX1_713 ( .A(w_mem_inst_w_mem_14__13_), .Y(w_mem_inst__abc_19396_new_n2712_));
INVX1 INVX1_714 ( .A(\block[45] ), .Y(w_mem_inst__abc_19396_new_n2713_));
INVX1 INVX1_715 ( .A(w_mem_inst_w_mem_14__14_), .Y(w_mem_inst__abc_19396_new_n2717_));
INVX1 INVX1_716 ( .A(\block[46] ), .Y(w_mem_inst__abc_19396_new_n2718_));
INVX1 INVX1_717 ( .A(w_mem_inst_w_mem_14__15_), .Y(w_mem_inst__abc_19396_new_n2722_));
INVX1 INVX1_718 ( .A(\block[47] ), .Y(w_mem_inst__abc_19396_new_n2723_));
INVX1 INVX1_719 ( .A(w_mem_inst_w_mem_14__16_), .Y(w_mem_inst__abc_19396_new_n2727_));
INVX1 INVX1_72 ( .A(_abc_15497_new_n970_), .Y(_abc_15497_new_n971_));
INVX1 INVX1_720 ( .A(\block[48] ), .Y(w_mem_inst__abc_19396_new_n2728_));
INVX1 INVX1_721 ( .A(w_mem_inst_w_mem_14__17_), .Y(w_mem_inst__abc_19396_new_n2732_));
INVX1 INVX1_722 ( .A(\block[49] ), .Y(w_mem_inst__abc_19396_new_n2733_));
INVX1 INVX1_723 ( .A(w_mem_inst_w_mem_14__18_), .Y(w_mem_inst__abc_19396_new_n2737_));
INVX1 INVX1_724 ( .A(\block[50] ), .Y(w_mem_inst__abc_19396_new_n2738_));
INVX1 INVX1_725 ( .A(w_mem_inst_w_mem_14__19_), .Y(w_mem_inst__abc_19396_new_n2742_));
INVX1 INVX1_726 ( .A(\block[51] ), .Y(w_mem_inst__abc_19396_new_n2743_));
INVX1 INVX1_727 ( .A(w_mem_inst_w_mem_14__20_), .Y(w_mem_inst__abc_19396_new_n2747_));
INVX1 INVX1_728 ( .A(\block[52] ), .Y(w_mem_inst__abc_19396_new_n2748_));
INVX1 INVX1_729 ( .A(w_mem_inst_w_mem_14__21_), .Y(w_mem_inst__abc_19396_new_n2752_));
INVX1 INVX1_73 ( .A(_abc_15497_new_n994_), .Y(_abc_15497_new_n995_));
INVX1 INVX1_730 ( .A(\block[53] ), .Y(w_mem_inst__abc_19396_new_n2753_));
INVX1 INVX1_731 ( .A(w_mem_inst_w_mem_14__22_), .Y(w_mem_inst__abc_19396_new_n2757_));
INVX1 INVX1_732 ( .A(\block[54] ), .Y(w_mem_inst__abc_19396_new_n2758_));
INVX1 INVX1_733 ( .A(w_mem_inst_w_mem_14__23_), .Y(w_mem_inst__abc_19396_new_n2762_));
INVX1 INVX1_734 ( .A(\block[55] ), .Y(w_mem_inst__abc_19396_new_n2763_));
INVX1 INVX1_735 ( .A(w_mem_inst_w_mem_14__24_), .Y(w_mem_inst__abc_19396_new_n2767_));
INVX1 INVX1_736 ( .A(\block[56] ), .Y(w_mem_inst__abc_19396_new_n2768_));
INVX1 INVX1_737 ( .A(w_mem_inst_w_mem_14__25_), .Y(w_mem_inst__abc_19396_new_n2772_));
INVX1 INVX1_738 ( .A(\block[57] ), .Y(w_mem_inst__abc_19396_new_n2773_));
INVX1 INVX1_739 ( .A(w_mem_inst_w_mem_14__26_), .Y(w_mem_inst__abc_19396_new_n2777_));
INVX1 INVX1_74 ( .A(_abc_15497_new_n997_), .Y(_abc_15497_new_n998_));
INVX1 INVX1_740 ( .A(\block[58] ), .Y(w_mem_inst__abc_19396_new_n2778_));
INVX1 INVX1_741 ( .A(w_mem_inst_w_mem_14__27_), .Y(w_mem_inst__abc_19396_new_n2782_));
INVX1 INVX1_742 ( .A(\block[59] ), .Y(w_mem_inst__abc_19396_new_n2783_));
INVX1 INVX1_743 ( .A(w_mem_inst_w_mem_14__28_), .Y(w_mem_inst__abc_19396_new_n2787_));
INVX1 INVX1_744 ( .A(\block[60] ), .Y(w_mem_inst__abc_19396_new_n2788_));
INVX1 INVX1_745 ( .A(w_mem_inst_w_mem_14__29_), .Y(w_mem_inst__abc_19396_new_n2792_));
INVX1 INVX1_746 ( .A(\block[61] ), .Y(w_mem_inst__abc_19396_new_n2793_));
INVX1 INVX1_747 ( .A(w_mem_inst_w_mem_14__30_), .Y(w_mem_inst__abc_19396_new_n2797_));
INVX1 INVX1_748 ( .A(\block[62] ), .Y(w_mem_inst__abc_19396_new_n2798_));
INVX1 INVX1_749 ( .A(w_mem_inst_w_mem_14__31_), .Y(w_mem_inst__abc_19396_new_n2802_));
INVX1 INVX1_75 ( .A(_abc_15497_new_n999_), .Y(_abc_15497_new_n1000_));
INVX1 INVX1_750 ( .A(\block[63] ), .Y(w_mem_inst__abc_19396_new_n2803_));
INVX1 INVX1_751 ( .A(w_mem_inst_w_mem_10__0_), .Y(w_mem_inst__abc_19396_new_n2807_));
INVX1 INVX1_752 ( .A(\block[160] ), .Y(w_mem_inst__abc_19396_new_n2808_));
INVX1 INVX1_753 ( .A(w_mem_inst_w_mem_10__1_), .Y(w_mem_inst__abc_19396_new_n2812_));
INVX1 INVX1_754 ( .A(\block[161] ), .Y(w_mem_inst__abc_19396_new_n2813_));
INVX1 INVX1_755 ( .A(w_mem_inst_w_mem_10__2_), .Y(w_mem_inst__abc_19396_new_n2817_));
INVX1 INVX1_756 ( .A(\block[162] ), .Y(w_mem_inst__abc_19396_new_n2818_));
INVX1 INVX1_757 ( .A(w_mem_inst_w_mem_10__3_), .Y(w_mem_inst__abc_19396_new_n2822_));
INVX1 INVX1_758 ( .A(\block[163] ), .Y(w_mem_inst__abc_19396_new_n2823_));
INVX1 INVX1_759 ( .A(w_mem_inst_w_mem_10__4_), .Y(w_mem_inst__abc_19396_new_n2827_));
INVX1 INVX1_76 ( .A(e_reg_8_), .Y(_abc_15497_new_n1006_));
INVX1 INVX1_760 ( .A(\block[164] ), .Y(w_mem_inst__abc_19396_new_n2828_));
INVX1 INVX1_761 ( .A(w_mem_inst_w_mem_10__5_), .Y(w_mem_inst__abc_19396_new_n2832_));
INVX1 INVX1_762 ( .A(\block[165] ), .Y(w_mem_inst__abc_19396_new_n2833_));
INVX1 INVX1_763 ( .A(w_mem_inst_w_mem_10__6_), .Y(w_mem_inst__abc_19396_new_n2837_));
INVX1 INVX1_764 ( .A(\block[166] ), .Y(w_mem_inst__abc_19396_new_n2838_));
INVX1 INVX1_765 ( .A(w_mem_inst_w_mem_10__7_), .Y(w_mem_inst__abc_19396_new_n2842_));
INVX1 INVX1_766 ( .A(\block[167] ), .Y(w_mem_inst__abc_19396_new_n2843_));
INVX1 INVX1_767 ( .A(w_mem_inst_w_mem_10__8_), .Y(w_mem_inst__abc_19396_new_n2847_));
INVX1 INVX1_768 ( .A(\block[168] ), .Y(w_mem_inst__abc_19396_new_n2848_));
INVX1 INVX1_769 ( .A(w_mem_inst_w_mem_10__9_), .Y(w_mem_inst__abc_19396_new_n2852_));
INVX1 INVX1_77 ( .A(_auto_iopadmap_cc_368_execute_22625_8_), .Y(_abc_15497_new_n1007_));
INVX1 INVX1_770 ( .A(\block[169] ), .Y(w_mem_inst__abc_19396_new_n2853_));
INVX1 INVX1_771 ( .A(w_mem_inst_w_mem_10__10_), .Y(w_mem_inst__abc_19396_new_n2857_));
INVX1 INVX1_772 ( .A(\block[170] ), .Y(w_mem_inst__abc_19396_new_n2858_));
INVX1 INVX1_773 ( .A(w_mem_inst_w_mem_10__11_), .Y(w_mem_inst__abc_19396_new_n2862_));
INVX1 INVX1_774 ( .A(\block[171] ), .Y(w_mem_inst__abc_19396_new_n2863_));
INVX1 INVX1_775 ( .A(w_mem_inst_w_mem_10__12_), .Y(w_mem_inst__abc_19396_new_n2867_));
INVX1 INVX1_776 ( .A(\block[172] ), .Y(w_mem_inst__abc_19396_new_n2868_));
INVX1 INVX1_777 ( .A(w_mem_inst_w_mem_10__13_), .Y(w_mem_inst__abc_19396_new_n2872_));
INVX1 INVX1_778 ( .A(\block[173] ), .Y(w_mem_inst__abc_19396_new_n2873_));
INVX1 INVX1_779 ( .A(w_mem_inst_w_mem_10__14_), .Y(w_mem_inst__abc_19396_new_n2877_));
INVX1 INVX1_78 ( .A(_auto_iopadmap_cc_368_execute_22625_9_), .Y(_abc_15497_new_n1024_));
INVX1 INVX1_780 ( .A(\block[174] ), .Y(w_mem_inst__abc_19396_new_n2878_));
INVX1 INVX1_781 ( .A(w_mem_inst_w_mem_10__15_), .Y(w_mem_inst__abc_19396_new_n2882_));
INVX1 INVX1_782 ( .A(\block[175] ), .Y(w_mem_inst__abc_19396_new_n2883_));
INVX1 INVX1_783 ( .A(w_mem_inst_w_mem_10__16_), .Y(w_mem_inst__abc_19396_new_n2887_));
INVX1 INVX1_784 ( .A(\block[176] ), .Y(w_mem_inst__abc_19396_new_n2888_));
INVX1 INVX1_785 ( .A(w_mem_inst_w_mem_10__17_), .Y(w_mem_inst__abc_19396_new_n2892_));
INVX1 INVX1_786 ( .A(\block[177] ), .Y(w_mem_inst__abc_19396_new_n2893_));
INVX1 INVX1_787 ( .A(w_mem_inst_w_mem_10__18_), .Y(w_mem_inst__abc_19396_new_n2897_));
INVX1 INVX1_788 ( .A(\block[178] ), .Y(w_mem_inst__abc_19396_new_n2898_));
INVX1 INVX1_789 ( .A(w_mem_inst_w_mem_10__19_), .Y(w_mem_inst__abc_19396_new_n2902_));
INVX1 INVX1_79 ( .A(_abc_15497_new_n1027_), .Y(_abc_15497_new_n1028_));
INVX1 INVX1_790 ( .A(\block[179] ), .Y(w_mem_inst__abc_19396_new_n2903_));
INVX1 INVX1_791 ( .A(w_mem_inst_w_mem_10__20_), .Y(w_mem_inst__abc_19396_new_n2907_));
INVX1 INVX1_792 ( .A(\block[180] ), .Y(w_mem_inst__abc_19396_new_n2908_));
INVX1 INVX1_793 ( .A(w_mem_inst_w_mem_10__21_), .Y(w_mem_inst__abc_19396_new_n2912_));
INVX1 INVX1_794 ( .A(\block[181] ), .Y(w_mem_inst__abc_19396_new_n2913_));
INVX1 INVX1_795 ( .A(w_mem_inst_w_mem_10__22_), .Y(w_mem_inst__abc_19396_new_n2917_));
INVX1 INVX1_796 ( .A(\block[182] ), .Y(w_mem_inst__abc_19396_new_n2918_));
INVX1 INVX1_797 ( .A(w_mem_inst_w_mem_10__23_), .Y(w_mem_inst__abc_19396_new_n2922_));
INVX1 INVX1_798 ( .A(\block[183] ), .Y(w_mem_inst__abc_19396_new_n2923_));
INVX1 INVX1_799 ( .A(w_mem_inst_w_mem_10__24_), .Y(w_mem_inst__abc_19396_new_n2927_));
INVX1 INVX1_8 ( .A(_abc_15497_new_n724_), .Y(_abc_15497_new_n725_));
INVX1 INVX1_80 ( .A(_auto_iopadmap_cc_368_execute_22625_10_), .Y(_abc_15497_new_n1033_));
INVX1 INVX1_800 ( .A(\block[184] ), .Y(w_mem_inst__abc_19396_new_n2928_));
INVX1 INVX1_801 ( .A(w_mem_inst_w_mem_10__25_), .Y(w_mem_inst__abc_19396_new_n2932_));
INVX1 INVX1_802 ( .A(\block[185] ), .Y(w_mem_inst__abc_19396_new_n2933_));
INVX1 INVX1_803 ( .A(w_mem_inst_w_mem_10__26_), .Y(w_mem_inst__abc_19396_new_n2937_));
INVX1 INVX1_804 ( .A(\block[186] ), .Y(w_mem_inst__abc_19396_new_n2938_));
INVX1 INVX1_805 ( .A(w_mem_inst_w_mem_10__27_), .Y(w_mem_inst__abc_19396_new_n2942_));
INVX1 INVX1_806 ( .A(\block[187] ), .Y(w_mem_inst__abc_19396_new_n2943_));
INVX1 INVX1_807 ( .A(w_mem_inst_w_mem_10__28_), .Y(w_mem_inst__abc_19396_new_n2947_));
INVX1 INVX1_808 ( .A(\block[188] ), .Y(w_mem_inst__abc_19396_new_n2948_));
INVX1 INVX1_809 ( .A(w_mem_inst_w_mem_10__29_), .Y(w_mem_inst__abc_19396_new_n2952_));
INVX1 INVX1_81 ( .A(e_reg_9_), .Y(_abc_15497_new_n1034_));
INVX1 INVX1_810 ( .A(\block[189] ), .Y(w_mem_inst__abc_19396_new_n2953_));
INVX1 INVX1_811 ( .A(w_mem_inst_w_mem_10__30_), .Y(w_mem_inst__abc_19396_new_n2957_));
INVX1 INVX1_812 ( .A(\block[190] ), .Y(w_mem_inst__abc_19396_new_n2958_));
INVX1 INVX1_813 ( .A(w_mem_inst_w_mem_10__31_), .Y(w_mem_inst__abc_19396_new_n2962_));
INVX1 INVX1_814 ( .A(\block[191] ), .Y(w_mem_inst__abc_19396_new_n2963_));
INVX1 INVX1_815 ( .A(w_mem_inst_w_mem_12__0_), .Y(w_mem_inst__abc_19396_new_n2967_));
INVX1 INVX1_816 ( .A(\block[96] ), .Y(w_mem_inst__abc_19396_new_n2968_));
INVX1 INVX1_817 ( .A(w_mem_inst_w_mem_12__1_), .Y(w_mem_inst__abc_19396_new_n2972_));
INVX1 INVX1_818 ( .A(\block[97] ), .Y(w_mem_inst__abc_19396_new_n2973_));
INVX1 INVX1_819 ( .A(w_mem_inst_w_mem_12__2_), .Y(w_mem_inst__abc_19396_new_n2977_));
INVX1 INVX1_82 ( .A(_abc_15497_new_n1036_), .Y(_abc_15497_new_n1037_));
INVX1 INVX1_820 ( .A(\block[98] ), .Y(w_mem_inst__abc_19396_new_n2978_));
INVX1 INVX1_821 ( .A(w_mem_inst_w_mem_12__3_), .Y(w_mem_inst__abc_19396_new_n2982_));
INVX1 INVX1_822 ( .A(\block[99] ), .Y(w_mem_inst__abc_19396_new_n2983_));
INVX1 INVX1_823 ( .A(w_mem_inst_w_mem_12__4_), .Y(w_mem_inst__abc_19396_new_n2987_));
INVX1 INVX1_824 ( .A(\block[100] ), .Y(w_mem_inst__abc_19396_new_n2988_));
INVX1 INVX1_825 ( .A(w_mem_inst_w_mem_12__5_), .Y(w_mem_inst__abc_19396_new_n2992_));
INVX1 INVX1_826 ( .A(\block[101] ), .Y(w_mem_inst__abc_19396_new_n2993_));
INVX1 INVX1_827 ( .A(w_mem_inst_w_mem_12__6_), .Y(w_mem_inst__abc_19396_new_n2997_));
INVX1 INVX1_828 ( .A(\block[102] ), .Y(w_mem_inst__abc_19396_new_n2998_));
INVX1 INVX1_829 ( .A(w_mem_inst_w_mem_12__7_), .Y(w_mem_inst__abc_19396_new_n3002_));
INVX1 INVX1_83 ( .A(_abc_15497_new_n1040_), .Y(_abc_15497_new_n1041_));
INVX1 INVX1_830 ( .A(\block[103] ), .Y(w_mem_inst__abc_19396_new_n3003_));
INVX1 INVX1_831 ( .A(w_mem_inst_w_mem_12__8_), .Y(w_mem_inst__abc_19396_new_n3007_));
INVX1 INVX1_832 ( .A(\block[104] ), .Y(w_mem_inst__abc_19396_new_n3008_));
INVX1 INVX1_833 ( .A(w_mem_inst_w_mem_12__9_), .Y(w_mem_inst__abc_19396_new_n3012_));
INVX1 INVX1_834 ( .A(\block[105] ), .Y(w_mem_inst__abc_19396_new_n3013_));
INVX1 INVX1_835 ( .A(w_mem_inst_w_mem_12__10_), .Y(w_mem_inst__abc_19396_new_n3017_));
INVX1 INVX1_836 ( .A(\block[106] ), .Y(w_mem_inst__abc_19396_new_n3018_));
INVX1 INVX1_837 ( .A(w_mem_inst_w_mem_12__11_), .Y(w_mem_inst__abc_19396_new_n3022_));
INVX1 INVX1_838 ( .A(\block[107] ), .Y(w_mem_inst__abc_19396_new_n3023_));
INVX1 INVX1_839 ( .A(w_mem_inst_w_mem_12__12_), .Y(w_mem_inst__abc_19396_new_n3027_));
INVX1 INVX1_84 ( .A(_abc_15497_new_n1042_), .Y(_abc_15497_new_n1043_));
INVX1 INVX1_840 ( .A(\block[108] ), .Y(w_mem_inst__abc_19396_new_n3028_));
INVX1 INVX1_841 ( .A(w_mem_inst_w_mem_12__13_), .Y(w_mem_inst__abc_19396_new_n3032_));
INVX1 INVX1_842 ( .A(\block[109] ), .Y(w_mem_inst__abc_19396_new_n3033_));
INVX1 INVX1_843 ( .A(w_mem_inst_w_mem_12__14_), .Y(w_mem_inst__abc_19396_new_n3037_));
INVX1 INVX1_844 ( .A(\block[110] ), .Y(w_mem_inst__abc_19396_new_n3038_));
INVX1 INVX1_845 ( .A(w_mem_inst_w_mem_12__15_), .Y(w_mem_inst__abc_19396_new_n3042_));
INVX1 INVX1_846 ( .A(\block[111] ), .Y(w_mem_inst__abc_19396_new_n3043_));
INVX1 INVX1_847 ( .A(w_mem_inst_w_mem_12__16_), .Y(w_mem_inst__abc_19396_new_n3047_));
INVX1 INVX1_848 ( .A(\block[112] ), .Y(w_mem_inst__abc_19396_new_n3048_));
INVX1 INVX1_849 ( .A(w_mem_inst_w_mem_12__17_), .Y(w_mem_inst__abc_19396_new_n3052_));
INVX1 INVX1_85 ( .A(_auto_iopadmap_cc_368_execute_22625_11_), .Y(_abc_15497_new_n1048_));
INVX1 INVX1_850 ( .A(\block[113] ), .Y(w_mem_inst__abc_19396_new_n3053_));
INVX1 INVX1_851 ( .A(w_mem_inst_w_mem_12__18_), .Y(w_mem_inst__abc_19396_new_n3057_));
INVX1 INVX1_852 ( .A(\block[114] ), .Y(w_mem_inst__abc_19396_new_n3058_));
INVX1 INVX1_853 ( .A(w_mem_inst_w_mem_12__19_), .Y(w_mem_inst__abc_19396_new_n3062_));
INVX1 INVX1_854 ( .A(\block[115] ), .Y(w_mem_inst__abc_19396_new_n3063_));
INVX1 INVX1_855 ( .A(w_mem_inst_w_mem_12__20_), .Y(w_mem_inst__abc_19396_new_n3067_));
INVX1 INVX1_856 ( .A(\block[116] ), .Y(w_mem_inst__abc_19396_new_n3068_));
INVX1 INVX1_857 ( .A(w_mem_inst_w_mem_12__21_), .Y(w_mem_inst__abc_19396_new_n3072_));
INVX1 INVX1_858 ( .A(\block[117] ), .Y(w_mem_inst__abc_19396_new_n3073_));
INVX1 INVX1_859 ( .A(w_mem_inst_w_mem_12__22_), .Y(w_mem_inst__abc_19396_new_n3077_));
INVX1 INVX1_86 ( .A(e_reg_10_), .Y(_abc_15497_new_n1049_));
INVX1 INVX1_860 ( .A(\block[118] ), .Y(w_mem_inst__abc_19396_new_n3078_));
INVX1 INVX1_861 ( .A(w_mem_inst_w_mem_12__23_), .Y(w_mem_inst__abc_19396_new_n3082_));
INVX1 INVX1_862 ( .A(\block[119] ), .Y(w_mem_inst__abc_19396_new_n3083_));
INVX1 INVX1_863 ( .A(w_mem_inst_w_mem_12__24_), .Y(w_mem_inst__abc_19396_new_n3087_));
INVX1 INVX1_864 ( .A(\block[120] ), .Y(w_mem_inst__abc_19396_new_n3088_));
INVX1 INVX1_865 ( .A(w_mem_inst_w_mem_12__25_), .Y(w_mem_inst__abc_19396_new_n3092_));
INVX1 INVX1_866 ( .A(\block[121] ), .Y(w_mem_inst__abc_19396_new_n3093_));
INVX1 INVX1_867 ( .A(w_mem_inst_w_mem_12__26_), .Y(w_mem_inst__abc_19396_new_n3097_));
INVX1 INVX1_868 ( .A(\block[122] ), .Y(w_mem_inst__abc_19396_new_n3098_));
INVX1 INVX1_869 ( .A(w_mem_inst_w_mem_12__27_), .Y(w_mem_inst__abc_19396_new_n3102_));
INVX1 INVX1_87 ( .A(_abc_15497_new_n1051_), .Y(_abc_15497_new_n1052_));
INVX1 INVX1_870 ( .A(\block[123] ), .Y(w_mem_inst__abc_19396_new_n3103_));
INVX1 INVX1_871 ( .A(w_mem_inst_w_mem_12__28_), .Y(w_mem_inst__abc_19396_new_n3107_));
INVX1 INVX1_872 ( .A(\block[124] ), .Y(w_mem_inst__abc_19396_new_n3108_));
INVX1 INVX1_873 ( .A(w_mem_inst_w_mem_12__29_), .Y(w_mem_inst__abc_19396_new_n3112_));
INVX1 INVX1_874 ( .A(\block[125] ), .Y(w_mem_inst__abc_19396_new_n3113_));
INVX1 INVX1_875 ( .A(w_mem_inst_w_mem_12__30_), .Y(w_mem_inst__abc_19396_new_n3117_));
INVX1 INVX1_876 ( .A(\block[126] ), .Y(w_mem_inst__abc_19396_new_n3118_));
INVX1 INVX1_877 ( .A(w_mem_inst_w_mem_12__31_), .Y(w_mem_inst__abc_19396_new_n3122_));
INVX1 INVX1_878 ( .A(\block[127] ), .Y(w_mem_inst__abc_19396_new_n3123_));
INVX1 INVX1_879 ( .A(w_mem_inst_w_mem_11__0_), .Y(w_mem_inst__abc_19396_new_n3127_));
INVX1 INVX1_88 ( .A(_abc_15497_new_n1058_), .Y(_abc_15497_new_n1059_));
INVX1 INVX1_880 ( .A(\block[128] ), .Y(w_mem_inst__abc_19396_new_n3128_));
INVX1 INVX1_881 ( .A(w_mem_inst_w_mem_11__1_), .Y(w_mem_inst__abc_19396_new_n3132_));
INVX1 INVX1_882 ( .A(\block[129] ), .Y(w_mem_inst__abc_19396_new_n3133_));
INVX1 INVX1_883 ( .A(w_mem_inst_w_mem_11__2_), .Y(w_mem_inst__abc_19396_new_n3137_));
INVX1 INVX1_884 ( .A(\block[130] ), .Y(w_mem_inst__abc_19396_new_n3138_));
INVX1 INVX1_885 ( .A(w_mem_inst_w_mem_11__3_), .Y(w_mem_inst__abc_19396_new_n3142_));
INVX1 INVX1_886 ( .A(\block[131] ), .Y(w_mem_inst__abc_19396_new_n3143_));
INVX1 INVX1_887 ( .A(w_mem_inst_w_mem_11__4_), .Y(w_mem_inst__abc_19396_new_n3147_));
INVX1 INVX1_888 ( .A(\block[132] ), .Y(w_mem_inst__abc_19396_new_n3148_));
INVX1 INVX1_889 ( .A(w_mem_inst_w_mem_11__5_), .Y(w_mem_inst__abc_19396_new_n3152_));
INVX1 INVX1_89 ( .A(_abc_15497_new_n1073_), .Y(_abc_15497_new_n1074_));
INVX1 INVX1_890 ( .A(\block[133] ), .Y(w_mem_inst__abc_19396_new_n3153_));
INVX1 INVX1_891 ( .A(w_mem_inst_w_mem_11__6_), .Y(w_mem_inst__abc_19396_new_n3157_));
INVX1 INVX1_892 ( .A(\block[134] ), .Y(w_mem_inst__abc_19396_new_n3158_));
INVX1 INVX1_893 ( .A(w_mem_inst_w_mem_11__7_), .Y(w_mem_inst__abc_19396_new_n3162_));
INVX1 INVX1_894 ( .A(\block[135] ), .Y(w_mem_inst__abc_19396_new_n3163_));
INVX1 INVX1_895 ( .A(w_mem_inst_w_mem_11__8_), .Y(w_mem_inst__abc_19396_new_n3167_));
INVX1 INVX1_896 ( .A(\block[136] ), .Y(w_mem_inst__abc_19396_new_n3168_));
INVX1 INVX1_897 ( .A(w_mem_inst_w_mem_11__9_), .Y(w_mem_inst__abc_19396_new_n3172_));
INVX1 INVX1_898 ( .A(\block[137] ), .Y(w_mem_inst__abc_19396_new_n3173_));
INVX1 INVX1_899 ( .A(w_mem_inst_w_mem_11__10_), .Y(w_mem_inst__abc_19396_new_n3177_));
INVX1 INVX1_9 ( .A(c_reg_10_), .Y(_abc_15497_new_n727_));
INVX1 INVX1_90 ( .A(_auto_iopadmap_cc_368_execute_22625_14_), .Y(_abc_15497_new_n1081_));
INVX1 INVX1_900 ( .A(\block[138] ), .Y(w_mem_inst__abc_19396_new_n3178_));
INVX1 INVX1_901 ( .A(w_mem_inst_w_mem_11__11_), .Y(w_mem_inst__abc_19396_new_n3182_));
INVX1 INVX1_902 ( .A(\block[139] ), .Y(w_mem_inst__abc_19396_new_n3183_));
INVX1 INVX1_903 ( .A(w_mem_inst_w_mem_11__12_), .Y(w_mem_inst__abc_19396_new_n3187_));
INVX1 INVX1_904 ( .A(\block[140] ), .Y(w_mem_inst__abc_19396_new_n3188_));
INVX1 INVX1_905 ( .A(w_mem_inst_w_mem_11__13_), .Y(w_mem_inst__abc_19396_new_n3192_));
INVX1 INVX1_906 ( .A(\block[141] ), .Y(w_mem_inst__abc_19396_new_n3193_));
INVX1 INVX1_907 ( .A(w_mem_inst_w_mem_11__14_), .Y(w_mem_inst__abc_19396_new_n3197_));
INVX1 INVX1_908 ( .A(\block[142] ), .Y(w_mem_inst__abc_19396_new_n3198_));
INVX1 INVX1_909 ( .A(w_mem_inst_w_mem_11__15_), .Y(w_mem_inst__abc_19396_new_n3202_));
INVX1 INVX1_91 ( .A(_abc_15497_new_n1062_), .Y(_abc_15497_new_n1084_));
INVX1 INVX1_910 ( .A(\block[143] ), .Y(w_mem_inst__abc_19396_new_n3203_));
INVX1 INVX1_911 ( .A(w_mem_inst_w_mem_11__16_), .Y(w_mem_inst__abc_19396_new_n3207_));
INVX1 INVX1_912 ( .A(\block[144] ), .Y(w_mem_inst__abc_19396_new_n3208_));
INVX1 INVX1_913 ( .A(w_mem_inst_w_mem_11__17_), .Y(w_mem_inst__abc_19396_new_n3212_));
INVX1 INVX1_914 ( .A(\block[145] ), .Y(w_mem_inst__abc_19396_new_n3213_));
INVX1 INVX1_915 ( .A(w_mem_inst_w_mem_11__18_), .Y(w_mem_inst__abc_19396_new_n3217_));
INVX1 INVX1_916 ( .A(\block[146] ), .Y(w_mem_inst__abc_19396_new_n3218_));
INVX1 INVX1_917 ( .A(w_mem_inst_w_mem_11__19_), .Y(w_mem_inst__abc_19396_new_n3222_));
INVX1 INVX1_918 ( .A(\block[147] ), .Y(w_mem_inst__abc_19396_new_n3223_));
INVX1 INVX1_919 ( .A(w_mem_inst_w_mem_11__20_), .Y(w_mem_inst__abc_19396_new_n3227_));
INVX1 INVX1_92 ( .A(_abc_15497_new_n1095_), .Y(_abc_15497_new_n1096_));
INVX1 INVX1_920 ( .A(\block[148] ), .Y(w_mem_inst__abc_19396_new_n3228_));
INVX1 INVX1_921 ( .A(w_mem_inst_w_mem_11__21_), .Y(w_mem_inst__abc_19396_new_n3232_));
INVX1 INVX1_922 ( .A(\block[149] ), .Y(w_mem_inst__abc_19396_new_n3233_));
INVX1 INVX1_923 ( .A(w_mem_inst_w_mem_11__22_), .Y(w_mem_inst__abc_19396_new_n3237_));
INVX1 INVX1_924 ( .A(\block[150] ), .Y(w_mem_inst__abc_19396_new_n3238_));
INVX1 INVX1_925 ( .A(w_mem_inst_w_mem_11__23_), .Y(w_mem_inst__abc_19396_new_n3242_));
INVX1 INVX1_926 ( .A(\block[151] ), .Y(w_mem_inst__abc_19396_new_n3243_));
INVX1 INVX1_927 ( .A(w_mem_inst_w_mem_11__24_), .Y(w_mem_inst__abc_19396_new_n3247_));
INVX1 INVX1_928 ( .A(\block[152] ), .Y(w_mem_inst__abc_19396_new_n3248_));
INVX1 INVX1_929 ( .A(w_mem_inst_w_mem_11__25_), .Y(w_mem_inst__abc_19396_new_n3252_));
INVX1 INVX1_93 ( .A(_abc_15497_new_n1061_), .Y(_abc_15497_new_n1102_));
INVX1 INVX1_930 ( .A(\block[153] ), .Y(w_mem_inst__abc_19396_new_n3253_));
INVX1 INVX1_931 ( .A(w_mem_inst_w_mem_11__26_), .Y(w_mem_inst__abc_19396_new_n3257_));
INVX1 INVX1_932 ( .A(\block[154] ), .Y(w_mem_inst__abc_19396_new_n3258_));
INVX1 INVX1_933 ( .A(w_mem_inst_w_mem_11__27_), .Y(w_mem_inst__abc_19396_new_n3262_));
INVX1 INVX1_934 ( .A(\block[155] ), .Y(w_mem_inst__abc_19396_new_n3263_));
INVX1 INVX1_935 ( .A(w_mem_inst_w_mem_11__28_), .Y(w_mem_inst__abc_19396_new_n3267_));
INVX1 INVX1_936 ( .A(\block[156] ), .Y(w_mem_inst__abc_19396_new_n3268_));
INVX1 INVX1_937 ( .A(w_mem_inst_w_mem_11__29_), .Y(w_mem_inst__abc_19396_new_n3272_));
INVX1 INVX1_938 ( .A(\block[157] ), .Y(w_mem_inst__abc_19396_new_n3273_));
INVX1 INVX1_939 ( .A(w_mem_inst_w_mem_11__30_), .Y(w_mem_inst__abc_19396_new_n3277_));
INVX1 INVX1_94 ( .A(_auto_iopadmap_cc_368_execute_22625_17_), .Y(_abc_15497_new_n1122_));
INVX1 INVX1_940 ( .A(\block[158] ), .Y(w_mem_inst__abc_19396_new_n3278_));
INVX1 INVX1_941 ( .A(w_mem_inst_w_mem_11__31_), .Y(w_mem_inst__abc_19396_new_n3282_));
INVX1 INVX1_942 ( .A(\block[159] ), .Y(w_mem_inst__abc_19396_new_n3283_));
INVX1 INVX1_943 ( .A(\block[256] ), .Y(w_mem_inst__abc_19396_new_n3287_));
INVX1 INVX1_944 ( .A(\block[257] ), .Y(w_mem_inst__abc_19396_new_n3291_));
INVX1 INVX1_945 ( .A(\block[258] ), .Y(w_mem_inst__abc_19396_new_n3295_));
INVX1 INVX1_946 ( .A(\block[259] ), .Y(w_mem_inst__abc_19396_new_n3299_));
INVX1 INVX1_947 ( .A(\block[260] ), .Y(w_mem_inst__abc_19396_new_n3303_));
INVX1 INVX1_948 ( .A(\block[261] ), .Y(w_mem_inst__abc_19396_new_n3307_));
INVX1 INVX1_949 ( .A(\block[262] ), .Y(w_mem_inst__abc_19396_new_n3311_));
INVX1 INVX1_95 ( .A(_auto_iopadmap_cc_368_execute_22625_18_), .Y(_abc_15497_new_n1128_));
INVX1 INVX1_950 ( .A(\block[263] ), .Y(w_mem_inst__abc_19396_new_n3315_));
INVX1 INVX1_951 ( .A(\block[264] ), .Y(w_mem_inst__abc_19396_new_n3319_));
INVX1 INVX1_952 ( .A(\block[265] ), .Y(w_mem_inst__abc_19396_new_n3323_));
INVX1 INVX1_953 ( .A(\block[266] ), .Y(w_mem_inst__abc_19396_new_n3327_));
INVX1 INVX1_954 ( .A(\block[267] ), .Y(w_mem_inst__abc_19396_new_n3331_));
INVX1 INVX1_955 ( .A(\block[268] ), .Y(w_mem_inst__abc_19396_new_n3335_));
INVX1 INVX1_956 ( .A(\block[269] ), .Y(w_mem_inst__abc_19396_new_n3339_));
INVX1 INVX1_957 ( .A(\block[270] ), .Y(w_mem_inst__abc_19396_new_n3343_));
INVX1 INVX1_958 ( .A(\block[271] ), .Y(w_mem_inst__abc_19396_new_n3347_));
INVX1 INVX1_959 ( .A(\block[272] ), .Y(w_mem_inst__abc_19396_new_n3351_));
INVX1 INVX1_96 ( .A(_abc_15497_new_n1132_), .Y(_abc_15497_new_n1133_));
INVX1 INVX1_960 ( .A(\block[273] ), .Y(w_mem_inst__abc_19396_new_n3355_));
INVX1 INVX1_961 ( .A(\block[274] ), .Y(w_mem_inst__abc_19396_new_n3359_));
INVX1 INVX1_962 ( .A(\block[275] ), .Y(w_mem_inst__abc_19396_new_n3363_));
INVX1 INVX1_963 ( .A(\block[276] ), .Y(w_mem_inst__abc_19396_new_n3367_));
INVX1 INVX1_964 ( .A(\block[277] ), .Y(w_mem_inst__abc_19396_new_n3371_));
INVX1 INVX1_965 ( .A(\block[278] ), .Y(w_mem_inst__abc_19396_new_n3375_));
INVX1 INVX1_966 ( .A(\block[279] ), .Y(w_mem_inst__abc_19396_new_n3379_));
INVX1 INVX1_967 ( .A(\block[280] ), .Y(w_mem_inst__abc_19396_new_n3383_));
INVX1 INVX1_968 ( .A(\block[281] ), .Y(w_mem_inst__abc_19396_new_n3387_));
INVX1 INVX1_969 ( .A(\block[282] ), .Y(w_mem_inst__abc_19396_new_n3391_));
INVX1 INVX1_97 ( .A(_abc_15497_new_n1116_), .Y(_abc_15497_new_n1134_));
INVX1 INVX1_970 ( .A(\block[283] ), .Y(w_mem_inst__abc_19396_new_n3395_));
INVX1 INVX1_971 ( .A(\block[284] ), .Y(w_mem_inst__abc_19396_new_n3399_));
INVX1 INVX1_972 ( .A(\block[285] ), .Y(w_mem_inst__abc_19396_new_n3403_));
INVX1 INVX1_973 ( .A(\block[286] ), .Y(w_mem_inst__abc_19396_new_n3407_));
INVX1 INVX1_974 ( .A(\block[287] ), .Y(w_mem_inst__abc_19396_new_n3411_));
INVX1 INVX1_975 ( .A(w_mem_inst_w_mem_9__0_), .Y(w_mem_inst__abc_19396_new_n3415_));
INVX1 INVX1_976 ( .A(\block[192] ), .Y(w_mem_inst__abc_19396_new_n3416_));
INVX1 INVX1_977 ( .A(w_mem_inst_w_mem_9__1_), .Y(w_mem_inst__abc_19396_new_n3420_));
INVX1 INVX1_978 ( .A(\block[193] ), .Y(w_mem_inst__abc_19396_new_n3421_));
INVX1 INVX1_979 ( .A(w_mem_inst_w_mem_9__2_), .Y(w_mem_inst__abc_19396_new_n3425_));
INVX1 INVX1_98 ( .A(_abc_15497_new_n1120_), .Y(_abc_15497_new_n1135_));
INVX1 INVX1_980 ( .A(\block[194] ), .Y(w_mem_inst__abc_19396_new_n3426_));
INVX1 INVX1_981 ( .A(w_mem_inst_w_mem_9__3_), .Y(w_mem_inst__abc_19396_new_n3430_));
INVX1 INVX1_982 ( .A(\block[195] ), .Y(w_mem_inst__abc_19396_new_n3431_));
INVX1 INVX1_983 ( .A(w_mem_inst_w_mem_9__4_), .Y(w_mem_inst__abc_19396_new_n3435_));
INVX1 INVX1_984 ( .A(\block[196] ), .Y(w_mem_inst__abc_19396_new_n3436_));
INVX1 INVX1_985 ( .A(w_mem_inst_w_mem_9__5_), .Y(w_mem_inst__abc_19396_new_n3440_));
INVX1 INVX1_986 ( .A(\block[197] ), .Y(w_mem_inst__abc_19396_new_n3441_));
INVX1 INVX1_987 ( .A(w_mem_inst_w_mem_9__6_), .Y(w_mem_inst__abc_19396_new_n3445_));
INVX1 INVX1_988 ( .A(\block[198] ), .Y(w_mem_inst__abc_19396_new_n3446_));
INVX1 INVX1_989 ( .A(w_mem_inst_w_mem_9__7_), .Y(w_mem_inst__abc_19396_new_n3450_));
INVX1 INVX1_99 ( .A(_abc_15497_new_n1113_), .Y(_abc_15497_new_n1136_));
INVX1 INVX1_990 ( .A(\block[199] ), .Y(w_mem_inst__abc_19396_new_n3451_));
INVX1 INVX1_991 ( .A(w_mem_inst_w_mem_9__8_), .Y(w_mem_inst__abc_19396_new_n3455_));
INVX1 INVX1_992 ( .A(\block[200] ), .Y(w_mem_inst__abc_19396_new_n3456_));
INVX1 INVX1_993 ( .A(w_mem_inst_w_mem_9__9_), .Y(w_mem_inst__abc_19396_new_n3460_));
INVX1 INVX1_994 ( .A(\block[201] ), .Y(w_mem_inst__abc_19396_new_n3461_));
INVX1 INVX1_995 ( .A(w_mem_inst_w_mem_9__10_), .Y(w_mem_inst__abc_19396_new_n3465_));
INVX1 INVX1_996 ( .A(\block[202] ), .Y(w_mem_inst__abc_19396_new_n3466_));
INVX1 INVX1_997 ( .A(w_mem_inst_w_mem_9__11_), .Y(w_mem_inst__abc_19396_new_n3470_));
INVX1 INVX1_998 ( .A(\block[203] ), .Y(w_mem_inst__abc_19396_new_n3471_));
INVX1 INVX1_999 ( .A(w_mem_inst_w_mem_9__12_), .Y(w_mem_inst__abc_19396_new_n3475_));
INVX2 INVX2_1 ( .A(_auto_iopadmap_cc_368_execute_22625_90_), .Y(_abc_15497_new_n698_));
INVX2 INVX2_10 ( .A(e_reg_12_), .Y(_abc_15497_new_n1064_));
INVX2 INVX2_11 ( .A(e_reg_14_), .Y(_abc_15497_new_n1080_));
INVX2 INVX2_12 ( .A(_auto_iopadmap_cc_368_execute_22625_16_), .Y(_abc_15497_new_n1101_));
INVX2 INVX2_13 ( .A(e_reg_16_), .Y(_abc_15497_new_n1112_));
INVX2 INVX2_14 ( .A(e_reg_17_), .Y(_abc_15497_new_n1121_));
INVX2 INVX2_15 ( .A(e_reg_18_), .Y(_abc_15497_new_n1130_));
INVX2 INVX2_16 ( .A(e_reg_19_), .Y(_abc_15497_new_n1146_));
INVX2 INVX2_17 ( .A(e_reg_20_), .Y(_abc_15497_new_n1162_));
INVX2 INVX2_18 ( .A(_auto_iopadmap_cc_368_execute_22625_21_), .Y(_abc_15497_new_n1171_));
INVX2 INVX2_19 ( .A(e_reg_21_), .Y(_abc_15497_new_n1173_));
INVX2 INVX2_2 ( .A(c_reg_14_), .Y(_abc_15497_new_n702_));
INVX2 INVX2_20 ( .A(_auto_iopadmap_cc_368_execute_22625_26_), .Y(_abc_15497_new_n1231_));
INVX2 INVX2_21 ( .A(e_reg_26_), .Y(_abc_15497_new_n1239_));
INVX2 INVX2_22 ( .A(_auto_iopadmap_cc_368_execute_22625_27_), .Y(_abc_15497_new_n1247_));
INVX2 INVX2_23 ( .A(e_reg_27_), .Y(_abc_15497_new_n1250_));
INVX2 INVX2_24 ( .A(e_reg_29_), .Y(_abc_15497_new_n1273_));
INVX2 INVX2_25 ( .A(d_reg_0_), .Y(_abc_15497_new_n1299_));
INVX2 INVX2_26 ( .A(d_reg_1_), .Y(_abc_15497_new_n1308_));
INVX2 INVX2_27 ( .A(d_reg_3_), .Y(_abc_15497_new_n1320_));
INVX2 INVX2_28 ( .A(d_reg_4_), .Y(_abc_15497_new_n1333_));
INVX2 INVX2_29 ( .A(d_reg_5_), .Y(_abc_15497_new_n1343_));
INVX2 INVX2_3 ( .A(c_reg_0_), .Y(_abc_15497_new_n769_));
INVX2 INVX2_30 ( .A(d_reg_7_), .Y(_abc_15497_new_n1353_));
INVX2 INVX2_31 ( .A(d_reg_6_), .Y(_abc_15497_new_n1357_));
INVX2 INVX2_32 ( .A(_auto_iopadmap_cc_368_execute_22625_40_), .Y(_abc_15497_new_n1361_));
INVX2 INVX2_33 ( .A(_abc_15497_new_n1366_), .Y(_abc_15497_new_n1367_));
INVX2 INVX2_34 ( .A(d_reg_9_), .Y(_abc_15497_new_n1374_));
INVX2 INVX2_35 ( .A(d_reg_11_), .Y(_abc_15497_new_n1398_));
INVX2 INVX2_36 ( .A(d_reg_12_), .Y(_abc_15497_new_n1414_));
INVX2 INVX2_37 ( .A(d_reg_13_), .Y(_abc_15497_new_n1425_));
INVX2 INVX2_38 ( .A(d_reg_15_), .Y(_abc_15497_new_n1447_));
INVX2 INVX2_39 ( .A(d_reg_16_), .Y(_abc_15497_new_n1462_));
INVX2 INVX2_4 ( .A(_auto_iopadmap_cc_368_execute_22625_64_), .Y(_abc_15497_new_n770_));
INVX2 INVX2_40 ( .A(d_reg_19_), .Y(_abc_15497_new_n1495_));
INVX2 INVX2_41 ( .A(d_reg_20_), .Y(_abc_15497_new_n1511_));
INVX2 INVX2_42 ( .A(_auto_iopadmap_cc_368_execute_22625_54_), .Y(_abc_15497_new_n1528_));
INVX2 INVX2_43 ( .A(d_reg_22_), .Y(_abc_15497_new_n1530_));
INVX2 INVX2_44 ( .A(_abc_15497_new_n1532_), .Y(_abc_15497_new_n1533_));
INVX2 INVX2_45 ( .A(d_reg_23_), .Y(_abc_15497_new_n1543_));
INVX2 INVX2_46 ( .A(_auto_iopadmap_cc_368_execute_22625_56_), .Y(_abc_15497_new_n1550_));
INVX2 INVX2_47 ( .A(d_reg_24_), .Y(_abc_15497_new_n1562_));
INVX2 INVX2_48 ( .A(d_reg_25_), .Y(_abc_15497_new_n1572_));
INVX2 INVX2_49 ( .A(_auto_iopadmap_cc_368_execute_22625_58_), .Y(_abc_15497_new_n1580_));
INVX2 INVX2_5 ( .A(_abc_15497_new_n859_), .Y(_abc_15497_new_n860_));
INVX2 INVX2_50 ( .A(d_reg_26_), .Y(_abc_15497_new_n1586_));
INVX2 INVX2_51 ( .A(_abc_15497_new_n1588_), .Y(_abc_15497_new_n1589_));
INVX2 INVX2_52 ( .A(d_reg_27_), .Y(_abc_15497_new_n1596_));
INVX2 INVX2_53 ( .A(b_reg_0_), .Y(_abc_15497_new_n1752_));
INVX2 INVX2_54 ( .A(_auto_iopadmap_cc_368_execute_22625_101_), .Y(_abc_15497_new_n1787_));
INVX2 INVX2_55 ( .A(_abc_15497_new_n1824_), .Y(_abc_15497_new_n1825_));
INVX2 INVX2_56 ( .A(_auto_iopadmap_cc_368_execute_22625_106_), .Y(_abc_15497_new_n1836_));
INVX2 INVX2_57 ( .A(b_reg_16_), .Y(_abc_15497_new_n1908_));
INVX2 INVX2_58 ( .A(_auto_iopadmap_cc_368_execute_22625_113_), .Y(_abc_15497_new_n1916_));
INVX2 INVX2_59 ( .A(b_reg_26_), .Y(_abc_15497_new_n2031_));
INVX2 INVX2_6 ( .A(c_reg_26_), .Y(_abc_15497_new_n866_));
INVX2 INVX2_60 ( .A(_auto_iopadmap_cc_368_execute_22625_131_), .Y(_abc_15497_new_n2112_));
INVX2 INVX2_61 ( .A(_auto_iopadmap_cc_368_execute_22625_133_), .Y(_abc_15497_new_n2129_));
INVX2 INVX2_62 ( .A(_auto_iopadmap_cc_368_execute_22625_134_), .Y(_abc_15497_new_n2141_));
INVX2 INVX2_63 ( .A(_auto_iopadmap_cc_368_execute_22625_140_), .Y(_abc_15497_new_n2203_));
INVX2 INVX2_64 ( .A(a_reg_12_), .Y(_abc_15497_new_n2214_));
INVX2 INVX2_65 ( .A(_auto_iopadmap_cc_368_execute_22625_142_), .Y(_abc_15497_new_n2228_));
INVX2 INVX2_66 ( .A(a_reg_14_), .Y(_abc_15497_new_n2230_));
INVX2 INVX2_67 ( .A(a_reg_16_), .Y(_abc_15497_new_n2258_));
INVX2 INVX2_68 ( .A(a_reg_24_), .Y(_abc_15497_new_n2360_));
INVX2 INVX2_69 ( .A(round_ctr_reg_6_), .Y(_abc_15497_new_n2735_));
INVX2 INVX2_7 ( .A(_auto_iopadmap_cc_368_execute_22625_94_), .Y(_abc_15497_new_n911_));
INVX2 INVX2_70 ( .A(round_ctr_reg_5_), .Y(_abc_15497_new_n2740_));
INVX2 INVX2_71 ( .A(d_reg_2_), .Y(_abc_15497_new_n2829_));
INVX2 INVX2_72 ( .A(d_reg_10_), .Y(_abc_15497_new_n3290_));
INVX2 INVX2_73 ( .A(d_reg_17_), .Y(_abc_15497_new_n3726_));
INVX2 INVX2_74 ( .A(round_ctr_reg_0_), .Y(_abc_15497_new_n4443_));
INVX2 INVX2_8 ( .A(c_reg_30_), .Y(_abc_15497_new_n912_));
INVX2 INVX2_9 ( .A(_auto_iopadmap_cc_368_execute_22625_12_), .Y(_abc_15497_new_n1057_));
INVX4 INVX4_1 ( .A(d_reg_8_), .Y(_abc_15497_new_n1364_));
INVX4 INVX4_2 ( .A(round_ctr_inc_bF_buf13), .Y(_abc_15497_new_n1646_));
INVX4 INVX4_3 ( .A(_abc_15497_new_n2738_), .Y(_abc_15497_new_n2739_));
INVX4 INVX4_4 ( .A(_abc_15497_new_n3678_), .Y(_abc_15497_new_n3679_));
INVX8 INVX8_1 ( .A(digest_update_bF_buf8), .Y(_abc_15497_new_n870_));
INVX8 INVX8_10 ( .A(w_mem_inst__abc_19396_new_n1627_), .Y(w_mem_inst__abc_19396_new_n1635_));
INVX8 INVX8_11 ( .A(round_ctr_rst_bF_buf6), .Y(w_mem_inst__abc_19396_new_n2420_));
INVX8 INVX8_12 ( .A(w_mem_inst__abc_19396_new_n2422__bF_buf32), .Y(w_mem_inst__abc_19396_new_n2582_));
INVX8 INVX8_2 ( .A(_auto_iopadmap_cc_368_execute_22788), .Y(_abc_15497_new_n871_));
INVX8 INVX8_3 ( .A(init), .Y(_abc_15497_new_n872_));
INVX8 INVX8_4 ( .A(_abc_15497_new_n1644_), .Y(round_ctr_rst));
INVX8 INVX8_5 ( .A(_abc_15497_new_n1648__bF_buf4), .Y(_abc_15497_new_n1663_));
INVX8 INVX8_6 ( .A(_abc_15497_new_n2742__bF_buf3), .Y(_abc_15497_new_n2743_));
INVX8 INVX8_7 ( .A(w_mem_inst__abc_19396_new_n1586__bF_buf4), .Y(w_mem_inst__abc_19396_new_n1587_));
INVX8 INVX8_8 ( .A(w_mem_inst__abc_19396_new_n1593_), .Y(w_mem_inst__abc_19396_new_n1594_));
INVX8 INVX8_9 ( .A(w_mem_inst__abc_19396_new_n1612_), .Y(w_mem_inst__abc_19396_new_n1617_));
MUX2X1 MUX2X1_1 ( .A(_abc_15497_new_n1304_), .B(_abc_15497_new_n1305_), .S(digest_update_bF_buf3), .Y(_0H3_reg_31_0__1_));
MUX2X1 MUX2X1_10 ( .A(\block[0] ), .B(w_mem_inst_w_mem_15__0_), .S(round_ctr_rst_bF_buf5), .Y(w_mem_inst__abc_19396_new_n2583_));
MUX2X1 MUX2X1_11 ( .A(w_mem_inst__abc_19396_new_n1590_), .B(w_mem_inst__abc_19396_new_n2583_), .S(w_mem_inst__abc_19396_new_n2582__bF_buf4), .Y(w_mem_inst__0w_mem_15__31_0__0_));
MUX2X1 MUX2X1_12 ( .A(\block[1] ), .B(w_mem_inst_w_mem_15__1_), .S(round_ctr_rst_bF_buf4), .Y(w_mem_inst__abc_19396_new_n2585_));
MUX2X1 MUX2X1_13 ( .A(w_mem_inst__abc_19396_new_n1645_), .B(w_mem_inst__abc_19396_new_n2585_), .S(w_mem_inst__abc_19396_new_n2582__bF_buf3), .Y(w_mem_inst__0w_mem_15__31_0__1_));
MUX2X1 MUX2X1_14 ( .A(\block[2] ), .B(w_mem_inst_w_mem_15__2_), .S(round_ctr_rst_bF_buf3), .Y(w_mem_inst__abc_19396_new_n2587_));
MUX2X1 MUX2X1_15 ( .A(w_mem_inst__abc_19396_new_n1670_), .B(w_mem_inst__abc_19396_new_n2587_), .S(w_mem_inst__abc_19396_new_n2582__bF_buf2), .Y(w_mem_inst__0w_mem_15__31_0__2_));
MUX2X1 MUX2X1_16 ( .A(\block[3] ), .B(w_mem_inst_w_mem_15__3_), .S(round_ctr_rst_bF_buf2), .Y(w_mem_inst__abc_19396_new_n2589_));
MUX2X1 MUX2X1_17 ( .A(w_mem_inst__abc_19396_new_n1695_), .B(w_mem_inst__abc_19396_new_n2589_), .S(w_mem_inst__abc_19396_new_n2582__bF_buf1), .Y(w_mem_inst__0w_mem_15__31_0__3_));
MUX2X1 MUX2X1_18 ( .A(\block[4] ), .B(w_mem_inst_w_mem_15__4_), .S(round_ctr_rst_bF_buf1), .Y(w_mem_inst__abc_19396_new_n2591_));
MUX2X1 MUX2X1_19 ( .A(w_mem_inst__abc_19396_new_n1720_), .B(w_mem_inst__abc_19396_new_n2591_), .S(w_mem_inst__abc_19396_new_n2582__bF_buf0), .Y(w_mem_inst__0w_mem_15__31_0__4_));
MUX2X1 MUX2X1_2 ( .A(_abc_15497_new_n1314_), .B(_abc_15497_new_n1315_), .S(digest_update_bF_buf2), .Y(_0H3_reg_31_0__2_));
MUX2X1 MUX2X1_20 ( .A(\block[5] ), .B(w_mem_inst_w_mem_15__5_), .S(round_ctr_rst_bF_buf0), .Y(w_mem_inst__abc_19396_new_n2593_));
MUX2X1 MUX2X1_21 ( .A(w_mem_inst__abc_19396_new_n1745_), .B(w_mem_inst__abc_19396_new_n2593_), .S(w_mem_inst__abc_19396_new_n2582__bF_buf4), .Y(w_mem_inst__0w_mem_15__31_0__5_));
MUX2X1 MUX2X1_22 ( .A(\block[6] ), .B(w_mem_inst_w_mem_15__6_), .S(round_ctr_rst_bF_buf8), .Y(w_mem_inst__abc_19396_new_n2595_));
MUX2X1 MUX2X1_23 ( .A(w_mem_inst__abc_19396_new_n1770_), .B(w_mem_inst__abc_19396_new_n2595_), .S(w_mem_inst__abc_19396_new_n2582__bF_buf3), .Y(w_mem_inst__0w_mem_15__31_0__6_));
MUX2X1 MUX2X1_24 ( .A(\block[7] ), .B(w_mem_inst_w_mem_15__7_), .S(round_ctr_rst_bF_buf7), .Y(w_mem_inst__abc_19396_new_n2597_));
MUX2X1 MUX2X1_25 ( .A(w_mem_inst__abc_19396_new_n1795_), .B(w_mem_inst__abc_19396_new_n2597_), .S(w_mem_inst__abc_19396_new_n2582__bF_buf2), .Y(w_mem_inst__0w_mem_15__31_0__7_));
MUX2X1 MUX2X1_26 ( .A(\block[8] ), .B(w_mem_inst_w_mem_15__8_), .S(round_ctr_rst_bF_buf6), .Y(w_mem_inst__abc_19396_new_n2599_));
MUX2X1 MUX2X1_27 ( .A(w_mem_inst__abc_19396_new_n1820_), .B(w_mem_inst__abc_19396_new_n2599_), .S(w_mem_inst__abc_19396_new_n2582__bF_buf1), .Y(w_mem_inst__0w_mem_15__31_0__8_));
MUX2X1 MUX2X1_28 ( .A(\block[9] ), .B(w_mem_inst_w_mem_15__9_), .S(round_ctr_rst_bF_buf5), .Y(w_mem_inst__abc_19396_new_n2601_));
MUX2X1 MUX2X1_29 ( .A(w_mem_inst__abc_19396_new_n1845_), .B(w_mem_inst__abc_19396_new_n2601_), .S(w_mem_inst__abc_19396_new_n2582__bF_buf0), .Y(w_mem_inst__0w_mem_15__31_0__9_));
MUX2X1 MUX2X1_3 ( .A(_abc_15497_new_n1329_), .B(_abc_15497_new_n1330_), .S(digest_update_bF_buf0), .Y(_0H3_reg_31_0__4_));
MUX2X1 MUX2X1_30 ( .A(\block[10] ), .B(w_mem_inst_w_mem_15__10_), .S(round_ctr_rst_bF_buf4), .Y(w_mem_inst__abc_19396_new_n2603_));
MUX2X1 MUX2X1_31 ( .A(w_mem_inst__abc_19396_new_n1870_), .B(w_mem_inst__abc_19396_new_n2603_), .S(w_mem_inst__abc_19396_new_n2582__bF_buf4), .Y(w_mem_inst__0w_mem_15__31_0__10_));
MUX2X1 MUX2X1_32 ( .A(\block[11] ), .B(w_mem_inst_w_mem_15__11_), .S(round_ctr_rst_bF_buf3), .Y(w_mem_inst__abc_19396_new_n2605_));
MUX2X1 MUX2X1_33 ( .A(w_mem_inst__abc_19396_new_n1895_), .B(w_mem_inst__abc_19396_new_n2605_), .S(w_mem_inst__abc_19396_new_n2582__bF_buf3), .Y(w_mem_inst__0w_mem_15__31_0__11_));
MUX2X1 MUX2X1_34 ( .A(\block[12] ), .B(w_mem_inst_w_mem_15__12_), .S(round_ctr_rst_bF_buf2), .Y(w_mem_inst__abc_19396_new_n2607_));
MUX2X1 MUX2X1_35 ( .A(w_mem_inst__abc_19396_new_n1920_), .B(w_mem_inst__abc_19396_new_n2607_), .S(w_mem_inst__abc_19396_new_n2582__bF_buf2), .Y(w_mem_inst__0w_mem_15__31_0__12_));
MUX2X1 MUX2X1_36 ( .A(\block[13] ), .B(w_mem_inst_w_mem_15__13_), .S(round_ctr_rst_bF_buf1), .Y(w_mem_inst__abc_19396_new_n2609_));
MUX2X1 MUX2X1_37 ( .A(w_mem_inst__abc_19396_new_n1945_), .B(w_mem_inst__abc_19396_new_n2609_), .S(w_mem_inst__abc_19396_new_n2582__bF_buf1), .Y(w_mem_inst__0w_mem_15__31_0__13_));
MUX2X1 MUX2X1_38 ( .A(\block[14] ), .B(w_mem_inst_w_mem_15__14_), .S(round_ctr_rst_bF_buf0), .Y(w_mem_inst__abc_19396_new_n2611_));
MUX2X1 MUX2X1_39 ( .A(w_mem_inst__abc_19396_new_n1970_), .B(w_mem_inst__abc_19396_new_n2611_), .S(w_mem_inst__abc_19396_new_n2582__bF_buf0), .Y(w_mem_inst__0w_mem_15__31_0__14_));
MUX2X1 MUX2X1_4 ( .A(c_reg_31_), .B(d_reg_31_), .S(b_reg_31_), .Y(_abc_15497_new_n4416_));
MUX2X1 MUX2X1_40 ( .A(\block[15] ), .B(w_mem_inst_w_mem_15__15_), .S(round_ctr_rst_bF_buf8), .Y(w_mem_inst__abc_19396_new_n2613_));
MUX2X1 MUX2X1_41 ( .A(w_mem_inst__abc_19396_new_n1995_), .B(w_mem_inst__abc_19396_new_n2613_), .S(w_mem_inst__abc_19396_new_n2582__bF_buf4), .Y(w_mem_inst__0w_mem_15__31_0__15_));
MUX2X1 MUX2X1_42 ( .A(\block[16] ), .B(w_mem_inst_w_mem_15__16_), .S(round_ctr_rst_bF_buf7), .Y(w_mem_inst__abc_19396_new_n2615_));
MUX2X1 MUX2X1_43 ( .A(w_mem_inst__abc_19396_new_n2020_), .B(w_mem_inst__abc_19396_new_n2615_), .S(w_mem_inst__abc_19396_new_n2582__bF_buf3), .Y(w_mem_inst__0w_mem_15__31_0__16_));
MUX2X1 MUX2X1_44 ( .A(\block[17] ), .B(w_mem_inst_w_mem_15__17_), .S(round_ctr_rst_bF_buf6), .Y(w_mem_inst__abc_19396_new_n2617_));
MUX2X1 MUX2X1_45 ( .A(w_mem_inst__abc_19396_new_n2045_), .B(w_mem_inst__abc_19396_new_n2617_), .S(w_mem_inst__abc_19396_new_n2582__bF_buf2), .Y(w_mem_inst__0w_mem_15__31_0__17_));
MUX2X1 MUX2X1_46 ( .A(\block[18] ), .B(w_mem_inst_w_mem_15__18_), .S(round_ctr_rst_bF_buf5), .Y(w_mem_inst__abc_19396_new_n2619_));
MUX2X1 MUX2X1_47 ( .A(w_mem_inst__abc_19396_new_n2070_), .B(w_mem_inst__abc_19396_new_n2619_), .S(w_mem_inst__abc_19396_new_n2582__bF_buf1), .Y(w_mem_inst__0w_mem_15__31_0__18_));
MUX2X1 MUX2X1_48 ( .A(\block[19] ), .B(w_mem_inst_w_mem_15__19_), .S(round_ctr_rst_bF_buf4), .Y(w_mem_inst__abc_19396_new_n2621_));
MUX2X1 MUX2X1_49 ( .A(w_mem_inst__abc_19396_new_n2095_), .B(w_mem_inst__abc_19396_new_n2621_), .S(w_mem_inst__abc_19396_new_n2582__bF_buf0), .Y(w_mem_inst__0w_mem_15__31_0__19_));
MUX2X1 MUX2X1_5 ( .A(round_ctr_reg_4_), .B(_abc_15497_new_n4466_), .S(_abc_15497_new_n4464_), .Y(_0round_ctr_reg_6_0__4_));
MUX2X1 MUX2X1_50 ( .A(\block[20] ), .B(w_mem_inst_w_mem_15__20_), .S(round_ctr_rst_bF_buf3), .Y(w_mem_inst__abc_19396_new_n2623_));
MUX2X1 MUX2X1_51 ( .A(w_mem_inst__abc_19396_new_n2120_), .B(w_mem_inst__abc_19396_new_n2623_), .S(w_mem_inst__abc_19396_new_n2582__bF_buf4), .Y(w_mem_inst__0w_mem_15__31_0__20_));
MUX2X1 MUX2X1_52 ( .A(\block[21] ), .B(w_mem_inst_w_mem_15__21_), .S(round_ctr_rst_bF_buf2), .Y(w_mem_inst__abc_19396_new_n2625_));
MUX2X1 MUX2X1_53 ( .A(w_mem_inst__abc_19396_new_n2145_), .B(w_mem_inst__abc_19396_new_n2625_), .S(w_mem_inst__abc_19396_new_n2582__bF_buf3), .Y(w_mem_inst__0w_mem_15__31_0__21_));
MUX2X1 MUX2X1_54 ( .A(\block[22] ), .B(w_mem_inst_w_mem_15__22_), .S(round_ctr_rst_bF_buf1), .Y(w_mem_inst__abc_19396_new_n2627_));
MUX2X1 MUX2X1_55 ( .A(w_mem_inst__abc_19396_new_n2170_), .B(w_mem_inst__abc_19396_new_n2627_), .S(w_mem_inst__abc_19396_new_n2582__bF_buf2), .Y(w_mem_inst__0w_mem_15__31_0__22_));
MUX2X1 MUX2X1_56 ( .A(\block[23] ), .B(w_mem_inst_w_mem_15__23_), .S(round_ctr_rst_bF_buf0), .Y(w_mem_inst__abc_19396_new_n2629_));
MUX2X1 MUX2X1_57 ( .A(w_mem_inst__abc_19396_new_n2195_), .B(w_mem_inst__abc_19396_new_n2629_), .S(w_mem_inst__abc_19396_new_n2582__bF_buf1), .Y(w_mem_inst__0w_mem_15__31_0__23_));
MUX2X1 MUX2X1_58 ( .A(\block[24] ), .B(w_mem_inst_w_mem_15__24_), .S(round_ctr_rst_bF_buf8), .Y(w_mem_inst__abc_19396_new_n2631_));
MUX2X1 MUX2X1_59 ( .A(w_mem_inst__abc_19396_new_n2220_), .B(w_mem_inst__abc_19396_new_n2631_), .S(w_mem_inst__abc_19396_new_n2582__bF_buf0), .Y(w_mem_inst__0w_mem_15__31_0__24_));
MUX2X1 MUX2X1_6 ( .A(round_ctr_reg_6_), .B(_abc_15497_new_n4472_), .S(_abc_15497_new_n4470_), .Y(_0round_ctr_reg_6_0__6_));
MUX2X1 MUX2X1_60 ( .A(\block[25] ), .B(w_mem_inst_w_mem_15__25_), .S(round_ctr_rst_bF_buf7), .Y(w_mem_inst__abc_19396_new_n2633_));
MUX2X1 MUX2X1_61 ( .A(w_mem_inst__abc_19396_new_n2245_), .B(w_mem_inst__abc_19396_new_n2633_), .S(w_mem_inst__abc_19396_new_n2582__bF_buf4), .Y(w_mem_inst__0w_mem_15__31_0__25_));
MUX2X1 MUX2X1_62 ( .A(\block[26] ), .B(w_mem_inst_w_mem_15__26_), .S(round_ctr_rst_bF_buf6), .Y(w_mem_inst__abc_19396_new_n2635_));
MUX2X1 MUX2X1_63 ( .A(w_mem_inst__abc_19396_new_n2270_), .B(w_mem_inst__abc_19396_new_n2635_), .S(w_mem_inst__abc_19396_new_n2582__bF_buf3), .Y(w_mem_inst__0w_mem_15__31_0__26_));
MUX2X1 MUX2X1_64 ( .A(\block[27] ), .B(w_mem_inst_w_mem_15__27_), .S(round_ctr_rst_bF_buf5), .Y(w_mem_inst__abc_19396_new_n2637_));
MUX2X1 MUX2X1_65 ( .A(w_mem_inst__abc_19396_new_n2295_), .B(w_mem_inst__abc_19396_new_n2637_), .S(w_mem_inst__abc_19396_new_n2582__bF_buf2), .Y(w_mem_inst__0w_mem_15__31_0__27_));
MUX2X1 MUX2X1_66 ( .A(\block[28] ), .B(w_mem_inst_w_mem_15__28_), .S(round_ctr_rst_bF_buf4), .Y(w_mem_inst__abc_19396_new_n2639_));
MUX2X1 MUX2X1_67 ( .A(w_mem_inst__abc_19396_new_n2320_), .B(w_mem_inst__abc_19396_new_n2639_), .S(w_mem_inst__abc_19396_new_n2582__bF_buf1), .Y(w_mem_inst__0w_mem_15__31_0__28_));
MUX2X1 MUX2X1_68 ( .A(\block[29] ), .B(w_mem_inst_w_mem_15__29_), .S(round_ctr_rst_bF_buf3), .Y(w_mem_inst__abc_19396_new_n2641_));
MUX2X1 MUX2X1_69 ( .A(w_mem_inst__abc_19396_new_n2345_), .B(w_mem_inst__abc_19396_new_n2641_), .S(w_mem_inst__abc_19396_new_n2582__bF_buf0), .Y(w_mem_inst__0w_mem_15__31_0__29_));
MUX2X1 MUX2X1_7 ( .A(_abc_15497_new_n4480_), .B(_abc_15497_new_n4479_), .S(digest_update_bF_buf2), .Y(_0H2_reg_31_0__1_));
MUX2X1 MUX2X1_70 ( .A(\block[30] ), .B(w_mem_inst_w_mem_15__30_), .S(round_ctr_rst_bF_buf2), .Y(w_mem_inst__abc_19396_new_n2643_));
MUX2X1 MUX2X1_71 ( .A(w_mem_inst__abc_19396_new_n2370_), .B(w_mem_inst__abc_19396_new_n2643_), .S(w_mem_inst__abc_19396_new_n2582__bF_buf4), .Y(w_mem_inst__0w_mem_15__31_0__30_));
MUX2X1 MUX2X1_72 ( .A(\block[31] ), .B(w_mem_inst_w_mem_15__31_), .S(round_ctr_rst_bF_buf1), .Y(w_mem_inst__abc_19396_new_n2645_));
MUX2X1 MUX2X1_73 ( .A(w_mem_inst__abc_19396_new_n2395_), .B(w_mem_inst__abc_19396_new_n2645_), .S(w_mem_inst__abc_19396_new_n2582__bF_buf3), .Y(w_mem_inst__0w_mem_15__31_0__31_));
MUX2X1 MUX2X1_74 ( .A(w_mem_inst__abc_19396_new_n4796_), .B(w_mem_inst_w_ctr_reg_2_), .S(w_mem_inst__abc_19396_new_n4797_), .Y(w_mem_inst__0w_ctr_reg_6_0__2_));
MUX2X1 MUX2X1_8 ( .A(_abc_15497_new_n4483_), .B(_abc_15497_new_n4482_), .S(digest_update_bF_buf1), .Y(_0H2_reg_31_0__2_));
MUX2X1 MUX2X1_9 ( .A(_abc_15497_new_n4491_), .B(_abc_15497_new_n4490_), .S(digest_update_bF_buf0), .Y(_0H2_reg_31_0__4_));
NAND2X1 NAND2X1_1 ( .A(_abc_15497_new_n701_), .B(_abc_15497_new_n706_), .Y(_abc_15497_new_n707_));
NAND2X1 NAND2X1_10 ( .A(c_reg_23_), .B(_auto_iopadmap_cc_368_execute_22625_87_), .Y(_abc_15497_new_n794_));
NAND2X1 NAND2X1_100 ( .A(_abc_15497_new_n1766_), .B(_abc_15497_new_n1765_), .Y(_abc_15497_new_n1767_));
NAND2X1 NAND2X1_101 ( .A(_abc_15497_new_n1780_), .B(_abc_15497_new_n1782_), .Y(_abc_15497_new_n1784_));
NAND2X1 NAND2X1_102 ( .A(digest_update_bF_buf7), .B(_abc_15497_new_n1784_), .Y(_abc_15497_new_n1785_));
NAND2X1 NAND2X1_103 ( .A(_abc_15497_new_n1796_), .B(_abc_15497_new_n1794_), .Y(_abc_15497_new_n1797_));
NAND2X1 NAND2X1_104 ( .A(_auto_iopadmap_cc_368_execute_22625_103_), .B(b_reg_7_), .Y(_abc_15497_new_n1809_));
NAND2X1 NAND2X1_105 ( .A(_abc_15497_new_n1811_), .B(_abc_15497_new_n1807_), .Y(_abc_15497_new_n1812_));
NAND2X1 NAND2X1_106 ( .A(_abc_15497_new_n1816_), .B(_abc_15497_new_n1815_), .Y(_0H1_reg_31_0__7_));
NAND2X1 NAND2X1_107 ( .A(_abc_15497_new_n1809_), .B(_abc_15497_new_n1807_), .Y(_abc_15497_new_n1823_));
NAND2X1 NAND2X1_108 ( .A(_abc_15497_new_n1832_), .B(_abc_15497_new_n1822_), .Y(_abc_15497_new_n1837_));
NAND2X1 NAND2X1_109 ( .A(_abc_15497_new_n1843_), .B(_abc_15497_new_n1839_), .Y(_abc_15497_new_n1845_));
NAND2X1 NAND2X1_11 ( .A(_abc_15497_new_n822_), .B(_abc_15497_new_n827_), .Y(_abc_15497_new_n828_));
NAND2X1 NAND2X1_110 ( .A(digest_update_bF_buf5), .B(_abc_15497_new_n1845_), .Y(_abc_15497_new_n1846_));
NAND2X1 NAND2X1_111 ( .A(_auto_iopadmap_cc_368_execute_22625_107_), .B(b_reg_11_), .Y(_abc_15497_new_n1850_));
NAND2X1 NAND2X1_112 ( .A(_abc_15497_new_n1852_), .B(_abc_15497_new_n1843_), .Y(_abc_15497_new_n1862_));
NAND2X1 NAND2X1_113 ( .A(_abc_15497_new_n1870_), .B(_abc_15497_new_n1860_), .Y(_abc_15497_new_n1884_));
NAND2X1 NAND2X1_114 ( .A(_auto_iopadmap_cc_368_execute_22625_111_), .B(b_reg_15_), .Y(_abc_15497_new_n1893_));
NAND2X1 NAND2X1_115 ( .A(_abc_15497_new_n1895_), .B(_abc_15497_new_n1878_), .Y(_abc_15497_new_n1900_));
NAND2X1 NAND2X1_116 ( .A(_abc_15497_new_n1864_), .B(_abc_15497_new_n1902_), .Y(_abc_15497_new_n1904_));
NAND2X1 NAND2X1_117 ( .A(_abc_15497_new_n1910_), .B(_abc_15497_new_n1905_), .Y(_abc_15497_new_n1912_));
NAND2X1 NAND2X1_118 ( .A(digest_update_bF_buf3), .B(_abc_15497_new_n1912_), .Y(_abc_15497_new_n1913_));
NAND2X1 NAND2X1_119 ( .A(_abc_15497_new_n1909_), .B(_abc_15497_new_n1920_), .Y(_abc_15497_new_n1926_));
NAND2X1 NAND2X1_12 ( .A(_abc_15497_new_n868_), .B(_abc_15497_new_n864_), .Y(_abc_15497_new_n874_));
NAND2X1 NAND2X1_120 ( .A(_auto_iopadmap_cc_368_execute_22625_114_), .B(b_reg_18_), .Y(_abc_15497_new_n1930_));
NAND2X1 NAND2X1_121 ( .A(digest_update_bF_buf2), .B(_abc_15497_new_n1934_), .Y(_abc_15497_new_n1935_));
NAND2X1 NAND2X1_122 ( .A(_abc_15497_new_n1930_), .B(_abc_15497_new_n1934_), .Y(_abc_15497_new_n1938_));
NAND2X1 NAND2X1_123 ( .A(_auto_iopadmap_cc_368_execute_22625_115_), .B(b_reg_19_), .Y(_abc_15497_new_n1940_));
NAND2X1 NAND2X1_124 ( .A(_abc_15497_new_n1947_), .B(_abc_15497_new_n1946_), .Y(_0H1_reg_31_0__19_));
NAND2X1 NAND2X1_125 ( .A(_abc_15497_new_n1932_), .B(_abc_15497_new_n1942_), .Y(_abc_15497_new_n1951_));
NAND2X1 NAND2X1_126 ( .A(_abc_15497_new_n1910_), .B(_abc_15497_new_n1920_), .Y(_abc_15497_new_n1954_));
NAND2X1 NAND2X1_127 ( .A(_auto_iopadmap_cc_368_execute_22625_118_), .B(b_reg_22_), .Y(_abc_15497_new_n1980_));
NAND2X1 NAND2X1_128 ( .A(_auto_iopadmap_cc_368_execute_22625_119_), .B(b_reg_23_), .Y(_abc_15497_new_n1988_));
NAND2X1 NAND2X1_129 ( .A(_abc_15497_new_n1982_), .B(_abc_15497_new_n1990_), .Y(_abc_15497_new_n1994_));
NAND2X1 NAND2X1_13 ( .A(digest_update_bF_buf7), .B(_abc_15497_new_n874_), .Y(_abc_15497_new_n875_));
NAND2X1 NAND2X1_130 ( .A(_abc_15497_new_n1953_), .B(_abc_15497_new_n1995_), .Y(_abc_15497_new_n1996_));
NAND2X1 NAND2X1_131 ( .A(_auto_iopadmap_cc_368_execute_22625_121_), .B(b_reg_25_), .Y(_abc_15497_new_n2017_));
NAND2X1 NAND2X1_132 ( .A(_abc_15497_new_n2033_), .B(_abc_15497_new_n2028_), .Y(_abc_15497_new_n2035_));
NAND2X1 NAND2X1_133 ( .A(digest_update_bF_buf7), .B(_abc_15497_new_n2035_), .Y(_abc_15497_new_n2036_));
NAND2X1 NAND2X1_134 ( .A(_auto_iopadmap_cc_368_execute_22625_123_), .B(b_reg_27_), .Y(_abc_15497_new_n2041_));
NAND2X1 NAND2X1_135 ( .A(_abc_15497_new_n2048_), .B(_abc_15497_new_n2024_), .Y(_abc_15497_new_n2049_));
NAND2X1 NAND2X1_136 ( .A(_abc_15497_new_n2047_), .B(_abc_15497_new_n2054_), .Y(_abc_15497_new_n2055_));
NAND2X1 NAND2X1_137 ( .A(_auto_iopadmap_cc_368_execute_22625_124_), .B(b_reg_28_), .Y(_abc_15497_new_n2056_));
NAND2X1 NAND2X1_138 ( .A(_abc_15497_new_n2056_), .B(_abc_15497_new_n2055_), .Y(_abc_15497_new_n2059_));
NAND2X1 NAND2X1_139 ( .A(_auto_iopadmap_cc_368_execute_22625_125_), .B(b_reg_29_), .Y(_abc_15497_new_n2065_));
NAND2X1 NAND2X1_14 ( .A(_auto_iopadmap_cc_368_execute_22625_91_), .B(c_reg_27_), .Y(_abc_15497_new_n879_));
NAND2X1 NAND2X1_140 ( .A(_abc_15497_new_n2073_), .B(_abc_15497_new_n2076_), .Y(_abc_15497_new_n2077_));
NAND2X1 NAND2X1_141 ( .A(_abc_15497_new_n2077_), .B(_abc_15497_new_n2078_), .Y(_abc_15497_new_n2079_));
NAND2X1 NAND2X1_142 ( .A(_auto_iopadmap_cc_368_execute_22625_126_), .B(b_reg_30_), .Y(_abc_15497_new_n2082_));
NAND2X1 NAND2X1_143 ( .A(_abc_15497_new_n2086_), .B(_abc_15497_new_n2085_), .Y(_abc_15497_new_n2087_));
NAND2X1 NAND2X1_144 ( .A(_abc_15497_new_n2089_), .B(_abc_15497_new_n2088_), .Y(_0H1_reg_31_0__31_));
NAND2X1 NAND2X1_145 ( .A(_abc_15497_new_n2098_), .B(_abc_15497_new_n2099_), .Y(_abc_15497_new_n2105_));
NAND2X1 NAND2X1_146 ( .A(_abc_15497_new_n2107_), .B(_abc_15497_new_n2106_), .Y(_abc_15497_new_n2108_));
NAND2X1 NAND2X1_147 ( .A(_abc_15497_new_n2112_), .B(_abc_15497_new_n2115_), .Y(_abc_15497_new_n2116_));
NAND2X1 NAND2X1_148 ( .A(_abc_15497_new_n2116_), .B(_abc_15497_new_n2118_), .Y(_abc_15497_new_n2119_));
NAND2X1 NAND2X1_149 ( .A(_abc_15497_new_n2123_), .B(_abc_15497_new_n2124_), .Y(_abc_15497_new_n2126_));
NAND2X1 NAND2X1_15 ( .A(_abc_15497_new_n886_), .B(_abc_15497_new_n861_), .Y(_abc_15497_new_n887_));
NAND2X1 NAND2X1_150 ( .A(digest_update_bF_buf2), .B(_abc_15497_new_n2126_), .Y(_abc_15497_new_n2127_));
NAND2X1 NAND2X1_151 ( .A(_abc_15497_new_n2138_), .B(_abc_15497_new_n2136_), .Y(_abc_15497_new_n2139_));
NAND2X1 NAND2X1_152 ( .A(_abc_15497_new_n2146_), .B(_abc_15497_new_n2142_), .Y(_abc_15497_new_n2148_));
NAND2X1 NAND2X1_153 ( .A(digest_update_bF_buf1), .B(_abc_15497_new_n2148_), .Y(_abc_15497_new_n2149_));
NAND2X1 NAND2X1_154 ( .A(_abc_15497_new_n2145_), .B(_abc_15497_new_n2152_), .Y(_abc_15497_new_n2160_));
NAND2X1 NAND2X1_155 ( .A(_abc_15497_new_n2176_), .B(_abc_15497_new_n2168_), .Y(_abc_15497_new_n2191_));
NAND2X1 NAND2X1_156 ( .A(_abc_15497_new_n2200_), .B(_abc_15497_new_n2184_), .Y(_abc_15497_new_n2204_));
NAND2X1 NAND2X1_157 ( .A(_abc_15497_new_n2216_), .B(_abc_15497_new_n2212_), .Y(_abc_15497_new_n2218_));
NAND2X1 NAND2X1_158 ( .A(digest_update_bF_buf7), .B(_abc_15497_new_n2218_), .Y(_abc_15497_new_n2219_));
NAND2X1 NAND2X1_159 ( .A(_abc_15497_new_n2224_), .B(_abc_15497_new_n2216_), .Y(_abc_15497_new_n2235_));
NAND2X1 NAND2X1_16 ( .A(_auto_iopadmap_cc_368_execute_22625_92_), .B(c_reg_28_), .Y(_abc_15497_new_n894_));
NAND2X1 NAND2X1_160 ( .A(_abc_15497_new_n2232_), .B(_abc_15497_new_n2236_), .Y(_abc_15497_new_n2238_));
NAND2X1 NAND2X1_161 ( .A(digest_update_bF_buf6), .B(_abc_15497_new_n2238_), .Y(_abc_15497_new_n2239_));
NAND2X1 NAND2X1_162 ( .A(_abc_15497_new_n2232_), .B(_abc_15497_new_n2246_), .Y(_abc_15497_new_n2250_));
NAND2X1 NAND2X1_163 ( .A(_abc_15497_new_n2205_), .B(_abc_15497_new_n2252_), .Y(_abc_15497_new_n2254_));
NAND2X1 NAND2X1_164 ( .A(_abc_15497_new_n2286_), .B(_abc_15497_new_n2298_), .Y(_abc_15497_new_n2304_));
NAND2X1 NAND2X1_165 ( .A(_abc_15497_new_n2328_), .B(_abc_15497_new_n2325_), .Y(_abc_15497_new_n2329_));
NAND2X1 NAND2X1_166 ( .A(_abc_15497_new_n2387_), .B(_abc_15497_new_n2382_), .Y(_abc_15497_new_n2389_));
NAND2X1 NAND2X1_167 ( .A(digest_update_bF_buf8), .B(_abc_15497_new_n2389_), .Y(_abc_15497_new_n2390_));
NAND2X1 NAND2X1_168 ( .A(_abc_15497_new_n2402_), .B(_abc_15497_new_n2379_), .Y(_abc_15497_new_n2403_));
NAND2X1 NAND2X1_169 ( .A(_abc_15497_new_n2409_), .B(_abc_15497_new_n2408_), .Y(_abc_15497_new_n2411_));
NAND2X1 NAND2X1_17 ( .A(_abc_15497_new_n899_), .B(_abc_15497_new_n898_), .Y(_0H2_reg_31_0__28_));
NAND2X1 NAND2X1_170 ( .A(digest_update_bF_buf7), .B(_abc_15497_new_n2411_), .Y(_abc_15497_new_n2412_));
NAND2X1 NAND2X1_171 ( .A(_abc_15497_new_n2425_), .B(_abc_15497_new_n2426_), .Y(_abc_15497_new_n2427_));
NAND2X1 NAND2X1_172 ( .A(_auto_iopadmap_cc_368_execute_22625_158_), .B(a_reg_30_), .Y(_abc_15497_new_n2428_));
NAND2X1 NAND2X1_173 ( .A(_abc_15497_new_n2428_), .B(_abc_15497_new_n2427_), .Y(_abc_15497_new_n2429_));
NAND2X1 NAND2X1_174 ( .A(d_reg_31_), .B(_abc_15497_new_n1663__bF_buf0), .Y(_abc_15497_new_n2636_));
NAND2X1 NAND2X1_175 ( .A(c_reg_31_), .B(round_ctr_inc_bF_buf12), .Y(_abc_15497_new_n2637_));
NAND2X1 NAND2X1_176 ( .A(round_ctr_reg_5_), .B(round_ctr_reg_4_), .Y(_abc_15497_new_n2736_));
NAND2X1 NAND2X1_177 ( .A(round_ctr_reg_5_), .B(round_ctr_reg_3_), .Y(_abc_15497_new_n2737_));
NAND2X1 NAND2X1_178 ( .A(_abc_15497_new_n1299_), .B(_abc_15497_new_n2746_), .Y(_abc_15497_new_n2747_));
NAND2X1 NAND2X1_179 ( .A(b_reg_0_), .B(c_reg_0_), .Y(_abc_15497_new_n2748_));
NAND2X1 NAND2X1_18 ( .A(_auto_iopadmap_cc_368_execute_22625_94_), .B(_abc_15497_new_n912_), .Y(_abc_15497_new_n913_));
NAND2X1 NAND2X1_180 ( .A(_abc_15497_new_n2735_), .B(_abc_15497_new_n2737_), .Y(_abc_15497_new_n2752_));
NAND2X1 NAND2X1_181 ( .A(round_ctr_reg_4_), .B(round_ctr_reg_2_), .Y(_abc_15497_new_n2753_));
NAND2X1 NAND2X1_182 ( .A(_abc_15497_new_n2735_), .B(_abc_15497_new_n2753_), .Y(_abc_15497_new_n2754_));
NAND2X1 NAND2X1_183 ( .A(_abc_15497_new_n2752_), .B(_abc_15497_new_n2754_), .Y(_abc_15497_new_n2755_));
NAND2X1 NAND2X1_184 ( .A(e_reg_0_), .B(a_reg_27_), .Y(_abc_15497_new_n2764_));
NAND2X1 NAND2X1_185 ( .A(_abc_15497_new_n2745_), .B(_abc_15497_new_n2743__bF_buf3), .Y(_abc_15497_new_n2769_));
NAND2X1 NAND2X1_186 ( .A(_abc_15497_new_n2760_), .B(_abc_15497_new_n2757_), .Y(_abc_15497_new_n2770_));
NAND2X1 NAND2X1_187 ( .A(b_reg_1_), .B(c_reg_1_), .Y(_abc_15497_new_n2783_));
NAND2X1 NAND2X1_188 ( .A(_abc_15497_new_n2789_), .B(_abc_15497_new_n2787_), .Y(_abc_15497_new_n2790_));
NAND2X1 NAND2X1_189 ( .A(e_reg_1_), .B(a_reg_28_), .Y(_abc_15497_new_n2794_));
NAND2X1 NAND2X1_19 ( .A(c_reg_30_), .B(_abc_15497_new_n911_), .Y(_abc_15497_new_n914_));
NAND2X1 NAND2X1_190 ( .A(_abc_15497_new_n2799_), .B(_abc_15497_new_n2803_), .Y(_abc_15497_new_n2804_));
NAND2X1 NAND2X1_191 ( .A(_abc_15497_new_n2804_), .B(_abc_15497_new_n2790_), .Y(_abc_15497_new_n2805_));
NAND2X1 NAND2X1_192 ( .A(_abc_15497_new_n2807_), .B(_abc_15497_new_n2806_), .Y(_abc_15497_new_n2808_));
NAND2X1 NAND2X1_193 ( .A(_abc_15497_new_n2790_), .B(_abc_15497_new_n2807_), .Y(_abc_15497_new_n2810_));
NAND2X1 NAND2X1_194 ( .A(_abc_15497_new_n2804_), .B(_abc_15497_new_n2806_), .Y(_abc_15497_new_n2811_));
NAND2X1 NAND2X1_195 ( .A(_abc_15497_new_n2816_), .B(_abc_15497_new_n2813_), .Y(_abc_15497_new_n2817_));
NAND2X1 NAND2X1_196 ( .A(round_ctr_inc_bF_buf5), .B(_abc_15497_new_n2821_), .Y(_abc_15497_new_n2822_));
NAND2X1 NAND2X1_197 ( .A(b_reg_2_), .B(c_reg_2_), .Y(_abc_15497_new_n2831_));
NAND2X1 NAND2X1_198 ( .A(_abc_15497_new_n2837_), .B(_abc_15497_new_n2835_), .Y(_abc_15497_new_n2838_));
NAND2X1 NAND2X1_199 ( .A(e_reg_2_), .B(a_reg_29_), .Y(_abc_15497_new_n2842_));
NAND2X1 NAND2X1_2 ( .A(_abc_15497_new_n731_), .B(_abc_15497_new_n735_), .Y(_abc_15497_new_n736_));
NAND2X1 NAND2X1_20 ( .A(_abc_15497_new_n918_), .B(_abc_15497_new_n892_), .Y(_abc_15497_new_n919_));
NAND2X1 NAND2X1_200 ( .A(_abc_15497_new_n2844_), .B(_abc_15497_new_n2846_), .Y(_abc_15497_new_n2849_));
NAND2X1 NAND2X1_201 ( .A(_abc_15497_new_n2848_), .B(_abc_15497_new_n2849_), .Y(_abc_15497_new_n2850_));
NAND2X1 NAND2X1_202 ( .A(_abc_15497_new_n2838_), .B(_abc_15497_new_n2851_), .Y(_abc_15497_new_n2852_));
NAND2X1 NAND2X1_203 ( .A(_abc_15497_new_n2847_), .B(_abc_15497_new_n2850_), .Y(_abc_15497_new_n2854_));
NAND2X1 NAND2X1_204 ( .A(_abc_15497_new_n2854_), .B(_abc_15497_new_n2853_), .Y(_abc_15497_new_n2855_));
NAND2X1 NAND2X1_205 ( .A(_abc_15497_new_n2838_), .B(_abc_15497_new_n2854_), .Y(_abc_15497_new_n2859_));
NAND2X1 NAND2X1_206 ( .A(_abc_15497_new_n2853_), .B(_abc_15497_new_n2851_), .Y(_abc_15497_new_n2860_));
NAND2X1 NAND2X1_207 ( .A(_abc_15497_new_n2739_), .B(_abc_15497_new_n2773_), .Y(_abc_15497_new_n2874_));
NAND2X1 NAND2X1_208 ( .A(_abc_15497_new_n2878_), .B(_abc_15497_new_n2873_), .Y(_abc_15497_new_n2879_));
NAND2X1 NAND2X1_209 ( .A(b_reg_3_), .B(c_reg_3_), .Y(_abc_15497_new_n2890_));
NAND2X1 NAND2X1_21 ( .A(_abc_15497_new_n913_), .B(_abc_15497_new_n914_), .Y(_abc_15497_new_n921_));
NAND2X1 NAND2X1_210 ( .A(_abc_15497_new_n2890_), .B(_abc_15497_new_n2891_), .Y(_abc_15497_new_n2893_));
NAND2X1 NAND2X1_211 ( .A(_abc_15497_new_n2896_), .B(_abc_15497_new_n2894_), .Y(_abc_15497_new_n2897_));
NAND2X1 NAND2X1_212 ( .A(_abc_15497_new_n960_), .B(_abc_15497_new_n2426_), .Y(_abc_15497_new_n2899_));
NAND2X1 NAND2X1_213 ( .A(e_reg_3_), .B(a_reg_30_), .Y(_abc_15497_new_n2900_));
NAND2X1 NAND2X1_214 ( .A(_abc_15497_new_n2900_), .B(_abc_15497_new_n2899_), .Y(_abc_15497_new_n2904_));
NAND2X1 NAND2X1_215 ( .A(_abc_15497_new_n2909_), .B(_abc_15497_new_n2906_), .Y(_abc_15497_new_n2910_));
NAND2X1 NAND2X1_216 ( .A(_abc_15497_new_n2897_), .B(_abc_15497_new_n2910_), .Y(_abc_15497_new_n2911_));
NAND2X1 NAND2X1_217 ( .A(_abc_15497_new_n2914_), .B(_abc_15497_new_n2913_), .Y(_abc_15497_new_n2915_));
NAND2X1 NAND2X1_218 ( .A(_abc_15497_new_n2915_), .B(_abc_15497_new_n2912_), .Y(_abc_15497_new_n2916_));
NAND2X1 NAND2X1_219 ( .A(_abc_15497_new_n2897_), .B(_abc_15497_new_n2915_), .Y(_abc_15497_new_n2919_));
NAND2X1 NAND2X1_22 ( .A(_abc_15497_new_n932_), .B(_abc_15497_new_n930_), .Y(_abc_15497_new_n933_));
NAND2X1 NAND2X1_220 ( .A(_abc_15497_new_n2910_), .B(_abc_15497_new_n2912_), .Y(_abc_15497_new_n2920_));
NAND2X1 NAND2X1_221 ( .A(_abc_15497_new_n2742__bF_buf2), .B(_abc_15497_new_n2924__bF_buf4), .Y(_abc_15497_new_n2925_));
NAND2X1 NAND2X1_222 ( .A(_abc_15497_new_n2934_), .B(_abc_15497_new_n2929_), .Y(_abc_15497_new_n2935_));
NAND2X1 NAND2X1_223 ( .A(_abc_15497_new_n1333_), .B(_abc_15497_new_n2946_), .Y(_abc_15497_new_n2947_));
NAND2X1 NAND2X1_224 ( .A(b_reg_4_), .B(c_reg_4_), .Y(_abc_15497_new_n2948_));
NAND2X1 NAND2X1_225 ( .A(_abc_15497_new_n2947_), .B(_abc_15497_new_n2950_), .Y(_abc_15497_new_n2951_));
NAND2X1 NAND2X1_226 ( .A(e_reg_4_), .B(a_reg_31_), .Y(_abc_15497_new_n2959_));
NAND2X1 NAND2X1_227 ( .A(_abc_15497_new_n2961_), .B(_abc_15497_new_n2963_), .Y(_abc_15497_new_n2967_));
NAND2X1 NAND2X1_228 ( .A(_abc_15497_new_n2966_), .B(_abc_15497_new_n2967_), .Y(_abc_15497_new_n2968_));
NAND2X1 NAND2X1_229 ( .A(_abc_15497_new_n2964_), .B(_abc_15497_new_n2968_), .Y(_abc_15497_new_n2982_));
NAND2X1 NAND2X1_23 ( .A(_abc_15497_new_n938_), .B(_abc_15497_new_n942_), .Y(_abc_15497_new_n948_));
NAND2X1 NAND2X1_230 ( .A(_abc_15497_new_n2989_), .B(_abc_15497_new_n2993_), .Y(_abc_15497_new_n2997_));
NAND2X1 NAND2X1_231 ( .A(_abc_15497_new_n2994_), .B(_abc_15497_new_n2942_), .Y(_abc_15497_new_n3002_));
NAND2X1 NAND2X1_232 ( .A(_abc_15497_new_n2982_), .B(_abc_15497_new_n2980_), .Y(_abc_15497_new_n3004_));
NAND2X1 NAND2X1_233 ( .A(b_reg_5_), .B(c_reg_5_), .Y(_abc_15497_new_n3009_));
NAND2X1 NAND2X1_234 ( .A(_abc_15497_new_n3015_), .B(_abc_15497_new_n3013_), .Y(_abc_15497_new_n3016_));
NAND2X1 NAND2X1_235 ( .A(e_reg_5_), .B(a_reg_0_), .Y(_abc_15497_new_n3020_));
NAND2X1 NAND2X1_236 ( .A(_abc_15497_new_n3016_), .B(_abc_15497_new_n3030_), .Y(_abc_15497_new_n3031_));
NAND2X1 NAND2X1_237 ( .A(_abc_15497_new_n3025_), .B(_abc_15497_new_n3029_), .Y(_abc_15497_new_n3033_));
NAND2X1 NAND2X1_238 ( .A(_abc_15497_new_n3033_), .B(_abc_15497_new_n3032_), .Y(_abc_15497_new_n3034_));
NAND2X1 NAND2X1_239 ( .A(_abc_15497_new_n3033_), .B(_abc_15497_new_n3016_), .Y(_abc_15497_new_n3038_));
NAND2X1 NAND2X1_24 ( .A(_abc_15497_new_n950_), .B(_abc_15497_new_n949_), .Y(_abc_15497_new_n951_));
NAND2X1 NAND2X1_240 ( .A(_abc_15497_new_n3030_), .B(_abc_15497_new_n3032_), .Y(_abc_15497_new_n3039_));
NAND2X1 NAND2X1_241 ( .A(_abc_15497_new_n2969_), .B(_abc_15497_new_n3004_), .Y(_abc_15497_new_n3046_));
NAND2X1 NAND2X1_242 ( .A(_abc_15497_new_n3045_), .B(_abc_15497_new_n3051_), .Y(_abc_15497_new_n3052_));
NAND2X1 NAND2X1_243 ( .A(_abc_15497_new_n3058_), .B(_abc_15497_new_n2942_), .Y(_abc_15497_new_n3059_));
NAND2X1 NAND2X1_244 ( .A(_abc_15497_new_n3062_), .B(_abc_15497_new_n3059_), .Y(_abc_15497_new_n3063_));
NAND2X1 NAND2X1_245 ( .A(b_reg_6_), .B(c_reg_6_), .Y(_abc_15497_new_n3067_));
NAND2X1 NAND2X1_246 ( .A(_abc_15497_new_n3073_), .B(_abc_15497_new_n3071_), .Y(_abc_15497_new_n3074_));
NAND2X1 NAND2X1_247 ( .A(e_reg_6_), .B(a_reg_1_), .Y(_abc_15497_new_n3078_));
NAND2X1 NAND2X1_248 ( .A(_abc_15497_new_n3074_), .B(_abc_15497_new_n3088_), .Y(_abc_15497_new_n3089_));
NAND2X1 NAND2X1_249 ( .A(_abc_15497_new_n3083_), .B(_abc_15497_new_n3087_), .Y(_abc_15497_new_n3091_));
NAND2X1 NAND2X1_25 ( .A(_abc_15497_new_n959_), .B(_abc_15497_new_n962_), .Y(_abc_15497_new_n963_));
NAND2X1 NAND2X1_250 ( .A(_abc_15497_new_n3091_), .B(_abc_15497_new_n3090_), .Y(_abc_15497_new_n3092_));
NAND2X1 NAND2X1_251 ( .A(_abc_15497_new_n3091_), .B(_abc_15497_new_n3074_), .Y(_abc_15497_new_n3096_));
NAND2X1 NAND2X1_252 ( .A(_abc_15497_new_n3088_), .B(_abc_15497_new_n3090_), .Y(_abc_15497_new_n3097_));
NAND2X1 NAND2X1_253 ( .A(_abc_15497_new_n3103_), .B(_abc_15497_new_n3107_), .Y(_abc_15497_new_n3108_));
NAND2X1 NAND2X1_254 ( .A(b_reg_7_), .B(c_reg_7_), .Y(_abc_15497_new_n3121_));
NAND2X1 NAND2X1_255 ( .A(e_reg_7_), .B(a_reg_2_), .Y(_abc_15497_new_n3133_));
NAND2X1 NAND2X1_256 ( .A(_abc_15497_new_n3138_), .B(_abc_15497_new_n3142_), .Y(_abc_15497_new_n3143_));
NAND2X1 NAND2X1_257 ( .A(_abc_15497_new_n3146_), .B(_abc_15497_new_n3145_), .Y(_abc_15497_new_n3147_));
NAND2X1 NAND2X1_258 ( .A(_abc_15497_new_n3148_), .B(_abc_15497_new_n3149_), .Y(_abc_15497_new_n3150_));
NAND2X1 NAND2X1_259 ( .A(_abc_15497_new_n3158_), .B(_abc_15497_new_n3118_), .Y(_abc_15497_new_n3159_));
NAND2X1 NAND2X1_26 ( .A(e_reg_4_), .B(_auto_iopadmap_cc_368_execute_22625_4_), .Y(_abc_15497_new_n967_));
NAND2X1 NAND2X1_260 ( .A(_abc_15497_new_n3157_), .B(_abc_15497_new_n3152_), .Y(_abc_15497_new_n3160_));
NAND2X1 NAND2X1_261 ( .A(_abc_15497_new_n3161_), .B(_abc_15497_new_n3159_), .Y(_abc_15497_new_n3162_));
NAND2X1 NAND2X1_262 ( .A(b_reg_8_), .B(c_reg_8_), .Y(_abc_15497_new_n3171_));
NAND2X1 NAND2X1_263 ( .A(e_reg_8_), .B(a_reg_3_), .Y(_abc_15497_new_n3181_));
NAND2X1 NAND2X1_264 ( .A(_abc_15497_new_n3183_), .B(_abc_15497_new_n3185_), .Y(_abc_15497_new_n3186_));
NAND2X1 NAND2X1_265 ( .A(_abc_15497_new_n3177_), .B(_abc_15497_new_n3175_), .Y(_abc_15497_new_n3190_));
NAND2X1 NAND2X1_266 ( .A(_abc_15497_new_n3192_), .B(_abc_15497_new_n3186_), .Y(_abc_15497_new_n3193_));
NAND2X1 NAND2X1_267 ( .A(_abc_15497_new_n3191_), .B(_abc_15497_new_n3193_), .Y(_abc_15497_new_n3200_));
NAND2X1 NAND2X1_268 ( .A(_abc_15497_new_n3200_), .B(_abc_15497_new_n3199_), .Y(_abc_15497_new_n3201_));
NAND2X1 NAND2X1_269 ( .A(_abc_15497_new_n3207_), .B(_abc_15497_new_n3210_), .Y(_abc_15497_new_n3211_));
NAND2X1 NAND2X1_27 ( .A(_abc_15497_new_n967_), .B(_abc_15497_new_n966_), .Y(_abc_15497_new_n968_));
NAND2X1 NAND2X1_270 ( .A(_abc_15497_new_n3232_), .B(_abc_15497_new_n738_), .Y(_abc_15497_new_n3233_));
NAND2X1 NAND2X1_271 ( .A(e_reg_9_), .B(a_reg_4_), .Y(_abc_15497_new_n3244_));
NAND2X1 NAND2X1_272 ( .A(_abc_15497_new_n1034_), .B(_abc_15497_new_n2130_), .Y(_abc_15497_new_n3247_));
NAND2X1 NAND2X1_273 ( .A(_abc_15497_new_n3248_), .B(_abc_15497_new_n3246_), .Y(_abc_15497_new_n3249_));
NAND2X1 NAND2X1_274 ( .A(b_reg_9_), .B(c_reg_9_), .Y(_abc_15497_new_n3254_));
NAND2X1 NAND2X1_275 ( .A(d_reg_9_), .B(_abc_15497_new_n3231_), .Y(_abc_15497_new_n3256_));
NAND2X1 NAND2X1_276 ( .A(_abc_15497_new_n3259_), .B(_abc_15497_new_n3262_), .Y(_abc_15497_new_n3263_));
NAND2X1 NAND2X1_277 ( .A(_abc_15497_new_n3263_), .B(_abc_15497_new_n3258_), .Y(_abc_15497_new_n3264_));
NAND2X1 NAND2X1_278 ( .A(_abc_15497_new_n3253_), .B(_abc_15497_new_n3264_), .Y(_abc_15497_new_n3270_));
NAND2X1 NAND2X1_279 ( .A(b_reg_10_), .B(c_reg_10_), .Y(_abc_15497_new_n3292_));
NAND2X1 NAND2X1_28 ( .A(_abc_15497_new_n968_), .B(_abc_15497_new_n969_), .Y(_abc_15497_new_n972_));
NAND2X1 NAND2X1_280 ( .A(_abc_15497_new_n3298_), .B(_abc_15497_new_n3296_), .Y(_abc_15497_new_n3299_));
NAND2X1 NAND2X1_281 ( .A(e_reg_10_), .B(a_reg_5_), .Y(_abc_15497_new_n3304_));
NAND2X1 NAND2X1_282 ( .A(_abc_15497_new_n3309_), .B(_abc_15497_new_n3312_), .Y(_abc_15497_new_n3313_));
NAND2X1 NAND2X1_283 ( .A(_abc_15497_new_n3313_), .B(_abc_15497_new_n3299_), .Y(_abc_15497_new_n3314_));
NAND2X1 NAND2X1_284 ( .A(_abc_15497_new_n3319_), .B(_abc_15497_new_n3320_), .Y(_abc_15497_new_n3321_));
NAND2X1 NAND2X1_285 ( .A(_abc_15497_new_n3321_), .B(_abc_15497_new_n3318_), .Y(_abc_15497_new_n3322_));
NAND2X1 NAND2X1_286 ( .A(_abc_15497_new_n3321_), .B(_abc_15497_new_n3299_), .Y(_abc_15497_new_n3324_));
NAND2X1 NAND2X1_287 ( .A(_abc_15497_new_n3313_), .B(_abc_15497_new_n3318_), .Y(_abc_15497_new_n3325_));
NAND2X1 NAND2X1_288 ( .A(_abc_15497_new_n3340_), .B(_abc_15497_new_n3336_), .Y(_abc_15497_new_n3341_));
NAND2X1 NAND2X1_289 ( .A(b_reg_11_), .B(c_reg_11_), .Y(_abc_15497_new_n3353_));
NAND2X1 NAND2X1_29 ( .A(e_reg_7_), .B(_auto_iopadmap_cc_368_execute_22625_7_), .Y(_abc_15497_new_n996_));
NAND2X1 NAND2X1_290 ( .A(_abc_15497_new_n1684_), .B(_abc_15497_new_n2144_), .Y(_abc_15497_new_n3365_));
NAND2X1 NAND2X1_291 ( .A(e_reg_11_), .B(a_reg_6_), .Y(_abc_15497_new_n3366_));
NAND2X1 NAND2X1_292 ( .A(_abc_15497_new_n3368_), .B(_abc_15497_new_n3372_), .Y(_abc_15497_new_n3373_));
NAND2X1 NAND2X1_293 ( .A(_abc_15497_new_n3359_), .B(_abc_15497_new_n3357_), .Y(_abc_15497_new_n3375_));
NAND2X1 NAND2X1_294 ( .A(_abc_15497_new_n3377_), .B(_abc_15497_new_n3376_), .Y(_abc_15497_new_n3378_));
NAND2X1 NAND2X1_295 ( .A(_abc_15497_new_n3390_), .B(_abc_15497_new_n3396_), .Y(_abc_15497_new_n3404_));
NAND2X1 NAND2X1_296 ( .A(_abc_15497_new_n3373_), .B(_abc_15497_new_n3375_), .Y(_abc_15497_new_n3410_));
NAND2X1 NAND2X1_297 ( .A(_abc_15497_new_n3378_), .B(_abc_15497_new_n3414_), .Y(_abc_15497_new_n3415_));
NAND2X1 NAND2X1_298 ( .A(b_reg_12_), .B(c_reg_12_), .Y(_abc_15497_new_n3420_));
NAND2X1 NAND2X1_299 ( .A(d_reg_12_), .B(_abc_15497_new_n3422_), .Y(_abc_15497_new_n3423_));
NAND2X1 NAND2X1_3 ( .A(_abc_15497_new_n752_), .B(_abc_15497_new_n756_), .Y(_abc_15497_new_n757_));
NAND2X1 NAND2X1_30 ( .A(_abc_15497_new_n996_), .B(_abc_15497_new_n995_), .Y(_abc_15497_new_n997_));
NAND2X1 NAND2X1_300 ( .A(_abc_15497_new_n3427_), .B(_abc_15497_new_n3425_), .Y(_abc_15497_new_n3428_));
NAND2X1 NAND2X1_301 ( .A(e_reg_12_), .B(a_reg_7_), .Y(_abc_15497_new_n3433_));
NAND2X1 NAND2X1_302 ( .A(_abc_15497_new_n1064_), .B(_abc_15497_new_n2159_), .Y(_abc_15497_new_n3436_));
NAND2X1 NAND2X1_303 ( .A(_abc_15497_new_n3438_), .B(_abc_15497_new_n3441_), .Y(_abc_15497_new_n3442_));
NAND2X1 NAND2X1_304 ( .A(_abc_15497_new_n3442_), .B(_abc_15497_new_n3428_), .Y(_abc_15497_new_n3443_));
NAND2X1 NAND2X1_305 ( .A(_abc_15497_new_n1414_), .B(_abc_15497_new_n3420_), .Y(_abc_15497_new_n3444_));
NAND2X1 NAND2X1_306 ( .A(_abc_15497_new_n3449_), .B(_abc_15497_new_n3450_), .Y(_abc_15497_new_n3451_));
NAND2X1 NAND2X1_307 ( .A(_abc_15497_new_n3451_), .B(_abc_15497_new_n3448_), .Y(_abc_15497_new_n3452_));
NAND2X1 NAND2X1_308 ( .A(_abc_15497_new_n3451_), .B(_abc_15497_new_n3428_), .Y(_abc_15497_new_n3456_));
NAND2X1 NAND2X1_309 ( .A(_abc_15497_new_n3442_), .B(_abc_15497_new_n3448_), .Y(_abc_15497_new_n3457_));
NAND2X1 NAND2X1_31 ( .A(_abc_15497_new_n998_), .B(_abc_15497_new_n993_), .Y(_abc_15497_new_n999_));
NAND2X1 NAND2X1_310 ( .A(_abc_15497_new_n3378_), .B(_abc_15497_new_n3375_), .Y(_abc_15497_new_n3464_));
NAND2X1 NAND2X1_311 ( .A(_abc_15497_new_n3373_), .B(_abc_15497_new_n3414_), .Y(_abc_15497_new_n3465_));
NAND2X1 NAND2X1_312 ( .A(_abc_15497_new_n3471_), .B(_abc_15497_new_n3409_), .Y(_abc_15497_new_n3473_));
NAND2X1 NAND2X1_313 ( .A(round_ctr_inc_bF_buf11), .B(_abc_15497_new_n3473_), .Y(_abc_15497_new_n3474_));
NAND2X1 NAND2X1_314 ( .A(_abc_15497_new_n3470_), .B(_abc_15497_new_n3473_), .Y(_abc_15497_new_n3478_));
NAND2X1 NAND2X1_315 ( .A(_abc_15497_new_n1881_), .B(_abc_15497_new_n708_), .Y(_abc_15497_new_n3484_));
NAND2X1 NAND2X1_316 ( .A(b_reg_13_), .B(c_reg_13_), .Y(_abc_15497_new_n3485_));
NAND2X1 NAND2X1_317 ( .A(_abc_15497_new_n3483_), .B(_abc_15497_new_n3486_), .Y(_abc_15497_new_n3487_));
NAND2X1 NAND2X1_318 ( .A(e_reg_13_), .B(a_reg_8_), .Y(_abc_15497_new_n3499_));
NAND2X1 NAND2X1_319 ( .A(_abc_15497_new_n3497_), .B(_abc_15497_new_n3500_), .Y(_abc_15497_new_n3501_));
NAND2X1 NAND2X1_32 ( .A(_abc_15497_new_n1003_), .B(_abc_15497_new_n1002_), .Y(_0H4_reg_31_0__7_));
NAND2X1 NAND2X1_320 ( .A(_abc_15497_new_n3503_), .B(_abc_15497_new_n3501_), .Y(_abc_15497_new_n3509_));
NAND2X1 NAND2X1_321 ( .A(_abc_15497_new_n3508_), .B(_abc_15497_new_n3509_), .Y(_abc_15497_new_n3510_));
NAND2X1 NAND2X1_322 ( .A(_abc_15497_new_n3510_), .B(_abc_15497_new_n3507_), .Y(_abc_15497_new_n3511_));
NAND2X1 NAND2X1_323 ( .A(_abc_15497_new_n3522_), .B(_abc_15497_new_n3526_), .Y(_abc_15497_new_n3527_));
NAND2X1 NAND2X1_324 ( .A(_abc_15497_new_n3535_), .B(_abc_15497_new_n3526_), .Y(_abc_15497_new_n3536_));
NAND2X1 NAND2X1_325 ( .A(_abc_15497_new_n3463_), .B(_abc_15497_new_n3470_), .Y(_abc_15497_new_n3537_));
NAND2X1 NAND2X1_326 ( .A(_abc_15497_new_n3538_), .B(_abc_15497_new_n3409_), .Y(_abc_15497_new_n3539_));
NAND2X1 NAND2X1_327 ( .A(_abc_15497_new_n1876_), .B(_abc_15497_new_n702_), .Y(_abc_15497_new_n3547_));
NAND2X1 NAND2X1_328 ( .A(b_reg_14_), .B(c_reg_14_), .Y(_abc_15497_new_n3548_));
NAND2X1 NAND2X1_329 ( .A(_abc_15497_new_n3546_), .B(_abc_15497_new_n3549_), .Y(_abc_15497_new_n3550_));
NAND2X1 NAND2X1_33 ( .A(_abc_15497_new_n1009_), .B(_abc_15497_new_n1010_), .Y(_abc_15497_new_n1011_));
NAND2X1 NAND2X1_330 ( .A(_abc_15497_new_n1080_), .B(_abc_15497_new_n2187_), .Y(_abc_15497_new_n3563_));
NAND2X1 NAND2X1_331 ( .A(e_reg_14_), .B(a_reg_9_), .Y(_abc_15497_new_n3564_));
NAND2X1 NAND2X1_332 ( .A(_abc_15497_new_n3569_), .B(_abc_15497_new_n3566_), .Y(_abc_15497_new_n3570_));
NAND2X1 NAND2X1_333 ( .A(_abc_15497_new_n3574_), .B(_abc_15497_new_n3575_), .Y(_abc_15497_new_n3576_));
NAND2X1 NAND2X1_334 ( .A(_abc_15497_new_n3576_), .B(_abc_15497_new_n3573_), .Y(_abc_15497_new_n3577_));
NAND2X1 NAND2X1_335 ( .A(_abc_15497_new_n3570_), .B(_abc_15497_new_n3573_), .Y(_abc_15497_new_n3580_));
NAND2X1 NAND2X1_336 ( .A(_abc_15497_new_n3591_), .B(_abc_15497_new_n3595_), .Y(_abc_15497_new_n3596_));
NAND2X1 NAND2X1_337 ( .A(_abc_15497_new_n3596_), .B(_abc_15497_new_n3540_), .Y(_abc_15497_new_n3598_));
NAND2X1 NAND2X1_338 ( .A(round_ctr_inc_bF_buf9), .B(_abc_15497_new_n3598_), .Y(_abc_15497_new_n3599_));
NAND2X1 NAND2X1_339 ( .A(_abc_15497_new_n3590_), .B(_abc_15497_new_n3582_), .Y(_abc_15497_new_n3603_));
NAND2X1 NAND2X1_34 ( .A(_abc_15497_new_n991_), .B(_abc_15497_new_n998_), .Y(_abc_15497_new_n1013_));
NAND2X1 NAND2X1_340 ( .A(_abc_15497_new_n3608_), .B(_abc_15497_new_n3609_), .Y(_abc_15497_new_n3610_));
NAND2X1 NAND2X1_341 ( .A(b_reg_15_), .B(c_reg_15_), .Y(_abc_15497_new_n3616_));
NAND2X1 NAND2X1_342 ( .A(_abc_15497_new_n3617_), .B(_abc_15497_new_n2743__bF_buf2), .Y(_abc_15497_new_n3618_));
NAND2X1 NAND2X1_343 ( .A(e_reg_15_), .B(a_reg_10_), .Y(_abc_15497_new_n3624_));
NAND2X1 NAND2X1_344 ( .A(_abc_15497_new_n3629_), .B(_abc_15497_new_n3632_), .Y(_abc_15497_new_n3633_));
NAND2X1 NAND2X1_345 ( .A(_abc_15497_new_n3639_), .B(_abc_15497_new_n3640_), .Y(_abc_15497_new_n3641_));
NAND2X1 NAND2X1_346 ( .A(_abc_15497_new_n3655_), .B(_abc_15497_new_n3659_), .Y(_abc_15497_new_n3660_));
NAND2X1 NAND2X1_347 ( .A(_abc_15497_new_n3668_), .B(_abc_15497_new_n3538_), .Y(_abc_15497_new_n3669_));
NAND2X1 NAND2X1_348 ( .A(_abc_15497_new_n3522_), .B(_abc_15497_new_n3536_), .Y(_abc_15497_new_n3670_));
NAND2X1 NAND2X1_349 ( .A(_abc_15497_new_n3639_), .B(_abc_15497_new_n3634_), .Y(_abc_15497_new_n3680_));
NAND2X1 NAND2X1_35 ( .A(_abc_15497_new_n1020_), .B(_abc_15497_new_n1018_), .Y(_abc_15497_new_n1021_));
NAND2X1 NAND2X1_350 ( .A(_abc_15497_new_n3689_), .B(_abc_15497_new_n3685_), .Y(_abc_15497_new_n3690_));
NAND2X1 NAND2X1_351 ( .A(_abc_15497_new_n3692_), .B(_abc_15497_new_n3693_), .Y(_abc_15497_new_n3694_));
NAND2X1 NAND2X1_352 ( .A(_abc_15497_new_n3694_), .B(_abc_15497_new_n3695_), .Y(_abc_15497_new_n3696_));
NAND2X1 NAND2X1_353 ( .A(_abc_15497_new_n3690_), .B(_abc_15497_new_n3697_), .Y(_abc_15497_new_n3698_));
NAND2X1 NAND2X1_354 ( .A(_abc_15497_new_n3699_), .B(_abc_15497_new_n3700_), .Y(_abc_15497_new_n3701_));
NAND2X1 NAND2X1_355 ( .A(_abc_15497_new_n3690_), .B(_abc_15497_new_n3700_), .Y(_abc_15497_new_n3703_));
NAND2X1 NAND2X1_356 ( .A(_abc_15497_new_n3699_), .B(_abc_15497_new_n3697_), .Y(_abc_15497_new_n3704_));
NAND2X1 NAND2X1_357 ( .A(_abc_15497_new_n3710_), .B(_abc_15497_new_n3712_), .Y(_abc_15497_new_n3714_));
NAND2X1 NAND2X1_358 ( .A(_abc_15497_new_n3726_), .B(_abc_15497_new_n3727_), .Y(_abc_15497_new_n3728_));
NAND2X1 NAND2X1_359 ( .A(b_reg_17_), .B(c_reg_17_), .Y(_abc_15497_new_n3729_));
NAND2X1 NAND2X1_36 ( .A(_abc_15497_new_n1025_), .B(_abc_15497_new_n1019_), .Y(_abc_15497_new_n1026_));
NAND2X1 NAND2X1_360 ( .A(_abc_15497_new_n3728_), .B(_abc_15497_new_n3731_), .Y(_abc_15497_new_n3732_));
NAND2X1 NAND2X1_361 ( .A(w_17_), .B(_abc_15497_new_n3742_), .Y(_abc_15497_new_n3743_));
NAND2X1 NAND2X1_362 ( .A(_abc_15497_new_n3741_), .B(_abc_15497_new_n3743_), .Y(_abc_15497_new_n3747_));
NAND2X1 NAND2X1_363 ( .A(_abc_15497_new_n3746_), .B(_abc_15497_new_n3747_), .Y(_abc_15497_new_n3748_));
NAND2X1 NAND2X1_364 ( .A(_abc_15497_new_n3735_), .B(_abc_15497_new_n3749_), .Y(_abc_15497_new_n3750_));
NAND2X1 NAND2X1_365 ( .A(_abc_15497_new_n3748_), .B(_abc_15497_new_n3745_), .Y(_abc_15497_new_n3752_));
NAND2X1 NAND2X1_366 ( .A(_abc_15497_new_n3751_), .B(_abc_15497_new_n3752_), .Y(_abc_15497_new_n3753_));
NAND2X1 NAND2X1_367 ( .A(_abc_15497_new_n3764_), .B(_abc_15497_new_n3768_), .Y(_abc_15497_new_n3769_));
NAND2X1 NAND2X1_368 ( .A(b_reg_18_), .B(_abc_15497_new_n823_), .Y(_abc_15497_new_n3784_));
NAND2X1 NAND2X1_369 ( .A(c_reg_18_), .B(_abc_15497_new_n3785_), .Y(_abc_15497_new_n3786_));
NAND2X1 NAND2X1_37 ( .A(_abc_15497_new_n1008_), .B(_abc_15497_new_n1025_), .Y(_abc_15497_new_n1035_));
NAND2X1 NAND2X1_370 ( .A(_abc_15497_new_n3784_), .B(_abc_15497_new_n3786_), .Y(_abc_15497_new_n3787_));
NAND2X1 NAND2X1_371 ( .A(_abc_15497_new_n3792_), .B(_abc_15497_new_n2759__bF_buf2), .Y(_abc_15497_new_n3793_));
NAND2X1 NAND2X1_372 ( .A(_abc_15497_new_n3797_), .B(_abc_15497_new_n3798_), .Y(_abc_15497_new_n3799_));
NAND2X1 NAND2X1_373 ( .A(_abc_15497_new_n3799_), .B(_abc_15497_new_n3800_), .Y(_abc_15497_new_n3801_));
NAND2X1 NAND2X1_374 ( .A(_abc_15497_new_n3795_), .B(_abc_15497_new_n3802_), .Y(_abc_15497_new_n3803_));
NAND2X1 NAND2X1_375 ( .A(_abc_15497_new_n3796_), .B(_abc_15497_new_n3805_), .Y(_abc_15497_new_n3806_));
NAND2X1 NAND2X1_376 ( .A(_abc_15497_new_n3783_), .B(_abc_15497_new_n3809_), .Y(_abc_15497_new_n3810_));
NAND2X1 NAND2X1_377 ( .A(_abc_15497_new_n3803_), .B(_abc_15497_new_n3808_), .Y(_abc_15497_new_n3812_));
NAND2X1 NAND2X1_378 ( .A(_abc_15497_new_n3811_), .B(_abc_15497_new_n3812_), .Y(_abc_15497_new_n3813_));
NAND2X1 NAND2X1_379 ( .A(_abc_15497_new_n3813_), .B(_abc_15497_new_n3810_), .Y(_abc_15497_new_n3814_));
NAND2X1 NAND2X1_38 ( .A(e_reg_10_), .B(_auto_iopadmap_cc_368_execute_22625_10_), .Y(_abc_15497_new_n1040_));
NAND2X1 NAND2X1_380 ( .A(_abc_15497_new_n3782_), .B(_abc_15497_new_n3814_), .Y(_abc_15497_new_n3815_));
NAND2X1 NAND2X1_381 ( .A(_abc_15497_new_n3815_), .B(_abc_15497_new_n3817_), .Y(_abc_15497_new_n3818_));
NAND2X1 NAND2X1_382 ( .A(_abc_15497_new_n1495_), .B(_abc_15497_new_n3833_), .Y(_abc_15497_new_n3834_));
NAND2X1 NAND2X1_383 ( .A(_abc_15497_new_n3837_), .B(_abc_15497_new_n2759__bF_buf1), .Y(_abc_15497_new_n3838_));
NAND2X1 NAND2X1_384 ( .A(_abc_15497_new_n3841_), .B(_abc_15497_new_n3842_), .Y(_abc_15497_new_n3843_));
NAND2X1 NAND2X1_385 ( .A(_abc_15497_new_n3843_), .B(_abc_15497_new_n3844_), .Y(_abc_15497_new_n3845_));
NAND2X1 NAND2X1_386 ( .A(_abc_15497_new_n3848_), .B(_abc_15497_new_n3849_), .Y(_abc_15497_new_n3850_));
NAND2X1 NAND2X1_387 ( .A(_abc_15497_new_n3848_), .B(_abc_15497_new_n3846_), .Y(_abc_15497_new_n3854_));
NAND2X1 NAND2X1_388 ( .A(_abc_15497_new_n3863_), .B(_abc_15497_new_n3860_), .Y(_abc_15497_new_n3864_));
NAND2X1 NAND2X1_389 ( .A(_abc_15497_new_n3811_), .B(_abc_15497_new_n3809_), .Y(_abc_15497_new_n3871_));
NAND2X1 NAND2X1_39 ( .A(digest_update_bF_buf8), .B(_abc_15497_new_n1045_), .Y(_abc_15497_new_n1046_));
NAND2X1 NAND2X1_390 ( .A(_abc_15497_new_n3783_), .B(_abc_15497_new_n3812_), .Y(_abc_15497_new_n3872_));
NAND2X1 NAND2X1_391 ( .A(_abc_15497_new_n3861_), .B(_abc_15497_new_n3862_), .Y(_abc_15497_new_n3878_));
NAND2X1 NAND2X1_392 ( .A(_abc_15497_new_n3901_), .B(_abc_15497_new_n3897_), .Y(_abc_15497_new_n3902_));
NAND2X1 NAND2X1_393 ( .A(_abc_15497_new_n3904_), .B(_abc_15497_new_n3905_), .Y(_abc_15497_new_n3906_));
NAND2X1 NAND2X1_394 ( .A(_abc_15497_new_n3906_), .B(_abc_15497_new_n3907_), .Y(_abc_15497_new_n3908_));
NAND2X1 NAND2X1_395 ( .A(_abc_15497_new_n3902_), .B(_abc_15497_new_n3909_), .Y(_abc_15497_new_n3910_));
NAND2X1 NAND2X1_396 ( .A(_abc_15497_new_n3911_), .B(_abc_15497_new_n3912_), .Y(_abc_15497_new_n3913_));
NAND2X1 NAND2X1_397 ( .A(_abc_15497_new_n3902_), .B(_abc_15497_new_n3912_), .Y(_abc_15497_new_n3916_));
NAND2X1 NAND2X1_398 ( .A(_abc_15497_new_n3911_), .B(_abc_15497_new_n3909_), .Y(_abc_15497_new_n3917_));
NAND2X1 NAND2X1_399 ( .A(_abc_15497_new_n3927_), .B(_abc_15497_new_n3923_), .Y(_abc_15497_new_n3928_));
NAND2X1 NAND2X1_4 ( .A(c_reg_4_), .B(_auto_iopadmap_cc_368_execute_22625_68_), .Y(_abc_15497_new_n764_));
NAND2X1 NAND2X1_40 ( .A(e_reg_11_), .B(_auto_iopadmap_cc_368_execute_22625_11_), .Y(_abc_15497_new_n1053_));
NAND2X1 NAND2X1_400 ( .A(_abc_15497_new_n3928_), .B(_abc_15497_new_n3885_), .Y(_abc_15497_new_n3930_));
NAND2X1 NAND2X1_401 ( .A(round_ctr_inc_bF_buf4), .B(_abc_15497_new_n3930_), .Y(_abc_15497_new_n3931_));
NAND2X1 NAND2X1_402 ( .A(_abc_15497_new_n3952_), .B(_abc_15497_new_n3947_), .Y(_abc_15497_new_n3953_));
NAND2X1 NAND2X1_403 ( .A(_abc_15497_new_n3955_), .B(_abc_15497_new_n3956_), .Y(_abc_15497_new_n3957_));
NAND2X1 NAND2X1_404 ( .A(_abc_15497_new_n3957_), .B(_abc_15497_new_n3958_), .Y(_abc_15497_new_n3959_));
NAND2X1 NAND2X1_405 ( .A(_abc_15497_new_n3953_), .B(_abc_15497_new_n3960_), .Y(_abc_15497_new_n3961_));
NAND2X1 NAND2X1_406 ( .A(_abc_15497_new_n3962_), .B(_abc_15497_new_n3963_), .Y(_abc_15497_new_n3964_));
NAND2X1 NAND2X1_407 ( .A(_abc_15497_new_n3953_), .B(_abc_15497_new_n3963_), .Y(_abc_15497_new_n3967_));
NAND2X1 NAND2X1_408 ( .A(_abc_15497_new_n3962_), .B(_abc_15497_new_n3960_), .Y(_abc_15497_new_n3968_));
NAND2X1 NAND2X1_409 ( .A(_abc_15497_new_n3974_), .B(_abc_15497_new_n3978_), .Y(_abc_15497_new_n3979_));
NAND2X1 NAND2X1_41 ( .A(_abc_15497_new_n1053_), .B(_abc_15497_new_n1052_), .Y(_abc_15497_new_n1054_));
NAND2X1 NAND2X1_410 ( .A(_abc_15497_new_n3986_), .B(_abc_15497_new_n3885_), .Y(_abc_15497_new_n3987_));
NAND2X1 NAND2X1_411 ( .A(_abc_15497_new_n4007_), .B(_abc_15497_new_n4002_), .Y(_abc_15497_new_n4008_));
NAND2X1 NAND2X1_412 ( .A(_abc_15497_new_n4010_), .B(_abc_15497_new_n4011_), .Y(_abc_15497_new_n4012_));
NAND2X1 NAND2X1_413 ( .A(_abc_15497_new_n4012_), .B(_abc_15497_new_n4013_), .Y(_abc_15497_new_n4014_));
NAND2X1 NAND2X1_414 ( .A(_abc_15497_new_n4008_), .B(_abc_15497_new_n4015_), .Y(_abc_15497_new_n4016_));
NAND2X1 NAND2X1_415 ( .A(_abc_15497_new_n4017_), .B(_abc_15497_new_n4018_), .Y(_abc_15497_new_n4019_));
NAND2X1 NAND2X1_416 ( .A(_abc_15497_new_n4008_), .B(_abc_15497_new_n4018_), .Y(_abc_15497_new_n4022_));
NAND2X1 NAND2X1_417 ( .A(_abc_15497_new_n4017_), .B(_abc_15497_new_n4015_), .Y(_abc_15497_new_n4023_));
NAND2X1 NAND2X1_418 ( .A(_abc_15497_new_n4029_), .B(_abc_15497_new_n4033_), .Y(_abc_15497_new_n4034_));
NAND2X1 NAND2X1_419 ( .A(_abc_15497_new_n1543_), .B(_abc_15497_new_n4050_), .Y(_abc_15497_new_n4051_));
NAND2X1 NAND2X1_42 ( .A(_abc_15497_new_n1066_), .B(_abc_15497_new_n1062_), .Y(_abc_15497_new_n1068_));
NAND2X1 NAND2X1_420 ( .A(b_reg_23_), .B(c_reg_23_), .Y(_abc_15497_new_n4052_));
NAND2X1 NAND2X1_421 ( .A(_abc_15497_new_n4051_), .B(_abc_15497_new_n4054_), .Y(_abc_15497_new_n4055_));
NAND2X1 NAND2X1_422 ( .A(_abc_15497_new_n4064_), .B(_abc_15497_new_n4065_), .Y(_abc_15497_new_n4066_));
NAND2X1 NAND2X1_423 ( .A(_abc_15497_new_n4066_), .B(_abc_15497_new_n4067_), .Y(_abc_15497_new_n4069_));
NAND2X1 NAND2X1_424 ( .A(_abc_15497_new_n4068_), .B(_abc_15497_new_n4070_), .Y(_abc_15497_new_n4071_));
NAND2X1 NAND2X1_425 ( .A(_abc_15497_new_n4059_), .B(_abc_15497_new_n4071_), .Y(_abc_15497_new_n4073_));
NAND2X1 NAND2X1_426 ( .A(_abc_15497_new_n4058_), .B(_abc_15497_new_n4071_), .Y(_abc_15497_new_n4077_));
NAND2X1 NAND2X1_427 ( .A(_abc_15497_new_n4084_), .B(_abc_15497_new_n4088_), .Y(_abc_15497_new_n4089_));
NAND2X1 NAND2X1_428 ( .A(round_ctr_inc_bF_buf1), .B(_abc_15497_new_n4092_), .Y(_abc_15497_new_n4093_));
NAND2X1 NAND2X1_429 ( .A(_abc_15497_new_n4034_), .B(_abc_15497_new_n4089_), .Y(_abc_15497_new_n4099_));
NAND2X1 NAND2X1_43 ( .A(digest_update_bF_buf7), .B(_abc_15497_new_n1068_), .Y(_abc_15497_new_n1069_));
NAND2X1 NAND2X1_430 ( .A(b_reg_24_), .B(c_reg_24_), .Y(_abc_15497_new_n4110_));
NAND2X1 NAND2X1_431 ( .A(_abc_15497_new_n4116_), .B(_abc_15497_new_n4114_), .Y(_abc_15497_new_n4117_));
NAND2X1 NAND2X1_432 ( .A(w_24_), .B(_abc_15497_new_n4126_), .Y(_abc_15497_new_n4127_));
NAND2X1 NAND2X1_433 ( .A(_abc_15497_new_n4125_), .B(_abc_15497_new_n4127_), .Y(_abc_15497_new_n4129_));
NAND2X1 NAND2X1_434 ( .A(_abc_15497_new_n4128_), .B(_abc_15497_new_n4130_), .Y(_abc_15497_new_n4131_));
NAND2X1 NAND2X1_435 ( .A(_abc_15497_new_n4108_), .B(_abc_15497_new_n4132_), .Y(_abc_15497_new_n4134_));
NAND2X1 NAND2X1_436 ( .A(_abc_15497_new_n2759__bF_buf1), .B(_abc_15497_new_n4136_), .Y(_abc_15497_new_n4137_));
NAND2X1 NAND2X1_437 ( .A(_abc_15497_new_n4138_), .B(_abc_15497_new_n4137_), .Y(_abc_15497_new_n4139_));
NAND2X1 NAND2X1_438 ( .A(_abc_15497_new_n4107_), .B(_abc_15497_new_n4139_), .Y(_abc_15497_new_n4140_));
NAND2X1 NAND2X1_439 ( .A(_abc_15497_new_n4142_), .B(_abc_15497_new_n4140_), .Y(_abc_15497_new_n4143_));
NAND2X1 NAND2X1_44 ( .A(e_reg_13_), .B(_auto_iopadmap_cc_368_execute_22625_13_), .Y(_abc_15497_new_n1073_));
NAND2X1 NAND2X1_440 ( .A(_abc_15497_new_n4143_), .B(_abc_15497_new_n4106_), .Y(_abc_15497_new_n4150_));
NAND2X1 NAND2X1_441 ( .A(b_reg_25_), .B(c_reg_25_), .Y(_abc_15497_new_n4156_));
NAND2X1 NAND2X1_442 ( .A(_abc_15497_new_n4163_), .B(_abc_15497_new_n4168_), .Y(_abc_15497_new_n4170_));
NAND2X1 NAND2X1_443 ( .A(_abc_15497_new_n4170_), .B(_abc_15497_new_n4169_), .Y(_abc_15497_new_n4171_));
NAND2X1 NAND2X1_444 ( .A(_abc_15497_new_n4153_), .B(_abc_15497_new_n4172_), .Y(_abc_15497_new_n4175_));
NAND2X1 NAND2X1_445 ( .A(_abc_15497_new_n4175_), .B(_abc_15497_new_n4174_), .Y(_abc_15497_new_n4176_));
NAND2X1 NAND2X1_446 ( .A(_abc_15497_new_n4151_), .B(_abc_15497_new_n4176_), .Y(_abc_15497_new_n4178_));
NAND2X1 NAND2X1_447 ( .A(_abc_15497_new_n4178_), .B(_abc_15497_new_n4177_), .Y(_abc_15497_new_n4179_));
NAND2X1 NAND2X1_448 ( .A(_abc_15497_new_n4189_), .B(_abc_15497_new_n4106_), .Y(_abc_15497_new_n4190_));
NAND2X1 NAND2X1_449 ( .A(_abc_15497_new_n4188_), .B(_abc_15497_new_n4190_), .Y(_abc_15497_new_n4191_));
NAND2X1 NAND2X1_45 ( .A(_abc_15497_new_n1075_), .B(_abc_15497_new_n1066_), .Y(_abc_15497_new_n1086_));
NAND2X1 NAND2X1_450 ( .A(c_reg_26_), .B(b_reg_26_), .Y(_abc_15497_new_n4194_));
NAND2X1 NAND2X1_451 ( .A(_abc_15497_new_n866_), .B(_abc_15497_new_n2031_), .Y(_abc_15497_new_n4195_));
NAND2X1 NAND2X1_452 ( .A(_abc_15497_new_n4194_), .B(_abc_15497_new_n4195_), .Y(_abc_15497_new_n4197_));
NAND2X1 NAND2X1_453 ( .A(_abc_15497_new_n4203_), .B(_abc_15497_new_n4199_), .Y(_abc_15497_new_n4204_));
NAND2X1 NAND2X1_454 ( .A(w_25_), .B(_abc_15497_new_n4167_), .Y(_abc_15497_new_n4205_));
NAND2X1 NAND2X1_455 ( .A(w_26_), .B(_abc_15497_new_n4211_), .Y(_abc_15497_new_n4212_));
NAND2X1 NAND2X1_456 ( .A(_abc_15497_new_n4210_), .B(_abc_15497_new_n4212_), .Y(_abc_15497_new_n4213_));
NAND2X1 NAND2X1_457 ( .A(_abc_15497_new_n4224_), .B(_abc_15497_new_n4222_), .Y(_abc_15497_new_n4225_));
NAND2X1 NAND2X1_458 ( .A(_abc_15497_new_n4220_), .B(_abc_15497_new_n4223_), .Y(_abc_15497_new_n4231_));
NAND2X1 NAND2X1_459 ( .A(_abc_15497_new_n4225_), .B(_abc_15497_new_n4191_), .Y(_abc_15497_new_n4232_));
NAND2X1 NAND2X1_46 ( .A(_abc_15497_new_n1083_), .B(_abc_15497_new_n1087_), .Y(_abc_15497_new_n1089_));
NAND2X1 NAND2X1_460 ( .A(c_reg_27_), .B(b_reg_27_), .Y(_abc_15497_new_n4243_));
NAND2X1 NAND2X1_461 ( .A(_abc_15497_new_n4239_), .B(_abc_15497_new_n4240_), .Y(_abc_15497_new_n4244_));
NAND2X1 NAND2X1_462 ( .A(_abc_15497_new_n4243_), .B(_abc_15497_new_n4244_), .Y(_abc_15497_new_n4245_));
NAND2X1 NAND2X1_463 ( .A(_abc_15497_new_n4250_), .B(_abc_15497_new_n4255_), .Y(_abc_15497_new_n4257_));
NAND2X1 NAND2X1_464 ( .A(_abc_15497_new_n4257_), .B(_abc_15497_new_n4256_), .Y(_abc_15497_new_n4258_));
NAND2X1 NAND2X1_465 ( .A(_abc_15497_new_n4182_), .B(_abc_15497_new_n4143_), .Y(_abc_15497_new_n4269_));
NAND2X1 NAND2X1_466 ( .A(_abc_15497_new_n4263_), .B(_abc_15497_new_n4225_), .Y(_abc_15497_new_n4270_));
NAND2X1 NAND2X1_467 ( .A(_abc_15497_new_n4276_), .B(_abc_15497_new_n4259_), .Y(_abc_15497_new_n4277_));
NAND2X1 NAND2X1_468 ( .A(c_reg_28_), .B(b_reg_28_), .Y(_abc_15497_new_n4280_));
NAND2X1 NAND2X1_469 ( .A(_abc_15497_new_n4295_), .B(_abc_15497_new_n4291_), .Y(_abc_15497_new_n4297_));
NAND2X1 NAND2X1_47 ( .A(digest_update_bF_buf6), .B(_abc_15497_new_n1089_), .Y(_abc_15497_new_n1090_));
NAND2X1 NAND2X1_470 ( .A(_abc_15497_new_n4297_), .B(_abc_15497_new_n4296_), .Y(_abc_15497_new_n4298_));
NAND2X1 NAND2X1_471 ( .A(_abc_15497_new_n3397_), .B(_abc_15497_new_n3341_), .Y(_abc_15497_new_n4306_));
NAND2X1 NAND2X1_472 ( .A(_abc_15497_new_n4307_), .B(_abc_15497_new_n4310_), .Y(_abc_15497_new_n4311_));
NAND2X1 NAND2X1_473 ( .A(_abc_15497_new_n3986_), .B(_abc_15497_new_n4097_), .Y(_abc_15497_new_n4313_));
NAND2X1 NAND2X1_474 ( .A(_abc_15497_new_n4304_), .B(_abc_15497_new_n4319_), .Y(_abc_15497_new_n4320_));
NAND2X1 NAND2X1_475 ( .A(_abc_15497_new_n4332_), .B(_abc_15497_new_n2743__bF_buf3), .Y(_abc_15497_new_n4333_));
NAND2X1 NAND2X1_476 ( .A(_abc_15497_new_n1622_), .B(_abc_15497_new_n4335_), .Y(_abc_15497_new_n4336_));
NAND2X1 NAND2X1_477 ( .A(_abc_15497_new_n4342_), .B(_abc_15497_new_n4349_), .Y(_abc_15497_new_n4351_));
NAND2X1 NAND2X1_478 ( .A(_abc_15497_new_n4351_), .B(_abc_15497_new_n4350_), .Y(_abc_15497_new_n4352_));
NAND2X1 NAND2X1_479 ( .A(_abc_15497_new_n4354_), .B(_abc_15497_new_n4355_), .Y(_abc_15497_new_n4356_));
NAND2X1 NAND2X1_48 ( .A(e_reg_15_), .B(_auto_iopadmap_cc_368_execute_22625_15_), .Y(_abc_15497_new_n1095_));
NAND2X1 NAND2X1_480 ( .A(_abc_15497_new_n4327_), .B(_abc_15497_new_n4356_), .Y(_abc_15497_new_n4357_));
NAND2X1 NAND2X1_481 ( .A(_abc_15497_new_n4318_), .B(_abc_15497_new_n4359_), .Y(_abc_15497_new_n4365_));
NAND2X1 NAND2X1_482 ( .A(_abc_15497_new_n4374_), .B(_abc_15497_new_n2743__bF_buf1), .Y(_abc_15497_new_n4375_));
NAND2X1 NAND2X1_483 ( .A(_abc_15497_new_n2630_), .B(_abc_15497_new_n4377_), .Y(_abc_15497_new_n4378_));
NAND2X1 NAND2X1_484 ( .A(w_29_), .B(_abc_15497_new_n4346_), .Y(_abc_15497_new_n4385_));
NAND2X1 NAND2X1_485 ( .A(w_30_), .B(_abc_15497_new_n4390_), .Y(_abc_15497_new_n4392_));
NAND2X1 NAND2X1_486 ( .A(_abc_15497_new_n4384_), .B(_abc_15497_new_n4395_), .Y(_abc_15497_new_n4397_));
NAND2X1 NAND2X1_487 ( .A(_abc_15497_new_n4397_), .B(_abc_15497_new_n4396_), .Y(_abc_15497_new_n4398_));
NAND2X1 NAND2X1_488 ( .A(_abc_15497_new_n4386_), .B(_abc_15497_new_n4393_), .Y(_abc_15497_new_n4414_));
NAND2X1 NAND2X1_489 ( .A(_abc_15497_new_n4416_), .B(_abc_15497_new_n2743__bF_buf0), .Y(_abc_15497_new_n4417_));
NAND2X1 NAND2X1_49 ( .A(_abc_15497_new_n1097_), .B(_abc_15497_new_n1083_), .Y(_abc_15497_new_n1103_));
NAND2X1 NAND2X1_490 ( .A(_abc_15497_new_n3392_), .B(_abc_15497_new_n4444_), .Y(_abc_15497_new_n4445_));
NAND2X1 NAND2X1_491 ( .A(round_ctr_inc_bF_buf9), .B(_abc_15497_new_n4443_), .Y(_abc_15497_new_n4453_));
NAND2X1 NAND2X1_492 ( .A(round_ctr_reg_1_), .B(_abc_15497_new_n1663__bF_buf0), .Y(_abc_15497_new_n4455_));
NAND2X1 NAND2X1_493 ( .A(round_ctr_reg_2_), .B(_abc_15497_new_n4444_), .Y(_abc_15497_new_n4459_));
NAND2X1 NAND2X1_494 ( .A(round_ctr_reg_4_), .B(_abc_15497_new_n4464_), .Y(_abc_15497_new_n4468_));
NAND2X1 NAND2X1_495 ( .A(_abc_15497_new_n4497_), .B(_abc_15497_new_n4496_), .Y(_0H2_reg_31_0__5_));
NAND2X1 NAND2X1_496 ( .A(_abc_15497_new_n764_), .B(_abc_15497_new_n780_), .Y(_abc_15497_new_n4500_));
NAND2X1 NAND2X1_497 ( .A(_abc_15497_new_n756_), .B(_abc_15497_new_n782_), .Y(_abc_15497_new_n4503_));
NAND2X1 NAND2X1_498 ( .A(_abc_15497_new_n4502_), .B(_abc_15497_new_n4503_), .Y(_abc_15497_new_n4504_));
NAND2X1 NAND2X1_499 ( .A(_abc_15497_new_n735_), .B(_abc_15497_new_n790_), .Y(_abc_15497_new_n4522_));
NAND2X1 NAND2X1_5 ( .A(c_reg_3_), .B(_auto_iopadmap_cc_368_execute_22625_67_), .Y(_abc_15497_new_n765_));
NAND2X1 NAND2X1_50 ( .A(_abc_15497_new_n1104_), .B(_abc_15497_new_n1108_), .Y(_abc_15497_new_n1109_));
NAND2X1 NAND2X1_500 ( .A(_abc_15497_new_n4521_), .B(_abc_15497_new_n4522_), .Y(_abc_15497_new_n4523_));
NAND2X1 NAND2X1_501 ( .A(_abc_15497_new_n706_), .B(_abc_15497_new_n4539_), .Y(_abc_15497_new_n4541_));
NAND2X1 NAND2X1_502 ( .A(digest_update_bF_buf3), .B(_abc_15497_new_n4541_), .Y(_abc_15497_new_n4542_));
NAND2X1 NAND2X1_503 ( .A(_abc_15497_new_n4575_), .B(_abc_15497_new_n4574_), .Y(_0H2_reg_31_0__21_));
NAND2X1 NAND2X1_504 ( .A(w_mem_inst_w_ctr_reg_0_), .B(w_mem_inst__abc_19396_new_n1592_), .Y(w_mem_inst__abc_19396_new_n1593_));
NAND2X1 NAND2X1_505 ( .A(w_mem_inst_w_ctr_reg_2_), .B(w_mem_inst__abc_19396_new_n1595_), .Y(w_mem_inst__abc_19396_new_n1596_));
NAND2X1 NAND2X1_506 ( .A(w_mem_inst__abc_19396_new_n1594__bF_buf7), .B(w_mem_inst__abc_19396_new_n1597_), .Y(w_mem_inst__abc_19396_new_n1598_));
NAND2X1 NAND2X1_507 ( .A(w_mem_inst_w_ctr_reg_3_), .B(w_mem_inst__abc_19396_new_n1602_), .Y(w_mem_inst__abc_19396_new_n1603_));
NAND2X1 NAND2X1_508 ( .A(w_mem_inst_w_ctr_reg_1_), .B(w_mem_inst_w_ctr_reg_0_), .Y(w_mem_inst__abc_19396_new_n1605_));
NAND2X1 NAND2X1_509 ( .A(w_mem_inst_w_mem_11__0_), .B(w_mem_inst__abc_19396_new_n1606__bF_buf4), .Y(w_mem_inst__abc_19396_new_n1607_));
NAND2X1 NAND2X1_51 ( .A(_abc_15497_new_n1114_), .B(_abc_15497_new_n1110_), .Y(_abc_15497_new_n1116_));
NAND2X1 NAND2X1_510 ( .A(w_mem_inst__abc_19396_new_n1610_), .B(w_mem_inst__abc_19396_new_n1597_), .Y(w_mem_inst__abc_19396_new_n1611_));
NAND2X1 NAND2X1_511 ( .A(w_mem_inst_w_ctr_reg_3_), .B(w_mem_inst_w_ctr_reg_2_), .Y(w_mem_inst__abc_19396_new_n1612_));
NAND2X1 NAND2X1_512 ( .A(w_mem_inst_w_mem_15__0_), .B(w_mem_inst__abc_19396_new_n1613__bF_buf4), .Y(w_mem_inst__abc_19396_new_n1614_));
NAND2X1 NAND2X1_513 ( .A(w_mem_inst_w_mem_0__0_), .B(w_mem_inst__abc_19396_new_n1621__bF_buf4), .Y(w_mem_inst__abc_19396_new_n1622_));
NAND2X1 NAND2X1_514 ( .A(w_mem_inst_w_ctr_reg_1_), .B(w_mem_inst__abc_19396_new_n1626_), .Y(w_mem_inst__abc_19396_new_n1627_));
NAND2X1 NAND2X1_515 ( .A(w_mem_inst__abc_19396_new_n1632_), .B(w_mem_inst__abc_19396_new_n1629_), .Y(w_mem_inst__abc_19396_new_n1633_));
NAND2X1 NAND2X1_516 ( .A(w_mem_inst_w_mem_11__1_), .B(w_mem_inst__abc_19396_new_n1606__bF_buf3), .Y(w_mem_inst__abc_19396_new_n1649_));
NAND2X1 NAND2X1_517 ( .A(w_mem_inst_w_mem_15__1_), .B(w_mem_inst__abc_19396_new_n1613__bF_buf3), .Y(w_mem_inst__abc_19396_new_n1652_));
NAND2X1 NAND2X1_518 ( .A(w_mem_inst_w_mem_0__1_), .B(w_mem_inst__abc_19396_new_n1621__bF_buf3), .Y(w_mem_inst__abc_19396_new_n1656_));
NAND2X1 NAND2X1_519 ( .A(w_mem_inst__abc_19396_new_n1660_), .B(w_mem_inst__abc_19396_new_n1659_), .Y(w_mem_inst__abc_19396_new_n1661_));
NAND2X1 NAND2X1_52 ( .A(digest_update_bF_buf5), .B(_abc_15497_new_n1116_), .Y(_abc_15497_new_n1117_));
NAND2X1 NAND2X1_520 ( .A(w_mem_inst_w_mem_11__2_), .B(w_mem_inst__abc_19396_new_n1606__bF_buf2), .Y(w_mem_inst__abc_19396_new_n1674_));
NAND2X1 NAND2X1_521 ( .A(w_mem_inst_w_mem_15__2_), .B(w_mem_inst__abc_19396_new_n1613__bF_buf2), .Y(w_mem_inst__abc_19396_new_n1677_));
NAND2X1 NAND2X1_522 ( .A(w_mem_inst_w_mem_0__2_), .B(w_mem_inst__abc_19396_new_n1621__bF_buf2), .Y(w_mem_inst__abc_19396_new_n1681_));
NAND2X1 NAND2X1_523 ( .A(w_mem_inst__abc_19396_new_n1685_), .B(w_mem_inst__abc_19396_new_n1684_), .Y(w_mem_inst__abc_19396_new_n1686_));
NAND2X1 NAND2X1_524 ( .A(w_mem_inst_w_mem_11__3_), .B(w_mem_inst__abc_19396_new_n1606__bF_buf1), .Y(w_mem_inst__abc_19396_new_n1699_));
NAND2X1 NAND2X1_525 ( .A(w_mem_inst_w_mem_15__3_), .B(w_mem_inst__abc_19396_new_n1613__bF_buf1), .Y(w_mem_inst__abc_19396_new_n1702_));
NAND2X1 NAND2X1_526 ( .A(w_mem_inst_w_mem_0__3_), .B(w_mem_inst__abc_19396_new_n1621__bF_buf1), .Y(w_mem_inst__abc_19396_new_n1706_));
NAND2X1 NAND2X1_527 ( .A(w_mem_inst__abc_19396_new_n1710_), .B(w_mem_inst__abc_19396_new_n1709_), .Y(w_mem_inst__abc_19396_new_n1711_));
NAND2X1 NAND2X1_528 ( .A(w_mem_inst_w_mem_11__4_), .B(w_mem_inst__abc_19396_new_n1606__bF_buf0), .Y(w_mem_inst__abc_19396_new_n1724_));
NAND2X1 NAND2X1_529 ( .A(w_mem_inst_w_mem_15__4_), .B(w_mem_inst__abc_19396_new_n1613__bF_buf0), .Y(w_mem_inst__abc_19396_new_n1727_));
NAND2X1 NAND2X1_53 ( .A(_abc_15497_new_n1132_), .B(_abc_15497_new_n1148_), .Y(_abc_15497_new_n1153_));
NAND2X1 NAND2X1_530 ( .A(w_mem_inst_w_mem_0__4_), .B(w_mem_inst__abc_19396_new_n1621__bF_buf0), .Y(w_mem_inst__abc_19396_new_n1731_));
NAND2X1 NAND2X1_531 ( .A(w_mem_inst__abc_19396_new_n1735_), .B(w_mem_inst__abc_19396_new_n1734_), .Y(w_mem_inst__abc_19396_new_n1736_));
NAND2X1 NAND2X1_532 ( .A(w_mem_inst_w_mem_11__5_), .B(w_mem_inst__abc_19396_new_n1606__bF_buf4), .Y(w_mem_inst__abc_19396_new_n1749_));
NAND2X1 NAND2X1_533 ( .A(w_mem_inst_w_mem_15__5_), .B(w_mem_inst__abc_19396_new_n1613__bF_buf4), .Y(w_mem_inst__abc_19396_new_n1752_));
NAND2X1 NAND2X1_534 ( .A(w_mem_inst_w_mem_0__5_), .B(w_mem_inst__abc_19396_new_n1621__bF_buf4), .Y(w_mem_inst__abc_19396_new_n1756_));
NAND2X1 NAND2X1_535 ( .A(w_mem_inst__abc_19396_new_n1760_), .B(w_mem_inst__abc_19396_new_n1759_), .Y(w_mem_inst__abc_19396_new_n1761_));
NAND2X1 NAND2X1_536 ( .A(w_mem_inst_w_mem_11__6_), .B(w_mem_inst__abc_19396_new_n1606__bF_buf3), .Y(w_mem_inst__abc_19396_new_n1774_));
NAND2X1 NAND2X1_537 ( .A(w_mem_inst_w_mem_15__6_), .B(w_mem_inst__abc_19396_new_n1613__bF_buf3), .Y(w_mem_inst__abc_19396_new_n1777_));
NAND2X1 NAND2X1_538 ( .A(w_mem_inst_w_mem_0__6_), .B(w_mem_inst__abc_19396_new_n1621__bF_buf3), .Y(w_mem_inst__abc_19396_new_n1781_));
NAND2X1 NAND2X1_539 ( .A(w_mem_inst__abc_19396_new_n1785_), .B(w_mem_inst__abc_19396_new_n1784_), .Y(w_mem_inst__abc_19396_new_n1786_));
NAND2X1 NAND2X1_54 ( .A(_abc_15497_new_n1114_), .B(_abc_15497_new_n1124_), .Y(_abc_15497_new_n1156_));
NAND2X1 NAND2X1_540 ( .A(w_mem_inst_w_mem_11__7_), .B(w_mem_inst__abc_19396_new_n1606__bF_buf2), .Y(w_mem_inst__abc_19396_new_n1799_));
NAND2X1 NAND2X1_541 ( .A(w_mem_inst_w_mem_15__7_), .B(w_mem_inst__abc_19396_new_n1613__bF_buf2), .Y(w_mem_inst__abc_19396_new_n1802_));
NAND2X1 NAND2X1_542 ( .A(w_mem_inst_w_mem_0__7_), .B(w_mem_inst__abc_19396_new_n1621__bF_buf2), .Y(w_mem_inst__abc_19396_new_n1806_));
NAND2X1 NAND2X1_543 ( .A(w_mem_inst__abc_19396_new_n1810_), .B(w_mem_inst__abc_19396_new_n1809_), .Y(w_mem_inst__abc_19396_new_n1811_));
NAND2X1 NAND2X1_544 ( .A(w_mem_inst_w_mem_11__8_), .B(w_mem_inst__abc_19396_new_n1606__bF_buf1), .Y(w_mem_inst__abc_19396_new_n1824_));
NAND2X1 NAND2X1_545 ( .A(w_mem_inst_w_mem_15__8_), .B(w_mem_inst__abc_19396_new_n1613__bF_buf1), .Y(w_mem_inst__abc_19396_new_n1827_));
NAND2X1 NAND2X1_546 ( .A(w_mem_inst_w_mem_0__8_), .B(w_mem_inst__abc_19396_new_n1621__bF_buf1), .Y(w_mem_inst__abc_19396_new_n1831_));
NAND2X1 NAND2X1_547 ( .A(w_mem_inst__abc_19396_new_n1835_), .B(w_mem_inst__abc_19396_new_n1834_), .Y(w_mem_inst__abc_19396_new_n1836_));
NAND2X1 NAND2X1_548 ( .A(w_mem_inst_w_mem_11__9_), .B(w_mem_inst__abc_19396_new_n1606__bF_buf0), .Y(w_mem_inst__abc_19396_new_n1849_));
NAND2X1 NAND2X1_549 ( .A(w_mem_inst_w_mem_15__9_), .B(w_mem_inst__abc_19396_new_n1613__bF_buf0), .Y(w_mem_inst__abc_19396_new_n1852_));
NAND2X1 NAND2X1_55 ( .A(_abc_15497_new_n1155_), .B(_abc_15497_new_n1159_), .Y(_abc_15497_new_n1160_));
NAND2X1 NAND2X1_550 ( .A(w_mem_inst_w_mem_0__9_), .B(w_mem_inst__abc_19396_new_n1621__bF_buf0), .Y(w_mem_inst__abc_19396_new_n1856_));
NAND2X1 NAND2X1_551 ( .A(w_mem_inst__abc_19396_new_n1860_), .B(w_mem_inst__abc_19396_new_n1859_), .Y(w_mem_inst__abc_19396_new_n1861_));
NAND2X1 NAND2X1_552 ( .A(w_mem_inst_w_mem_11__10_), .B(w_mem_inst__abc_19396_new_n1606__bF_buf4), .Y(w_mem_inst__abc_19396_new_n1874_));
NAND2X1 NAND2X1_553 ( .A(w_mem_inst_w_mem_15__10_), .B(w_mem_inst__abc_19396_new_n1613__bF_buf4), .Y(w_mem_inst__abc_19396_new_n1877_));
NAND2X1 NAND2X1_554 ( .A(w_mem_inst_w_mem_0__10_), .B(w_mem_inst__abc_19396_new_n1621__bF_buf4), .Y(w_mem_inst__abc_19396_new_n1881_));
NAND2X1 NAND2X1_555 ( .A(w_mem_inst__abc_19396_new_n1885_), .B(w_mem_inst__abc_19396_new_n1884_), .Y(w_mem_inst__abc_19396_new_n1886_));
NAND2X1 NAND2X1_556 ( .A(w_mem_inst_w_mem_11__11_), .B(w_mem_inst__abc_19396_new_n1606__bF_buf3), .Y(w_mem_inst__abc_19396_new_n1899_));
NAND2X1 NAND2X1_557 ( .A(w_mem_inst_w_mem_15__11_), .B(w_mem_inst__abc_19396_new_n1613__bF_buf3), .Y(w_mem_inst__abc_19396_new_n1902_));
NAND2X1 NAND2X1_558 ( .A(w_mem_inst_w_mem_0__11_), .B(w_mem_inst__abc_19396_new_n1621__bF_buf3), .Y(w_mem_inst__abc_19396_new_n1906_));
NAND2X1 NAND2X1_559 ( .A(w_mem_inst__abc_19396_new_n1910_), .B(w_mem_inst__abc_19396_new_n1909_), .Y(w_mem_inst__abc_19396_new_n1911_));
NAND2X1 NAND2X1_56 ( .A(digest_update_bF_buf3), .B(_abc_15497_new_n1167_), .Y(_abc_15497_new_n1168_));
NAND2X1 NAND2X1_560 ( .A(w_mem_inst_w_mem_11__12_), .B(w_mem_inst__abc_19396_new_n1606__bF_buf2), .Y(w_mem_inst__abc_19396_new_n1924_));
NAND2X1 NAND2X1_561 ( .A(w_mem_inst_w_mem_15__12_), .B(w_mem_inst__abc_19396_new_n1613__bF_buf2), .Y(w_mem_inst__abc_19396_new_n1927_));
NAND2X1 NAND2X1_562 ( .A(w_mem_inst_w_mem_0__12_), .B(w_mem_inst__abc_19396_new_n1621__bF_buf2), .Y(w_mem_inst__abc_19396_new_n1931_));
NAND2X1 NAND2X1_563 ( .A(w_mem_inst__abc_19396_new_n1935_), .B(w_mem_inst__abc_19396_new_n1934_), .Y(w_mem_inst__abc_19396_new_n1936_));
NAND2X1 NAND2X1_564 ( .A(w_mem_inst_w_mem_11__13_), .B(w_mem_inst__abc_19396_new_n1606__bF_buf1), .Y(w_mem_inst__abc_19396_new_n1949_));
NAND2X1 NAND2X1_565 ( .A(w_mem_inst_w_mem_15__13_), .B(w_mem_inst__abc_19396_new_n1613__bF_buf1), .Y(w_mem_inst__abc_19396_new_n1952_));
NAND2X1 NAND2X1_566 ( .A(w_mem_inst_w_mem_0__13_), .B(w_mem_inst__abc_19396_new_n1621__bF_buf1), .Y(w_mem_inst__abc_19396_new_n1956_));
NAND2X1 NAND2X1_567 ( .A(w_mem_inst__abc_19396_new_n1960_), .B(w_mem_inst__abc_19396_new_n1959_), .Y(w_mem_inst__abc_19396_new_n1961_));
NAND2X1 NAND2X1_568 ( .A(w_mem_inst_w_mem_11__14_), .B(w_mem_inst__abc_19396_new_n1606__bF_buf0), .Y(w_mem_inst__abc_19396_new_n1974_));
NAND2X1 NAND2X1_569 ( .A(w_mem_inst_w_mem_15__14_), .B(w_mem_inst__abc_19396_new_n1613__bF_buf0), .Y(w_mem_inst__abc_19396_new_n1977_));
NAND2X1 NAND2X1_57 ( .A(_abc_15497_new_n1165_), .B(_abc_15497_new_n1175_), .Y(_abc_15497_new_n1179_));
NAND2X1 NAND2X1_570 ( .A(w_mem_inst_w_mem_0__14_), .B(w_mem_inst__abc_19396_new_n1621__bF_buf0), .Y(w_mem_inst__abc_19396_new_n1981_));
NAND2X1 NAND2X1_571 ( .A(w_mem_inst__abc_19396_new_n1985_), .B(w_mem_inst__abc_19396_new_n1984_), .Y(w_mem_inst__abc_19396_new_n1986_));
NAND2X1 NAND2X1_572 ( .A(w_mem_inst_w_mem_11__15_), .B(w_mem_inst__abc_19396_new_n1606__bF_buf4), .Y(w_mem_inst__abc_19396_new_n1999_));
NAND2X1 NAND2X1_573 ( .A(w_mem_inst_w_mem_15__15_), .B(w_mem_inst__abc_19396_new_n1613__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2002_));
NAND2X1 NAND2X1_574 ( .A(w_mem_inst_w_mem_0__15_), .B(w_mem_inst__abc_19396_new_n1621__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2006_));
NAND2X1 NAND2X1_575 ( .A(w_mem_inst__abc_19396_new_n2010_), .B(w_mem_inst__abc_19396_new_n2009_), .Y(w_mem_inst__abc_19396_new_n2011_));
NAND2X1 NAND2X1_576 ( .A(w_mem_inst_w_mem_11__16_), .B(w_mem_inst__abc_19396_new_n1606__bF_buf3), .Y(w_mem_inst__abc_19396_new_n2024_));
NAND2X1 NAND2X1_577 ( .A(w_mem_inst_w_mem_15__16_), .B(w_mem_inst__abc_19396_new_n1613__bF_buf3), .Y(w_mem_inst__abc_19396_new_n2027_));
NAND2X1 NAND2X1_578 ( .A(w_mem_inst_w_mem_0__16_), .B(w_mem_inst__abc_19396_new_n1621__bF_buf3), .Y(w_mem_inst__abc_19396_new_n2031_));
NAND2X1 NAND2X1_579 ( .A(w_mem_inst__abc_19396_new_n2035_), .B(w_mem_inst__abc_19396_new_n2034_), .Y(w_mem_inst__abc_19396_new_n2036_));
NAND2X1 NAND2X1_58 ( .A(_abc_15497_new_n1164_), .B(_abc_15497_new_n1175_), .Y(_abc_15497_new_n1181_));
NAND2X1 NAND2X1_580 ( .A(w_mem_inst_w_mem_11__17_), .B(w_mem_inst__abc_19396_new_n1606__bF_buf2), .Y(w_mem_inst__abc_19396_new_n2049_));
NAND2X1 NAND2X1_581 ( .A(w_mem_inst_w_mem_15__17_), .B(w_mem_inst__abc_19396_new_n1613__bF_buf2), .Y(w_mem_inst__abc_19396_new_n2052_));
NAND2X1 NAND2X1_582 ( .A(w_mem_inst_w_mem_0__17_), .B(w_mem_inst__abc_19396_new_n1621__bF_buf2), .Y(w_mem_inst__abc_19396_new_n2056_));
NAND2X1 NAND2X1_583 ( .A(w_mem_inst__abc_19396_new_n2060_), .B(w_mem_inst__abc_19396_new_n2059_), .Y(w_mem_inst__abc_19396_new_n2061_));
NAND2X1 NAND2X1_584 ( .A(w_mem_inst_w_mem_11__18_), .B(w_mem_inst__abc_19396_new_n1606__bF_buf1), .Y(w_mem_inst__abc_19396_new_n2074_));
NAND2X1 NAND2X1_585 ( .A(w_mem_inst_w_mem_15__18_), .B(w_mem_inst__abc_19396_new_n1613__bF_buf1), .Y(w_mem_inst__abc_19396_new_n2077_));
NAND2X1 NAND2X1_586 ( .A(w_mem_inst_w_mem_0__18_), .B(w_mem_inst__abc_19396_new_n1621__bF_buf1), .Y(w_mem_inst__abc_19396_new_n2081_));
NAND2X1 NAND2X1_587 ( .A(w_mem_inst__abc_19396_new_n2085_), .B(w_mem_inst__abc_19396_new_n2084_), .Y(w_mem_inst__abc_19396_new_n2086_));
NAND2X1 NAND2X1_588 ( .A(w_mem_inst_w_mem_11__19_), .B(w_mem_inst__abc_19396_new_n1606__bF_buf0), .Y(w_mem_inst__abc_19396_new_n2099_));
NAND2X1 NAND2X1_589 ( .A(w_mem_inst_w_mem_15__19_), .B(w_mem_inst__abc_19396_new_n1613__bF_buf0), .Y(w_mem_inst__abc_19396_new_n2102_));
NAND2X1 NAND2X1_59 ( .A(e_reg_22_), .B(_auto_iopadmap_cc_368_execute_22625_22_), .Y(_abc_15497_new_n1185_));
NAND2X1 NAND2X1_590 ( .A(w_mem_inst_w_mem_0__19_), .B(w_mem_inst__abc_19396_new_n1621__bF_buf0), .Y(w_mem_inst__abc_19396_new_n2106_));
NAND2X1 NAND2X1_591 ( .A(w_mem_inst__abc_19396_new_n2110_), .B(w_mem_inst__abc_19396_new_n2109_), .Y(w_mem_inst__abc_19396_new_n2111_));
NAND2X1 NAND2X1_592 ( .A(w_mem_inst_w_mem_11__20_), .B(w_mem_inst__abc_19396_new_n1606__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2124_));
NAND2X1 NAND2X1_593 ( .A(w_mem_inst_w_mem_15__20_), .B(w_mem_inst__abc_19396_new_n1613__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2127_));
NAND2X1 NAND2X1_594 ( .A(w_mem_inst_w_mem_0__20_), .B(w_mem_inst__abc_19396_new_n1621__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2131_));
NAND2X1 NAND2X1_595 ( .A(w_mem_inst__abc_19396_new_n2135_), .B(w_mem_inst__abc_19396_new_n2134_), .Y(w_mem_inst__abc_19396_new_n2136_));
NAND2X1 NAND2X1_596 ( .A(w_mem_inst_w_mem_11__21_), .B(w_mem_inst__abc_19396_new_n1606__bF_buf3), .Y(w_mem_inst__abc_19396_new_n2149_));
NAND2X1 NAND2X1_597 ( .A(w_mem_inst_w_mem_15__21_), .B(w_mem_inst__abc_19396_new_n1613__bF_buf3), .Y(w_mem_inst__abc_19396_new_n2152_));
NAND2X1 NAND2X1_598 ( .A(w_mem_inst_w_mem_0__21_), .B(w_mem_inst__abc_19396_new_n1621__bF_buf3), .Y(w_mem_inst__abc_19396_new_n2156_));
NAND2X1 NAND2X1_599 ( .A(w_mem_inst__abc_19396_new_n2160_), .B(w_mem_inst__abc_19396_new_n2159_), .Y(w_mem_inst__abc_19396_new_n2161_));
NAND2X1 NAND2X1_6 ( .A(c_reg_1_), .B(_auto_iopadmap_cc_368_execute_22625_65_), .Y(_abc_15497_new_n768_));
NAND2X1 NAND2X1_60 ( .A(e_reg_23_), .B(_auto_iopadmap_cc_368_execute_22625_23_), .Y(_abc_15497_new_n1195_));
NAND2X1 NAND2X1_600 ( .A(w_mem_inst_w_mem_11__22_), .B(w_mem_inst__abc_19396_new_n1606__bF_buf2), .Y(w_mem_inst__abc_19396_new_n2174_));
NAND2X1 NAND2X1_601 ( .A(w_mem_inst_w_mem_15__22_), .B(w_mem_inst__abc_19396_new_n1613__bF_buf2), .Y(w_mem_inst__abc_19396_new_n2177_));
NAND2X1 NAND2X1_602 ( .A(w_mem_inst_w_mem_0__22_), .B(w_mem_inst__abc_19396_new_n1621__bF_buf2), .Y(w_mem_inst__abc_19396_new_n2181_));
NAND2X1 NAND2X1_603 ( .A(w_mem_inst__abc_19396_new_n2185_), .B(w_mem_inst__abc_19396_new_n2184_), .Y(w_mem_inst__abc_19396_new_n2186_));
NAND2X1 NAND2X1_604 ( .A(w_mem_inst_w_mem_11__23_), .B(w_mem_inst__abc_19396_new_n1606__bF_buf1), .Y(w_mem_inst__abc_19396_new_n2199_));
NAND2X1 NAND2X1_605 ( .A(w_mem_inst_w_mem_15__23_), .B(w_mem_inst__abc_19396_new_n1613__bF_buf1), .Y(w_mem_inst__abc_19396_new_n2202_));
NAND2X1 NAND2X1_606 ( .A(w_mem_inst_w_mem_0__23_), .B(w_mem_inst__abc_19396_new_n1621__bF_buf1), .Y(w_mem_inst__abc_19396_new_n2206_));
NAND2X1 NAND2X1_607 ( .A(w_mem_inst__abc_19396_new_n2210_), .B(w_mem_inst__abc_19396_new_n2209_), .Y(w_mem_inst__abc_19396_new_n2211_));
NAND2X1 NAND2X1_608 ( .A(w_mem_inst_w_mem_11__24_), .B(w_mem_inst__abc_19396_new_n1606__bF_buf0), .Y(w_mem_inst__abc_19396_new_n2224_));
NAND2X1 NAND2X1_609 ( .A(w_mem_inst_w_mem_15__24_), .B(w_mem_inst__abc_19396_new_n1613__bF_buf0), .Y(w_mem_inst__abc_19396_new_n2227_));
NAND2X1 NAND2X1_61 ( .A(_abc_15497_new_n1187_), .B(_abc_15497_new_n1197_), .Y(_abc_15497_new_n1201_));
NAND2X1 NAND2X1_610 ( .A(w_mem_inst_w_mem_0__24_), .B(w_mem_inst__abc_19396_new_n1621__bF_buf0), .Y(w_mem_inst__abc_19396_new_n2231_));
NAND2X1 NAND2X1_611 ( .A(w_mem_inst__abc_19396_new_n2235_), .B(w_mem_inst__abc_19396_new_n2234_), .Y(w_mem_inst__abc_19396_new_n2236_));
NAND2X1 NAND2X1_612 ( .A(w_mem_inst_w_mem_11__25_), .B(w_mem_inst__abc_19396_new_n1606__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2249_));
NAND2X1 NAND2X1_613 ( .A(w_mem_inst_w_mem_15__25_), .B(w_mem_inst__abc_19396_new_n1613__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2252_));
NAND2X1 NAND2X1_614 ( .A(w_mem_inst_w_mem_0__25_), .B(w_mem_inst__abc_19396_new_n1621__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2256_));
NAND2X1 NAND2X1_615 ( .A(w_mem_inst__abc_19396_new_n2260_), .B(w_mem_inst__abc_19396_new_n2259_), .Y(w_mem_inst__abc_19396_new_n2261_));
NAND2X1 NAND2X1_616 ( .A(w_mem_inst_w_mem_11__26_), .B(w_mem_inst__abc_19396_new_n1606__bF_buf3), .Y(w_mem_inst__abc_19396_new_n2274_));
NAND2X1 NAND2X1_617 ( .A(w_mem_inst_w_mem_15__26_), .B(w_mem_inst__abc_19396_new_n1613__bF_buf3), .Y(w_mem_inst__abc_19396_new_n2277_));
NAND2X1 NAND2X1_618 ( .A(w_mem_inst_w_mem_0__26_), .B(w_mem_inst__abc_19396_new_n1621__bF_buf3), .Y(w_mem_inst__abc_19396_new_n2281_));
NAND2X1 NAND2X1_619 ( .A(w_mem_inst__abc_19396_new_n2285_), .B(w_mem_inst__abc_19396_new_n2284_), .Y(w_mem_inst__abc_19396_new_n2286_));
NAND2X1 NAND2X1_62 ( .A(e_reg_25_), .B(_auto_iopadmap_cc_368_execute_22625_25_), .Y(_abc_15497_new_n1225_));
NAND2X1 NAND2X1_620 ( .A(w_mem_inst_w_mem_11__27_), .B(w_mem_inst__abc_19396_new_n1606__bF_buf2), .Y(w_mem_inst__abc_19396_new_n2299_));
NAND2X1 NAND2X1_621 ( .A(w_mem_inst_w_mem_15__27_), .B(w_mem_inst__abc_19396_new_n1613__bF_buf2), .Y(w_mem_inst__abc_19396_new_n2302_));
NAND2X1 NAND2X1_622 ( .A(w_mem_inst_w_mem_0__27_), .B(w_mem_inst__abc_19396_new_n1621__bF_buf2), .Y(w_mem_inst__abc_19396_new_n2306_));
NAND2X1 NAND2X1_623 ( .A(w_mem_inst__abc_19396_new_n2310_), .B(w_mem_inst__abc_19396_new_n2309_), .Y(w_mem_inst__abc_19396_new_n2311_));
NAND2X1 NAND2X1_624 ( .A(w_mem_inst_w_mem_11__28_), .B(w_mem_inst__abc_19396_new_n1606__bF_buf1), .Y(w_mem_inst__abc_19396_new_n2324_));
NAND2X1 NAND2X1_625 ( .A(w_mem_inst_w_mem_15__28_), .B(w_mem_inst__abc_19396_new_n1613__bF_buf1), .Y(w_mem_inst__abc_19396_new_n2327_));
NAND2X1 NAND2X1_626 ( .A(w_mem_inst_w_mem_0__28_), .B(w_mem_inst__abc_19396_new_n1621__bF_buf1), .Y(w_mem_inst__abc_19396_new_n2331_));
NAND2X1 NAND2X1_627 ( .A(w_mem_inst__abc_19396_new_n2335_), .B(w_mem_inst__abc_19396_new_n2334_), .Y(w_mem_inst__abc_19396_new_n2336_));
NAND2X1 NAND2X1_628 ( .A(w_mem_inst_w_mem_11__29_), .B(w_mem_inst__abc_19396_new_n1606__bF_buf0), .Y(w_mem_inst__abc_19396_new_n2349_));
NAND2X1 NAND2X1_629 ( .A(w_mem_inst_w_mem_15__29_), .B(w_mem_inst__abc_19396_new_n1613__bF_buf0), .Y(w_mem_inst__abc_19396_new_n2352_));
NAND2X1 NAND2X1_63 ( .A(_abc_15497_new_n1240_), .B(_abc_15497_new_n1252_), .Y(_abc_15497_new_n1261_));
NAND2X1 NAND2X1_630 ( .A(w_mem_inst_w_mem_0__29_), .B(w_mem_inst__abc_19396_new_n1621__bF_buf0), .Y(w_mem_inst__abc_19396_new_n2356_));
NAND2X1 NAND2X1_631 ( .A(w_mem_inst__abc_19396_new_n2360_), .B(w_mem_inst__abc_19396_new_n2359_), .Y(w_mem_inst__abc_19396_new_n2361_));
NAND2X1 NAND2X1_632 ( .A(w_mem_inst_w_mem_11__30_), .B(w_mem_inst__abc_19396_new_n1606__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2374_));
NAND2X1 NAND2X1_633 ( .A(w_mem_inst_w_mem_15__30_), .B(w_mem_inst__abc_19396_new_n1613__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2377_));
NAND2X1 NAND2X1_634 ( .A(w_mem_inst_w_mem_0__30_), .B(w_mem_inst__abc_19396_new_n1621__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2381_));
NAND2X1 NAND2X1_635 ( .A(w_mem_inst__abc_19396_new_n2385_), .B(w_mem_inst__abc_19396_new_n2384_), .Y(w_mem_inst__abc_19396_new_n2386_));
NAND2X1 NAND2X1_636 ( .A(w_mem_inst_w_mem_11__31_), .B(w_mem_inst__abc_19396_new_n1606__bF_buf3), .Y(w_mem_inst__abc_19396_new_n2399_));
NAND2X1 NAND2X1_637 ( .A(w_mem_inst_w_mem_15__31_), .B(w_mem_inst__abc_19396_new_n1613__bF_buf3), .Y(w_mem_inst__abc_19396_new_n2402_));
NAND2X1 NAND2X1_638 ( .A(w_mem_inst_w_mem_0__31_), .B(w_mem_inst__abc_19396_new_n1621__bF_buf3), .Y(w_mem_inst__abc_19396_new_n2406_));
NAND2X1 NAND2X1_639 ( .A(w_mem_inst__abc_19396_new_n2410_), .B(w_mem_inst__abc_19396_new_n2409_), .Y(w_mem_inst__abc_19396_new_n2411_));
NAND2X1 NAND2X1_64 ( .A(digest_update_bF_buf8), .B(_abc_15497_new_n1266_), .Y(_abc_15497_new_n1267_));
NAND2X1 NAND2X1_640 ( .A(w_mem_inst__abc_19396_new_n2419_), .B(w_mem_inst__abc_19396_new_n2420__bF_buf6), .Y(w_mem_inst__abc_19396_new_n4791_));
NAND2X1 NAND2X1_641 ( .A(round_ctr_inc_bF_buf0), .B(w_mem_inst__abc_19396_new_n1626_), .Y(w_mem_inst__abc_19396_new_n4792_));
NAND2X1 NAND2X1_642 ( .A(round_ctr_inc_bF_buf11), .B(w_mem_inst__abc_19396_new_n1610_), .Y(w_mem_inst__abc_19396_new_n4797_));
NAND2X1 NAND2X1_643 ( .A(round_ctr_inc_bF_buf9), .B(w_mem_inst__abc_19396_new_n1613__bF_buf2), .Y(w_mem_inst__abc_19396_new_n4801_));
NAND2X1 NAND2X1_644 ( .A(round_ctr_rst_bF_buf0), .B(w_mem_inst__abc_19396_new_n2419_), .Y(w_mem_inst__abc_19396_new_n4807_));
NAND2X1 NAND2X1_65 ( .A(e_reg_28_), .B(_auto_iopadmap_cc_368_execute_22625_28_), .Y(_abc_15497_new_n1270_));
NAND2X1 NAND2X1_66 ( .A(e_reg_30_), .B(_auto_iopadmap_cc_368_execute_22625_30_), .Y(_abc_15497_new_n1290_));
NAND2X1 NAND2X1_67 ( .A(_abc_15497_new_n1296_), .B(_abc_15497_new_n1295_), .Y(_0H4_reg_31_0__31_));
NAND2X1 NAND2X1_68 ( .A(_abc_15497_new_n1300_), .B(_abc_15497_new_n1303_), .Y(_abc_15497_new_n1309_));
NAND2X1 NAND2X1_69 ( .A(_abc_15497_new_n1326_), .B(_abc_15497_new_n1328_), .Y(_abc_15497_new_n1334_));
NAND2X1 NAND2X1_7 ( .A(_abc_15497_new_n771_), .B(_abc_15497_new_n772_), .Y(_abc_15497_new_n773_));
NAND2X1 NAND2X1_70 ( .A(_abc_15497_new_n1336_), .B(_abc_15497_new_n1335_), .Y(_abc_15497_new_n1338_));
NAND2X1 NAND2X1_71 ( .A(digest_update_bF_buf8), .B(_abc_15497_new_n1338_), .Y(_abc_15497_new_n1339_));
NAND2X1 NAND2X1_72 ( .A(_abc_15497_new_n1345_), .B(_abc_15497_new_n1344_), .Y(_abc_15497_new_n1347_));
NAND2X1 NAND2X1_73 ( .A(digest_update_bF_buf7), .B(_abc_15497_new_n1347_), .Y(_abc_15497_new_n1348_));
NAND2X1 NAND2X1_74 ( .A(_auto_iopadmap_cc_368_execute_22625_42_), .B(d_reg_10_), .Y(_abc_15497_new_n1387_));
NAND2X1 NAND2X1_75 ( .A(_abc_15497_new_n1393_), .B(_abc_15497_new_n1392_), .Y(_0H3_reg_31_0__10_));
NAND2X1 NAND2X1_76 ( .A(_abc_15497_new_n1389_), .B(_abc_15497_new_n1400_), .Y(_abc_15497_new_n1405_));
NAND2X1 NAND2X1_77 ( .A(_abc_15497_new_n1416_), .B(_abc_15497_new_n1411_), .Y(_abc_15497_new_n1418_));
NAND2X1 NAND2X1_78 ( .A(digest_update_bF_buf4), .B(_abc_15497_new_n1418_), .Y(_abc_15497_new_n1419_));
NAND2X1 NAND2X1_79 ( .A(_auto_iopadmap_cc_368_execute_22625_46_), .B(d_reg_14_), .Y(_abc_15497_new_n1436_));
NAND2X1 NAND2X1_8 ( .A(_abc_15497_new_n768_), .B(_abc_15497_new_n773_), .Y(_abc_15497_new_n774_));
NAND2X1 NAND2X1_80 ( .A(_abc_15497_new_n1438_), .B(_abc_15497_new_n1449_), .Y(_abc_15497_new_n1453_));
NAND2X1 NAND2X1_81 ( .A(_abc_15497_new_n1416_), .B(_abc_15497_new_n1427_), .Y(_abc_15497_new_n1456_));
NAND2X1 NAND2X1_82 ( .A(_abc_15497_new_n1457_), .B(_abc_15497_new_n1406_), .Y(_abc_15497_new_n1459_));
NAND2X1 NAND2X1_83 ( .A(_auto_iopadmap_cc_368_execute_22625_49_), .B(d_reg_17_), .Y(_abc_15497_new_n1469_));
NAND2X1 NAND2X1_84 ( .A(_abc_15497_new_n1475_), .B(_abc_15497_new_n1474_), .Y(_0H3_reg_31_0__17_));
NAND2X1 NAND2X1_85 ( .A(_abc_15497_new_n1471_), .B(_abc_15497_new_n1464_), .Y(_abc_15497_new_n1480_));
NAND2X1 NAND2X1_86 ( .A(_auto_iopadmap_cc_368_execute_22625_53_), .B(d_reg_21_), .Y(_abc_15497_new_n1523_));
NAND2X1 NAND2X1_87 ( .A(_abc_15497_new_n1523_), .B(_abc_15497_new_n1522_), .Y(_abc_15497_new_n1524_));
NAND2X1 NAND2X1_88 ( .A(_abc_15497_new_n1540_), .B(_abc_15497_new_n1543_), .Y(_abc_15497_new_n1544_));
NAND2X1 NAND2X1_89 ( .A(_auto_iopadmap_cc_368_execute_22625_55_), .B(d_reg_23_), .Y(_abc_15497_new_n1545_));
NAND2X1 NAND2X1_9 ( .A(_abc_15497_new_n779_), .B(_abc_15497_new_n778_), .Y(_abc_15497_new_n780_));
NAND2X1 NAND2X1_90 ( .A(_abc_15497_new_n1545_), .B(_abc_15497_new_n1544_), .Y(_abc_15497_new_n1546_));
NAND2X1 NAND2X1_91 ( .A(_abc_15497_new_n1535_), .B(_abc_15497_new_n1553_), .Y(_abc_15497_new_n1555_));
NAND2X1 NAND2X1_92 ( .A(_abc_15497_new_n1581_), .B(_abc_15497_new_n1604_), .Y(_abc_15497_new_n1605_));
NAND2X1 NAND2X1_93 ( .A(_abc_15497_new_n1611_), .B(_abc_15497_new_n1610_), .Y(_abc_15497_new_n1613_));
NAND2X1 NAND2X1_94 ( .A(digest_update_bF_buf3), .B(_abc_15497_new_n1613_), .Y(_abc_15497_new_n1614_));
NAND2X1 NAND2X1_95 ( .A(_auto_iopadmap_cc_368_execute_22625_60_), .B(d_reg_28_), .Y(_abc_15497_new_n1618_));
NAND2X1 NAND2X1_96 ( .A(_auto_iopadmap_cc_368_execute_22625_62_), .B(d_reg_30_), .Y(_abc_15497_new_n1638_));
NAND2X1 NAND2X1_97 ( .A(e_reg_31_), .B(_abc_15497_new_n1663__bF_buf5), .Y(_abc_15497_new_n1747_));
NAND2X1 NAND2X1_98 ( .A(d_reg_31_), .B(round_ctr_inc_bF_buf12), .Y(_abc_15497_new_n1748_));
NAND2X1 NAND2X1_99 ( .A(_abc_15497_new_n1757_), .B(_abc_15497_new_n1758_), .Y(_abc_15497_new_n1764_));
NAND3X1 NAND3X1_1 ( .A(_abc_15497_new_n926_), .B(_abc_15497_new_n929_), .C(_abc_15497_new_n928_), .Y(_abc_15497_new_n930_));
NAND3X1 NAND3X1_10 ( .A(_abc_15497_new_n2735_), .B(_abc_15497_new_n2736_), .C(_abc_15497_new_n2737_), .Y(_abc_15497_new_n2738_));
NAND3X1 NAND3X1_100 ( .A(w_12_), .B(_abc_15497_new_n3433_), .C(_abc_15497_new_n3436_), .Y(_abc_15497_new_n3437_));
NAND3X1 NAND3X1_101 ( .A(_abc_15497_new_n3435_), .B(_abc_15497_new_n3437_), .C(_abc_15497_new_n3430_), .Y(_abc_15497_new_n3438_));
NAND3X1 NAND3X1_102 ( .A(_abc_15497_new_n3429_), .B(_abc_15497_new_n3437_), .C(_abc_15497_new_n3435_), .Y(_abc_15497_new_n3449_));
NAND3X1 NAND3X1_103 ( .A(_abc_15497_new_n3456_), .B(_abc_15497_new_n3457_), .C(_abc_15497_new_n3455_), .Y(_abc_15497_new_n3460_));
NAND3X1 NAND3X1_104 ( .A(_abc_15497_new_n3443_), .B(_abc_15497_new_n3452_), .C(_abc_15497_new_n3418_), .Y(_abc_15497_new_n3461_));
NAND3X1 NAND3X1_105 ( .A(_abc_15497_new_n2756__bF_buf3), .B(_abc_15497_new_n3460_), .C(_abc_15497_new_n3461_), .Y(_abc_15497_new_n3462_));
NAND3X1 NAND3X1_106 ( .A(_abc_15497_new_n3462_), .B(_abc_15497_new_n3417_), .C(_abc_15497_new_n3459_), .Y(_abc_15497_new_n3463_));
NAND3X1 NAND3X1_107 ( .A(_abc_15497_new_n2925__bF_buf1), .B(_abc_15497_new_n3460_), .C(_abc_15497_new_n3461_), .Y(_abc_15497_new_n3468_));
NAND3X1 NAND3X1_108 ( .A(_abc_15497_new_n3468_), .B(_abc_15497_new_n3467_), .C(_abc_15497_new_n3469_), .Y(_abc_15497_new_n3470_));
NAND3X1 NAND3X1_109 ( .A(d_reg_13_), .B(_abc_15497_new_n3485_), .C(_abc_15497_new_n3484_), .Y(_abc_15497_new_n3486_));
NAND3X1 NAND3X1_11 ( .A(_abc_15497_new_n2740_), .B(_abc_15497_new_n2735_), .C(_abc_15497_new_n2741_), .Y(_abc_15497_new_n2742_));
NAND3X1 NAND3X1_110 ( .A(w_13_), .B(_abc_15497_new_n3499_), .C(_abc_15497_new_n3498_), .Y(_abc_15497_new_n3500_));
NAND3X1 NAND3X1_111 ( .A(_abc_15497_new_n3493_), .B(_abc_15497_new_n3497_), .C(_abc_15497_new_n3500_), .Y(_abc_15497_new_n3508_));
NAND3X1 NAND3X1_112 ( .A(_abc_15497_new_n3513_), .B(_abc_15497_new_n3514_), .C(_abc_15497_new_n3518_), .Y(_abc_15497_new_n3519_));
NAND3X1 NAND3X1_113 ( .A(_abc_15497_new_n3505_), .B(_abc_15497_new_n3511_), .C(_abc_15497_new_n3480_), .Y(_abc_15497_new_n3520_));
NAND3X1 NAND3X1_114 ( .A(_abc_15497_new_n2755_), .B(_abc_15497_new_n3519_), .C(_abc_15497_new_n3520_), .Y(_abc_15497_new_n3521_));
NAND3X1 NAND3X1_115 ( .A(_abc_15497_new_n3521_), .B(_abc_15497_new_n3516_), .C(_abc_15497_new_n3479_), .Y(_abc_15497_new_n3522_));
NAND3X1 NAND3X1_116 ( .A(_abc_15497_new_n3522_), .B(_abc_15497_new_n3536_), .C(_abc_15497_new_n3539_), .Y(_abc_15497_new_n3540_));
NAND3X1 NAND3X1_117 ( .A(d_reg_14_), .B(_abc_15497_new_n3548_), .C(_abc_15497_new_n3547_), .Y(_abc_15497_new_n3549_));
NAND3X1 NAND3X1_118 ( .A(w_14_), .B(_abc_15497_new_n3564_), .C(_abc_15497_new_n3563_), .Y(_abc_15497_new_n3565_));
NAND3X1 NAND3X1_119 ( .A(_abc_15497_new_n3562_), .B(_abc_15497_new_n3565_), .C(_abc_15497_new_n3558_), .Y(_abc_15497_new_n3566_));
NAND3X1 NAND3X1_12 ( .A(_abc_15497_new_n2747_), .B(_abc_15497_new_n2750_), .C(_abc_15497_new_n2756__bF_buf4), .Y(_abc_15497_new_n2757_));
NAND3X1 NAND3X1_120 ( .A(_abc_15497_new_n3557_), .B(_abc_15497_new_n3562_), .C(_abc_15497_new_n3565_), .Y(_abc_15497_new_n3574_));
NAND3X1 NAND3X1_121 ( .A(_abc_15497_new_n3579_), .B(_abc_15497_new_n3580_), .C(_abc_15497_new_n3587_), .Y(_abc_15497_new_n3588_));
NAND3X1 NAND3X1_122 ( .A(_abc_15497_new_n3571_), .B(_abc_15497_new_n3577_), .C(_abc_15497_new_n3542_), .Y(_abc_15497_new_n3589_));
NAND3X1 NAND3X1_123 ( .A(_abc_15497_new_n2924__bF_buf0), .B(_abc_15497_new_n3589_), .C(_abc_15497_new_n3588_), .Y(_abc_15497_new_n3590_));
NAND3X1 NAND3X1_124 ( .A(_abc_15497_new_n3590_), .B(_abc_15497_new_n3582_), .C(_abc_15497_new_n3541_), .Y(_abc_15497_new_n3591_));
NAND3X1 NAND3X1_125 ( .A(w_15_), .B(_abc_15497_new_n3624_), .C(_abc_15497_new_n3627_), .Y(_abc_15497_new_n3628_));
NAND3X1 NAND3X1_126 ( .A(_abc_15497_new_n3626_), .B(_abc_15497_new_n3628_), .C(_abc_15497_new_n3621_), .Y(_abc_15497_new_n3629_));
NAND3X1 NAND3X1_127 ( .A(_abc_15497_new_n3613_), .B(_abc_15497_new_n3636_), .C(_abc_15497_new_n2756__bF_buf3), .Y(_abc_15497_new_n3637_));
NAND3X1 NAND3X1_128 ( .A(_abc_15497_new_n3620_), .B(_abc_15497_new_n3628_), .C(_abc_15497_new_n3626_), .Y(_abc_15497_new_n3639_));
NAND3X1 NAND3X1_129 ( .A(_abc_15497_new_n3637_), .B(_abc_15497_new_n3638_), .C(_abc_15497_new_n3641_), .Y(_abc_15497_new_n3642_));
NAND3X1 NAND3X1_13 ( .A(_abc_15497_new_n2769_), .B(_abc_15497_new_n2767_), .C(_abc_15497_new_n2770_), .Y(_abc_15497_new_n2771_));
NAND3X1 NAND3X1_130 ( .A(_abc_15497_new_n3637_), .B(_abc_15497_new_n3638_), .C(_abc_15497_new_n3633_), .Y(_abc_15497_new_n3645_));
NAND3X1 NAND3X1_131 ( .A(_abc_15497_new_n3644_), .B(_abc_15497_new_n3645_), .C(_abc_15497_new_n3651_), .Y(_abc_15497_new_n3652_));
NAND3X1 NAND3X1_132 ( .A(_abc_15497_new_n3634_), .B(_abc_15497_new_n3642_), .C(_abc_15497_new_n3606_), .Y(_abc_15497_new_n3653_));
NAND3X1 NAND3X1_133 ( .A(_abc_15497_new_n2742__bF_buf3), .B(_abc_15497_new_n3652_), .C(_abc_15497_new_n3653_), .Y(_abc_15497_new_n3654_));
NAND3X1 NAND3X1_134 ( .A(_abc_15497_new_n3654_), .B(_abc_15497_new_n3605_), .C(_abc_15497_new_n3647_), .Y(_abc_15497_new_n3655_));
NAND3X1 NAND3X1_135 ( .A(_abc_15497_new_n3698_), .B(_abc_15497_new_n3701_), .C(_abc_15497_new_n3681_), .Y(_abc_15497_new_n3702_));
NAND3X1 NAND3X1_136 ( .A(_abc_15497_new_n3680_), .B(_abc_15497_new_n3703_), .C(_abc_15497_new_n3704_), .Y(_abc_15497_new_n3705_));
NAND3X1 NAND3X1_137 ( .A(_abc_15497_new_n3679_), .B(_abc_15497_new_n3705_), .C(_abc_15497_new_n3702_), .Y(_abc_15497_new_n3706_));
NAND3X1 NAND3X1_138 ( .A(_abc_15497_new_n3706_), .B(_abc_15497_new_n3709_), .C(_abc_15497_new_n3677_), .Y(_abc_15497_new_n3710_));
NAND3X1 NAND3X1_139 ( .A(_abc_15497_new_n3753_), .B(_abc_15497_new_n3750_), .C(_abc_15497_new_n3725_), .Y(_abc_15497_new_n3762_));
NAND3X1 NAND3X1_14 ( .A(w_1_), .B(_abc_15497_new_n2794_), .C(_abc_15497_new_n2797_), .Y(_abc_15497_new_n2798_));
NAND3X1 NAND3X1_140 ( .A(_abc_15497_new_n2781__bF_buf1), .B(_abc_15497_new_n3762_), .C(_abc_15497_new_n3761_), .Y(_abc_15497_new_n3763_));
NAND3X1 NAND3X1_141 ( .A(_abc_15497_new_n3722_), .B(_abc_15497_new_n3763_), .C(_abc_15497_new_n3760_), .Y(_abc_15497_new_n3764_));
NAND3X1 NAND3X1_142 ( .A(_abc_15497_new_n2944_), .B(_abc_15497_new_n3762_), .C(_abc_15497_new_n3761_), .Y(_abc_15497_new_n3766_));
NAND3X1 NAND3X1_143 ( .A(_abc_15497_new_n3765_), .B(_abc_15497_new_n3766_), .C(_abc_15497_new_n3767_), .Y(_abc_15497_new_n3768_));
NAND3X1 NAND3X1_144 ( .A(_abc_15497_new_n3765_), .B(_abc_15497_new_n3763_), .C(_abc_15497_new_n3760_), .Y(_abc_15497_new_n3778_));
NAND3X1 NAND3X1_145 ( .A(_abc_15497_new_n3806_), .B(_abc_15497_new_n3807_), .C(_abc_15497_new_n3804_), .Y(_abc_15497_new_n3808_));
NAND3X1 NAND3X1_146 ( .A(_abc_15497_new_n3810_), .B(_abc_15497_new_n3813_), .C(_abc_15497_new_n3816_), .Y(_abc_15497_new_n3817_));
NAND3X1 NAND3X1_147 ( .A(_abc_15497_new_n3847_), .B(_abc_15497_new_n3850_), .C(_abc_15497_new_n3829_), .Y(_abc_15497_new_n3851_));
NAND3X1 NAND3X1_148 ( .A(_abc_15497_new_n3853_), .B(_abc_15497_new_n3854_), .C(_abc_15497_new_n3852_), .Y(_abc_15497_new_n3855_));
NAND3X1 NAND3X1_149 ( .A(_abc_15497_new_n3679_), .B(_abc_15497_new_n3851_), .C(_abc_15497_new_n3855_), .Y(_abc_15497_new_n3856_));
NAND3X1 NAND3X1_15 ( .A(_abc_15497_new_n2791_), .B(_abc_15497_new_n2796_), .C(_abc_15497_new_n2798_), .Y(_abc_15497_new_n2799_));
NAND3X1 NAND3X1_150 ( .A(_abc_15497_new_n3856_), .B(_abc_15497_new_n3859_), .C(_abc_15497_new_n3827_), .Y(_abc_15497_new_n3860_));
NAND3X1 NAND3X1_151 ( .A(_abc_15497_new_n3678_), .B(_abc_15497_new_n3851_), .C(_abc_15497_new_n3855_), .Y(_abc_15497_new_n3861_));
NAND3X1 NAND3X1_152 ( .A(_abc_15497_new_n3810_), .B(_abc_15497_new_n3861_), .C(_abc_15497_new_n3862_), .Y(_abc_15497_new_n3863_));
NAND3X1 NAND3X1_153 ( .A(_abc_15497_new_n3769_), .B(_abc_15497_new_n3883_), .C(_abc_15497_new_n3713_), .Y(_abc_15497_new_n3884_));
NAND3X1 NAND3X1_154 ( .A(_abc_15497_new_n3910_), .B(_abc_15497_new_n3913_), .C(_abc_15497_new_n3893_), .Y(_abc_15497_new_n3914_));
NAND3X1 NAND3X1_155 ( .A(_abc_15497_new_n3916_), .B(_abc_15497_new_n3917_), .C(_abc_15497_new_n3915_), .Y(_abc_15497_new_n3918_));
NAND3X1 NAND3X1_156 ( .A(_abc_15497_new_n3679_), .B(_abc_15497_new_n3918_), .C(_abc_15497_new_n3914_), .Y(_abc_15497_new_n3919_));
NAND3X1 NAND3X1_157 ( .A(_abc_15497_new_n3919_), .B(_abc_15497_new_n3886_), .C(_abc_15497_new_n3922_), .Y(_abc_15497_new_n3923_));
NAND3X1 NAND3X1_158 ( .A(_abc_15497_new_n3678_), .B(_abc_15497_new_n3918_), .C(_abc_15497_new_n3914_), .Y(_abc_15497_new_n3925_));
NAND3X1 NAND3X1_159 ( .A(_abc_15497_new_n3925_), .B(_abc_15497_new_n3924_), .C(_abc_15497_new_n3926_), .Y(_abc_15497_new_n3927_));
NAND3X1 NAND3X1_16 ( .A(_abc_15497_new_n2774_), .B(_abc_15497_new_n2819_), .C(_abc_15497_new_n2820_), .Y(_abc_15497_new_n2821_));
NAND3X1 NAND3X1_160 ( .A(_abc_15497_new_n3961_), .B(_abc_15497_new_n3964_), .C(_abc_15497_new_n3943_), .Y(_abc_15497_new_n3965_));
NAND3X1 NAND3X1_161 ( .A(_abc_15497_new_n3967_), .B(_abc_15497_new_n3968_), .C(_abc_15497_new_n3966_), .Y(_abc_15497_new_n3969_));
NAND3X1 NAND3X1_162 ( .A(_abc_15497_new_n2755_), .B(_abc_15497_new_n3969_), .C(_abc_15497_new_n3965_), .Y(_abc_15497_new_n3970_));
NAND3X1 NAND3X1_163 ( .A(_abc_15497_new_n3970_), .B(_abc_15497_new_n3937_), .C(_abc_15497_new_n3973_), .Y(_abc_15497_new_n3974_));
NAND3X1 NAND3X1_164 ( .A(_abc_15497_new_n2780__bF_buf1), .B(_abc_15497_new_n3969_), .C(_abc_15497_new_n3965_), .Y(_abc_15497_new_n3976_));
NAND3X1 NAND3X1_165 ( .A(_abc_15497_new_n3976_), .B(_abc_15497_new_n3977_), .C(_abc_15497_new_n3975_), .Y(_abc_15497_new_n3978_));
NAND3X1 NAND3X1_166 ( .A(_abc_15497_new_n3970_), .B(_abc_15497_new_n3973_), .C(_abc_15497_new_n3975_), .Y(_abc_15497_new_n3989_));
NAND3X1 NAND3X1_167 ( .A(_abc_15497_new_n4016_), .B(_abc_15497_new_n4019_), .C(_abc_15497_new_n3998_), .Y(_abc_15497_new_n4020_));
NAND3X1 NAND3X1_168 ( .A(_abc_15497_new_n4022_), .B(_abc_15497_new_n4023_), .C(_abc_15497_new_n4021_), .Y(_abc_15497_new_n4024_));
NAND3X1 NAND3X1_169 ( .A(_abc_15497_new_n2925__bF_buf1), .B(_abc_15497_new_n4024_), .C(_abc_15497_new_n4020_), .Y(_abc_15497_new_n4025_));
NAND3X1 NAND3X1_17 ( .A(_abc_15497_new_n2805_), .B(_abc_15497_new_n2808_), .C(_abc_15497_new_n2771_), .Y(_abc_15497_new_n2826_));
NAND3X1 NAND3X1_170 ( .A(_abc_15497_new_n4025_), .B(_abc_15497_new_n3992_), .C(_abc_15497_new_n4028_), .Y(_abc_15497_new_n4029_));
NAND3X1 NAND3X1_171 ( .A(_abc_15497_new_n2756__bF_buf2), .B(_abc_15497_new_n4024_), .C(_abc_15497_new_n4020_), .Y(_abc_15497_new_n4031_));
NAND3X1 NAND3X1_172 ( .A(_abc_15497_new_n4031_), .B(_abc_15497_new_n4032_), .C(_abc_15497_new_n4030_), .Y(_abc_15497_new_n4033_));
NAND3X1 NAND3X1_173 ( .A(_abc_15497_new_n4066_), .B(_abc_15497_new_n4063_), .C(_abc_15497_new_n4067_), .Y(_abc_15497_new_n4068_));
NAND3X1 NAND3X1_174 ( .A(_abc_15497_new_n4062_), .B(_abc_15497_new_n4013_), .C(_abc_15497_new_n4069_), .Y(_abc_15497_new_n4070_));
NAND3X1 NAND3X1_175 ( .A(_abc_15497_new_n4077_), .B(_abc_15497_new_n4078_), .C(_abc_15497_new_n4076_), .Y(_abc_15497_new_n4081_));
NAND3X1 NAND3X1_176 ( .A(_abc_15497_new_n4073_), .B(_abc_15497_new_n4072_), .C(_abc_15497_new_n4049_), .Y(_abc_15497_new_n4082_));
NAND3X1 NAND3X1_177 ( .A(_abc_15497_new_n2738_), .B(_abc_15497_new_n4082_), .C(_abc_15497_new_n4081_), .Y(_abc_15497_new_n4083_));
NAND3X1 NAND3X1_178 ( .A(_abc_15497_new_n4083_), .B(_abc_15497_new_n4044_), .C(_abc_15497_new_n4080_), .Y(_abc_15497_new_n4084_));
NAND3X1 NAND3X1_179 ( .A(_abc_15497_new_n2739_), .B(_abc_15497_new_n4082_), .C(_abc_15497_new_n4081_), .Y(_abc_15497_new_n4086_));
NAND3X1 NAND3X1_18 ( .A(w_2_), .B(_abc_15497_new_n2842_), .C(_abc_15497_new_n2845_), .Y(_abc_15497_new_n2846_));
NAND3X1 NAND3X1_180 ( .A(_abc_15497_new_n4086_), .B(_abc_15497_new_n4087_), .C(_abc_15497_new_n4085_), .Y(_abc_15497_new_n4088_));
NAND3X1 NAND3X1_181 ( .A(_abc_15497_new_n4083_), .B(_abc_15497_new_n4080_), .C(_abc_15497_new_n4085_), .Y(_abc_15497_new_n4101_));
NAND3X1 NAND3X1_182 ( .A(_abc_15497_new_n3776_), .B(_abc_15497_new_n3883_), .C(_abc_15497_new_n4098_), .Y(_abc_15497_new_n4105_));
NAND3X1 NAND3X1_183 ( .A(_abc_15497_new_n4112_), .B(_abc_15497_new_n4113_), .C(_abc_15497_new_n2756__bF_buf0), .Y(_abc_15497_new_n4114_));
NAND3X1 NAND3X1_184 ( .A(_abc_15497_new_n4125_), .B(_abc_15497_new_n4127_), .C(_abc_15497_new_n4121_), .Y(_abc_15497_new_n4128_));
NAND3X1 NAND3X1_185 ( .A(_abc_15497_new_n4120_), .B(_abc_15497_new_n4067_), .C(_abc_15497_new_n4129_), .Y(_abc_15497_new_n4130_));
NAND3X1 NAND3X1_186 ( .A(_abc_15497_new_n4141_), .B(_abc_15497_new_n4138_), .C(_abc_15497_new_n4137_), .Y(_abc_15497_new_n4142_));
NAND3X1 NAND3X1_187 ( .A(_abc_15497_new_n4107_), .B(_abc_15497_new_n4138_), .C(_abc_15497_new_n4137_), .Y(_abc_15497_new_n4149_));
NAND3X1 NAND3X1_188 ( .A(_abc_15497_new_n4162_), .B(_abc_15497_new_n4170_), .C(_abc_15497_new_n4169_), .Y(_abc_15497_new_n4192_));
NAND3X1 NAND3X1_189 ( .A(_abc_15497_new_n4173_), .B(_abc_15497_new_n4220_), .C(_abc_15497_new_n4223_), .Y(_abc_15497_new_n4224_));
NAND3X1 NAND3X1_19 ( .A(_abc_15497_new_n2839_), .B(_abc_15497_new_n2844_), .C(_abc_15497_new_n2846_), .Y(_abc_15497_new_n2847_));
NAND3X1 NAND3X1_190 ( .A(_abc_15497_new_n4210_), .B(_abc_15497_new_n4212_), .C(_abc_15497_new_n4206_), .Y(_abc_15497_new_n4237_));
NAND3X1 NAND3X1_191 ( .A(_abc_15497_new_n4257_), .B(_abc_15497_new_n4249_), .C(_abc_15497_new_n4256_), .Y(_abc_15497_new_n4278_));
NAND3X1 NAND3X1_192 ( .A(_abc_15497_new_n3058_), .B(_abc_15497_new_n3213_), .C(_abc_15497_new_n2942_), .Y(_abc_15497_new_n4305_));
NAND3X1 NAND3X1_193 ( .A(_abc_15497_new_n3522_), .B(_abc_15497_new_n3526_), .C(_abc_15497_new_n3471_), .Y(_abc_15497_new_n4308_));
NAND3X1 NAND3X1_194 ( .A(_abc_15497_new_n3655_), .B(_abc_15497_new_n3659_), .C(_abc_15497_new_n3596_), .Y(_abc_15497_new_n4309_));
NAND3X1 NAND3X1_195 ( .A(_abc_15497_new_n4225_), .B(_abc_15497_new_n4263_), .C(_abc_15497_new_n4189_), .Y(_abc_15497_new_n4316_));
NAND3X1 NAND3X1_196 ( .A(_abc_15497_new_n4289_), .B(_abc_15497_new_n4297_), .C(_abc_15497_new_n4296_), .Y(_abc_15497_new_n4328_));
NAND3X1 NAND3X1_197 ( .A(_abc_15497_new_n4329_), .B(_abc_15497_new_n4351_), .C(_abc_15497_new_n4350_), .Y(_abc_15497_new_n4369_));
NAND3X1 NAND3X1_198 ( .A(_abc_15497_new_n4396_), .B(_abc_15497_new_n4397_), .C(_abc_15497_new_n4371_), .Y(_abc_15497_new_n4411_));
NAND3X1 NAND3X1_199 ( .A(round_ctr_reg_6_), .B(_abc_15497_new_n4441_), .C(_abc_15497_new_n4446_), .Y(_abc_15497_new_n4447_));
NAND3X1 NAND3X1_2 ( .A(_abc_15497_new_n996_), .B(_abc_15497_new_n1013_), .C(_abc_15497_new_n1015_), .Y(_abc_15497_new_n1016_));
NAND3X1 NAND3X1_20 ( .A(_abc_15497_new_n2855_), .B(_abc_15497_new_n2852_), .C(_abc_15497_new_n2828_), .Y(_abc_15497_new_n2856_));
NAND3X1 NAND3X1_200 ( .A(w_mem_inst_w_mem_13__0_), .B(w_mem_inst__abc_19396_new_n1617__bF_buf7), .C(w_mem_inst__abc_19396_new_n1594__bF_buf6), .Y(w_mem_inst__abc_19396_new_n1618_));
NAND3X1 NAND3X1_201 ( .A(w_mem_inst_w_mem_12__0_), .B(w_mem_inst__abc_19396_new_n1619__bF_buf3), .C(w_mem_inst__abc_19396_new_n1617__bF_buf6), .Y(w_mem_inst__abc_19396_new_n1623_));
NAND3X1 NAND3X1_202 ( .A(w_mem_inst__abc_19396_new_n1623_), .B(w_mem_inst__abc_19396_new_n1622_), .C(w_mem_inst__abc_19396_new_n1618_), .Y(w_mem_inst__abc_19396_new_n1624_));
NAND3X1 NAND3X1_203 ( .A(w_mem_inst_w_mem_1__0_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf6), .C(w_mem_inst__abc_19396_new_n1594__bF_buf5), .Y(w_mem_inst__abc_19396_new_n1634_));
NAND3X1 NAND3X1_204 ( .A(w_mem_inst_w_mem_2__0_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf5), .C(w_mem_inst__abc_19396_new_n1635__bF_buf4), .Y(w_mem_inst__abc_19396_new_n1636_));
NAND3X1 NAND3X1_205 ( .A(w_mem_inst__abc_19396_new_n1634_), .B(w_mem_inst__abc_19396_new_n1636_), .C(w_mem_inst__abc_19396_new_n1639_), .Y(w_mem_inst__abc_19396_new_n1640_));
NAND3X1 NAND3X1_206 ( .A(w_mem_inst_w_mem_13__1_), .B(w_mem_inst__abc_19396_new_n1617__bF_buf5), .C(w_mem_inst__abc_19396_new_n1594__bF_buf4), .Y(w_mem_inst__abc_19396_new_n1655_));
NAND3X1 NAND3X1_207 ( .A(w_mem_inst_w_mem_12__1_), .B(w_mem_inst__abc_19396_new_n1619__bF_buf2), .C(w_mem_inst__abc_19396_new_n1617__bF_buf4), .Y(w_mem_inst__abc_19396_new_n1657_));
NAND3X1 NAND3X1_208 ( .A(w_mem_inst__abc_19396_new_n1657_), .B(w_mem_inst__abc_19396_new_n1656_), .C(w_mem_inst__abc_19396_new_n1655_), .Y(w_mem_inst__abc_19396_new_n1658_));
NAND3X1 NAND3X1_209 ( .A(w_mem_inst_w_mem_1__1_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf4), .C(w_mem_inst__abc_19396_new_n1594__bF_buf3), .Y(w_mem_inst__abc_19396_new_n1662_));
NAND3X1 NAND3X1_21 ( .A(_abc_15497_new_n2858_), .B(_abc_15497_new_n2859_), .C(_abc_15497_new_n2860_), .Y(_abc_15497_new_n2861_));
NAND3X1 NAND3X1_210 ( .A(w_mem_inst_w_mem_2__1_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf3), .C(w_mem_inst__abc_19396_new_n1635__bF_buf3), .Y(w_mem_inst__abc_19396_new_n1663_));
NAND3X1 NAND3X1_211 ( .A(w_mem_inst__abc_19396_new_n1662_), .B(w_mem_inst__abc_19396_new_n1663_), .C(w_mem_inst__abc_19396_new_n1664_), .Y(w_mem_inst__abc_19396_new_n1665_));
NAND3X1 NAND3X1_212 ( .A(w_mem_inst_w_mem_13__2_), .B(w_mem_inst__abc_19396_new_n1617__bF_buf3), .C(w_mem_inst__abc_19396_new_n1594__bF_buf2), .Y(w_mem_inst__abc_19396_new_n1680_));
NAND3X1 NAND3X1_213 ( .A(w_mem_inst_w_mem_12__2_), .B(w_mem_inst__abc_19396_new_n1619__bF_buf1), .C(w_mem_inst__abc_19396_new_n1617__bF_buf2), .Y(w_mem_inst__abc_19396_new_n1682_));
NAND3X1 NAND3X1_214 ( .A(w_mem_inst__abc_19396_new_n1682_), .B(w_mem_inst__abc_19396_new_n1681_), .C(w_mem_inst__abc_19396_new_n1680_), .Y(w_mem_inst__abc_19396_new_n1683_));
NAND3X1 NAND3X1_215 ( .A(w_mem_inst_w_mem_1__2_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf2), .C(w_mem_inst__abc_19396_new_n1594__bF_buf1), .Y(w_mem_inst__abc_19396_new_n1687_));
NAND3X1 NAND3X1_216 ( .A(w_mem_inst_w_mem_2__2_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf1), .C(w_mem_inst__abc_19396_new_n1635__bF_buf2), .Y(w_mem_inst__abc_19396_new_n1688_));
NAND3X1 NAND3X1_217 ( .A(w_mem_inst__abc_19396_new_n1687_), .B(w_mem_inst__abc_19396_new_n1688_), .C(w_mem_inst__abc_19396_new_n1689_), .Y(w_mem_inst__abc_19396_new_n1690_));
NAND3X1 NAND3X1_218 ( .A(w_mem_inst_w_mem_13__3_), .B(w_mem_inst__abc_19396_new_n1617__bF_buf1), .C(w_mem_inst__abc_19396_new_n1594__bF_buf0), .Y(w_mem_inst__abc_19396_new_n1705_));
NAND3X1 NAND3X1_219 ( .A(w_mem_inst_w_mem_12__3_), .B(w_mem_inst__abc_19396_new_n1619__bF_buf0), .C(w_mem_inst__abc_19396_new_n1617__bF_buf0), .Y(w_mem_inst__abc_19396_new_n1707_));
NAND3X1 NAND3X1_22 ( .A(_abc_15497_new_n2859_), .B(_abc_15497_new_n2860_), .C(_abc_15497_new_n2828_), .Y(_abc_15497_new_n2864_));
NAND3X1 NAND3X1_220 ( .A(w_mem_inst__abc_19396_new_n1707_), .B(w_mem_inst__abc_19396_new_n1706_), .C(w_mem_inst__abc_19396_new_n1705_), .Y(w_mem_inst__abc_19396_new_n1708_));
NAND3X1 NAND3X1_221 ( .A(w_mem_inst_w_mem_1__3_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf0), .C(w_mem_inst__abc_19396_new_n1594__bF_buf7), .Y(w_mem_inst__abc_19396_new_n1712_));
NAND3X1 NAND3X1_222 ( .A(w_mem_inst_w_mem_2__3_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf7), .C(w_mem_inst__abc_19396_new_n1635__bF_buf1), .Y(w_mem_inst__abc_19396_new_n1713_));
NAND3X1 NAND3X1_223 ( .A(w_mem_inst__abc_19396_new_n1712_), .B(w_mem_inst__abc_19396_new_n1713_), .C(w_mem_inst__abc_19396_new_n1714_), .Y(w_mem_inst__abc_19396_new_n1715_));
NAND3X1 NAND3X1_224 ( .A(w_mem_inst_w_mem_13__4_), .B(w_mem_inst__abc_19396_new_n1617__bF_buf7), .C(w_mem_inst__abc_19396_new_n1594__bF_buf6), .Y(w_mem_inst__abc_19396_new_n1730_));
NAND3X1 NAND3X1_225 ( .A(w_mem_inst_w_mem_12__4_), .B(w_mem_inst__abc_19396_new_n1619__bF_buf4), .C(w_mem_inst__abc_19396_new_n1617__bF_buf6), .Y(w_mem_inst__abc_19396_new_n1732_));
NAND3X1 NAND3X1_226 ( .A(w_mem_inst__abc_19396_new_n1732_), .B(w_mem_inst__abc_19396_new_n1731_), .C(w_mem_inst__abc_19396_new_n1730_), .Y(w_mem_inst__abc_19396_new_n1733_));
NAND3X1 NAND3X1_227 ( .A(w_mem_inst_w_mem_1__4_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf6), .C(w_mem_inst__abc_19396_new_n1594__bF_buf5), .Y(w_mem_inst__abc_19396_new_n1737_));
NAND3X1 NAND3X1_228 ( .A(w_mem_inst_w_mem_2__4_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf5), .C(w_mem_inst__abc_19396_new_n1635__bF_buf0), .Y(w_mem_inst__abc_19396_new_n1738_));
NAND3X1 NAND3X1_229 ( .A(w_mem_inst__abc_19396_new_n1737_), .B(w_mem_inst__abc_19396_new_n1738_), .C(w_mem_inst__abc_19396_new_n1739_), .Y(w_mem_inst__abc_19396_new_n1740_));
NAND3X1 NAND3X1_23 ( .A(_abc_15497_new_n2858_), .B(_abc_15497_new_n2855_), .C(_abc_15497_new_n2852_), .Y(_abc_15497_new_n2865_));
NAND3X1 NAND3X1_230 ( .A(w_mem_inst_w_mem_13__5_), .B(w_mem_inst__abc_19396_new_n1617__bF_buf5), .C(w_mem_inst__abc_19396_new_n1594__bF_buf4), .Y(w_mem_inst__abc_19396_new_n1755_));
NAND3X1 NAND3X1_231 ( .A(w_mem_inst_w_mem_12__5_), .B(w_mem_inst__abc_19396_new_n1619__bF_buf3), .C(w_mem_inst__abc_19396_new_n1617__bF_buf4), .Y(w_mem_inst__abc_19396_new_n1757_));
NAND3X1 NAND3X1_232 ( .A(w_mem_inst__abc_19396_new_n1757_), .B(w_mem_inst__abc_19396_new_n1756_), .C(w_mem_inst__abc_19396_new_n1755_), .Y(w_mem_inst__abc_19396_new_n1758_));
NAND3X1 NAND3X1_233 ( .A(w_mem_inst_w_mem_1__5_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf4), .C(w_mem_inst__abc_19396_new_n1594__bF_buf3), .Y(w_mem_inst__abc_19396_new_n1762_));
NAND3X1 NAND3X1_234 ( .A(w_mem_inst_w_mem_2__5_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf3), .C(w_mem_inst__abc_19396_new_n1635__bF_buf4), .Y(w_mem_inst__abc_19396_new_n1763_));
NAND3X1 NAND3X1_235 ( .A(w_mem_inst__abc_19396_new_n1762_), .B(w_mem_inst__abc_19396_new_n1763_), .C(w_mem_inst__abc_19396_new_n1764_), .Y(w_mem_inst__abc_19396_new_n1765_));
NAND3X1 NAND3X1_236 ( .A(w_mem_inst_w_mem_13__6_), .B(w_mem_inst__abc_19396_new_n1617__bF_buf3), .C(w_mem_inst__abc_19396_new_n1594__bF_buf2), .Y(w_mem_inst__abc_19396_new_n1780_));
NAND3X1 NAND3X1_237 ( .A(w_mem_inst_w_mem_12__6_), .B(w_mem_inst__abc_19396_new_n1619__bF_buf2), .C(w_mem_inst__abc_19396_new_n1617__bF_buf2), .Y(w_mem_inst__abc_19396_new_n1782_));
NAND3X1 NAND3X1_238 ( .A(w_mem_inst__abc_19396_new_n1782_), .B(w_mem_inst__abc_19396_new_n1781_), .C(w_mem_inst__abc_19396_new_n1780_), .Y(w_mem_inst__abc_19396_new_n1783_));
NAND3X1 NAND3X1_239 ( .A(w_mem_inst_w_mem_1__6_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf2), .C(w_mem_inst__abc_19396_new_n1594__bF_buf1), .Y(w_mem_inst__abc_19396_new_n1787_));
NAND3X1 NAND3X1_24 ( .A(_abc_15497_new_n2810_), .B(_abc_15497_new_n2811_), .C(_abc_15497_new_n2772_), .Y(_abc_15497_new_n2868_));
NAND3X1 NAND3X1_240 ( .A(w_mem_inst_w_mem_2__6_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf1), .C(w_mem_inst__abc_19396_new_n1635__bF_buf3), .Y(w_mem_inst__abc_19396_new_n1788_));
NAND3X1 NAND3X1_241 ( .A(w_mem_inst__abc_19396_new_n1787_), .B(w_mem_inst__abc_19396_new_n1788_), .C(w_mem_inst__abc_19396_new_n1789_), .Y(w_mem_inst__abc_19396_new_n1790_));
NAND3X1 NAND3X1_242 ( .A(w_mem_inst_w_mem_13__7_), .B(w_mem_inst__abc_19396_new_n1617__bF_buf1), .C(w_mem_inst__abc_19396_new_n1594__bF_buf0), .Y(w_mem_inst__abc_19396_new_n1805_));
NAND3X1 NAND3X1_243 ( .A(w_mem_inst_w_mem_12__7_), .B(w_mem_inst__abc_19396_new_n1619__bF_buf1), .C(w_mem_inst__abc_19396_new_n1617__bF_buf0), .Y(w_mem_inst__abc_19396_new_n1807_));
NAND3X1 NAND3X1_244 ( .A(w_mem_inst__abc_19396_new_n1807_), .B(w_mem_inst__abc_19396_new_n1806_), .C(w_mem_inst__abc_19396_new_n1805_), .Y(w_mem_inst__abc_19396_new_n1808_));
NAND3X1 NAND3X1_245 ( .A(w_mem_inst_w_mem_1__7_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf0), .C(w_mem_inst__abc_19396_new_n1594__bF_buf7), .Y(w_mem_inst__abc_19396_new_n1812_));
NAND3X1 NAND3X1_246 ( .A(w_mem_inst_w_mem_2__7_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf7), .C(w_mem_inst__abc_19396_new_n1635__bF_buf2), .Y(w_mem_inst__abc_19396_new_n1813_));
NAND3X1 NAND3X1_247 ( .A(w_mem_inst__abc_19396_new_n1812_), .B(w_mem_inst__abc_19396_new_n1813_), .C(w_mem_inst__abc_19396_new_n1814_), .Y(w_mem_inst__abc_19396_new_n1815_));
NAND3X1 NAND3X1_248 ( .A(w_mem_inst_w_mem_13__8_), .B(w_mem_inst__abc_19396_new_n1617__bF_buf7), .C(w_mem_inst__abc_19396_new_n1594__bF_buf6), .Y(w_mem_inst__abc_19396_new_n1830_));
NAND3X1 NAND3X1_249 ( .A(w_mem_inst_w_mem_12__8_), .B(w_mem_inst__abc_19396_new_n1619__bF_buf0), .C(w_mem_inst__abc_19396_new_n1617__bF_buf6), .Y(w_mem_inst__abc_19396_new_n1832_));
NAND3X1 NAND3X1_25 ( .A(_abc_15497_new_n2739_), .B(_abc_15497_new_n2865_), .C(_abc_15497_new_n2864_), .Y(_abc_15497_new_n2870_));
NAND3X1 NAND3X1_250 ( .A(w_mem_inst__abc_19396_new_n1832_), .B(w_mem_inst__abc_19396_new_n1831_), .C(w_mem_inst__abc_19396_new_n1830_), .Y(w_mem_inst__abc_19396_new_n1833_));
NAND3X1 NAND3X1_251 ( .A(w_mem_inst_w_mem_1__8_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf6), .C(w_mem_inst__abc_19396_new_n1594__bF_buf5), .Y(w_mem_inst__abc_19396_new_n1837_));
NAND3X1 NAND3X1_252 ( .A(w_mem_inst_w_mem_2__8_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf5), .C(w_mem_inst__abc_19396_new_n1635__bF_buf1), .Y(w_mem_inst__abc_19396_new_n1838_));
NAND3X1 NAND3X1_253 ( .A(w_mem_inst__abc_19396_new_n1837_), .B(w_mem_inst__abc_19396_new_n1838_), .C(w_mem_inst__abc_19396_new_n1839_), .Y(w_mem_inst__abc_19396_new_n1840_));
NAND3X1 NAND3X1_254 ( .A(w_mem_inst_w_mem_13__9_), .B(w_mem_inst__abc_19396_new_n1617__bF_buf5), .C(w_mem_inst__abc_19396_new_n1594__bF_buf4), .Y(w_mem_inst__abc_19396_new_n1855_));
NAND3X1 NAND3X1_255 ( .A(w_mem_inst_w_mem_12__9_), .B(w_mem_inst__abc_19396_new_n1619__bF_buf4), .C(w_mem_inst__abc_19396_new_n1617__bF_buf4), .Y(w_mem_inst__abc_19396_new_n1857_));
NAND3X1 NAND3X1_256 ( .A(w_mem_inst__abc_19396_new_n1857_), .B(w_mem_inst__abc_19396_new_n1856_), .C(w_mem_inst__abc_19396_new_n1855_), .Y(w_mem_inst__abc_19396_new_n1858_));
NAND3X1 NAND3X1_257 ( .A(w_mem_inst_w_mem_1__9_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf4), .C(w_mem_inst__abc_19396_new_n1594__bF_buf3), .Y(w_mem_inst__abc_19396_new_n1862_));
NAND3X1 NAND3X1_258 ( .A(w_mem_inst_w_mem_2__9_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf3), .C(w_mem_inst__abc_19396_new_n1635__bF_buf0), .Y(w_mem_inst__abc_19396_new_n1863_));
NAND3X1 NAND3X1_259 ( .A(w_mem_inst__abc_19396_new_n1862_), .B(w_mem_inst__abc_19396_new_n1863_), .C(w_mem_inst__abc_19396_new_n1864_), .Y(w_mem_inst__abc_19396_new_n1865_));
NAND3X1 NAND3X1_26 ( .A(_abc_15497_new_n2738_), .B(_abc_15497_new_n2861_), .C(_abc_15497_new_n2856_), .Y(_abc_15497_new_n2871_));
NAND3X1 NAND3X1_260 ( .A(w_mem_inst_w_mem_13__10_), .B(w_mem_inst__abc_19396_new_n1617__bF_buf3), .C(w_mem_inst__abc_19396_new_n1594__bF_buf2), .Y(w_mem_inst__abc_19396_new_n1880_));
NAND3X1 NAND3X1_261 ( .A(w_mem_inst_w_mem_12__10_), .B(w_mem_inst__abc_19396_new_n1619__bF_buf3), .C(w_mem_inst__abc_19396_new_n1617__bF_buf2), .Y(w_mem_inst__abc_19396_new_n1882_));
NAND3X1 NAND3X1_262 ( .A(w_mem_inst__abc_19396_new_n1882_), .B(w_mem_inst__abc_19396_new_n1881_), .C(w_mem_inst__abc_19396_new_n1880_), .Y(w_mem_inst__abc_19396_new_n1883_));
NAND3X1 NAND3X1_263 ( .A(w_mem_inst_w_mem_1__10_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf2), .C(w_mem_inst__abc_19396_new_n1594__bF_buf1), .Y(w_mem_inst__abc_19396_new_n1887_));
NAND3X1 NAND3X1_264 ( .A(w_mem_inst_w_mem_2__10_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf1), .C(w_mem_inst__abc_19396_new_n1635__bF_buf4), .Y(w_mem_inst__abc_19396_new_n1888_));
NAND3X1 NAND3X1_265 ( .A(w_mem_inst__abc_19396_new_n1887_), .B(w_mem_inst__abc_19396_new_n1888_), .C(w_mem_inst__abc_19396_new_n1889_), .Y(w_mem_inst__abc_19396_new_n1890_));
NAND3X1 NAND3X1_266 ( .A(w_mem_inst_w_mem_13__11_), .B(w_mem_inst__abc_19396_new_n1617__bF_buf1), .C(w_mem_inst__abc_19396_new_n1594__bF_buf0), .Y(w_mem_inst__abc_19396_new_n1905_));
NAND3X1 NAND3X1_267 ( .A(w_mem_inst_w_mem_12__11_), .B(w_mem_inst__abc_19396_new_n1619__bF_buf2), .C(w_mem_inst__abc_19396_new_n1617__bF_buf0), .Y(w_mem_inst__abc_19396_new_n1907_));
NAND3X1 NAND3X1_268 ( .A(w_mem_inst__abc_19396_new_n1907_), .B(w_mem_inst__abc_19396_new_n1906_), .C(w_mem_inst__abc_19396_new_n1905_), .Y(w_mem_inst__abc_19396_new_n1908_));
NAND3X1 NAND3X1_269 ( .A(w_mem_inst_w_mem_1__11_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf0), .C(w_mem_inst__abc_19396_new_n1594__bF_buf7), .Y(w_mem_inst__abc_19396_new_n1912_));
NAND3X1 NAND3X1_27 ( .A(_abc_15497_new_n2871_), .B(_abc_15497_new_n2870_), .C(_abc_15497_new_n2869_), .Y(_abc_15497_new_n2876_));
NAND3X1 NAND3X1_270 ( .A(w_mem_inst_w_mem_2__11_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf7), .C(w_mem_inst__abc_19396_new_n1635__bF_buf3), .Y(w_mem_inst__abc_19396_new_n1913_));
NAND3X1 NAND3X1_271 ( .A(w_mem_inst__abc_19396_new_n1912_), .B(w_mem_inst__abc_19396_new_n1913_), .C(w_mem_inst__abc_19396_new_n1914_), .Y(w_mem_inst__abc_19396_new_n1915_));
NAND3X1 NAND3X1_272 ( .A(w_mem_inst_w_mem_13__12_), .B(w_mem_inst__abc_19396_new_n1617__bF_buf7), .C(w_mem_inst__abc_19396_new_n1594__bF_buf6), .Y(w_mem_inst__abc_19396_new_n1930_));
NAND3X1 NAND3X1_273 ( .A(w_mem_inst_w_mem_12__12_), .B(w_mem_inst__abc_19396_new_n1619__bF_buf1), .C(w_mem_inst__abc_19396_new_n1617__bF_buf6), .Y(w_mem_inst__abc_19396_new_n1932_));
NAND3X1 NAND3X1_274 ( .A(w_mem_inst__abc_19396_new_n1932_), .B(w_mem_inst__abc_19396_new_n1931_), .C(w_mem_inst__abc_19396_new_n1930_), .Y(w_mem_inst__abc_19396_new_n1933_));
NAND3X1 NAND3X1_275 ( .A(w_mem_inst_w_mem_1__12_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf6), .C(w_mem_inst__abc_19396_new_n1594__bF_buf5), .Y(w_mem_inst__abc_19396_new_n1937_));
NAND3X1 NAND3X1_276 ( .A(w_mem_inst_w_mem_2__12_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf5), .C(w_mem_inst__abc_19396_new_n1635__bF_buf2), .Y(w_mem_inst__abc_19396_new_n1938_));
NAND3X1 NAND3X1_277 ( .A(w_mem_inst__abc_19396_new_n1937_), .B(w_mem_inst__abc_19396_new_n1938_), .C(w_mem_inst__abc_19396_new_n1939_), .Y(w_mem_inst__abc_19396_new_n1940_));
NAND3X1 NAND3X1_278 ( .A(w_mem_inst_w_mem_13__13_), .B(w_mem_inst__abc_19396_new_n1617__bF_buf5), .C(w_mem_inst__abc_19396_new_n1594__bF_buf4), .Y(w_mem_inst__abc_19396_new_n1955_));
NAND3X1 NAND3X1_279 ( .A(w_mem_inst_w_mem_12__13_), .B(w_mem_inst__abc_19396_new_n1619__bF_buf0), .C(w_mem_inst__abc_19396_new_n1617__bF_buf4), .Y(w_mem_inst__abc_19396_new_n1957_));
NAND3X1 NAND3X1_28 ( .A(_abc_15497_new_n2876_), .B(_abc_15497_new_n2875_), .C(_abc_15497_new_n2877_), .Y(_abc_15497_new_n2878_));
NAND3X1 NAND3X1_280 ( .A(w_mem_inst__abc_19396_new_n1957_), .B(w_mem_inst__abc_19396_new_n1956_), .C(w_mem_inst__abc_19396_new_n1955_), .Y(w_mem_inst__abc_19396_new_n1958_));
NAND3X1 NAND3X1_281 ( .A(w_mem_inst_w_mem_1__13_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf4), .C(w_mem_inst__abc_19396_new_n1594__bF_buf3), .Y(w_mem_inst__abc_19396_new_n1962_));
NAND3X1 NAND3X1_282 ( .A(w_mem_inst_w_mem_2__13_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf3), .C(w_mem_inst__abc_19396_new_n1635__bF_buf1), .Y(w_mem_inst__abc_19396_new_n1963_));
NAND3X1 NAND3X1_283 ( .A(w_mem_inst__abc_19396_new_n1962_), .B(w_mem_inst__abc_19396_new_n1963_), .C(w_mem_inst__abc_19396_new_n1964_), .Y(w_mem_inst__abc_19396_new_n1965_));
NAND3X1 NAND3X1_284 ( .A(w_mem_inst_w_mem_13__14_), .B(w_mem_inst__abc_19396_new_n1617__bF_buf3), .C(w_mem_inst__abc_19396_new_n1594__bF_buf2), .Y(w_mem_inst__abc_19396_new_n1980_));
NAND3X1 NAND3X1_285 ( .A(w_mem_inst_w_mem_12__14_), .B(w_mem_inst__abc_19396_new_n1619__bF_buf4), .C(w_mem_inst__abc_19396_new_n1617__bF_buf2), .Y(w_mem_inst__abc_19396_new_n1982_));
NAND3X1 NAND3X1_286 ( .A(w_mem_inst__abc_19396_new_n1982_), .B(w_mem_inst__abc_19396_new_n1981_), .C(w_mem_inst__abc_19396_new_n1980_), .Y(w_mem_inst__abc_19396_new_n1983_));
NAND3X1 NAND3X1_287 ( .A(w_mem_inst_w_mem_1__14_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf2), .C(w_mem_inst__abc_19396_new_n1594__bF_buf1), .Y(w_mem_inst__abc_19396_new_n1987_));
NAND3X1 NAND3X1_288 ( .A(w_mem_inst_w_mem_2__14_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf1), .C(w_mem_inst__abc_19396_new_n1635__bF_buf0), .Y(w_mem_inst__abc_19396_new_n1988_));
NAND3X1 NAND3X1_289 ( .A(w_mem_inst__abc_19396_new_n1987_), .B(w_mem_inst__abc_19396_new_n1988_), .C(w_mem_inst__abc_19396_new_n1989_), .Y(w_mem_inst__abc_19396_new_n1990_));
NAND3X1 NAND3X1_29 ( .A(_abc_15497_new_n2892_), .B(_abc_15497_new_n2893_), .C(_abc_15497_new_n2756__bF_buf3), .Y(_abc_15497_new_n2894_));
NAND3X1 NAND3X1_290 ( .A(w_mem_inst_w_mem_13__15_), .B(w_mem_inst__abc_19396_new_n1617__bF_buf1), .C(w_mem_inst__abc_19396_new_n1594__bF_buf0), .Y(w_mem_inst__abc_19396_new_n2005_));
NAND3X1 NAND3X1_291 ( .A(w_mem_inst_w_mem_12__15_), .B(w_mem_inst__abc_19396_new_n1619__bF_buf3), .C(w_mem_inst__abc_19396_new_n1617__bF_buf0), .Y(w_mem_inst__abc_19396_new_n2007_));
NAND3X1 NAND3X1_292 ( .A(w_mem_inst__abc_19396_new_n2007_), .B(w_mem_inst__abc_19396_new_n2006_), .C(w_mem_inst__abc_19396_new_n2005_), .Y(w_mem_inst__abc_19396_new_n2008_));
NAND3X1 NAND3X1_293 ( .A(w_mem_inst_w_mem_1__15_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf0), .C(w_mem_inst__abc_19396_new_n1594__bF_buf7), .Y(w_mem_inst__abc_19396_new_n2012_));
NAND3X1 NAND3X1_294 ( .A(w_mem_inst_w_mem_2__15_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf7), .C(w_mem_inst__abc_19396_new_n1635__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2013_));
NAND3X1 NAND3X1_295 ( .A(w_mem_inst__abc_19396_new_n2012_), .B(w_mem_inst__abc_19396_new_n2013_), .C(w_mem_inst__abc_19396_new_n2014_), .Y(w_mem_inst__abc_19396_new_n2015_));
NAND3X1 NAND3X1_296 ( .A(w_mem_inst_w_mem_13__16_), .B(w_mem_inst__abc_19396_new_n1617__bF_buf7), .C(w_mem_inst__abc_19396_new_n1594__bF_buf6), .Y(w_mem_inst__abc_19396_new_n2030_));
NAND3X1 NAND3X1_297 ( .A(w_mem_inst_w_mem_12__16_), .B(w_mem_inst__abc_19396_new_n1619__bF_buf2), .C(w_mem_inst__abc_19396_new_n1617__bF_buf6), .Y(w_mem_inst__abc_19396_new_n2032_));
NAND3X1 NAND3X1_298 ( .A(w_mem_inst__abc_19396_new_n2032_), .B(w_mem_inst__abc_19396_new_n2031_), .C(w_mem_inst__abc_19396_new_n2030_), .Y(w_mem_inst__abc_19396_new_n2033_));
NAND3X1 NAND3X1_299 ( .A(w_mem_inst_w_mem_1__16_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf6), .C(w_mem_inst__abc_19396_new_n1594__bF_buf5), .Y(w_mem_inst__abc_19396_new_n2037_));
NAND3X1 NAND3X1_3 ( .A(_abc_15497_new_n1746_), .B(_abc_15497_new_n1748_), .C(_abc_15497_new_n1747_), .Y(_0e_reg_31_0__31_));
NAND3X1 NAND3X1_30 ( .A(_abc_15497_new_n2898_), .B(_abc_15497_new_n2902_), .C(_abc_15497_new_n2905_), .Y(_abc_15497_new_n2906_));
NAND3X1 NAND3X1_300 ( .A(w_mem_inst_w_mem_2__16_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf5), .C(w_mem_inst__abc_19396_new_n1635__bF_buf3), .Y(w_mem_inst__abc_19396_new_n2038_));
NAND3X1 NAND3X1_301 ( .A(w_mem_inst__abc_19396_new_n2037_), .B(w_mem_inst__abc_19396_new_n2038_), .C(w_mem_inst__abc_19396_new_n2039_), .Y(w_mem_inst__abc_19396_new_n2040_));
NAND3X1 NAND3X1_302 ( .A(w_mem_inst_w_mem_13__17_), .B(w_mem_inst__abc_19396_new_n1617__bF_buf5), .C(w_mem_inst__abc_19396_new_n1594__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2055_));
NAND3X1 NAND3X1_303 ( .A(w_mem_inst_w_mem_12__17_), .B(w_mem_inst__abc_19396_new_n1619__bF_buf1), .C(w_mem_inst__abc_19396_new_n1617__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2057_));
NAND3X1 NAND3X1_304 ( .A(w_mem_inst__abc_19396_new_n2057_), .B(w_mem_inst__abc_19396_new_n2056_), .C(w_mem_inst__abc_19396_new_n2055_), .Y(w_mem_inst__abc_19396_new_n2058_));
NAND3X1 NAND3X1_305 ( .A(w_mem_inst_w_mem_1__17_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf4), .C(w_mem_inst__abc_19396_new_n1594__bF_buf3), .Y(w_mem_inst__abc_19396_new_n2062_));
NAND3X1 NAND3X1_306 ( .A(w_mem_inst_w_mem_2__17_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf3), .C(w_mem_inst__abc_19396_new_n1635__bF_buf2), .Y(w_mem_inst__abc_19396_new_n2063_));
NAND3X1 NAND3X1_307 ( .A(w_mem_inst__abc_19396_new_n2062_), .B(w_mem_inst__abc_19396_new_n2063_), .C(w_mem_inst__abc_19396_new_n2064_), .Y(w_mem_inst__abc_19396_new_n2065_));
NAND3X1 NAND3X1_308 ( .A(w_mem_inst_w_mem_13__18_), .B(w_mem_inst__abc_19396_new_n1617__bF_buf3), .C(w_mem_inst__abc_19396_new_n1594__bF_buf2), .Y(w_mem_inst__abc_19396_new_n2080_));
NAND3X1 NAND3X1_309 ( .A(w_mem_inst_w_mem_12__18_), .B(w_mem_inst__abc_19396_new_n1619__bF_buf0), .C(w_mem_inst__abc_19396_new_n1617__bF_buf2), .Y(w_mem_inst__abc_19396_new_n2082_));
NAND3X1 NAND3X1_31 ( .A(_abc_15497_new_n2907_), .B(_abc_15497_new_n2902_), .C(_abc_15497_new_n2905_), .Y(_abc_15497_new_n2913_));
NAND3X1 NAND3X1_310 ( .A(w_mem_inst__abc_19396_new_n2082_), .B(w_mem_inst__abc_19396_new_n2081_), .C(w_mem_inst__abc_19396_new_n2080_), .Y(w_mem_inst__abc_19396_new_n2083_));
NAND3X1 NAND3X1_311 ( .A(w_mem_inst_w_mem_1__18_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf2), .C(w_mem_inst__abc_19396_new_n1594__bF_buf1), .Y(w_mem_inst__abc_19396_new_n2087_));
NAND3X1 NAND3X1_312 ( .A(w_mem_inst_w_mem_2__18_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf1), .C(w_mem_inst__abc_19396_new_n1635__bF_buf1), .Y(w_mem_inst__abc_19396_new_n2088_));
NAND3X1 NAND3X1_313 ( .A(w_mem_inst__abc_19396_new_n2087_), .B(w_mem_inst__abc_19396_new_n2088_), .C(w_mem_inst__abc_19396_new_n2089_), .Y(w_mem_inst__abc_19396_new_n2090_));
NAND3X1 NAND3X1_314 ( .A(w_mem_inst_w_mem_13__19_), .B(w_mem_inst__abc_19396_new_n1617__bF_buf1), .C(w_mem_inst__abc_19396_new_n1594__bF_buf0), .Y(w_mem_inst__abc_19396_new_n2105_));
NAND3X1 NAND3X1_315 ( .A(w_mem_inst_w_mem_12__19_), .B(w_mem_inst__abc_19396_new_n1619__bF_buf4), .C(w_mem_inst__abc_19396_new_n1617__bF_buf0), .Y(w_mem_inst__abc_19396_new_n2107_));
NAND3X1 NAND3X1_316 ( .A(w_mem_inst__abc_19396_new_n2107_), .B(w_mem_inst__abc_19396_new_n2106_), .C(w_mem_inst__abc_19396_new_n2105_), .Y(w_mem_inst__abc_19396_new_n2108_));
NAND3X1 NAND3X1_317 ( .A(w_mem_inst_w_mem_1__19_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf0), .C(w_mem_inst__abc_19396_new_n1594__bF_buf7), .Y(w_mem_inst__abc_19396_new_n2112_));
NAND3X1 NAND3X1_318 ( .A(w_mem_inst_w_mem_2__19_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf7), .C(w_mem_inst__abc_19396_new_n1635__bF_buf0), .Y(w_mem_inst__abc_19396_new_n2113_));
NAND3X1 NAND3X1_319 ( .A(w_mem_inst__abc_19396_new_n2112_), .B(w_mem_inst__abc_19396_new_n2113_), .C(w_mem_inst__abc_19396_new_n2114_), .Y(w_mem_inst__abc_19396_new_n2115_));
NAND3X1 NAND3X1_32 ( .A(_abc_15497_new_n2919_), .B(_abc_15497_new_n2920_), .C(_abc_15497_new_n2918_), .Y(_abc_15497_new_n2926_));
NAND3X1 NAND3X1_320 ( .A(w_mem_inst_w_mem_13__20_), .B(w_mem_inst__abc_19396_new_n1617__bF_buf7), .C(w_mem_inst__abc_19396_new_n1594__bF_buf6), .Y(w_mem_inst__abc_19396_new_n2130_));
NAND3X1 NAND3X1_321 ( .A(w_mem_inst_w_mem_12__20_), .B(w_mem_inst__abc_19396_new_n1619__bF_buf3), .C(w_mem_inst__abc_19396_new_n1617__bF_buf6), .Y(w_mem_inst__abc_19396_new_n2132_));
NAND3X1 NAND3X1_322 ( .A(w_mem_inst__abc_19396_new_n2132_), .B(w_mem_inst__abc_19396_new_n2131_), .C(w_mem_inst__abc_19396_new_n2130_), .Y(w_mem_inst__abc_19396_new_n2133_));
NAND3X1 NAND3X1_323 ( .A(w_mem_inst_w_mem_1__20_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf6), .C(w_mem_inst__abc_19396_new_n1594__bF_buf5), .Y(w_mem_inst__abc_19396_new_n2137_));
NAND3X1 NAND3X1_324 ( .A(w_mem_inst_w_mem_2__20_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf5), .C(w_mem_inst__abc_19396_new_n1635__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2138_));
NAND3X1 NAND3X1_325 ( .A(w_mem_inst__abc_19396_new_n2137_), .B(w_mem_inst__abc_19396_new_n2138_), .C(w_mem_inst__abc_19396_new_n2139_), .Y(w_mem_inst__abc_19396_new_n2140_));
NAND3X1 NAND3X1_326 ( .A(w_mem_inst_w_mem_13__21_), .B(w_mem_inst__abc_19396_new_n1617__bF_buf5), .C(w_mem_inst__abc_19396_new_n1594__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2155_));
NAND3X1 NAND3X1_327 ( .A(w_mem_inst_w_mem_12__21_), .B(w_mem_inst__abc_19396_new_n1619__bF_buf2), .C(w_mem_inst__abc_19396_new_n1617__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2157_));
NAND3X1 NAND3X1_328 ( .A(w_mem_inst__abc_19396_new_n2157_), .B(w_mem_inst__abc_19396_new_n2156_), .C(w_mem_inst__abc_19396_new_n2155_), .Y(w_mem_inst__abc_19396_new_n2158_));
NAND3X1 NAND3X1_329 ( .A(w_mem_inst_w_mem_1__21_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf4), .C(w_mem_inst__abc_19396_new_n1594__bF_buf3), .Y(w_mem_inst__abc_19396_new_n2162_));
NAND3X1 NAND3X1_33 ( .A(_abc_15497_new_n2888_), .B(_abc_15497_new_n2911_), .C(_abc_15497_new_n2916_), .Y(_abc_15497_new_n2927_));
NAND3X1 NAND3X1_330 ( .A(w_mem_inst_w_mem_2__21_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf3), .C(w_mem_inst__abc_19396_new_n1635__bF_buf3), .Y(w_mem_inst__abc_19396_new_n2163_));
NAND3X1 NAND3X1_331 ( .A(w_mem_inst__abc_19396_new_n2162_), .B(w_mem_inst__abc_19396_new_n2163_), .C(w_mem_inst__abc_19396_new_n2164_), .Y(w_mem_inst__abc_19396_new_n2165_));
NAND3X1 NAND3X1_332 ( .A(w_mem_inst_w_mem_13__22_), .B(w_mem_inst__abc_19396_new_n1617__bF_buf3), .C(w_mem_inst__abc_19396_new_n1594__bF_buf2), .Y(w_mem_inst__abc_19396_new_n2180_));
NAND3X1 NAND3X1_333 ( .A(w_mem_inst_w_mem_12__22_), .B(w_mem_inst__abc_19396_new_n1619__bF_buf1), .C(w_mem_inst__abc_19396_new_n1617__bF_buf2), .Y(w_mem_inst__abc_19396_new_n2182_));
NAND3X1 NAND3X1_334 ( .A(w_mem_inst__abc_19396_new_n2182_), .B(w_mem_inst__abc_19396_new_n2181_), .C(w_mem_inst__abc_19396_new_n2180_), .Y(w_mem_inst__abc_19396_new_n2183_));
NAND3X1 NAND3X1_335 ( .A(w_mem_inst_w_mem_1__22_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf2), .C(w_mem_inst__abc_19396_new_n1594__bF_buf1), .Y(w_mem_inst__abc_19396_new_n2187_));
NAND3X1 NAND3X1_336 ( .A(w_mem_inst_w_mem_2__22_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf1), .C(w_mem_inst__abc_19396_new_n1635__bF_buf2), .Y(w_mem_inst__abc_19396_new_n2188_));
NAND3X1 NAND3X1_337 ( .A(w_mem_inst__abc_19396_new_n2187_), .B(w_mem_inst__abc_19396_new_n2188_), .C(w_mem_inst__abc_19396_new_n2189_), .Y(w_mem_inst__abc_19396_new_n2190_));
NAND3X1 NAND3X1_338 ( .A(w_mem_inst_w_mem_13__23_), .B(w_mem_inst__abc_19396_new_n1617__bF_buf1), .C(w_mem_inst__abc_19396_new_n1594__bF_buf0), .Y(w_mem_inst__abc_19396_new_n2205_));
NAND3X1 NAND3X1_339 ( .A(w_mem_inst_w_mem_12__23_), .B(w_mem_inst__abc_19396_new_n1619__bF_buf0), .C(w_mem_inst__abc_19396_new_n1617__bF_buf0), .Y(w_mem_inst__abc_19396_new_n2207_));
NAND3X1 NAND3X1_34 ( .A(_abc_15497_new_n2925__bF_buf3), .B(_abc_15497_new_n2927_), .C(_abc_15497_new_n2926_), .Y(_abc_15497_new_n2928_));
NAND3X1 NAND3X1_340 ( .A(w_mem_inst__abc_19396_new_n2207_), .B(w_mem_inst__abc_19396_new_n2206_), .C(w_mem_inst__abc_19396_new_n2205_), .Y(w_mem_inst__abc_19396_new_n2208_));
NAND3X1 NAND3X1_341 ( .A(w_mem_inst_w_mem_1__23_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf0), .C(w_mem_inst__abc_19396_new_n1594__bF_buf7), .Y(w_mem_inst__abc_19396_new_n2212_));
NAND3X1 NAND3X1_342 ( .A(w_mem_inst_w_mem_2__23_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf7), .C(w_mem_inst__abc_19396_new_n1635__bF_buf1), .Y(w_mem_inst__abc_19396_new_n2213_));
NAND3X1 NAND3X1_343 ( .A(w_mem_inst__abc_19396_new_n2212_), .B(w_mem_inst__abc_19396_new_n2213_), .C(w_mem_inst__abc_19396_new_n2214_), .Y(w_mem_inst__abc_19396_new_n2215_));
NAND3X1 NAND3X1_344 ( .A(w_mem_inst_w_mem_13__24_), .B(w_mem_inst__abc_19396_new_n1617__bF_buf7), .C(w_mem_inst__abc_19396_new_n1594__bF_buf6), .Y(w_mem_inst__abc_19396_new_n2230_));
NAND3X1 NAND3X1_345 ( .A(w_mem_inst_w_mem_12__24_), .B(w_mem_inst__abc_19396_new_n1619__bF_buf4), .C(w_mem_inst__abc_19396_new_n1617__bF_buf6), .Y(w_mem_inst__abc_19396_new_n2232_));
NAND3X1 NAND3X1_346 ( .A(w_mem_inst__abc_19396_new_n2232_), .B(w_mem_inst__abc_19396_new_n2231_), .C(w_mem_inst__abc_19396_new_n2230_), .Y(w_mem_inst__abc_19396_new_n2233_));
NAND3X1 NAND3X1_347 ( .A(w_mem_inst_w_mem_1__24_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf6), .C(w_mem_inst__abc_19396_new_n1594__bF_buf5), .Y(w_mem_inst__abc_19396_new_n2237_));
NAND3X1 NAND3X1_348 ( .A(w_mem_inst_w_mem_2__24_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf5), .C(w_mem_inst__abc_19396_new_n1635__bF_buf0), .Y(w_mem_inst__abc_19396_new_n2238_));
NAND3X1 NAND3X1_349 ( .A(w_mem_inst__abc_19396_new_n2237_), .B(w_mem_inst__abc_19396_new_n2238_), .C(w_mem_inst__abc_19396_new_n2239_), .Y(w_mem_inst__abc_19396_new_n2240_));
NAND3X1 NAND3X1_35 ( .A(_abc_15497_new_n2928_), .B(_abc_15497_new_n2922_), .C(_abc_15497_new_n2886_), .Y(_abc_15497_new_n2929_));
NAND3X1 NAND3X1_350 ( .A(w_mem_inst_w_mem_13__25_), .B(w_mem_inst__abc_19396_new_n1617__bF_buf5), .C(w_mem_inst__abc_19396_new_n1594__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2255_));
NAND3X1 NAND3X1_351 ( .A(w_mem_inst_w_mem_12__25_), .B(w_mem_inst__abc_19396_new_n1619__bF_buf3), .C(w_mem_inst__abc_19396_new_n1617__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2257_));
NAND3X1 NAND3X1_352 ( .A(w_mem_inst__abc_19396_new_n2257_), .B(w_mem_inst__abc_19396_new_n2256_), .C(w_mem_inst__abc_19396_new_n2255_), .Y(w_mem_inst__abc_19396_new_n2258_));
NAND3X1 NAND3X1_353 ( .A(w_mem_inst_w_mem_1__25_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf4), .C(w_mem_inst__abc_19396_new_n1594__bF_buf3), .Y(w_mem_inst__abc_19396_new_n2262_));
NAND3X1 NAND3X1_354 ( .A(w_mem_inst_w_mem_2__25_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf3), .C(w_mem_inst__abc_19396_new_n1635__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2263_));
NAND3X1 NAND3X1_355 ( .A(w_mem_inst__abc_19396_new_n2262_), .B(w_mem_inst__abc_19396_new_n2263_), .C(w_mem_inst__abc_19396_new_n2264_), .Y(w_mem_inst__abc_19396_new_n2265_));
NAND3X1 NAND3X1_356 ( .A(w_mem_inst_w_mem_13__26_), .B(w_mem_inst__abc_19396_new_n1617__bF_buf3), .C(w_mem_inst__abc_19396_new_n1594__bF_buf2), .Y(w_mem_inst__abc_19396_new_n2280_));
NAND3X1 NAND3X1_357 ( .A(w_mem_inst_w_mem_12__26_), .B(w_mem_inst__abc_19396_new_n1619__bF_buf2), .C(w_mem_inst__abc_19396_new_n1617__bF_buf2), .Y(w_mem_inst__abc_19396_new_n2282_));
NAND3X1 NAND3X1_358 ( .A(w_mem_inst__abc_19396_new_n2282_), .B(w_mem_inst__abc_19396_new_n2281_), .C(w_mem_inst__abc_19396_new_n2280_), .Y(w_mem_inst__abc_19396_new_n2283_));
NAND3X1 NAND3X1_359 ( .A(w_mem_inst_w_mem_1__26_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf2), .C(w_mem_inst__abc_19396_new_n1594__bF_buf1), .Y(w_mem_inst__abc_19396_new_n2287_));
NAND3X1 NAND3X1_36 ( .A(_abc_15497_new_n2911_), .B(_abc_15497_new_n2916_), .C(_abc_15497_new_n2918_), .Y(_abc_15497_new_n2931_));
NAND3X1 NAND3X1_360 ( .A(w_mem_inst_w_mem_2__26_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf1), .C(w_mem_inst__abc_19396_new_n1635__bF_buf3), .Y(w_mem_inst__abc_19396_new_n2288_));
NAND3X1 NAND3X1_361 ( .A(w_mem_inst__abc_19396_new_n2287_), .B(w_mem_inst__abc_19396_new_n2288_), .C(w_mem_inst__abc_19396_new_n2289_), .Y(w_mem_inst__abc_19396_new_n2290_));
NAND3X1 NAND3X1_362 ( .A(w_mem_inst_w_mem_13__27_), .B(w_mem_inst__abc_19396_new_n1617__bF_buf1), .C(w_mem_inst__abc_19396_new_n1594__bF_buf0), .Y(w_mem_inst__abc_19396_new_n2305_));
NAND3X1 NAND3X1_363 ( .A(w_mem_inst_w_mem_12__27_), .B(w_mem_inst__abc_19396_new_n1619__bF_buf1), .C(w_mem_inst__abc_19396_new_n1617__bF_buf0), .Y(w_mem_inst__abc_19396_new_n2307_));
NAND3X1 NAND3X1_364 ( .A(w_mem_inst__abc_19396_new_n2307_), .B(w_mem_inst__abc_19396_new_n2306_), .C(w_mem_inst__abc_19396_new_n2305_), .Y(w_mem_inst__abc_19396_new_n2308_));
NAND3X1 NAND3X1_365 ( .A(w_mem_inst_w_mem_1__27_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf0), .C(w_mem_inst__abc_19396_new_n1594__bF_buf7), .Y(w_mem_inst__abc_19396_new_n2312_));
NAND3X1 NAND3X1_366 ( .A(w_mem_inst_w_mem_2__27_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf7), .C(w_mem_inst__abc_19396_new_n1635__bF_buf2), .Y(w_mem_inst__abc_19396_new_n2313_));
NAND3X1 NAND3X1_367 ( .A(w_mem_inst__abc_19396_new_n2312_), .B(w_mem_inst__abc_19396_new_n2313_), .C(w_mem_inst__abc_19396_new_n2314_), .Y(w_mem_inst__abc_19396_new_n2315_));
NAND3X1 NAND3X1_368 ( .A(w_mem_inst_w_mem_13__28_), .B(w_mem_inst__abc_19396_new_n1617__bF_buf7), .C(w_mem_inst__abc_19396_new_n1594__bF_buf6), .Y(w_mem_inst__abc_19396_new_n2330_));
NAND3X1 NAND3X1_369 ( .A(w_mem_inst_w_mem_12__28_), .B(w_mem_inst__abc_19396_new_n1619__bF_buf0), .C(w_mem_inst__abc_19396_new_n1617__bF_buf6), .Y(w_mem_inst__abc_19396_new_n2332_));
NAND3X1 NAND3X1_37 ( .A(_abc_15497_new_n2888_), .B(_abc_15497_new_n2919_), .C(_abc_15497_new_n2920_), .Y(_abc_15497_new_n2932_));
NAND3X1 NAND3X1_370 ( .A(w_mem_inst__abc_19396_new_n2332_), .B(w_mem_inst__abc_19396_new_n2331_), .C(w_mem_inst__abc_19396_new_n2330_), .Y(w_mem_inst__abc_19396_new_n2333_));
NAND3X1 NAND3X1_371 ( .A(w_mem_inst_w_mem_1__28_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf6), .C(w_mem_inst__abc_19396_new_n1594__bF_buf5), .Y(w_mem_inst__abc_19396_new_n2337_));
NAND3X1 NAND3X1_372 ( .A(w_mem_inst_w_mem_2__28_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf5), .C(w_mem_inst__abc_19396_new_n1635__bF_buf1), .Y(w_mem_inst__abc_19396_new_n2338_));
NAND3X1 NAND3X1_373 ( .A(w_mem_inst__abc_19396_new_n2337_), .B(w_mem_inst__abc_19396_new_n2338_), .C(w_mem_inst__abc_19396_new_n2339_), .Y(w_mem_inst__abc_19396_new_n2340_));
NAND3X1 NAND3X1_374 ( .A(w_mem_inst_w_mem_13__29_), .B(w_mem_inst__abc_19396_new_n1617__bF_buf5), .C(w_mem_inst__abc_19396_new_n1594__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2355_));
NAND3X1 NAND3X1_375 ( .A(w_mem_inst_w_mem_12__29_), .B(w_mem_inst__abc_19396_new_n1619__bF_buf4), .C(w_mem_inst__abc_19396_new_n1617__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2357_));
NAND3X1 NAND3X1_376 ( .A(w_mem_inst__abc_19396_new_n2357_), .B(w_mem_inst__abc_19396_new_n2356_), .C(w_mem_inst__abc_19396_new_n2355_), .Y(w_mem_inst__abc_19396_new_n2358_));
NAND3X1 NAND3X1_377 ( .A(w_mem_inst_w_mem_1__29_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf4), .C(w_mem_inst__abc_19396_new_n1594__bF_buf3), .Y(w_mem_inst__abc_19396_new_n2362_));
NAND3X1 NAND3X1_378 ( .A(w_mem_inst_w_mem_2__29_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf3), .C(w_mem_inst__abc_19396_new_n1635__bF_buf0), .Y(w_mem_inst__abc_19396_new_n2363_));
NAND3X1 NAND3X1_379 ( .A(w_mem_inst__abc_19396_new_n2362_), .B(w_mem_inst__abc_19396_new_n2363_), .C(w_mem_inst__abc_19396_new_n2364_), .Y(w_mem_inst__abc_19396_new_n2365_));
NAND3X1 NAND3X1_38 ( .A(_abc_15497_new_n2736_), .B(_abc_15497_new_n2863_), .C(_abc_15497_new_n2742__bF_buf1), .Y(_abc_15497_new_n2944_));
NAND3X1 NAND3X1_380 ( .A(w_mem_inst_w_mem_13__30_), .B(w_mem_inst__abc_19396_new_n1617__bF_buf3), .C(w_mem_inst__abc_19396_new_n1594__bF_buf2), .Y(w_mem_inst__abc_19396_new_n2380_));
NAND3X1 NAND3X1_381 ( .A(w_mem_inst_w_mem_12__30_), .B(w_mem_inst__abc_19396_new_n1619__bF_buf3), .C(w_mem_inst__abc_19396_new_n1617__bF_buf2), .Y(w_mem_inst__abc_19396_new_n2382_));
NAND3X1 NAND3X1_382 ( .A(w_mem_inst__abc_19396_new_n2382_), .B(w_mem_inst__abc_19396_new_n2381_), .C(w_mem_inst__abc_19396_new_n2380_), .Y(w_mem_inst__abc_19396_new_n2383_));
NAND3X1 NAND3X1_383 ( .A(w_mem_inst_w_mem_1__30_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf2), .C(w_mem_inst__abc_19396_new_n1594__bF_buf1), .Y(w_mem_inst__abc_19396_new_n2387_));
NAND3X1 NAND3X1_384 ( .A(w_mem_inst_w_mem_2__30_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf1), .C(w_mem_inst__abc_19396_new_n1635__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2388_));
NAND3X1 NAND3X1_385 ( .A(w_mem_inst__abc_19396_new_n2387_), .B(w_mem_inst__abc_19396_new_n2388_), .C(w_mem_inst__abc_19396_new_n2389_), .Y(w_mem_inst__abc_19396_new_n2390_));
NAND3X1 NAND3X1_386 ( .A(w_mem_inst_w_mem_13__31_), .B(w_mem_inst__abc_19396_new_n1617__bF_buf1), .C(w_mem_inst__abc_19396_new_n1594__bF_buf0), .Y(w_mem_inst__abc_19396_new_n2405_));
NAND3X1 NAND3X1_387 ( .A(w_mem_inst_w_mem_12__31_), .B(w_mem_inst__abc_19396_new_n1619__bF_buf2), .C(w_mem_inst__abc_19396_new_n1617__bF_buf0), .Y(w_mem_inst__abc_19396_new_n2407_));
NAND3X1 NAND3X1_388 ( .A(w_mem_inst__abc_19396_new_n2407_), .B(w_mem_inst__abc_19396_new_n2406_), .C(w_mem_inst__abc_19396_new_n2405_), .Y(w_mem_inst__abc_19396_new_n2408_));
NAND3X1 NAND3X1_389 ( .A(w_mem_inst_w_mem_1__31_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf0), .C(w_mem_inst__abc_19396_new_n1594__bF_buf7), .Y(w_mem_inst__abc_19396_new_n2412_));
NAND3X1 NAND3X1_39 ( .A(w_4_), .B(_abc_15497_new_n2959_), .C(_abc_15497_new_n2962_), .Y(_abc_15497_new_n2963_));
NAND3X1 NAND3X1_390 ( .A(w_mem_inst_w_mem_2__31_), .B(w_mem_inst__abc_19396_new_n1620__bF_buf7), .C(w_mem_inst__abc_19396_new_n1635__bF_buf3), .Y(w_mem_inst__abc_19396_new_n2413_));
NAND3X1 NAND3X1_391 ( .A(w_mem_inst__abc_19396_new_n2412_), .B(w_mem_inst__abc_19396_new_n2413_), .C(w_mem_inst__abc_19396_new_n2414_), .Y(w_mem_inst__abc_19396_new_n2415_));
NAND3X1 NAND3X1_4 ( .A(_abc_15497_new_n2082_), .B(_abc_15497_new_n2083_), .C(_abc_15497_new_n2078_), .Y(_abc_15497_new_n2084_));
NAND3X1 NAND3X1_40 ( .A(_abc_15497_new_n2961_), .B(_abc_15497_new_n2963_), .C(_abc_15497_new_n2956_), .Y(_abc_15497_new_n2964_));
NAND3X1 NAND3X1_41 ( .A(_abc_15497_new_n2964_), .B(_abc_15497_new_n2968_), .C(_abc_15497_new_n2954_), .Y(_abc_15497_new_n2969_));
NAND3X1 NAND3X1_42 ( .A(_abc_15497_new_n2944_), .B(_abc_15497_new_n2984_), .C(_abc_15497_new_n2973_), .Y(_abc_15497_new_n2985_));
NAND3X1 NAND3X1_43 ( .A(_abc_15497_new_n2781__bF_buf1), .B(_abc_15497_new_n2986_), .C(_abc_15497_new_n2987_), .Y(_abc_15497_new_n2988_));
NAND3X1 NAND3X1_44 ( .A(_abc_15497_new_n2943_), .B(_abc_15497_new_n2985_), .C(_abc_15497_new_n2988_), .Y(_abc_15497_new_n2989_));
NAND3X1 NAND3X1_45 ( .A(_abc_15497_new_n2944_), .B(_abc_15497_new_n2986_), .C(_abc_15497_new_n2987_), .Y(_abc_15497_new_n2991_));
NAND3X1 NAND3X1_46 ( .A(_abc_15497_new_n2781__bF_buf0), .B(_abc_15497_new_n2984_), .C(_abc_15497_new_n2973_), .Y(_abc_15497_new_n2992_));
NAND3X1 NAND3X1_47 ( .A(_abc_15497_new_n2990_), .B(_abc_15497_new_n2991_), .C(_abc_15497_new_n2992_), .Y(_abc_15497_new_n2993_));
NAND3X1 NAND3X1_48 ( .A(w_5_), .B(_abc_15497_new_n3020_), .C(_abc_15497_new_n3023_), .Y(_abc_15497_new_n3024_));
NAND3X1 NAND3X1_49 ( .A(_abc_15497_new_n3017_), .B(_abc_15497_new_n3022_), .C(_abc_15497_new_n3024_), .Y(_abc_15497_new_n3025_));
NAND3X1 NAND3X1_5 ( .A(digest_update_bF_buf5), .B(_abc_15497_new_n2087_), .C(_abc_15497_new_n2084_), .Y(_abc_15497_new_n2088_));
NAND3X1 NAND3X1_50 ( .A(_abc_15497_new_n3038_), .B(_abc_15497_new_n3039_), .C(_abc_15497_new_n3037_), .Y(_abc_15497_new_n3042_));
NAND3X1 NAND3X1_51 ( .A(_abc_15497_new_n3031_), .B(_abc_15497_new_n3034_), .C(_abc_15497_new_n3007_), .Y(_abc_15497_new_n3043_));
NAND3X1 NAND3X1_52 ( .A(_abc_15497_new_n2781__bF_buf1), .B(_abc_15497_new_n3042_), .C(_abc_15497_new_n3043_), .Y(_abc_15497_new_n3044_));
NAND3X1 NAND3X1_53 ( .A(_abc_15497_new_n3044_), .B(_abc_15497_new_n3041_), .C(_abc_15497_new_n3006_), .Y(_abc_15497_new_n3045_));
NAND3X1 NAND3X1_54 ( .A(w_6_), .B(_abc_15497_new_n3078_), .C(_abc_15497_new_n3081_), .Y(_abc_15497_new_n3082_));
NAND3X1 NAND3X1_55 ( .A(_abc_15497_new_n3075_), .B(_abc_15497_new_n3080_), .C(_abc_15497_new_n3082_), .Y(_abc_15497_new_n3083_));
NAND3X1 NAND3X1_56 ( .A(_abc_15497_new_n3096_), .B(_abc_15497_new_n3097_), .C(_abc_15497_new_n3095_), .Y(_abc_15497_new_n3100_));
NAND3X1 NAND3X1_57 ( .A(_abc_15497_new_n3089_), .B(_abc_15497_new_n3092_), .C(_abc_15497_new_n3065_), .Y(_abc_15497_new_n3101_));
NAND3X1 NAND3X1_58 ( .A(_abc_15497_new_n2738_), .B(_abc_15497_new_n3100_), .C(_abc_15497_new_n3101_), .Y(_abc_15497_new_n3102_));
NAND3X1 NAND3X1_59 ( .A(_abc_15497_new_n3064_), .B(_abc_15497_new_n3102_), .C(_abc_15497_new_n3099_), .Y(_abc_15497_new_n3103_));
NAND3X1 NAND3X1_6 ( .A(_abc_15497_new_n2312_), .B(_abc_15497_new_n2324_), .C(_abc_15497_new_n2348_), .Y(_abc_15497_new_n2353_));
NAND3X1 NAND3X1_60 ( .A(_abc_15497_new_n3102_), .B(_abc_15497_new_n3099_), .C(_abc_15497_new_n3104_), .Y(_abc_15497_new_n3116_));
NAND3X1 NAND3X1_61 ( .A(d_reg_7_), .B(b_reg_7_), .C(c_reg_7_), .Y(_abc_15497_new_n3123_));
NAND3X1 NAND3X1_62 ( .A(w_7_), .B(_abc_15497_new_n3133_), .C(_abc_15497_new_n3136_), .Y(_abc_15497_new_n3137_));
NAND3X1 NAND3X1_63 ( .A(_abc_15497_new_n3130_), .B(_abc_15497_new_n3135_), .C(_abc_15497_new_n3137_), .Y(_abc_15497_new_n3138_));
NAND3X1 NAND3X1_64 ( .A(_abc_15497_new_n3135_), .B(_abc_15497_new_n3137_), .C(_abc_15497_new_n3139_), .Y(_abc_15497_new_n3148_));
NAND3X1 NAND3X1_65 ( .A(_abc_15497_new_n3101_), .B(_abc_15497_new_n3160_), .C(_abc_15497_new_n3102_), .Y(_abc_15497_new_n3161_));
NAND3X1 NAND3X1_66 ( .A(w_8_), .B(_abc_15497_new_n3181_), .C(_abc_15497_new_n3184_), .Y(_abc_15497_new_n3185_));
NAND3X1 NAND3X1_67 ( .A(_abc_15497_new_n3178_), .B(_abc_15497_new_n3183_), .C(_abc_15497_new_n3185_), .Y(_abc_15497_new_n3191_));
NAND3X1 NAND3X1_68 ( .A(_abc_15497_new_n3191_), .B(_abc_15497_new_n3193_), .C(_abc_15497_new_n3190_), .Y(_abc_15497_new_n3198_));
NAND3X1 NAND3X1_69 ( .A(_abc_15497_new_n3198_), .B(_abc_15497_new_n3201_), .C(_abc_15497_new_n3197_), .Y(_abc_15497_new_n3202_));
NAND3X1 NAND3X1_7 ( .A(_auto_iopadmap_cc_368_execute_22625_156_), .B(a_reg_28_), .C(_abc_15497_new_n2420_), .Y(_abc_15497_new_n2430_));
NAND3X1 NAND3X1_70 ( .A(_abc_15497_new_n2759__bF_buf2), .B(_abc_15497_new_n3202_), .C(_abc_15497_new_n3195_), .Y(_abc_15497_new_n3203_));
NAND3X1 NAND3X1_71 ( .A(_abc_15497_new_n3198_), .B(_abc_15497_new_n3201_), .C(_abc_15497_new_n3169_), .Y(_abc_15497_new_n3204_));
NAND3X1 NAND3X1_72 ( .A(_abc_15497_new_n2924__bF_buf1), .B(_abc_15497_new_n3204_), .C(_abc_15497_new_n3205_), .Y(_abc_15497_new_n3206_));
NAND3X1 NAND3X1_73 ( .A(_abc_15497_new_n3168_), .B(_abc_15497_new_n3203_), .C(_abc_15497_new_n3206_), .Y(_abc_15497_new_n3207_));
NAND3X1 NAND3X1_74 ( .A(_abc_15497_new_n2994_), .B(_abc_15497_new_n3212_), .C(_abc_15497_new_n3213_), .Y(_abc_15497_new_n3214_));
NAND3X1 NAND3X1_75 ( .A(_abc_15497_new_n3167_), .B(_abc_15497_new_n3203_), .C(_abc_15497_new_n3206_), .Y(_abc_15497_new_n3225_));
NAND3X1 NAND3X1_76 ( .A(w_9_), .B(_abc_15497_new_n3244_), .C(_abc_15497_new_n3247_), .Y(_abc_15497_new_n3248_));
NAND3X1 NAND3X1_77 ( .A(_abc_15497_new_n3241_), .B(_abc_15497_new_n3248_), .C(_abc_15497_new_n3246_), .Y(_abc_15497_new_n3259_));
NAND3X1 NAND3X1_78 ( .A(_abc_15497_new_n3191_), .B(_abc_15497_new_n3198_), .C(_abc_15497_new_n3270_), .Y(_abc_15497_new_n3271_));
NAND3X1 NAND3X1_79 ( .A(_abc_15497_new_n3253_), .B(_abc_15497_new_n3264_), .C(_abc_15497_new_n3230_), .Y(_abc_15497_new_n3272_));
NAND3X1 NAND3X1_8 ( .A(_auto_iopadmap_cc_368_execute_22625_63_), .B(_abc_15497_new_n1650__bF_buf4), .C(_abc_15497_new_n2634_), .Y(_abc_15497_new_n2635_));
NAND3X1 NAND3X1_80 ( .A(_abc_15497_new_n2781__bF_buf3), .B(_abc_15497_new_n3272_), .C(_abc_15497_new_n3271_), .Y(_abc_15497_new_n3273_));
NAND3X1 NAND3X1_81 ( .A(_abc_15497_new_n3229_), .B(_abc_15497_new_n3273_), .C(_abc_15497_new_n3269_), .Y(_abc_15497_new_n3274_));
NAND3X1 NAND3X1_82 ( .A(_abc_15497_new_n3274_), .B(_abc_15497_new_n3278_), .C(_abc_15497_new_n3211_), .Y(_abc_15497_new_n3285_));
NAND3X1 NAND3X1_83 ( .A(w_10_), .B(_abc_15497_new_n3304_), .C(_abc_15497_new_n3307_), .Y(_abc_15497_new_n3308_));
NAND3X1 NAND3X1_84 ( .A(_abc_15497_new_n3306_), .B(_abc_15497_new_n3308_), .C(_abc_15497_new_n3301_), .Y(_abc_15497_new_n3309_));
NAND3X1 NAND3X1_85 ( .A(_abc_15497_new_n3300_), .B(_abc_15497_new_n3306_), .C(_abc_15497_new_n3308_), .Y(_abc_15497_new_n3319_));
NAND3X1 NAND3X1_86 ( .A(_abc_15497_new_n3324_), .B(_abc_15497_new_n3325_), .C(_abc_15497_new_n3332_), .Y(_abc_15497_new_n3333_));
NAND3X1 NAND3X1_87 ( .A(_abc_15497_new_n3314_), .B(_abc_15497_new_n3322_), .C(_abc_15497_new_n3289_), .Y(_abc_15497_new_n3334_));
NAND3X1 NAND3X1_88 ( .A(_abc_15497_new_n2759__bF_buf3), .B(_abc_15497_new_n3334_), .C(_abc_15497_new_n3333_), .Y(_abc_15497_new_n3335_));
NAND3X1 NAND3X1_89 ( .A(_abc_15497_new_n3327_), .B(_abc_15497_new_n3335_), .C(_abc_15497_new_n3288_), .Y(_abc_15497_new_n3336_));
NAND3X1 NAND3X1_9 ( .A(_abc_15497_new_n2637_), .B(_abc_15497_new_n2635_), .C(_abc_15497_new_n2636_), .Y(_0d_reg_31_0__31_));
NAND3X1 NAND3X1_90 ( .A(_abc_15497_new_n3327_), .B(_abc_15497_new_n3335_), .C(_abc_15497_new_n3337_), .Y(_abc_15497_new_n3348_));
NAND3X1 NAND3X1_91 ( .A(d_reg_11_), .B(b_reg_11_), .C(c_reg_11_), .Y(_abc_15497_new_n3355_));
NAND3X1 NAND3X1_92 ( .A(w_11_), .B(_abc_15497_new_n3366_), .C(_abc_15497_new_n3365_), .Y(_abc_15497_new_n3367_));
NAND3X1 NAND3X1_93 ( .A(_abc_15497_new_n3360_), .B(_abc_15497_new_n3364_), .C(_abc_15497_new_n3367_), .Y(_abc_15497_new_n3368_));
NAND3X1 NAND3X1_94 ( .A(_abc_15497_new_n3364_), .B(_abc_15497_new_n3367_), .C(_abc_15497_new_n3369_), .Y(_abc_15497_new_n3376_));
NAND3X1 NAND3X1_95 ( .A(_abc_15497_new_n2780__bF_buf0), .B(_abc_15497_new_n3385_), .C(_abc_15497_new_n3380_), .Y(_abc_15497_new_n3386_));
NAND3X1 NAND3X1_96 ( .A(_abc_15497_new_n2755_), .B(_abc_15497_new_n3387_), .C(_abc_15497_new_n3388_), .Y(_abc_15497_new_n3389_));
NAND3X1 NAND3X1_97 ( .A(_abc_15497_new_n3386_), .B(_abc_15497_new_n3389_), .C(_abc_15497_new_n3350_), .Y(_abc_15497_new_n3390_));
NAND3X1 NAND3X1_98 ( .A(round_ctr_reg_5_), .B(round_ctr_reg_4_), .C(_abc_15497_new_n3392_), .Y(_abc_15497_new_n3393_));
NAND3X1 NAND3X1_99 ( .A(_abc_15497_new_n3211_), .B(_abc_15497_new_n3279_), .C(_abc_15497_new_n3405_), .Y(_abc_15497_new_n3408_));
NOR2X1 NOR2X1_1 ( .A(c_reg_15_), .B(_auto_iopadmap_cc_368_execute_22625_79_), .Y(_abc_15497_new_n700_));
NOR2X1 NOR2X1_10 ( .A(_abc_15497_new_n719_), .B(_abc_15497_new_n711_), .Y(_abc_15497_new_n720_));
NOR2X1 NOR2X1_100 ( .A(e_reg_10_), .B(_auto_iopadmap_cc_368_execute_22625_10_), .Y(_abc_15497_new_n1039_));
NOR2X1 NOR2X1_101 ( .A(_abc_15497_new_n1043_), .B(_abc_15497_new_n1038_), .Y(_abc_15497_new_n1044_));
NOR2X1 NOR2X1_102 ( .A(e_reg_11_), .B(_auto_iopadmap_cc_368_execute_22625_11_), .Y(_abc_15497_new_n1051_));
NOR2X1 NOR2X1_103 ( .A(_abc_15497_new_n1054_), .B(_abc_15497_new_n1042_), .Y(_abc_15497_new_n1058_));
NOR2X1 NOR2X1_104 ( .A(e_reg_12_), .B(_auto_iopadmap_cc_368_execute_22625_12_), .Y(_abc_15497_new_n1063_));
NOR2X1 NOR2X1_105 ( .A(_abc_15497_new_n1064_), .B(_abc_15497_new_n1057_), .Y(_abc_15497_new_n1065_));
NOR2X1 NOR2X1_106 ( .A(_abc_15497_new_n1063_), .B(_abc_15497_new_n1065_), .Y(_abc_15497_new_n1066_));
NOR2X1 NOR2X1_107 ( .A(_abc_15497_new_n1066_), .B(_abc_15497_new_n1062_), .Y(_abc_15497_new_n1067_));
NOR2X1 NOR2X1_108 ( .A(e_reg_13_), .B(_auto_iopadmap_cc_368_execute_22625_13_), .Y(_abc_15497_new_n1072_));
NOR2X1 NOR2X1_109 ( .A(_abc_15497_new_n1072_), .B(_abc_15497_new_n1074_), .Y(_abc_15497_new_n1075_));
NOR2X1 NOR2X1_11 ( .A(_abc_15497_new_n721_), .B(_abc_15497_new_n718_), .Y(_abc_15497_new_n722_));
NOR2X1 NOR2X1_110 ( .A(e_reg_14_), .B(_auto_iopadmap_cc_368_execute_22625_14_), .Y(_abc_15497_new_n1079_));
NOR2X1 NOR2X1_111 ( .A(_abc_15497_new_n1080_), .B(_abc_15497_new_n1081_), .Y(_abc_15497_new_n1082_));
NOR2X1 NOR2X1_112 ( .A(_abc_15497_new_n1079_), .B(_abc_15497_new_n1082_), .Y(_abc_15497_new_n1083_));
NOR2X1 NOR2X1_113 ( .A(_abc_15497_new_n1083_), .B(_abc_15497_new_n1087_), .Y(_abc_15497_new_n1088_));
NOR2X1 NOR2X1_114 ( .A(e_reg_15_), .B(_auto_iopadmap_cc_368_execute_22625_15_), .Y(_abc_15497_new_n1094_));
NOR2X1 NOR2X1_115 ( .A(_abc_15497_new_n1094_), .B(_abc_15497_new_n1096_), .Y(_abc_15497_new_n1097_));
NOR2X1 NOR2X1_116 ( .A(_abc_15497_new_n1086_), .B(_abc_15497_new_n1103_), .Y(_abc_15497_new_n1104_));
NOR2X1 NOR2X1_117 ( .A(_abc_15497_new_n1026_), .B(_abc_15497_new_n1059_), .Y(_abc_15497_new_n1108_));
NOR2X1 NOR2X1_118 ( .A(e_reg_16_), .B(_auto_iopadmap_cc_368_execute_22625_16_), .Y(_abc_15497_new_n1111_));
NOR2X1 NOR2X1_119 ( .A(_abc_15497_new_n1112_), .B(_abc_15497_new_n1101_), .Y(_abc_15497_new_n1113_));
NOR2X1 NOR2X1_12 ( .A(_abc_15497_new_n707_), .B(_abc_15497_new_n723_), .Y(_abc_15497_new_n724_));
NOR2X1 NOR2X1_120 ( .A(_abc_15497_new_n1111_), .B(_abc_15497_new_n1113_), .Y(_abc_15497_new_n1114_));
NOR2X1 NOR2X1_121 ( .A(_abc_15497_new_n1114_), .B(_abc_15497_new_n1110_), .Y(_abc_15497_new_n1115_));
NOR2X1 NOR2X1_122 ( .A(e_reg_17_), .B(_auto_iopadmap_cc_368_execute_22625_17_), .Y(_abc_15497_new_n1120_));
NOR2X1 NOR2X1_123 ( .A(_abc_15497_new_n1121_), .B(_abc_15497_new_n1122_), .Y(_abc_15497_new_n1123_));
NOR2X1 NOR2X1_124 ( .A(_abc_15497_new_n1120_), .B(_abc_15497_new_n1123_), .Y(_abc_15497_new_n1124_));
NOR2X1 NOR2X1_125 ( .A(e_reg_18_), .B(_auto_iopadmap_cc_368_execute_22625_18_), .Y(_abc_15497_new_n1129_));
NOR2X1 NOR2X1_126 ( .A(_abc_15497_new_n1130_), .B(_abc_15497_new_n1128_), .Y(_abc_15497_new_n1131_));
NOR2X1 NOR2X1_127 ( .A(_abc_15497_new_n1129_), .B(_abc_15497_new_n1131_), .Y(_abc_15497_new_n1132_));
NOR2X1 NOR2X1_128 ( .A(e_reg_19_), .B(_auto_iopadmap_cc_368_execute_22625_19_), .Y(_abc_15497_new_n1145_));
NOR2X1 NOR2X1_129 ( .A(_abc_15497_new_n1146_), .B(_abc_15497_new_n1142_), .Y(_abc_15497_new_n1147_));
NOR2X1 NOR2X1_13 ( .A(_abc_15497_new_n727_), .B(_abc_15497_new_n728_), .Y(_abc_15497_new_n729_));
NOR2X1 NOR2X1_130 ( .A(_abc_15497_new_n1145_), .B(_abc_15497_new_n1147_), .Y(_abc_15497_new_n1148_));
NOR2X1 NOR2X1_131 ( .A(_abc_15497_new_n1156_), .B(_abc_15497_new_n1153_), .Y(_abc_15497_new_n1157_));
NOR2X1 NOR2X1_132 ( .A(e_reg_20_), .B(_auto_iopadmap_cc_368_execute_22625_20_), .Y(_abc_15497_new_n1161_));
NOR2X1 NOR2X1_133 ( .A(_abc_15497_new_n1162_), .B(_abc_15497_new_n1163_), .Y(_abc_15497_new_n1164_));
NOR2X1 NOR2X1_134 ( .A(_abc_15497_new_n1161_), .B(_abc_15497_new_n1164_), .Y(_abc_15497_new_n1165_));
NOR2X1 NOR2X1_135 ( .A(_abc_15497_new_n1165_), .B(_abc_15497_new_n1160_), .Y(_abc_15497_new_n1166_));
NOR2X1 NOR2X1_136 ( .A(e_reg_21_), .B(_auto_iopadmap_cc_368_execute_22625_21_), .Y(_abc_15497_new_n1172_));
NOR2X1 NOR2X1_137 ( .A(_abc_15497_new_n1173_), .B(_abc_15497_new_n1171_), .Y(_abc_15497_new_n1174_));
NOR2X1 NOR2X1_138 ( .A(_abc_15497_new_n1172_), .B(_abc_15497_new_n1174_), .Y(_abc_15497_new_n1175_));
NOR2X1 NOR2X1_139 ( .A(e_reg_22_), .B(_auto_iopadmap_cc_368_execute_22625_22_), .Y(_abc_15497_new_n1184_));
NOR2X1 NOR2X1_14 ( .A(c_reg_11_), .B(_auto_iopadmap_cc_368_execute_22625_75_), .Y(_abc_15497_new_n730_));
NOR2X1 NOR2X1_140 ( .A(_abc_15497_new_n1184_), .B(_abc_15497_new_n1186_), .Y(_abc_15497_new_n1187_));
NOR2X1 NOR2X1_141 ( .A(e_reg_23_), .B(_auto_iopadmap_cc_368_execute_22625_23_), .Y(_abc_15497_new_n1194_));
NOR2X1 NOR2X1_142 ( .A(_abc_15497_new_n1194_), .B(_abc_15497_new_n1196_), .Y(_abc_15497_new_n1197_));
NOR2X1 NOR2X1_143 ( .A(_abc_15497_new_n1201_), .B(_abc_15497_new_n1179_), .Y(_abc_15497_new_n1202_));
NOR2X1 NOR2X1_144 ( .A(_abc_15497_new_n1203_), .B(_abc_15497_new_n1155_), .Y(_abc_15497_new_n1204_));
NOR2X1 NOR2X1_145 ( .A(_abc_15497_new_n1207_), .B(_abc_15497_new_n1204_), .Y(_abc_15497_new_n1208_));
NOR2X1 NOR2X1_146 ( .A(e_reg_24_), .B(_auto_iopadmap_cc_368_execute_22625_24_), .Y(_abc_15497_new_n1212_));
NOR2X1 NOR2X1_147 ( .A(_abc_15497_new_n1213_), .B(_abc_15497_new_n1214_), .Y(_abc_15497_new_n1215_));
NOR2X1 NOR2X1_148 ( .A(_abc_15497_new_n1212_), .B(_abc_15497_new_n1215_), .Y(_abc_15497_new_n1216_));
NOR2X1 NOR2X1_149 ( .A(_abc_15497_new_n1216_), .B(_abc_15497_new_n1211_), .Y(_abc_15497_new_n1217_));
NOR2X1 NOR2X1_15 ( .A(_abc_15497_new_n730_), .B(_abc_15497_new_n726_), .Y(_abc_15497_new_n731_));
NOR2X1 NOR2X1_150 ( .A(e_reg_25_), .B(_auto_iopadmap_cc_368_execute_22625_25_), .Y(_abc_15497_new_n1224_));
NOR2X1 NOR2X1_151 ( .A(_abc_15497_new_n1224_), .B(_abc_15497_new_n1226_), .Y(_abc_15497_new_n1227_));
NOR2X1 NOR2X1_152 ( .A(_abc_15497_new_n1232_), .B(_abc_15497_new_n1218_), .Y(_abc_15497_new_n1233_));
NOR2X1 NOR2X1_153 ( .A(e_reg_26_), .B(_auto_iopadmap_cc_368_execute_22625_26_), .Y(_abc_15497_new_n1238_));
NOR2X1 NOR2X1_154 ( .A(_abc_15497_new_n1239_), .B(_abc_15497_new_n1231_), .Y(_abc_15497_new_n1240_));
NOR2X1 NOR2X1_155 ( .A(_abc_15497_new_n1238_), .B(_abc_15497_new_n1240_), .Y(_abc_15497_new_n1241_));
NOR2X1 NOR2X1_156 ( .A(_abc_15497_new_n1241_), .B(_abc_15497_new_n1237_), .Y(_abc_15497_new_n1242_));
NOR2X1 NOR2X1_157 ( .A(_abc_15497_new_n1244_), .B(_abc_15497_new_n1243_), .Y(_abc_15497_new_n1248_));
NOR2X1 NOR2X1_158 ( .A(e_reg_27_), .B(_auto_iopadmap_cc_368_execute_22625_27_), .Y(_abc_15497_new_n1249_));
NOR2X1 NOR2X1_159 ( .A(_abc_15497_new_n1250_), .B(_abc_15497_new_n1247_), .Y(_abc_15497_new_n1251_));
NOR2X1 NOR2X1_16 ( .A(c_reg_10_), .B(_auto_iopadmap_cc_368_execute_22625_74_), .Y(_abc_15497_new_n734_));
NOR2X1 NOR2X1_160 ( .A(_abc_15497_new_n1249_), .B(_abc_15497_new_n1251_), .Y(_abc_15497_new_n1252_));
NOR2X1 NOR2X1_161 ( .A(_abc_15497_new_n1253_), .B(_abc_15497_new_n1244_), .Y(_abc_15497_new_n1259_));
NOR2X1 NOR2X1_162 ( .A(_abc_15497_new_n1264_), .B(_abc_15497_new_n1263_), .Y(_abc_15497_new_n1265_));
NOR2X1 NOR2X1_163 ( .A(e_reg_29_), .B(_auto_iopadmap_cc_368_execute_22625_29_), .Y(_abc_15497_new_n1272_));
NOR2X1 NOR2X1_164 ( .A(_abc_15497_new_n1273_), .B(_abc_15497_new_n1274_), .Y(_abc_15497_new_n1275_));
NOR2X1 NOR2X1_165 ( .A(_abc_15497_new_n1272_), .B(_abc_15497_new_n1275_), .Y(_abc_15497_new_n1276_));
NOR2X1 NOR2X1_166 ( .A(_abc_15497_new_n1292_), .B(_abc_15497_new_n1291_), .Y(_abc_15497_new_n1293_));
NOR2X1 NOR2X1_167 ( .A(_abc_15497_new_n1298_), .B(_abc_15497_new_n1299_), .Y(_abc_15497_new_n1300_));
NOR2X1 NOR2X1_168 ( .A(_auto_iopadmap_cc_368_execute_22625_33_), .B(_abc_15497_new_n883__bF_buf8), .Y(_abc_15497_new_n1305_));
NOR2X1 NOR2X1_169 ( .A(_auto_iopadmap_cc_368_execute_22625_34_), .B(d_reg_2_), .Y(_abc_15497_new_n1311_));
NOR2X1 NOR2X1_17 ( .A(_abc_15497_new_n734_), .B(_abc_15497_new_n729_), .Y(_abc_15497_new_n735_));
NOR2X1 NOR2X1_170 ( .A(_abc_15497_new_n1311_), .B(_abc_15497_new_n1312_), .Y(_abc_15497_new_n1313_));
NOR2X1 NOR2X1_171 ( .A(_auto_iopadmap_cc_368_execute_22625_34_), .B(_abc_15497_new_n883__bF_buf7), .Y(_abc_15497_new_n1315_));
NOR2X1 NOR2X1_172 ( .A(_auto_iopadmap_cc_368_execute_22625_35_), .B(d_reg_3_), .Y(_abc_15497_new_n1319_));
NOR2X1 NOR2X1_173 ( .A(_abc_15497_new_n1317_), .B(_abc_15497_new_n1320_), .Y(_abc_15497_new_n1321_));
NOR2X1 NOR2X1_174 ( .A(_auto_iopadmap_cc_368_execute_22625_36_), .B(_abc_15497_new_n883__bF_buf6), .Y(_abc_15497_new_n1330_));
NOR2X1 NOR2X1_175 ( .A(_abc_15497_new_n1336_), .B(_abc_15497_new_n1335_), .Y(_abc_15497_new_n1337_));
NOR2X1 NOR2X1_176 ( .A(_abc_15497_new_n1345_), .B(_abc_15497_new_n1344_), .Y(_abc_15497_new_n1346_));
NOR2X1 NOR2X1_177 ( .A(_auto_iopadmap_cc_368_execute_22625_39_), .B(d_reg_7_), .Y(_abc_15497_new_n1352_));
NOR2X1 NOR2X1_178 ( .A(_abc_15497_new_n1351_), .B(_abc_15497_new_n1353_), .Y(_abc_15497_new_n1354_));
NOR2X1 NOR2X1_179 ( .A(_abc_15497_new_n1352_), .B(_abc_15497_new_n1354_), .Y(_abc_15497_new_n1355_));
NOR2X1 NOR2X1_18 ( .A(_abc_15497_new_n738_), .B(_abc_15497_new_n739_), .Y(_abc_15497_new_n740_));
NOR2X1 NOR2X1_180 ( .A(_auto_iopadmap_cc_368_execute_22625_40_), .B(d_reg_8_), .Y(_abc_15497_new_n1363_));
NOR2X1 NOR2X1_181 ( .A(_abc_15497_new_n1361_), .B(_abc_15497_new_n1364_), .Y(_abc_15497_new_n1365_));
NOR2X1 NOR2X1_182 ( .A(_abc_15497_new_n1363_), .B(_abc_15497_new_n1365_), .Y(_abc_15497_new_n1366_));
NOR2X1 NOR2X1_183 ( .A(_abc_15497_new_n1367_), .B(_abc_15497_new_n1362_), .Y(_abc_15497_new_n1372_));
NOR2X1 NOR2X1_184 ( .A(_auto_iopadmap_cc_368_execute_22625_41_), .B(d_reg_9_), .Y(_abc_15497_new_n1373_));
NOR2X1 NOR2X1_185 ( .A(_abc_15497_new_n1371_), .B(_abc_15497_new_n1374_), .Y(_abc_15497_new_n1375_));
NOR2X1 NOR2X1_186 ( .A(_abc_15497_new_n1373_), .B(_abc_15497_new_n1375_), .Y(_abc_15497_new_n1376_));
NOR2X1 NOR2X1_187 ( .A(_abc_15497_new_n1367_), .B(_abc_15497_new_n1377_), .Y(_abc_15497_new_n1382_));
NOR2X1 NOR2X1_188 ( .A(_auto_iopadmap_cc_368_execute_22625_42_), .B(d_reg_10_), .Y(_abc_15497_new_n1386_));
NOR2X1 NOR2X1_189 ( .A(_abc_15497_new_n1386_), .B(_abc_15497_new_n1388_), .Y(_abc_15497_new_n1389_));
NOR2X1 NOR2X1_19 ( .A(_abc_15497_new_n741_), .B(_abc_15497_new_n742_), .Y(_abc_15497_new_n743_));
NOR2X1 NOR2X1_190 ( .A(_abc_15497_new_n870__bF_buf5), .B(_abc_15497_new_n1390_), .Y(_abc_15497_new_n1391_));
NOR2X1 NOR2X1_191 ( .A(_abc_15497_new_n1388_), .B(_abc_15497_new_n1390_), .Y(_abc_15497_new_n1396_));
NOR2X1 NOR2X1_192 ( .A(_auto_iopadmap_cc_368_execute_22625_43_), .B(d_reg_11_), .Y(_abc_15497_new_n1397_));
NOR2X1 NOR2X1_193 ( .A(_abc_15497_new_n1395_), .B(_abc_15497_new_n1398_), .Y(_abc_15497_new_n1399_));
NOR2X1 NOR2X1_194 ( .A(_abc_15497_new_n1397_), .B(_abc_15497_new_n1399_), .Y(_abc_15497_new_n1400_));
NOR2X1 NOR2X1_195 ( .A(_abc_15497_new_n1405_), .B(_abc_15497_new_n1383_), .Y(_abc_15497_new_n1406_));
NOR2X1 NOR2X1_196 ( .A(_auto_iopadmap_cc_368_execute_22625_44_), .B(d_reg_12_), .Y(_abc_15497_new_n1412_));
NOR2X1 NOR2X1_197 ( .A(_abc_15497_new_n1413_), .B(_abc_15497_new_n1414_), .Y(_abc_15497_new_n1415_));
NOR2X1 NOR2X1_198 ( .A(_abc_15497_new_n1412_), .B(_abc_15497_new_n1415_), .Y(_abc_15497_new_n1416_));
NOR2X1 NOR2X1_199 ( .A(_abc_15497_new_n1416_), .B(_abc_15497_new_n1411_), .Y(_abc_15497_new_n1417_));
NOR2X1 NOR2X1_2 ( .A(_abc_15497_new_n700_), .B(_abc_15497_new_n699_), .Y(_abc_15497_new_n701_));
NOR2X1 NOR2X1_20 ( .A(c_reg_9_), .B(_auto_iopadmap_cc_368_execute_22625_73_), .Y(_abc_15497_new_n744_));
NOR2X1 NOR2X1_200 ( .A(_auto_iopadmap_cc_368_execute_22625_45_), .B(d_reg_13_), .Y(_abc_15497_new_n1424_));
NOR2X1 NOR2X1_201 ( .A(_abc_15497_new_n1422_), .B(_abc_15497_new_n1425_), .Y(_abc_15497_new_n1426_));
NOR2X1 NOR2X1_202 ( .A(_abc_15497_new_n1424_), .B(_abc_15497_new_n1426_), .Y(_abc_15497_new_n1427_));
NOR2X1 NOR2X1_203 ( .A(_auto_iopadmap_cc_368_execute_22625_46_), .B(d_reg_14_), .Y(_abc_15497_new_n1435_));
NOR2X1 NOR2X1_204 ( .A(_abc_15497_new_n1435_), .B(_abc_15497_new_n1437_), .Y(_abc_15497_new_n1438_));
NOR2X1 NOR2X1_205 ( .A(_auto_iopadmap_cc_368_execute_22625_47_), .B(d_reg_15_), .Y(_abc_15497_new_n1446_));
NOR2X1 NOR2X1_206 ( .A(_abc_15497_new_n1444_), .B(_abc_15497_new_n1447_), .Y(_abc_15497_new_n1448_));
NOR2X1 NOR2X1_207 ( .A(_abc_15497_new_n1446_), .B(_abc_15497_new_n1448_), .Y(_abc_15497_new_n1449_));
NOR2X1 NOR2X1_208 ( .A(_abc_15497_new_n1453_), .B(_abc_15497_new_n1456_), .Y(_abc_15497_new_n1457_));
NOR2X1 NOR2X1_209 ( .A(_auto_iopadmap_cc_368_execute_22625_48_), .B(d_reg_16_), .Y(_abc_15497_new_n1461_));
NOR2X1 NOR2X1_21 ( .A(_abc_15497_new_n744_), .B(_abc_15497_new_n740_), .Y(_abc_15497_new_n745_));
NOR2X1 NOR2X1_210 ( .A(_abc_15497_new_n1452_), .B(_abc_15497_new_n1462_), .Y(_abc_15497_new_n1463_));
NOR2X1 NOR2X1_211 ( .A(_abc_15497_new_n1461_), .B(_abc_15497_new_n1463_), .Y(_abc_15497_new_n1464_));
NOR2X1 NOR2X1_212 ( .A(_auto_iopadmap_cc_368_execute_22625_49_), .B(d_reg_17_), .Y(_abc_15497_new_n1468_));
NOR2X1 NOR2X1_213 ( .A(_abc_15497_new_n1468_), .B(_abc_15497_new_n1470_), .Y(_abc_15497_new_n1471_));
NOR2X1 NOR2X1_214 ( .A(_abc_15497_new_n1471_), .B(_abc_15497_new_n1467_), .Y(_abc_15497_new_n1473_));
NOR2X1 NOR2X1_215 ( .A(_auto_iopadmap_cc_368_execute_22625_50_), .B(d_reg_18_), .Y(_abc_15497_new_n1484_));
NOR2X1 NOR2X1_216 ( .A(_abc_15497_new_n1477_), .B(_abc_15497_new_n1485_), .Y(_abc_15497_new_n1486_));
NOR2X1 NOR2X1_217 ( .A(_abc_15497_new_n1484_), .B(_abc_15497_new_n1486_), .Y(_abc_15497_new_n1487_));
NOR2X1 NOR2X1_218 ( .A(_abc_15497_new_n1487_), .B(_abc_15497_new_n1483_), .Y(_abc_15497_new_n1488_));
NOR2X1 NOR2X1_219 ( .A(_auto_iopadmap_cc_368_execute_22625_51_), .B(d_reg_19_), .Y(_abc_15497_new_n1494_));
NOR2X1 NOR2X1_22 ( .A(_abc_15497_new_n748_), .B(_abc_15497_new_n749_), .Y(_abc_15497_new_n750_));
NOR2X1 NOR2X1_220 ( .A(_abc_15497_new_n1492_), .B(_abc_15497_new_n1495_), .Y(_abc_15497_new_n1496_));
NOR2X1 NOR2X1_221 ( .A(_abc_15497_new_n1494_), .B(_abc_15497_new_n1496_), .Y(_abc_15497_new_n1497_));
NOR2X1 NOR2X1_222 ( .A(_abc_15497_new_n1489_), .B(_abc_15497_new_n1498_), .Y(_abc_15497_new_n1502_));
NOR2X1 NOR2X1_223 ( .A(_abc_15497_new_n1480_), .B(_abc_15497_new_n1503_), .Y(_abc_15497_new_n1504_));
NOR2X1 NOR2X1_224 ( .A(_auto_iopadmap_cc_368_execute_22625_52_), .B(d_reg_20_), .Y(_abc_15497_new_n1509_));
NOR2X1 NOR2X1_225 ( .A(_abc_15497_new_n1510_), .B(_abc_15497_new_n1511_), .Y(_abc_15497_new_n1512_));
NOR2X1 NOR2X1_226 ( .A(_abc_15497_new_n1509_), .B(_abc_15497_new_n1512_), .Y(_abc_15497_new_n1513_));
NOR2X1 NOR2X1_227 ( .A(_abc_15497_new_n1513_), .B(_abc_15497_new_n1508_), .Y(_abc_15497_new_n1514_));
NOR2X1 NOR2X1_228 ( .A(_auto_iopadmap_cc_368_execute_22625_53_), .B(d_reg_21_), .Y(_abc_15497_new_n1521_));
NOR2X1 NOR2X1_229 ( .A(_auto_iopadmap_cc_368_execute_22625_54_), .B(d_reg_22_), .Y(_abc_15497_new_n1529_));
NOR2X1 NOR2X1_23 ( .A(c_reg_7_), .B(_auto_iopadmap_cc_368_execute_22625_71_), .Y(_abc_15497_new_n751_));
NOR2X1 NOR2X1_230 ( .A(_abc_15497_new_n1528_), .B(_abc_15497_new_n1530_), .Y(_abc_15497_new_n1531_));
NOR2X1 NOR2X1_231 ( .A(_abc_15497_new_n1529_), .B(_abc_15497_new_n1531_), .Y(_abc_15497_new_n1532_));
NOR2X1 NOR2X1_232 ( .A(_abc_15497_new_n1524_), .B(_abc_15497_new_n1515_), .Y(_abc_15497_new_n1535_));
NOR2X1 NOR2X1_233 ( .A(_abc_15497_new_n1533_), .B(_abc_15497_new_n1536_), .Y(_abc_15497_new_n1541_));
NOR2X1 NOR2X1_234 ( .A(_abc_15497_new_n1531_), .B(_abc_15497_new_n1541_), .Y(_abc_15497_new_n1542_));
NOR2X1 NOR2X1_235 ( .A(_abc_15497_new_n1546_), .B(_abc_15497_new_n1533_), .Y(_abc_15497_new_n1553_));
NOR2X1 NOR2X1_236 ( .A(_abc_15497_new_n1555_), .B(_abc_15497_new_n1557_), .Y(_abc_15497_new_n1558_));
NOR2X1 NOR2X1_237 ( .A(_auto_iopadmap_cc_368_execute_22625_56_), .B(d_reg_24_), .Y(_abc_15497_new_n1561_));
NOR2X1 NOR2X1_238 ( .A(_abc_15497_new_n1550_), .B(_abc_15497_new_n1562_), .Y(_abc_15497_new_n1563_));
NOR2X1 NOR2X1_239 ( .A(_abc_15497_new_n1561_), .B(_abc_15497_new_n1563_), .Y(_abc_15497_new_n1564_));
NOR2X1 NOR2X1_24 ( .A(_abc_15497_new_n751_), .B(_abc_15497_new_n747_), .Y(_abc_15497_new_n752_));
NOR2X1 NOR2X1_240 ( .A(_abc_15497_new_n1564_), .B(_abc_15497_new_n1560_), .Y(_abc_15497_new_n1565_));
NOR2X1 NOR2X1_241 ( .A(_abc_15497_new_n1566_), .B(_abc_15497_new_n1559_), .Y(_abc_15497_new_n1570_));
NOR2X1 NOR2X1_242 ( .A(_auto_iopadmap_cc_368_execute_22625_57_), .B(d_reg_25_), .Y(_abc_15497_new_n1571_));
NOR2X1 NOR2X1_243 ( .A(_abc_15497_new_n1569_), .B(_abc_15497_new_n1572_), .Y(_abc_15497_new_n1573_));
NOR2X1 NOR2X1_244 ( .A(_abc_15497_new_n1571_), .B(_abc_15497_new_n1573_), .Y(_abc_15497_new_n1574_));
NOR2X1 NOR2X1_245 ( .A(_abc_15497_new_n1566_), .B(_abc_15497_new_n1575_), .Y(_abc_15497_new_n1581_));
NOR2X1 NOR2X1_246 ( .A(_auto_iopadmap_cc_368_execute_22625_58_), .B(d_reg_26_), .Y(_abc_15497_new_n1585_));
NOR2X1 NOR2X1_247 ( .A(_abc_15497_new_n1580_), .B(_abc_15497_new_n1586_), .Y(_abc_15497_new_n1587_));
NOR2X1 NOR2X1_248 ( .A(_abc_15497_new_n1585_), .B(_abc_15497_new_n1587_), .Y(_abc_15497_new_n1588_));
NOR2X1 NOR2X1_249 ( .A(_abc_15497_new_n1589_), .B(_abc_15497_new_n1584_), .Y(_abc_15497_new_n1594_));
NOR2X1 NOR2X1_25 ( .A(c_reg_6_), .B(_auto_iopadmap_cc_368_execute_22625_70_), .Y(_abc_15497_new_n755_));
NOR2X1 NOR2X1_250 ( .A(_auto_iopadmap_cc_368_execute_22625_59_), .B(d_reg_27_), .Y(_abc_15497_new_n1595_));
NOR2X1 NOR2X1_251 ( .A(_abc_15497_new_n1593_), .B(_abc_15497_new_n1596_), .Y(_abc_15497_new_n1597_));
NOR2X1 NOR2X1_252 ( .A(_abc_15497_new_n1595_), .B(_abc_15497_new_n1597_), .Y(_abc_15497_new_n1598_));
NOR2X1 NOR2X1_253 ( .A(_abc_15497_new_n1599_), .B(_abc_15497_new_n1589_), .Y(_abc_15497_new_n1604_));
NOR2X1 NOR2X1_254 ( .A(_abc_15497_new_n1611_), .B(_abc_15497_new_n1610_), .Y(_abc_15497_new_n1612_));
NOR2X1 NOR2X1_255 ( .A(_auto_iopadmap_cc_368_execute_22625_61_), .B(d_reg_29_), .Y(_abc_15497_new_n1620_));
NOR2X1 NOR2X1_256 ( .A(_abc_15497_new_n1621_), .B(_abc_15497_new_n1622_), .Y(_abc_15497_new_n1623_));
NOR2X1 NOR2X1_257 ( .A(_abc_15497_new_n1620_), .B(_abc_15497_new_n1623_), .Y(_abc_15497_new_n1624_));
NOR2X1 NOR2X1_258 ( .A(next), .B(init), .Y(_abc_15497_new_n1647_));
NOR2X1 NOR2X1_259 ( .A(_abc_15497_new_n936_), .B(_abc_15497_new_n883__bF_buf10), .Y(_abc_15497_new_n1649_));
NOR2X1 NOR2X1_26 ( .A(_abc_15497_new_n755_), .B(_abc_15497_new_n750_), .Y(_abc_15497_new_n756_));
NOR2X1 NOR2X1_260 ( .A(round_ctr_inc_bF_buf12), .B(_abc_15497_new_n1644_), .Y(_abc_15497_new_n1650_));
NOR2X1 NOR2X1_261 ( .A(_abc_15497_new_n941_), .B(_abc_15497_new_n883__bF_buf9), .Y(_abc_15497_new_n1653_));
NOR2X1 NOR2X1_262 ( .A(_abc_15497_new_n946_), .B(_abc_15497_new_n883__bF_buf8), .Y(_abc_15497_new_n1656_));
NOR2X1 NOR2X1_263 ( .A(_abc_15497_new_n955_), .B(_abc_15497_new_n883__bF_buf7), .Y(_abc_15497_new_n1659_));
NOR2X1 NOR2X1_264 ( .A(_abc_15497_new_n1024_), .B(_abc_15497_new_n883__bF_buf2), .Y(_abc_15497_new_n1678_));
NOR2X1 NOR2X1_265 ( .A(_abc_15497_new_n1033_), .B(_abc_15497_new_n883__bF_buf1), .Y(_abc_15497_new_n1681_));
NOR2X1 NOR2X1_266 ( .A(_abc_15497_new_n1048_), .B(_abc_15497_new_n883__bF_buf0), .Y(_abc_15497_new_n1685_));
NOR2X1 NOR2X1_267 ( .A(_abc_15497_new_n1057_), .B(_abc_15497_new_n883__bF_buf13), .Y(_abc_15497_new_n1688_));
NOR2X1 NOR2X1_268 ( .A(_abc_15497_new_n1101_), .B(_abc_15497_new_n883__bF_buf10), .Y(_abc_15497_new_n1700_));
NOR2X1 NOR2X1_269 ( .A(_abc_15497_new_n1128_), .B(_abc_15497_new_n883__bF_buf9), .Y(_abc_15497_new_n1706_));
NOR2X1 NOR2X1_27 ( .A(_abc_15497_new_n759_), .B(_abc_15497_new_n760_), .Y(_abc_15497_new_n761_));
NOR2X1 NOR2X1_270 ( .A(_abc_15497_new_n1142_), .B(_abc_15497_new_n883__bF_buf8), .Y(_abc_15497_new_n1709_));
NOR2X1 NOR2X1_271 ( .A(_abc_15497_new_n1171_), .B(_abc_15497_new_n883__bF_buf7), .Y(_abc_15497_new_n1715_));
NOR2X1 NOR2X1_272 ( .A(_abc_15497_new_n1231_), .B(_abc_15497_new_n883__bF_buf3), .Y(_abc_15497_new_n1730_));
NOR2X1 NOR2X1_273 ( .A(_abc_15497_new_n1247_), .B(_abc_15497_new_n883__bF_buf2), .Y(_abc_15497_new_n1733_));
NOR2X1 NOR2X1_274 ( .A(_abc_15497_new_n1258_), .B(_abc_15497_new_n883__bF_buf1), .Y(_abc_15497_new_n1737_));
NOR2X1 NOR2X1_275 ( .A(_abc_15497_new_n1274_), .B(_abc_15497_new_n883__bF_buf0), .Y(_abc_15497_new_n1740_));
NOR2X1 NOR2X1_276 ( .A(_auto_iopadmap_cc_368_execute_22625_96_), .B(b_reg_0_), .Y(_abc_15497_new_n1750_));
NOR2X1 NOR2X1_277 ( .A(_abc_15497_new_n1751_), .B(_abc_15497_new_n1752_), .Y(_abc_15497_new_n1757_));
NOR2X1 NOR2X1_278 ( .A(_auto_iopadmap_cc_368_execute_22625_99_), .B(b_reg_3_), .Y(_abc_15497_new_n1773_));
NOR2X1 NOR2X1_279 ( .A(_abc_15497_new_n1773_), .B(_abc_15497_new_n1774_), .Y(_abc_15497_new_n1775_));
NOR2X1 NOR2X1_28 ( .A(c_reg_5_), .B(_auto_iopadmap_cc_368_execute_22625_69_), .Y(_abc_15497_new_n763_));
NOR2X1 NOR2X1_280 ( .A(_abc_15497_new_n1780_), .B(_abc_15497_new_n1782_), .Y(_abc_15497_new_n1783_));
NOR2X1 NOR2X1_281 ( .A(_abc_15497_new_n1779_), .B(_abc_15497_new_n1788_), .Y(_abc_15497_new_n1789_));
NOR2X1 NOR2X1_282 ( .A(_abc_15497_new_n1789_), .B(_abc_15497_new_n1783_), .Y(_abc_15497_new_n1790_));
NOR2X1 NOR2X1_283 ( .A(_auto_iopadmap_cc_368_execute_22625_101_), .B(b_reg_5_), .Y(_abc_15497_new_n1791_));
NOR2X1 NOR2X1_284 ( .A(_abc_15497_new_n1787_), .B(_abc_15497_new_n1792_), .Y(_abc_15497_new_n1793_));
NOR2X1 NOR2X1_285 ( .A(_abc_15497_new_n1791_), .B(_abc_15497_new_n1793_), .Y(_abc_15497_new_n1795_));
NOR2X1 NOR2X1_286 ( .A(_auto_iopadmap_cc_368_execute_22625_102_), .B(b_reg_6_), .Y(_abc_15497_new_n1801_));
NOR2X1 NOR2X1_287 ( .A(_abc_15497_new_n1799_), .B(_abc_15497_new_n1802_), .Y(_abc_15497_new_n1803_));
NOR2X1 NOR2X1_288 ( .A(_abc_15497_new_n1801_), .B(_abc_15497_new_n1803_), .Y(_abc_15497_new_n1804_));
NOR2X1 NOR2X1_289 ( .A(_auto_iopadmap_cc_368_execute_22625_103_), .B(b_reg_7_), .Y(_abc_15497_new_n1808_));
NOR2X1 NOR2X1_29 ( .A(c_reg_3_), .B(_auto_iopadmap_cc_368_execute_22625_67_), .Y(_abc_15497_new_n766_));
NOR2X1 NOR2X1_290 ( .A(_abc_15497_new_n1808_), .B(_abc_15497_new_n1810_), .Y(_abc_15497_new_n1811_));
NOR2X1 NOR2X1_291 ( .A(_abc_15497_new_n1811_), .B(_abc_15497_new_n1807_), .Y(_abc_15497_new_n1814_));
NOR2X1 NOR2X1_292 ( .A(_auto_iopadmap_cc_368_execute_22625_104_), .B(b_reg_8_), .Y(_abc_15497_new_n1818_));
NOR2X1 NOR2X1_293 ( .A(_abc_15497_new_n1819_), .B(_abc_15497_new_n1820_), .Y(_abc_15497_new_n1821_));
NOR2X1 NOR2X1_294 ( .A(_abc_15497_new_n1818_), .B(_abc_15497_new_n1821_), .Y(_abc_15497_new_n1822_));
NOR2X1 NOR2X1_295 ( .A(_auto_iopadmap_cc_368_execute_22625_105_), .B(b_reg_9_), .Y(_abc_15497_new_n1830_));
NOR2X1 NOR2X1_296 ( .A(_abc_15497_new_n1830_), .B(_abc_15497_new_n1831_), .Y(_abc_15497_new_n1832_));
NOR2X1 NOR2X1_297 ( .A(_auto_iopadmap_cc_368_execute_22625_106_), .B(b_reg_10_), .Y(_abc_15497_new_n1840_));
NOR2X1 NOR2X1_298 ( .A(_abc_15497_new_n1836_), .B(_abc_15497_new_n1841_), .Y(_abc_15497_new_n1842_));
NOR2X1 NOR2X1_299 ( .A(_abc_15497_new_n1840_), .B(_abc_15497_new_n1842_), .Y(_abc_15497_new_n1843_));
NOR2X1 NOR2X1_3 ( .A(_abc_15497_new_n702_), .B(_abc_15497_new_n703_), .Y(_abc_15497_new_n704_));
NOR2X1 NOR2X1_30 ( .A(_abc_15497_new_n769_), .B(_abc_15497_new_n770_), .Y(_abc_15497_new_n771_));
NOR2X1 NOR2X1_300 ( .A(_abc_15497_new_n1843_), .B(_abc_15497_new_n1839_), .Y(_abc_15497_new_n1844_));
NOR2X1 NOR2X1_301 ( .A(_auto_iopadmap_cc_368_execute_22625_107_), .B(b_reg_11_), .Y(_abc_15497_new_n1849_));
NOR2X1 NOR2X1_302 ( .A(_abc_15497_new_n1849_), .B(_abc_15497_new_n1851_), .Y(_abc_15497_new_n1852_));
NOR2X1 NOR2X1_303 ( .A(_auto_iopadmap_cc_368_execute_22625_108_), .B(b_reg_12_), .Y(_abc_15497_new_n1857_));
NOR2X1 NOR2X1_304 ( .A(_abc_15497_new_n1856_), .B(_abc_15497_new_n1858_), .Y(_abc_15497_new_n1859_));
NOR2X1 NOR2X1_305 ( .A(_abc_15497_new_n1857_), .B(_abc_15497_new_n1859_), .Y(_abc_15497_new_n1860_));
NOR2X1 NOR2X1_306 ( .A(_abc_15497_new_n1862_), .B(_abc_15497_new_n1837_), .Y(_abc_15497_new_n1864_));
NOR2X1 NOR2X1_307 ( .A(_auto_iopadmap_cc_368_execute_22625_110_), .B(b_reg_14_), .Y(_abc_15497_new_n1875_));
NOR2X1 NOR2X1_308 ( .A(_abc_15497_new_n1874_), .B(_abc_15497_new_n1876_), .Y(_abc_15497_new_n1877_));
NOR2X1 NOR2X1_309 ( .A(_abc_15497_new_n1875_), .B(_abc_15497_new_n1877_), .Y(_abc_15497_new_n1878_));
NOR2X1 NOR2X1_31 ( .A(c_reg_2_), .B(_auto_iopadmap_cc_368_execute_22625_66_), .Y(_abc_15497_new_n775_));
NOR2X1 NOR2X1_310 ( .A(_auto_iopadmap_cc_368_execute_22625_111_), .B(b_reg_15_), .Y(_abc_15497_new_n1892_));
NOR2X1 NOR2X1_311 ( .A(_abc_15497_new_n1892_), .B(_abc_15497_new_n1894_), .Y(_abc_15497_new_n1895_));
NOR2X1 NOR2X1_312 ( .A(_abc_15497_new_n1900_), .B(_abc_15497_new_n1884_), .Y(_abc_15497_new_n1902_));
NOR2X1 NOR2X1_313 ( .A(_auto_iopadmap_cc_368_execute_22625_112_), .B(b_reg_16_), .Y(_abc_15497_new_n1906_));
NOR2X1 NOR2X1_314 ( .A(_abc_15497_new_n1907_), .B(_abc_15497_new_n1908_), .Y(_abc_15497_new_n1909_));
NOR2X1 NOR2X1_315 ( .A(_abc_15497_new_n1906_), .B(_abc_15497_new_n1909_), .Y(_abc_15497_new_n1910_));
NOR2X1 NOR2X1_316 ( .A(_abc_15497_new_n1910_), .B(_abc_15497_new_n1905_), .Y(_abc_15497_new_n1911_));
NOR2X1 NOR2X1_317 ( .A(_auto_iopadmap_cc_368_execute_22625_113_), .B(b_reg_17_), .Y(_abc_15497_new_n1917_));
NOR2X1 NOR2X1_318 ( .A(_abc_15497_new_n1916_), .B(_abc_15497_new_n1918_), .Y(_abc_15497_new_n1919_));
NOR2X1 NOR2X1_319 ( .A(_abc_15497_new_n1917_), .B(_abc_15497_new_n1919_), .Y(_abc_15497_new_n1920_));
NOR2X1 NOR2X1_32 ( .A(_abc_15497_new_n775_), .B(_abc_15497_new_n767_), .Y(_abc_15497_new_n776_));
NOR2X1 NOR2X1_320 ( .A(_abc_15497_new_n1924_), .B(_abc_15497_new_n1912_), .Y(_abc_15497_new_n1925_));
NOR2X1 NOR2X1_321 ( .A(_auto_iopadmap_cc_368_execute_22625_114_), .B(b_reg_18_), .Y(_abc_15497_new_n1929_));
NOR2X1 NOR2X1_322 ( .A(_abc_15497_new_n1929_), .B(_abc_15497_new_n1931_), .Y(_abc_15497_new_n1932_));
NOR2X1 NOR2X1_323 ( .A(_abc_15497_new_n1932_), .B(_abc_15497_new_n1928_), .Y(_abc_15497_new_n1933_));
NOR2X1 NOR2X1_324 ( .A(_auto_iopadmap_cc_368_execute_22625_115_), .B(b_reg_19_), .Y(_abc_15497_new_n1939_));
NOR2X1 NOR2X1_325 ( .A(_abc_15497_new_n1939_), .B(_abc_15497_new_n1941_), .Y(_abc_15497_new_n1942_));
NOR2X1 NOR2X1_326 ( .A(_abc_15497_new_n1943_), .B(_abc_15497_new_n1938_), .Y(_abc_15497_new_n1944_));
NOR2X1 NOR2X1_327 ( .A(_abc_15497_new_n1951_), .B(_abc_15497_new_n1954_), .Y(_abc_15497_new_n1955_));
NOR2X1 NOR2X1_328 ( .A(_auto_iopadmap_cc_368_execute_22625_116_), .B(b_reg_20_), .Y(_abc_15497_new_n1957_));
NOR2X1 NOR2X1_329 ( .A(_abc_15497_new_n1949_), .B(_abc_15497_new_n1958_), .Y(_abc_15497_new_n1959_));
NOR2X1 NOR2X1_33 ( .A(c_reg_8_), .B(_auto_iopadmap_cc_368_execute_22625_72_), .Y(_abc_15497_new_n785_));
NOR2X1 NOR2X1_330 ( .A(_abc_15497_new_n1957_), .B(_abc_15497_new_n1959_), .Y(_abc_15497_new_n1960_));
NOR2X1 NOR2X1_331 ( .A(_auto_iopadmap_cc_368_execute_22625_117_), .B(b_reg_21_), .Y(_abc_15497_new_n1966_));
NOR2X1 NOR2X1_332 ( .A(_abc_15497_new_n1965_), .B(_abc_15497_new_n1967_), .Y(_abc_15497_new_n1968_));
NOR2X1 NOR2X1_333 ( .A(_abc_15497_new_n1966_), .B(_abc_15497_new_n1968_), .Y(_abc_15497_new_n1969_));
NOR2X1 NOR2X1_334 ( .A(_abc_15497_new_n1961_), .B(_abc_15497_new_n1974_), .Y(_abc_15497_new_n1975_));
NOR2X1 NOR2X1_335 ( .A(_auto_iopadmap_cc_368_execute_22625_118_), .B(b_reg_22_), .Y(_abc_15497_new_n1979_));
NOR2X1 NOR2X1_336 ( .A(_abc_15497_new_n1979_), .B(_abc_15497_new_n1981_), .Y(_abc_15497_new_n1982_));
NOR2X1 NOR2X1_337 ( .A(_auto_iopadmap_cc_368_execute_22625_119_), .B(b_reg_23_), .Y(_abc_15497_new_n1987_));
NOR2X1 NOR2X1_338 ( .A(_abc_15497_new_n1987_), .B(_abc_15497_new_n1989_), .Y(_abc_15497_new_n1990_));
NOR2X1 NOR2X1_339 ( .A(_abc_15497_new_n1994_), .B(_abc_15497_new_n1976_), .Y(_abc_15497_new_n1995_));
NOR2X1 NOR2X1_34 ( .A(_abc_15497_new_n785_), .B(_abc_15497_new_n743_), .Y(_abc_15497_new_n786_));
NOR2X1 NOR2X1_340 ( .A(_abc_15497_new_n1999_), .B(_abc_15497_new_n1997_), .Y(_abc_15497_new_n2000_));
NOR2X1 NOR2X1_341 ( .A(_auto_iopadmap_cc_368_execute_22625_120_), .B(b_reg_24_), .Y(_abc_15497_new_n2004_));
NOR2X1 NOR2X1_342 ( .A(_abc_15497_new_n2005_), .B(_abc_15497_new_n2006_), .Y(_abc_15497_new_n2007_));
NOR2X1 NOR2X1_343 ( .A(_abc_15497_new_n2004_), .B(_abc_15497_new_n2007_), .Y(_abc_15497_new_n2008_));
NOR2X1 NOR2X1_344 ( .A(_auto_iopadmap_cc_368_execute_22625_121_), .B(b_reg_25_), .Y(_abc_15497_new_n2016_));
NOR2X1 NOR2X1_345 ( .A(_abc_15497_new_n2016_), .B(_abc_15497_new_n2018_), .Y(_abc_15497_new_n2019_));
NOR2X1 NOR2X1_346 ( .A(_abc_15497_new_n2023_), .B(_abc_15497_new_n2009_), .Y(_abc_15497_new_n2024_));
NOR2X1 NOR2X1_347 ( .A(_auto_iopadmap_cc_368_execute_22625_122_), .B(b_reg_26_), .Y(_abc_15497_new_n2029_));
NOR2X1 NOR2X1_348 ( .A(_abc_15497_new_n2030_), .B(_abc_15497_new_n2031_), .Y(_abc_15497_new_n2032_));
NOR2X1 NOR2X1_349 ( .A(_abc_15497_new_n2029_), .B(_abc_15497_new_n2032_), .Y(_abc_15497_new_n2033_));
NOR2X1 NOR2X1_35 ( .A(_abc_15497_new_n784_), .B(_abc_15497_new_n787_), .Y(_abc_15497_new_n788_));
NOR2X1 NOR2X1_350 ( .A(_abc_15497_new_n2033_), .B(_abc_15497_new_n2028_), .Y(_abc_15497_new_n2034_));
NOR2X1 NOR2X1_351 ( .A(_auto_iopadmap_cc_368_execute_22625_123_), .B(b_reg_27_), .Y(_abc_15497_new_n2040_));
NOR2X1 NOR2X1_352 ( .A(_abc_15497_new_n2040_), .B(_abc_15497_new_n2042_), .Y(_abc_15497_new_n2043_));
NOR2X1 NOR2X1_353 ( .A(_auto_iopadmap_cc_368_execute_22625_125_), .B(_abc_15497_new_n883__bF_buf8), .Y(_abc_15497_new_n2062_));
NOR2X1 NOR2X1_354 ( .A(_auto_iopadmap_cc_368_execute_22625_125_), .B(b_reg_29_), .Y(_abc_15497_new_n2064_));
NOR2X1 NOR2X1_355 ( .A(_abc_15497_new_n2064_), .B(_abc_15497_new_n2066_), .Y(_abc_15497_new_n2067_));
NOR2X1 NOR2X1_356 ( .A(_abc_15497_new_n2059_), .B(_abc_15497_new_n2068_), .Y(_abc_15497_new_n2075_));
NOR2X1 NOR2X1_357 ( .A(_auto_iopadmap_cc_368_execute_22625_128_), .B(a_reg_0_), .Y(_abc_15497_new_n2091_));
NOR2X1 NOR2X1_358 ( .A(_abc_15497_new_n2092_), .B(_abc_15497_new_n2093_), .Y(_abc_15497_new_n2098_));
NOR2X1 NOR2X1_359 ( .A(_abc_15497_new_n2112_), .B(_abc_15497_new_n2115_), .Y(_abc_15497_new_n2117_));
NOR2X1 NOR2X1_36 ( .A(c_reg_23_), .B(_auto_iopadmap_cc_368_execute_22625_87_), .Y(_abc_15497_new_n793_));
NOR2X1 NOR2X1_360 ( .A(_abc_15497_new_n2123_), .B(_abc_15497_new_n2124_), .Y(_abc_15497_new_n2125_));
NOR2X1 NOR2X1_361 ( .A(_abc_15497_new_n2122_), .B(_abc_15497_new_n2130_), .Y(_abc_15497_new_n2131_));
NOR2X1 NOR2X1_362 ( .A(_abc_15497_new_n2131_), .B(_abc_15497_new_n2125_), .Y(_abc_15497_new_n2132_));
NOR2X1 NOR2X1_363 ( .A(_auto_iopadmap_cc_368_execute_22625_133_), .B(a_reg_5_), .Y(_abc_15497_new_n2133_));
NOR2X1 NOR2X1_364 ( .A(_abc_15497_new_n2129_), .B(_abc_15497_new_n2134_), .Y(_abc_15497_new_n2135_));
NOR2X1 NOR2X1_365 ( .A(_abc_15497_new_n2133_), .B(_abc_15497_new_n2135_), .Y(_abc_15497_new_n2137_));
NOR2X1 NOR2X1_366 ( .A(_auto_iopadmap_cc_368_execute_22625_134_), .B(a_reg_6_), .Y(_abc_15497_new_n2143_));
NOR2X1 NOR2X1_367 ( .A(_abc_15497_new_n2141_), .B(_abc_15497_new_n2144_), .Y(_abc_15497_new_n2145_));
NOR2X1 NOR2X1_368 ( .A(_abc_15497_new_n2143_), .B(_abc_15497_new_n2145_), .Y(_abc_15497_new_n2146_));
NOR2X1 NOR2X1_369 ( .A(_abc_15497_new_n2146_), .B(_abc_15497_new_n2142_), .Y(_abc_15497_new_n2147_));
NOR2X1 NOR2X1_37 ( .A(_abc_15497_new_n793_), .B(_abc_15497_new_n795_), .Y(_abc_15497_new_n796_));
NOR2X1 NOR2X1_370 ( .A(_abc_15497_new_n2153_), .B(_abc_15497_new_n2148_), .Y(_abc_15497_new_n2154_));
NOR2X1 NOR2X1_371 ( .A(_abc_15497_new_n2161_), .B(_abc_15497_new_n2154_), .Y(_abc_15497_new_n2162_));
NOR2X1 NOR2X1_372 ( .A(_auto_iopadmap_cc_368_execute_22625_136_), .B(a_reg_8_), .Y(_abc_15497_new_n2164_));
NOR2X1 NOR2X1_373 ( .A(_abc_15497_new_n2165_), .B(_abc_15497_new_n2166_), .Y(_abc_15497_new_n2167_));
NOR2X1 NOR2X1_374 ( .A(_abc_15497_new_n2164_), .B(_abc_15497_new_n2167_), .Y(_abc_15497_new_n2168_));
NOR2X1 NOR2X1_375 ( .A(_abc_15497_new_n2168_), .B(_abc_15497_new_n2163_), .Y(_abc_15497_new_n2169_));
NOR2X1 NOR2X1_376 ( .A(_auto_iopadmap_cc_368_execute_22625_138_), .B(a_reg_10_), .Y(_abc_15497_new_n2181_));
NOR2X1 NOR2X1_377 ( .A(_abc_15497_new_n2180_), .B(_abc_15497_new_n2182_), .Y(_abc_15497_new_n2183_));
NOR2X1 NOR2X1_378 ( .A(_abc_15497_new_n2181_), .B(_abc_15497_new_n2183_), .Y(_abc_15497_new_n2184_));
NOR2X1 NOR2X1_379 ( .A(_abc_15497_new_n2191_), .B(_abc_15497_new_n2204_), .Y(_abc_15497_new_n2205_));
NOR2X1 NOR2X1_38 ( .A(_abc_15497_new_n798_), .B(_abc_15497_new_n799_), .Y(_abc_15497_new_n800_));
NOR2X1 NOR2X1_380 ( .A(_auto_iopadmap_cc_368_execute_22625_140_), .B(a_reg_12_), .Y(_abc_15497_new_n2213_));
NOR2X1 NOR2X1_381 ( .A(_abc_15497_new_n2203_), .B(_abc_15497_new_n2214_), .Y(_abc_15497_new_n2215_));
NOR2X1 NOR2X1_382 ( .A(_abc_15497_new_n2213_), .B(_abc_15497_new_n2215_), .Y(_abc_15497_new_n2216_));
NOR2X1 NOR2X1_383 ( .A(_abc_15497_new_n2216_), .B(_abc_15497_new_n2212_), .Y(_abc_15497_new_n2217_));
NOR2X1 NOR2X1_384 ( .A(_auto_iopadmap_cc_368_execute_22625_141_), .B(a_reg_13_), .Y(_abc_15497_new_n2222_));
NOR2X1 NOR2X1_385 ( .A(_abc_15497_new_n2222_), .B(_abc_15497_new_n2223_), .Y(_abc_15497_new_n2224_));
NOR2X1 NOR2X1_386 ( .A(_auto_iopadmap_cc_368_execute_22625_142_), .B(a_reg_14_), .Y(_abc_15497_new_n2229_));
NOR2X1 NOR2X1_387 ( .A(_abc_15497_new_n2228_), .B(_abc_15497_new_n2230_), .Y(_abc_15497_new_n2231_));
NOR2X1 NOR2X1_388 ( .A(_abc_15497_new_n2229_), .B(_abc_15497_new_n2231_), .Y(_abc_15497_new_n2232_));
NOR2X1 NOR2X1_389 ( .A(_abc_15497_new_n2232_), .B(_abc_15497_new_n2236_), .Y(_abc_15497_new_n2237_));
NOR2X1 NOR2X1_39 ( .A(c_reg_22_), .B(_auto_iopadmap_cc_368_execute_22625_86_), .Y(_abc_15497_new_n801_));
NOR2X1 NOR2X1_390 ( .A(_auto_iopadmap_cc_368_execute_22625_143_), .B(a_reg_15_), .Y(_abc_15497_new_n2243_));
NOR2X1 NOR2X1_391 ( .A(_abc_15497_new_n2241_), .B(_abc_15497_new_n2244_), .Y(_abc_15497_new_n2245_));
NOR2X1 NOR2X1_392 ( .A(_abc_15497_new_n2243_), .B(_abc_15497_new_n2245_), .Y(_abc_15497_new_n2246_));
NOR2X1 NOR2X1_393 ( .A(_abc_15497_new_n2235_), .B(_abc_15497_new_n2250_), .Y(_abc_15497_new_n2252_));
NOR2X1 NOR2X1_394 ( .A(_auto_iopadmap_cc_368_execute_22625_144_), .B(a_reg_16_), .Y(_abc_15497_new_n2256_));
NOR2X1 NOR2X1_395 ( .A(_abc_15497_new_n2257_), .B(_abc_15497_new_n2258_), .Y(_abc_15497_new_n2259_));
NOR2X1 NOR2X1_396 ( .A(_abc_15497_new_n2256_), .B(_abc_15497_new_n2259_), .Y(_abc_15497_new_n2260_));
NOR2X1 NOR2X1_397 ( .A(_abc_15497_new_n2260_), .B(_abc_15497_new_n2255_), .Y(_abc_15497_new_n2261_));
NOR2X1 NOR2X1_398 ( .A(_abc_15497_new_n2263_), .B(_abc_15497_new_n2262_), .Y(_abc_15497_new_n2268_));
NOR2X1 NOR2X1_399 ( .A(_auto_iopadmap_cc_368_execute_22625_145_), .B(a_reg_17_), .Y(_abc_15497_new_n2269_));
NOR2X1 NOR2X1_4 ( .A(c_reg_14_), .B(_auto_iopadmap_cc_368_execute_22625_78_), .Y(_abc_15497_new_n705_));
NOR2X1 NOR2X1_40 ( .A(_abc_15497_new_n801_), .B(_abc_15497_new_n800_), .Y(_abc_15497_new_n802_));
NOR2X1 NOR2X1_400 ( .A(_abc_15497_new_n2267_), .B(_abc_15497_new_n2270_), .Y(_abc_15497_new_n2271_));
NOR2X1 NOR2X1_401 ( .A(_abc_15497_new_n2269_), .B(_abc_15497_new_n2271_), .Y(_abc_15497_new_n2272_));
NOR2X1 NOR2X1_402 ( .A(_abc_15497_new_n2263_), .B(_abc_15497_new_n2273_), .Y(_abc_15497_new_n2278_));
NOR2X1 NOR2X1_403 ( .A(_auto_iopadmap_cc_368_execute_22625_146_), .B(a_reg_18_), .Y(_abc_15497_new_n2282_));
NOR2X1 NOR2X1_404 ( .A(_abc_15497_new_n2283_), .B(_abc_15497_new_n2284_), .Y(_abc_15497_new_n2285_));
NOR2X1 NOR2X1_405 ( .A(_abc_15497_new_n2282_), .B(_abc_15497_new_n2285_), .Y(_abc_15497_new_n2286_));
NOR2X1 NOR2X1_406 ( .A(_abc_15497_new_n870__bF_buf9), .B(_abc_15497_new_n2287_), .Y(_abc_15497_new_n2288_));
NOR2X1 NOR2X1_407 ( .A(_abc_15497_new_n2285_), .B(_abc_15497_new_n2287_), .Y(_abc_15497_new_n2294_));
NOR2X1 NOR2X1_408 ( .A(_auto_iopadmap_cc_368_execute_22625_147_), .B(a_reg_19_), .Y(_abc_15497_new_n2295_));
NOR2X1 NOR2X1_409 ( .A(_abc_15497_new_n2293_), .B(_abc_15497_new_n2296_), .Y(_abc_15497_new_n2297_));
NOR2X1 NOR2X1_41 ( .A(_abc_15497_new_n797_), .B(_abc_15497_new_n803_), .Y(_abc_15497_new_n804_));
NOR2X1 NOR2X1_410 ( .A(_abc_15497_new_n2295_), .B(_abc_15497_new_n2297_), .Y(_abc_15497_new_n2298_));
NOR2X1 NOR2X1_411 ( .A(_abc_15497_new_n2304_), .B(_abc_15497_new_n2279_), .Y(_abc_15497_new_n2305_));
NOR2X1 NOR2X1_412 ( .A(_auto_iopadmap_cc_368_execute_22625_148_), .B(a_reg_20_), .Y(_abc_15497_new_n2309_));
NOR2X1 NOR2X1_413 ( .A(_abc_15497_new_n2303_), .B(_abc_15497_new_n2310_), .Y(_abc_15497_new_n2311_));
NOR2X1 NOR2X1_414 ( .A(_abc_15497_new_n2309_), .B(_abc_15497_new_n2311_), .Y(_abc_15497_new_n2312_));
NOR2X1 NOR2X1_415 ( .A(_abc_15497_new_n2313_), .B(_abc_15497_new_n2308_), .Y(_abc_15497_new_n2318_));
NOR2X1 NOR2X1_416 ( .A(_auto_iopadmap_cc_368_execute_22625_149_), .B(a_reg_21_), .Y(_abc_15497_new_n2320_));
NOR2X1 NOR2X1_417 ( .A(_abc_15497_new_n2317_), .B(_abc_15497_new_n2321_), .Y(_abc_15497_new_n2322_));
NOR2X1 NOR2X1_418 ( .A(_abc_15497_new_n2320_), .B(_abc_15497_new_n2322_), .Y(_abc_15497_new_n2324_));
NOR2X1 NOR2X1_419 ( .A(_auto_iopadmap_cc_368_execute_22625_150_), .B(a_reg_22_), .Y(_abc_15497_new_n2330_));
NOR2X1 NOR2X1_42 ( .A(c_reg_21_), .B(_auto_iopadmap_cc_368_execute_22625_85_), .Y(_abc_15497_new_n808_));
NOR2X1 NOR2X1_420 ( .A(_abc_15497_new_n2331_), .B(_abc_15497_new_n2332_), .Y(_abc_15497_new_n2333_));
NOR2X1 NOR2X1_421 ( .A(_abc_15497_new_n2330_), .B(_abc_15497_new_n2333_), .Y(_abc_15497_new_n2334_));
NOR2X1 NOR2X1_422 ( .A(_abc_15497_new_n2339_), .B(_abc_15497_new_n2347_), .Y(_abc_15497_new_n2348_));
NOR2X1 NOR2X1_423 ( .A(_abc_15497_new_n2353_), .B(_abc_15497_new_n2355_), .Y(_abc_15497_new_n2356_));
NOR2X1 NOR2X1_424 ( .A(_auto_iopadmap_cc_368_execute_22625_152_), .B(a_reg_24_), .Y(_abc_15497_new_n2358_));
NOR2X1 NOR2X1_425 ( .A(_abc_15497_new_n2359_), .B(_abc_15497_new_n2360_), .Y(_abc_15497_new_n2361_));
NOR2X1 NOR2X1_426 ( .A(_abc_15497_new_n2358_), .B(_abc_15497_new_n2361_), .Y(_abc_15497_new_n2362_));
NOR2X1 NOR2X1_427 ( .A(_auto_iopadmap_cc_368_execute_22625_153_), .B(a_reg_25_), .Y(_abc_15497_new_n2370_));
NOR2X1 NOR2X1_428 ( .A(_abc_15497_new_n2371_), .B(_abc_15497_new_n2372_), .Y(_abc_15497_new_n2373_));
NOR2X1 NOR2X1_429 ( .A(_abc_15497_new_n2370_), .B(_abc_15497_new_n2373_), .Y(_abc_15497_new_n2374_));
NOR2X1 NOR2X1_43 ( .A(_abc_15497_new_n808_), .B(_abc_15497_new_n806_), .Y(_abc_15497_new_n809_));
NOR2X1 NOR2X1_430 ( .A(_abc_15497_new_n2363_), .B(_abc_15497_new_n2378_), .Y(_abc_15497_new_n2379_));
NOR2X1 NOR2X1_431 ( .A(_auto_iopadmap_cc_368_execute_22625_154_), .B(a_reg_26_), .Y(_abc_15497_new_n2383_));
NOR2X1 NOR2X1_432 ( .A(_abc_15497_new_n2384_), .B(_abc_15497_new_n2385_), .Y(_abc_15497_new_n2386_));
NOR2X1 NOR2X1_433 ( .A(_abc_15497_new_n2383_), .B(_abc_15497_new_n2386_), .Y(_abc_15497_new_n2387_));
NOR2X1 NOR2X1_434 ( .A(_abc_15497_new_n2387_), .B(_abc_15497_new_n2382_), .Y(_abc_15497_new_n2388_));
NOR2X1 NOR2X1_435 ( .A(_auto_iopadmap_cc_368_execute_22625_155_), .B(a_reg_27_), .Y(_abc_15497_new_n2394_));
NOR2X1 NOR2X1_436 ( .A(_abc_15497_new_n2393_), .B(_abc_15497_new_n2395_), .Y(_abc_15497_new_n2396_));
NOR2X1 NOR2X1_437 ( .A(_abc_15497_new_n2394_), .B(_abc_15497_new_n2396_), .Y(_abc_15497_new_n2397_));
NOR2X1 NOR2X1_438 ( .A(_abc_15497_new_n2409_), .B(_abc_15497_new_n2408_), .Y(_abc_15497_new_n2410_));
NOR2X1 NOR2X1_439 ( .A(_auto_iopadmap_cc_368_execute_22625_157_), .B(a_reg_29_), .Y(_abc_15497_new_n2416_));
NOR2X1 NOR2X1_44 ( .A(c_reg_20_), .B(_auto_iopadmap_cc_368_execute_22625_84_), .Y(_abc_15497_new_n814_));
NOR2X1 NOR2X1_440 ( .A(_abc_15497_new_n2417_), .B(_abc_15497_new_n2418_), .Y(_abc_15497_new_n2419_));
NOR2X1 NOR2X1_441 ( .A(_abc_15497_new_n2416_), .B(_abc_15497_new_n2419_), .Y(_abc_15497_new_n2420_));
NOR2X1 NOR2X1_442 ( .A(_abc_15497_new_n1756_), .B(_abc_15497_new_n883__bF_buf8), .Y(_abc_15497_new_n2447_));
NOR2X1 NOR2X1_443 ( .A(_abc_15497_new_n1762_), .B(_abc_15497_new_n883__bF_buf7), .Y(_abc_15497_new_n2450_));
NOR2X1 NOR2X1_444 ( .A(_abc_15497_new_n1779_), .B(_abc_15497_new_n883__bF_buf5), .Y(_abc_15497_new_n2456_));
NOR2X1 NOR2X1_445 ( .A(_abc_15497_new_n1787_), .B(_abc_15497_new_n883__bF_buf4), .Y(_abc_15497_new_n2459_));
NOR2X1 NOR2X1_446 ( .A(_abc_15497_new_n1799_), .B(_abc_15497_new_n883__bF_buf3), .Y(_abc_15497_new_n2462_));
NOR2X1 NOR2X1_447 ( .A(_abc_15497_new_n1836_), .B(_abc_15497_new_n883__bF_buf0), .Y(_abc_15497_new_n2474_));
NOR2X1 NOR2X1_448 ( .A(_abc_15497_new_n1856_), .B(_abc_15497_new_n883__bF_buf12), .Y(_abc_15497_new_n2480_));
NOR2X1 NOR2X1_449 ( .A(_abc_15497_new_n1874_), .B(_abc_15497_new_n883__bF_buf11), .Y(_abc_15497_new_n2486_));
NOR2X1 NOR2X1_45 ( .A(_abc_15497_new_n814_), .B(_abc_15497_new_n807_), .Y(_abc_15497_new_n815_));
NOR2X1 NOR2X1_450 ( .A(_abc_15497_new_n1916_), .B(_abc_15497_new_n883__bF_buf9), .Y(_abc_15497_new_n2495_));
NOR2X1 NOR2X1_451 ( .A(_abc_15497_new_n1949_), .B(_abc_15497_new_n883__bF_buf6), .Y(_abc_15497_new_n2504_));
NOR2X1 NOR2X1_452 ( .A(_abc_15497_new_n1965_), .B(_abc_15497_new_n883__bF_buf5), .Y(_abc_15497_new_n2507_));
NOR2X1 NOR2X1_453 ( .A(_abc_15497_new_n2047_), .B(_abc_15497_new_n883__bF_buf0), .Y(_abc_15497_new_n2528_));
NOR2X1 NOR2X1_454 ( .A(_abc_15497_new_n1298_), .B(_abc_15497_new_n883__bF_buf10), .Y(_abc_15497_new_n2540_));
NOR2X1 NOR2X1_455 ( .A(_abc_15497_new_n1317_), .B(_abc_15497_new_n883__bF_buf8), .Y(_abc_15497_new_n2549_));
NOR2X1 NOR2X1_456 ( .A(_abc_15497_new_n1351_), .B(_abc_15497_new_n883__bF_buf7), .Y(_abc_15497_new_n2561_));
NOR2X1 NOR2X1_457 ( .A(_abc_15497_new_n1361_), .B(_abc_15497_new_n883__bF_buf6), .Y(_abc_15497_new_n2564_));
NOR2X1 NOR2X1_458 ( .A(_abc_15497_new_n1371_), .B(_abc_15497_new_n883__bF_buf5), .Y(_abc_15497_new_n2567_));
NOR2X1 NOR2X1_459 ( .A(_abc_15497_new_n1395_), .B(_abc_15497_new_n883__bF_buf3), .Y(_abc_15497_new_n2573_));
NOR2X1 NOR2X1_46 ( .A(_abc_15497_new_n813_), .B(_abc_15497_new_n816_), .Y(_abc_15497_new_n817_));
NOR2X1 NOR2X1_460 ( .A(_abc_15497_new_n1422_), .B(_abc_15497_new_n883__bF_buf2), .Y(_abc_15497_new_n2579_));
NOR2X1 NOR2X1_461 ( .A(_abc_15497_new_n1444_), .B(_abc_15497_new_n883__bF_buf0), .Y(_abc_15497_new_n2585_));
NOR2X1 NOR2X1_462 ( .A(_abc_15497_new_n1452_), .B(_abc_15497_new_n883__bF_buf13), .Y(_abc_15497_new_n2588_));
NOR2X1 NOR2X1_463 ( .A(_abc_15497_new_n1477_), .B(_abc_15497_new_n883__bF_buf11), .Y(_abc_15497_new_n2594_));
NOR2X1 NOR2X1_464 ( .A(_abc_15497_new_n1492_), .B(_abc_15497_new_n883__bF_buf10), .Y(_abc_15497_new_n2597_));
NOR2X1 NOR2X1_465 ( .A(_abc_15497_new_n1528_), .B(_abc_15497_new_n883__bF_buf8), .Y(_abc_15497_new_n2606_));
NOR2X1 NOR2X1_466 ( .A(_abc_15497_new_n1540_), .B(_abc_15497_new_n883__bF_buf7), .Y(_abc_15497_new_n2609_));
NOR2X1 NOR2X1_467 ( .A(_abc_15497_new_n1550_), .B(_abc_15497_new_n883__bF_buf6), .Y(_abc_15497_new_n2612_));
NOR2X1 NOR2X1_468 ( .A(_abc_15497_new_n1569_), .B(_abc_15497_new_n883__bF_buf5), .Y(_abc_15497_new_n2615_));
NOR2X1 NOR2X1_469 ( .A(_abc_15497_new_n1580_), .B(_abc_15497_new_n883__bF_buf4), .Y(_abc_15497_new_n2618_));
NOR2X1 NOR2X1_47 ( .A(_abc_15497_new_n818_), .B(_abc_15497_new_n805_), .Y(_abc_15497_new_n819_));
NOR2X1 NOR2X1_470 ( .A(_abc_15497_new_n1593_), .B(_abc_15497_new_n883__bF_buf3), .Y(_abc_15497_new_n2621_));
NOR2X1 NOR2X1_471 ( .A(_abc_15497_new_n1621_), .B(_abc_15497_new_n883__bF_buf1), .Y(_abc_15497_new_n2627_));
NOR2X1 NOR2X1_472 ( .A(_abc_15497_new_n1628_), .B(_abc_15497_new_n883__bF_buf0), .Y(_abc_15497_new_n2631_));
NOR2X1 NOR2X1_473 ( .A(_abc_15497_new_n770_), .B(_abc_15497_new_n883__bF_buf12), .Y(_abc_15497_new_n2639_));
NOR2X1 NOR2X1_474 ( .A(_abc_15497_new_n742_), .B(_abc_15497_new_n883__bF_buf6), .Y(_abc_15497_new_n2663_));
NOR2X1 NOR2X1_475 ( .A(_abc_15497_new_n739_), .B(_abc_15497_new_n883__bF_buf5), .Y(_abc_15497_new_n2666_));
NOR2X1 NOR2X1_476 ( .A(_abc_15497_new_n709_), .B(_abc_15497_new_n883__bF_buf2), .Y(_abc_15497_new_n2678_));
NOR2X1 NOR2X1_477 ( .A(_abc_15497_new_n833_), .B(_abc_15497_new_n883__bF_buf0), .Y(_abc_15497_new_n2687_));
NOR2X1 NOR2X1_478 ( .A(_abc_15497_new_n824_), .B(_abc_15497_new_n883__bF_buf12), .Y(_abc_15497_new_n2693_));
NOR2X1 NOR2X1_479 ( .A(_abc_15497_new_n799_), .B(_abc_15497_new_n883__bF_buf8), .Y(_abc_15497_new_n2705_));
NOR2X1 NOR2X1_48 ( .A(c_reg_19_), .B(_auto_iopadmap_cc_368_execute_22625_83_), .Y(_abc_15497_new_n821_));
NOR2X1 NOR2X1_480 ( .A(_abc_15497_new_n856_), .B(_abc_15497_new_n883__bF_buf6), .Y(_abc_15497_new_n2711_));
NOR2X1 NOR2X1_481 ( .A(_abc_15497_new_n850_), .B(_abc_15497_new_n883__bF_buf5), .Y(_abc_15497_new_n2714_));
NOR2X1 NOR2X1_482 ( .A(_abc_15497_new_n698_), .B(_abc_15497_new_n883__bF_buf4), .Y(_abc_15497_new_n2717_));
NOR2X1 NOR2X1_483 ( .A(_abc_15497_new_n901_), .B(_abc_15497_new_n883__bF_buf1), .Y(_abc_15497_new_n2726_));
NOR2X1 NOR2X1_484 ( .A(_abc_15497_new_n911_), .B(_abc_15497_new_n883__bF_buf0), .Y(_abc_15497_new_n2729_));
NOR2X1 NOR2X1_485 ( .A(b_reg_0_), .B(c_reg_0_), .Y(_abc_15497_new_n2746_));
NOR2X1 NOR2X1_486 ( .A(e_reg_0_), .B(a_reg_27_), .Y(_abc_15497_new_n2763_));
NOR2X1 NOR2X1_487 ( .A(_abc_15497_new_n2763_), .B(_abc_15497_new_n2765_), .Y(_abc_15497_new_n2766_));
NOR2X1 NOR2X1_488 ( .A(_abc_15497_new_n2767_), .B(_abc_15497_new_n2761_), .Y(_abc_15497_new_n2768_));
NOR2X1 NOR2X1_489 ( .A(_abc_15497_new_n2768_), .B(_abc_15497_new_n2772_), .Y(_abc_15497_new_n2773_));
NOR2X1 NOR2X1_49 ( .A(_abc_15497_new_n821_), .B(_abc_15497_new_n820_), .Y(_abc_15497_new_n822_));
NOR2X1 NOR2X1_490 ( .A(_abc_15497_new_n1646_), .B(_abc_15497_new_n2774_), .Y(_abc_15497_new_n2775_));
NOR2X1 NOR2X1_491 ( .A(b_reg_1_), .B(c_reg_1_), .Y(_abc_15497_new_n2782_));
NOR2X1 NOR2X1_492 ( .A(e_reg_1_), .B(a_reg_28_), .Y(_abc_15497_new_n2793_));
NOR2X1 NOR2X1_493 ( .A(_abc_15497_new_n2774_), .B(_abc_15497_new_n2817_), .Y(_abc_15497_new_n2818_));
NOR2X1 NOR2X1_494 ( .A(_abc_15497_new_n2097_), .B(_abc_15497_new_n883__bF_buf11), .Y(_abc_15497_new_n2823_));
NOR2X1 NOR2X1_495 ( .A(b_reg_2_), .B(c_reg_2_), .Y(_abc_15497_new_n2830_));
NOR2X1 NOR2X1_496 ( .A(e_reg_2_), .B(a_reg_29_), .Y(_abc_15497_new_n2841_));
NOR2X1 NOR2X1_497 ( .A(_abc_15497_new_n2103_), .B(_abc_15497_new_n883__bF_buf10), .Y(_abc_15497_new_n2880_));
NOR2X1 NOR2X1_498 ( .A(b_reg_3_), .B(c_reg_3_), .Y(_abc_15497_new_n2889_));
NOR2X1 NOR2X1_499 ( .A(_abc_15497_new_n2903_), .B(_abc_15497_new_n2904_), .Y(_abc_15497_new_n2908_));
NOR2X1 NOR2X1_5 ( .A(_abc_15497_new_n705_), .B(_abc_15497_new_n704_), .Y(_abc_15497_new_n706_));
NOR2X1 NOR2X1_50 ( .A(_abc_15497_new_n823_), .B(_abc_15497_new_n824_), .Y(_abc_15497_new_n825_));
NOR2X1 NOR2X1_500 ( .A(_abc_15497_new_n2112_), .B(_abc_15497_new_n883__bF_buf9), .Y(_abc_15497_new_n2937_));
NOR2X1 NOR2X1_501 ( .A(b_reg_4_), .B(c_reg_4_), .Y(_abc_15497_new_n2946_));
NOR2X1 NOR2X1_502 ( .A(e_reg_4_), .B(a_reg_31_), .Y(_abc_15497_new_n2958_));
NOR2X1 NOR2X1_503 ( .A(_abc_15497_new_n2954_), .B(_abc_15497_new_n2971_), .Y(_abc_15497_new_n2972_));
NOR2X1 NOR2X1_504 ( .A(_abc_15497_new_n2980_), .B(_abc_15497_new_n2971_), .Y(_abc_15497_new_n2981_));
NOR2X1 NOR2X1_505 ( .A(_abc_15497_new_n2954_), .B(_abc_15497_new_n2982_), .Y(_abc_15497_new_n2983_));
NOR2X1 NOR2X1_506 ( .A(_abc_15497_new_n2994_), .B(_abc_15497_new_n2942_), .Y(_abc_15497_new_n2995_));
NOR2X1 NOR2X1_507 ( .A(_abc_15497_new_n2122_), .B(_abc_15497_new_n883__bF_buf8), .Y(_abc_15497_new_n2999_));
NOR2X1 NOR2X1_508 ( .A(b_reg_5_), .B(c_reg_5_), .Y(_abc_15497_new_n3008_));
NOR2X1 NOR2X1_509 ( .A(e_reg_5_), .B(a_reg_0_), .Y(_abc_15497_new_n3019_));
NOR2X1 NOR2X1_51 ( .A(c_reg_18_), .B(_auto_iopadmap_cc_368_execute_22625_82_), .Y(_abc_15497_new_n826_));
NOR2X1 NOR2X1_510 ( .A(_abc_15497_new_n2975_), .B(_abc_15497_new_n3046_), .Y(_abc_15497_new_n3047_));
NOR2X1 NOR2X1_511 ( .A(_abc_15497_new_n2129_), .B(_abc_15497_new_n883__bF_buf7), .Y(_abc_15497_new_n3055_));
NOR2X1 NOR2X1_512 ( .A(_abc_15497_new_n2997_), .B(_abc_15497_new_n3052_), .Y(_abc_15497_new_n3058_));
NOR2X1 NOR2X1_513 ( .A(b_reg_6_), .B(c_reg_6_), .Y(_abc_15497_new_n3066_));
NOR2X1 NOR2X1_514 ( .A(e_reg_6_), .B(a_reg_1_), .Y(_abc_15497_new_n3077_));
NOR2X1 NOR2X1_515 ( .A(_abc_15497_new_n3108_), .B(_abc_15497_new_n3063_), .Y(_abc_15497_new_n3109_));
NOR2X1 NOR2X1_516 ( .A(_abc_15497_new_n2141_), .B(_abc_15497_new_n883__bF_buf6), .Y(_abc_15497_new_n3113_));
NOR2X1 NOR2X1_517 ( .A(b_reg_7_), .B(c_reg_7_), .Y(_abc_15497_new_n3120_));
NOR2X1 NOR2X1_518 ( .A(e_reg_7_), .B(a_reg_2_), .Y(_abc_15497_new_n3132_));
NOR2X1 NOR2X1_519 ( .A(_abc_15497_new_n3143_), .B(_abc_15497_new_n3129_), .Y(_abc_15497_new_n3144_));
NOR2X1 NOR2X1_52 ( .A(_abc_15497_new_n826_), .B(_abc_15497_new_n825_), .Y(_abc_15497_new_n827_));
NOR2X1 NOR2X1_520 ( .A(_abc_15497_new_n3147_), .B(_abc_15497_new_n3150_), .Y(_abc_15497_new_n3151_));
NOR2X1 NOR2X1_521 ( .A(_abc_15497_new_n3150_), .B(_abc_15497_new_n3129_), .Y(_abc_15497_new_n3155_));
NOR2X1 NOR2X1_522 ( .A(_abc_15497_new_n3147_), .B(_abc_15497_new_n3143_), .Y(_abc_15497_new_n3156_));
NOR2X1 NOR2X1_523 ( .A(_abc_15497_new_n2151_), .B(_abc_15497_new_n883__bF_buf5), .Y(_abc_15497_new_n3164_));
NOR2X1 NOR2X1_524 ( .A(b_reg_8_), .B(c_reg_8_), .Y(_abc_15497_new_n3170_));
NOR2X1 NOR2X1_525 ( .A(e_reg_8_), .B(a_reg_3_), .Y(_abc_15497_new_n3180_));
NOR2X1 NOR2X1_526 ( .A(_abc_15497_new_n1646_), .B(_abc_15497_new_n3218_), .Y(_abc_15497_new_n3219_));
NOR2X1 NOR2X1_527 ( .A(_abc_15497_new_n3226_), .B(_abc_15497_new_n3218_), .Y(_abc_15497_new_n3227_));
NOR2X1 NOR2X1_528 ( .A(b_reg_9_), .B(c_reg_9_), .Y(_abc_15497_new_n3235_));
NOR2X1 NOR2X1_529 ( .A(e_reg_9_), .B(a_reg_4_), .Y(_abc_15497_new_n3243_));
NOR2X1 NOR2X1_53 ( .A(c_reg_17_), .B(_auto_iopadmap_cc_368_execute_22625_81_), .Y(_abc_15497_new_n830_));
NOR2X1 NOR2X1_530 ( .A(_abc_15497_new_n3241_), .B(_abc_15497_new_n3249_), .Y(_abc_15497_new_n3250_));
NOR2X1 NOR2X1_531 ( .A(b_reg_10_), .B(c_reg_10_), .Y(_abc_15497_new_n3291_));
NOR2X1 NOR2X1_532 ( .A(e_reg_10_), .B(a_reg_5_), .Y(_abc_15497_new_n3303_));
NOR2X1 NOR2X1_533 ( .A(_abc_15497_new_n2742__bF_buf0), .B(_abc_15497_new_n3239_), .Y(_abc_15497_new_n3328_));
NOR2X1 NOR2X1_534 ( .A(_abc_15497_new_n2180_), .B(_abc_15497_new_n883__bF_buf3), .Y(_abc_15497_new_n3345_));
NOR2X1 NOR2X1_535 ( .A(b_reg_11_), .B(c_reg_11_), .Y(_abc_15497_new_n3352_));
NOR2X1 NOR2X1_536 ( .A(e_reg_11_), .B(a_reg_6_), .Y(_abc_15497_new_n3362_));
NOR2X1 NOR2X1_537 ( .A(_abc_15497_new_n3378_), .B(_abc_15497_new_n3375_), .Y(_abc_15497_new_n3379_));
NOR2X1 NOR2X1_538 ( .A(_abc_15497_new_n2197_), .B(_abc_15497_new_n883__bF_buf2), .Y(_abc_15497_new_n3400_));
NOR2X1 NOR2X1_539 ( .A(b_reg_12_), .B(c_reg_12_), .Y(_abc_15497_new_n3419_));
NOR2X1 NOR2X1_54 ( .A(_abc_15497_new_n830_), .B(_abc_15497_new_n829_), .Y(_abc_15497_new_n831_));
NOR2X1 NOR2X1_540 ( .A(e_reg_12_), .B(a_reg_7_), .Y(_abc_15497_new_n3432_));
NOR2X1 NOR2X1_541 ( .A(_abc_15497_new_n3471_), .B(_abc_15497_new_n3409_), .Y(_abc_15497_new_n3472_));
NOR2X1 NOR2X1_542 ( .A(_abc_15497_new_n2203_), .B(_abc_15497_new_n883__bF_buf1), .Y(_abc_15497_new_n3475_));
NOR2X1 NOR2X1_543 ( .A(b_reg_13_), .B(c_reg_13_), .Y(_abc_15497_new_n3481_));
NOR2X1 NOR2X1_544 ( .A(e_reg_13_), .B(a_reg_8_), .Y(_abc_15497_new_n3495_));
NOR2X1 NOR2X1_545 ( .A(_abc_15497_new_n3493_), .B(_abc_15497_new_n3501_), .Y(_abc_15497_new_n3502_));
NOR2X1 NOR2X1_546 ( .A(_abc_15497_new_n3537_), .B(_abc_15497_new_n3527_), .Y(_abc_15497_new_n3538_));
NOR2X1 NOR2X1_547 ( .A(b_reg_14_), .B(c_reg_14_), .Y(_abc_15497_new_n3544_));
NOR2X1 NOR2X1_548 ( .A(e_reg_14_), .B(a_reg_9_), .Y(_abc_15497_new_n3560_));
NOR2X1 NOR2X1_549 ( .A(_abc_15497_new_n3596_), .B(_abc_15497_new_n3540_), .Y(_abc_15497_new_n3597_));
NOR2X1 NOR2X1_55 ( .A(_abc_15497_new_n832_), .B(_abc_15497_new_n833_), .Y(_abc_15497_new_n834_));
NOR2X1 NOR2X1_550 ( .A(_abc_15497_new_n2228_), .B(_abc_15497_new_n883__bF_buf13), .Y(_abc_15497_new_n3600_));
NOR2X1 NOR2X1_551 ( .A(b_reg_15_), .B(c_reg_15_), .Y(_abc_15497_new_n3612_));
NOR2X1 NOR2X1_552 ( .A(_abc_15497_new_n3614_), .B(_abc_15497_new_n2925__bF_buf2), .Y(_abc_15497_new_n3615_));
NOR2X1 NOR2X1_553 ( .A(e_reg_15_), .B(a_reg_10_), .Y(_abc_15497_new_n3623_));
NOR2X1 NOR2X1_554 ( .A(_abc_15497_new_n2241_), .B(_abc_15497_new_n883__bF_buf12), .Y(_abc_15497_new_n3665_));
NOR2X1 NOR2X1_555 ( .A(_abc_15497_new_n3408_), .B(_abc_15497_new_n3669_), .Y(_abc_15497_new_n3674_));
NOR2X1 NOR2X1_556 ( .A(_abc_15497_new_n3646_), .B(_abc_15497_new_n3658_), .Y(_abc_15497_new_n3677_));
NOR2X1 NOR2X1_557 ( .A(c_reg_16_), .B(_abc_15497_new_n3682_), .Y(_abc_15497_new_n3684_));
NOR2X1 NOR2X1_558 ( .A(_abc_15497_new_n3714_), .B(_abc_15497_new_n3675_), .Y(_abc_15497_new_n3715_));
NOR2X1 NOR2X1_559 ( .A(_abc_15497_new_n1646_), .B(_abc_15497_new_n3715_), .Y(_abc_15497_new_n3716_));
NOR2X1 NOR2X1_56 ( .A(c_reg_16_), .B(_auto_iopadmap_cc_368_execute_22625_80_), .Y(_abc_15497_new_n841_));
NOR2X1 NOR2X1_560 ( .A(_abc_15497_new_n3711_), .B(_abc_15497_new_n3715_), .Y(_abc_15497_new_n3721_));
NOR2X1 NOR2X1_561 ( .A(b_reg_17_), .B(c_reg_17_), .Y(_abc_15497_new_n3727_));
NOR2X1 NOR2X1_562 ( .A(_abc_15497_new_n1112_), .B(_abc_15497_new_n2207_), .Y(_abc_15497_new_n3736_));
NOR2X1 NOR2X1_563 ( .A(_abc_15497_new_n3692_), .B(_abc_15497_new_n3693_), .Y(_abc_15497_new_n3737_));
NOR2X1 NOR2X1_564 ( .A(e_reg_17_), .B(a_reg_12_), .Y(_abc_15497_new_n3739_));
NOR2X1 NOR2X1_565 ( .A(_abc_15497_new_n1121_), .B(_abc_15497_new_n2214_), .Y(_abc_15497_new_n3740_));
NOR2X1 NOR2X1_566 ( .A(_abc_15497_new_n3739_), .B(_abc_15497_new_n3740_), .Y(_abc_15497_new_n3742_));
NOR2X1 NOR2X1_567 ( .A(_abc_15497_new_n3736_), .B(_abc_15497_new_n3737_), .Y(_abc_15497_new_n3746_));
NOR2X1 NOR2X1_568 ( .A(_abc_15497_new_n3751_), .B(_abc_15497_new_n3752_), .Y(_abc_15497_new_n3757_));
NOR2X1 NOR2X1_569 ( .A(_abc_15497_new_n3735_), .B(_abc_15497_new_n3749_), .Y(_abc_15497_new_n3758_));
NOR2X1 NOR2X1_57 ( .A(_abc_15497_new_n841_), .B(_abc_15497_new_n834_), .Y(_abc_15497_new_n842_));
NOR2X1 NOR2X1_570 ( .A(_abc_15497_new_n2267_), .B(_abc_15497_new_n883__bF_buf10), .Y(_abc_15497_new_n3773_));
NOR2X1 NOR2X1_571 ( .A(_abc_15497_new_n2925__bF_buf3), .B(_abc_15497_new_n3788_), .Y(_abc_15497_new_n3789_));
NOR2X1 NOR2X1_572 ( .A(_abc_15497_new_n3794_), .B(_abc_15497_new_n3789_), .Y(_abc_15497_new_n3795_));
NOR2X1 NOR2X1_573 ( .A(_abc_15497_new_n3816_), .B(_abc_15497_new_n3814_), .Y(_abc_15497_new_n3824_));
NOR2X1 NOR2X1_574 ( .A(_abc_15497_new_n2925__bF_buf2), .B(_abc_15497_new_n3831_), .Y(_abc_15497_new_n3832_));
NOR2X1 NOR2X1_575 ( .A(_abc_15497_new_n3839_), .B(_abc_15497_new_n3832_), .Y(_abc_15497_new_n3848_));
NOR2X1 NOR2X1_576 ( .A(_abc_15497_new_n2293_), .B(_abc_15497_new_n883__bF_buf9), .Y(_abc_15497_new_n3867_));
NOR2X1 NOR2X1_577 ( .A(_abc_15497_new_n1130_), .B(_abc_15497_new_n3531_), .Y(_abc_15497_new_n3888_));
NOR2X1 NOR2X1_578 ( .A(c_reg_20_), .B(_abc_15497_new_n3894_), .Y(_abc_15497_new_n3896_));
NOR2X1 NOR2X1_579 ( .A(_abc_15497_new_n3928_), .B(_abc_15497_new_n3885_), .Y(_abc_15497_new_n3929_));
NOR2X1 NOR2X1_58 ( .A(_abc_15497_new_n840_), .B(_abc_15497_new_n843_), .Y(_abc_15497_new_n844_));
NOR2X1 NOR2X1_580 ( .A(_abc_15497_new_n2303_), .B(_abc_15497_new_n883__bF_buf8), .Y(_abc_15497_new_n3932_));
NOR2X1 NOR2X1_581 ( .A(_abc_15497_new_n1146_), .B(_abc_15497_new_n2230_), .Y(_abc_15497_new_n3938_));
NOR2X1 NOR2X1_582 ( .A(c_reg_21_), .B(_abc_15497_new_n3944_), .Y(_abc_15497_new_n3946_));
NOR2X1 NOR2X1_583 ( .A(_abc_15497_new_n2317_), .B(_abc_15497_new_n883__bF_buf7), .Y(_abc_15497_new_n3983_));
NOR2X1 NOR2X1_584 ( .A(_abc_15497_new_n1162_), .B(_abc_15497_new_n2244_), .Y(_abc_15497_new_n3993_));
NOR2X1 NOR2X1_585 ( .A(c_reg_22_), .B(_abc_15497_new_n3999_), .Y(_abc_15497_new_n4001_));
NOR2X1 NOR2X1_586 ( .A(_abc_15497_new_n4041_), .B(_abc_15497_new_n4042_), .Y(_abc_15497_new_n4043_));
NOR2X1 NOR2X1_587 ( .A(_abc_15497_new_n1173_), .B(_abc_15497_new_n2258_), .Y(_abc_15497_new_n4045_));
NOR2X1 NOR2X1_588 ( .A(b_reg_23_), .B(c_reg_23_), .Y(_abc_15497_new_n4050_));
NOR2X1 NOR2X1_589 ( .A(_abc_15497_new_n4060_), .B(_abc_15497_new_n2270_), .Y(_abc_15497_new_n4061_));
NOR2X1 NOR2X1_59 ( .A(_abc_15497_new_n828_), .B(_abc_15497_new_n845_), .Y(_abc_15497_new_n846_));
NOR2X1 NOR2X1_590 ( .A(_abc_15497_new_n2341_), .B(_abc_15497_new_n883__bF_buf6), .Y(_abc_15497_new_n4094_));
NOR2X1 NOR2X1_591 ( .A(b_reg_24_), .B(c_reg_24_), .Y(_abc_15497_new_n4109_));
NOR2X1 NOR2X1_592 ( .A(_abc_15497_new_n4118_), .B(_abc_15497_new_n2284_), .Y(_abc_15497_new_n4119_));
NOR2X1 NOR2X1_593 ( .A(e_reg_24_), .B(a_reg_19_), .Y(_abc_15497_new_n4123_));
NOR2X1 NOR2X1_594 ( .A(_abc_15497_new_n1213_), .B(_abc_15497_new_n2296_), .Y(_abc_15497_new_n4124_));
NOR2X1 NOR2X1_595 ( .A(_abc_15497_new_n4123_), .B(_abc_15497_new_n4124_), .Y(_abc_15497_new_n4126_));
NOR2X1 NOR2X1_596 ( .A(_abc_15497_new_n4108_), .B(_abc_15497_new_n4132_), .Y(_abc_15497_new_n4133_));
NOR2X1 NOR2X1_597 ( .A(_abc_15497_new_n4133_), .B(_abc_15497_new_n4135_), .Y(_abc_15497_new_n4136_));
NOR2X1 NOR2X1_598 ( .A(b_reg_25_), .B(c_reg_25_), .Y(_abc_15497_new_n4154_));
NOR2X1 NOR2X1_599 ( .A(e_reg_25_), .B(a_reg_20_), .Y(_abc_15497_new_n4164_));
NOR2X1 NOR2X1_6 ( .A(_abc_15497_new_n708_), .B(_abc_15497_new_n709_), .Y(_abc_15497_new_n710_));
NOR2X1 NOR2X1_60 ( .A(_abc_15497_new_n849_), .B(_abc_15497_new_n850_), .Y(_abc_15497_new_n851_));
NOR2X1 NOR2X1_600 ( .A(_abc_15497_new_n4165_), .B(_abc_15497_new_n2310_), .Y(_abc_15497_new_n4166_));
NOR2X1 NOR2X1_601 ( .A(_abc_15497_new_n4164_), .B(_abc_15497_new_n4166_), .Y(_abc_15497_new_n4167_));
NOR2X1 NOR2X1_602 ( .A(_abc_15497_new_n4153_), .B(_abc_15497_new_n4172_), .Y(_abc_15497_new_n4173_));
NOR2X1 NOR2X1_603 ( .A(d_reg_26_), .B(_abc_15497_new_n4197_), .Y(_abc_15497_new_n4198_));
NOR2X1 NOR2X1_604 ( .A(e_reg_26_), .B(a_reg_21_), .Y(_abc_15497_new_n4208_));
NOR2X1 NOR2X1_605 ( .A(_abc_15497_new_n1239_), .B(_abc_15497_new_n2321_), .Y(_abc_15497_new_n4209_));
NOR2X1 NOR2X1_606 ( .A(_abc_15497_new_n4208_), .B(_abc_15497_new_n4209_), .Y(_abc_15497_new_n4211_));
NOR2X1 NOR2X1_607 ( .A(_abc_15497_new_n4193_), .B(_abc_15497_new_n4215_), .Y(_abc_15497_new_n4216_));
NOR2X1 NOR2X1_608 ( .A(_abc_15497_new_n4216_), .B(_abc_15497_new_n4217_), .Y(_abc_15497_new_n4218_));
NOR2X1 NOR2X1_609 ( .A(e_reg_27_), .B(a_reg_22_), .Y(_abc_15497_new_n4252_));
NOR2X1 NOR2X1_61 ( .A(c_reg_25_), .B(_auto_iopadmap_cc_368_execute_22625_89_), .Y(_abc_15497_new_n852_));
NOR2X1 NOR2X1_610 ( .A(_abc_15497_new_n1250_), .B(_abc_15497_new_n2332_), .Y(_abc_15497_new_n4253_));
NOR2X1 NOR2X1_611 ( .A(_abc_15497_new_n4260_), .B(_abc_15497_new_n4235_), .Y(_abc_15497_new_n4261_));
NOR2X1 NOR2X1_612 ( .A(_abc_15497_new_n4261_), .B(_abc_15497_new_n4262_), .Y(_abc_15497_new_n4263_));
NOR2X1 NOR2X1_613 ( .A(_abc_15497_new_n2393_), .B(_abc_15497_new_n883__bF_buf3), .Y(_abc_15497_new_n4266_));
NOR2X1 NOR2X1_614 ( .A(_abc_15497_new_n4270_), .B(_abc_15497_new_n4269_), .Y(_abc_15497_new_n4271_));
NOR2X1 NOR2X1_615 ( .A(_abc_15497_new_n4173_), .B(_abc_15497_new_n4231_), .Y(_abc_15497_new_n4272_));
NOR2X1 NOR2X1_616 ( .A(c_reg_28_), .B(b_reg_28_), .Y(_abc_15497_new_n4282_));
NOR2X1 NOR2X1_617 ( .A(_abc_15497_new_n4282_), .B(_abc_15497_new_n4281_), .Y(_abc_15497_new_n4283_));
NOR2X1 NOR2X1_618 ( .A(d_reg_28_), .B(_abc_15497_new_n4281_), .Y(_abc_15497_new_n4285_));
NOR2X1 NOR2X1_619 ( .A(_abc_15497_new_n4282_), .B(_abc_15497_new_n4285_), .Y(_abc_15497_new_n4287_));
NOR2X1 NOR2X1_62 ( .A(_abc_15497_new_n852_), .B(_abc_15497_new_n851_), .Y(_abc_15497_new_n853_));
NOR2X1 NOR2X1_620 ( .A(_abc_15497_new_n4251_), .B(_abc_15497_new_n4254_), .Y(_abc_15497_new_n4290_));
NOR2X1 NOR2X1_621 ( .A(_abc_15497_new_n4253_), .B(_abc_15497_new_n4290_), .Y(_abc_15497_new_n4291_));
NOR2X1 NOR2X1_622 ( .A(e_reg_28_), .B(a_reg_23_), .Y(_abc_15497_new_n4292_));
NOR2X1 NOR2X1_623 ( .A(_abc_15497_new_n1736_), .B(_abc_15497_new_n2349_), .Y(_abc_15497_new_n4293_));
NOR2X1 NOR2X1_624 ( .A(_abc_15497_new_n4292_), .B(_abc_15497_new_n4293_), .Y(_abc_15497_new_n4294_));
NOR2X1 NOR2X1_625 ( .A(_abc_15497_new_n4277_), .B(_abc_15497_new_n4301_), .Y(_abc_15497_new_n4302_));
NOR2X1 NOR2X1_626 ( .A(_abc_15497_new_n3285_), .B(_abc_15497_new_n4306_), .Y(_abc_15497_new_n4307_));
NOR2X1 NOR2X1_627 ( .A(_abc_15497_new_n4309_), .B(_abc_15497_new_n4308_), .Y(_abc_15497_new_n4310_));
NOR2X1 NOR2X1_628 ( .A(_abc_15497_new_n4313_), .B(_abc_15497_new_n3884_), .Y(_abc_15497_new_n4314_));
NOR2X1 NOR2X1_629 ( .A(_abc_15497_new_n4302_), .B(_abc_15497_new_n4303_), .Y(_abc_15497_new_n4318_));
NOR2X1 NOR2X1_63 ( .A(_abc_15497_new_n855_), .B(_abc_15497_new_n856_), .Y(_abc_15497_new_n857_));
NOR2X1 NOR2X1_630 ( .A(_abc_15497_new_n2401_), .B(_abc_15497_new_n883__bF_buf2), .Y(_abc_15497_new_n4321_));
NOR2X1 NOR2X1_631 ( .A(_abc_15497_new_n904_), .B(_abc_15497_new_n4330_), .Y(_abc_15497_new_n4331_));
NOR2X1 NOR2X1_632 ( .A(c_reg_29_), .B(b_reg_29_), .Y(_abc_15497_new_n4334_));
NOR2X1 NOR2X1_633 ( .A(_abc_15497_new_n4334_), .B(_abc_15497_new_n4331_), .Y(_abc_15497_new_n4335_));
NOR2X1 NOR2X1_634 ( .A(e_reg_29_), .B(a_reg_24_), .Y(_abc_15497_new_n4344_));
NOR2X1 NOR2X1_635 ( .A(_abc_15497_new_n1273_), .B(_abc_15497_new_n2360_), .Y(_abc_15497_new_n4345_));
NOR2X1 NOR2X1_636 ( .A(_abc_15497_new_n4344_), .B(_abc_15497_new_n4345_), .Y(_abc_15497_new_n4346_));
NOR2X1 NOR2X1_637 ( .A(_abc_15497_new_n912_), .B(_abc_15497_new_n4372_), .Y(_abc_15497_new_n4373_));
NOR2X1 NOR2X1_638 ( .A(c_reg_30_), .B(b_reg_30_), .Y(_abc_15497_new_n4376_));
NOR2X1 NOR2X1_639 ( .A(_abc_15497_new_n4376_), .B(_abc_15497_new_n4373_), .Y(_abc_15497_new_n4377_));
NOR2X1 NOR2X1_64 ( .A(c_reg_24_), .B(_auto_iopadmap_cc_368_execute_22625_88_), .Y(_abc_15497_new_n858_));
NOR2X1 NOR2X1_640 ( .A(e_reg_30_), .B(a_reg_25_), .Y(_abc_15497_new_n4387_));
NOR2X1 NOR2X1_641 ( .A(_abc_15497_new_n4388_), .B(_abc_15497_new_n2372_), .Y(_abc_15497_new_n4389_));
NOR2X1 NOR2X1_642 ( .A(_abc_15497_new_n4387_), .B(_abc_15497_new_n4389_), .Y(_abc_15497_new_n4390_));
NOR2X1 NOR2X1_643 ( .A(c_reg_31_), .B(b_reg_31_), .Y(_abc_15497_new_n4419_));
NOR2X1 NOR2X1_644 ( .A(_abc_15497_new_n4419_), .B(_abc_15497_new_n4418_), .Y(_abc_15497_new_n4420_));
NOR2X1 NOR2X1_645 ( .A(_abc_15497_new_n2438_), .B(_abc_15497_new_n883__bF_buf1), .Y(_abc_15497_new_n4438_));
NOR2X1 NOR2X1_646 ( .A(round_ctr_reg_5_), .B(round_ctr_reg_4_), .Y(_abc_15497_new_n4441_));
NOR2X1 NOR2X1_647 ( .A(_abc_15497_new_n4442_), .B(_abc_15497_new_n4443_), .Y(_abc_15497_new_n4444_));
NOR2X1 NOR2X1_648 ( .A(_abc_15497_new_n1646_), .B(_abc_15497_new_n4447_), .Y(_abc_15497_abc_9717_auto_fsm_map_cc_118_implement_pattern_cache_863));
NOR2X1 NOR2X1_649 ( .A(round_ctr_reg_2_), .B(_abc_15497_new_n4444_), .Y(_abc_15497_new_n4458_));
NOR2X1 NOR2X1_65 ( .A(_abc_15497_new_n858_), .B(_abc_15497_new_n857_), .Y(_abc_15497_new_n859_));
NOR2X1 NOR2X1_650 ( .A(_abc_15497_new_n4458_), .B(_abc_15497_new_n4460_), .Y(_0round_ctr_reg_6_0__2_));
NOR2X1 NOR2X1_651 ( .A(_abc_15497_new_n1646_), .B(_abc_15497_new_n4445_), .Y(_abc_15497_new_n4464_));
NOR2X1 NOR2X1_652 ( .A(_abc_15497_new_n2740_), .B(_abc_15497_new_n4468_), .Y(_abc_15497_new_n4470_));
NOR2X1 NOR2X1_653 ( .A(c_reg_0_), .B(_auto_iopadmap_cc_368_execute_22625_64_), .Y(_abc_15497_new_n4476_));
NOR2X1 NOR2X1_654 ( .A(_auto_iopadmap_cc_368_execute_22625_65_), .B(_abc_15497_new_n883__bF_buf0), .Y(_abc_15497_new_n4479_));
NOR2X1 NOR2X1_655 ( .A(_auto_iopadmap_cc_368_execute_22625_66_), .B(_abc_15497_new_n883__bF_buf13), .Y(_abc_15497_new_n4482_));
NOR2X1 NOR2X1_656 ( .A(_abc_15497_new_n766_), .B(_abc_15497_new_n4485_), .Y(_abc_15497_new_n4486_));
NOR2X1 NOR2X1_657 ( .A(_auto_iopadmap_cc_368_execute_22625_68_), .B(_abc_15497_new_n883__bF_buf11), .Y(_abc_15497_new_n4490_));
NOR2X1 NOR2X1_658 ( .A(_abc_15497_new_n763_), .B(_abc_15497_new_n761_), .Y(_abc_15497_new_n4493_));
NOR2X1 NOR2X1_659 ( .A(_abc_15497_new_n4493_), .B(_abc_15497_new_n781_), .Y(_abc_15497_new_n4495_));
NOR2X1 NOR2X1_66 ( .A(_abc_15497_new_n854_), .B(_abc_15497_new_n860_), .Y(_abc_15497_new_n861_));
NOR2X1 NOR2X1_660 ( .A(_abc_15497_new_n786_), .B(_abc_15497_new_n4511_), .Y(_abc_15497_new_n4512_));
NOR2X1 NOR2X1_661 ( .A(_abc_15497_new_n720_), .B(_abc_15497_new_n4530_), .Y(_abc_15497_new_n4531_));
NOR2X1 NOR2X1_662 ( .A(_abc_15497_new_n706_), .B(_abc_15497_new_n4539_), .Y(_abc_15497_new_n4540_));
NOR2X1 NOR2X1_663 ( .A(_abc_15497_new_n842_), .B(_abc_15497_new_n792_), .Y(_abc_15497_new_n4549_));
NOR2X1 NOR2X1_664 ( .A(_abc_15497_new_n815_), .B(_abc_15497_new_n4565_), .Y(_abc_15497_new_n4566_));
NOR2X1 NOR2X1_665 ( .A(_abc_15497_new_n837_), .B(_abc_15497_new_n4564_), .Y(_abc_15497_new_n4567_));
NOR2X1 NOR2X1_666 ( .A(_abc_15497_new_n809_), .B(_abc_15497_new_n4571_), .Y(_abc_15497_new_n4573_));
NOR2X1 NOR2X1_667 ( .A(_abc_15497_new_n802_), .B(_abc_15497_new_n4577_), .Y(_abc_15497_new_n4578_));
NOR2X1 NOR2X1_668 ( .A(_auto_iopadmap_cc_368_execute_22625_87_), .B(_abc_15497_new_n883__bF_buf12), .Y(_abc_15497_new_n4582_));
NOR2X1 NOR2X1_669 ( .A(_abc_15497_new_n860_), .B(_abc_15497_new_n848_), .Y(_abc_15497_new_n4591_));
NOR2X1 NOR2X1_67 ( .A(_auto_iopadmap_cc_368_execute_22625_90_), .B(c_reg_26_), .Y(_abc_15497_new_n865_));
NOR2X1 NOR2X1_670 ( .A(_abc_15497_new_n857_), .B(_abc_15497_new_n4591_), .Y(_abc_15497_new_n4592_));
NOR2X1 NOR2X1_671 ( .A(w_mem_inst_w_ctr_reg_5_), .B(w_mem_inst__abc_19396_new_n1585_), .Y(w_mem_inst__abc_19396_new_n1586_));
NOR2X1 NOR2X1_672 ( .A(w_mem_inst__abc_19396_new_n1605_), .B(w_mem_inst__abc_19396_new_n1603_), .Y(w_mem_inst__abc_19396_new_n1606_));
NOR2X1 NOR2X1_673 ( .A(w_mem_inst__abc_19396_new_n1605_), .B(w_mem_inst__abc_19396_new_n1612_), .Y(w_mem_inst__abc_19396_new_n1613_));
NOR2X1 NOR2X1_674 ( .A(w_mem_inst_w_ctr_reg_1_), .B(w_mem_inst_w_ctr_reg_0_), .Y(w_mem_inst__abc_19396_new_n1619_));
NOR2X1 NOR2X1_675 ( .A(w_mem_inst_w_ctr_reg_3_), .B(w_mem_inst_w_ctr_reg_2_), .Y(w_mem_inst__abc_19396_new_n1620_));
NOR2X1 NOR2X1_676 ( .A(w_mem_inst__abc_19396_new_n1593_), .B(w_mem_inst__abc_19396_new_n1603_), .Y(w_mem_inst__abc_19396_new_n1625_));
NOR2X1 NOR2X1_677 ( .A(w_mem_inst__abc_19396_new_n1603_), .B(w_mem_inst__abc_19396_new_n1627_), .Y(w_mem_inst__abc_19396_new_n1628_));
NOR2X1 NOR2X1_678 ( .A(w_mem_inst__abc_19396_new_n1601_), .B(w_mem_inst__abc_19396_new_n1596_), .Y(w_mem_inst__abc_19396_new_n1630_));
NOR2X1 NOR2X1_679 ( .A(w_mem_inst__abc_19396_new_n1596_), .B(w_mem_inst__abc_19396_new_n1627_), .Y(w_mem_inst__abc_19396_new_n1631_));
NOR2X1 NOR2X1_68 ( .A(_abc_15497_new_n698_), .B(_abc_15497_new_n866_), .Y(_abc_15497_new_n867_));
NOR2X1 NOR2X1_680 ( .A(w_mem_inst__abc_19396_new_n4804_), .B(w_mem_inst__abc_19396_new_n4801_), .Y(w_mem_inst__abc_19396_new_n4805_));
NOR2X1 NOR2X1_681 ( .A(w_mem_inst__abc_19396_new_n4808_), .B(w_mem_inst__abc_19396_new_n4809_), .Y(w_mem_inst__0w_ctr_reg_6_0__5_));
NOR2X1 NOR2X1_69 ( .A(_abc_15497_new_n865_), .B(_abc_15497_new_n867_), .Y(_abc_15497_new_n868_));
NOR2X1 NOR2X1_7 ( .A(c_reg_13_), .B(_auto_iopadmap_cc_368_execute_22625_77_), .Y(_abc_15497_new_n712_));
NOR2X1 NOR2X1_70 ( .A(_abc_15497_new_n868_), .B(_abc_15497_new_n864_), .Y(_abc_15497_new_n869_));
NOR2X1 NOR2X1_71 ( .A(_auto_iopadmap_cc_368_execute_22625_91_), .B(c_reg_27_), .Y(_abc_15497_new_n878_));
NOR2X1 NOR2X1_72 ( .A(_abc_15497_new_n878_), .B(_abc_15497_new_n880_), .Y(_abc_15497_new_n881_));
NOR2X1 NOR2X1_73 ( .A(_abc_15497_new_n871__bF_buf3), .B(_abc_15497_new_n872__bF_buf3), .Y(_abc_15497_new_n883_));
NOR2X1 NOR2X1_74 ( .A(_auto_iopadmap_cc_368_execute_22625_92_), .B(c_reg_28_), .Y(_abc_15497_new_n893_));
NOR2X1 NOR2X1_75 ( .A(_abc_15497_new_n893_), .B(_abc_15497_new_n895_), .Y(_abc_15497_new_n896_));
NOR2X1 NOR2X1_76 ( .A(_auto_iopadmap_cc_368_execute_22625_93_), .B(c_reg_29_), .Y(_abc_15497_new_n903_));
NOR2X1 NOR2X1_77 ( .A(_abc_15497_new_n901_), .B(_abc_15497_new_n904_), .Y(_abc_15497_new_n905_));
NOR2X1 NOR2X1_78 ( .A(_abc_15497_new_n903_), .B(_abc_15497_new_n905_), .Y(_abc_15497_new_n906_));
NOR2X1 NOR2X1_79 ( .A(_abc_15497_new_n911_), .B(_abc_15497_new_n912_), .Y(_abc_15497_new_n925_));
NOR2X1 NOR2X1_8 ( .A(_abc_15497_new_n712_), .B(_abc_15497_new_n710_), .Y(_abc_15497_new_n713_));
NOR2X1 NOR2X1_80 ( .A(_abc_15497_new_n937_), .B(_abc_15497_new_n936_), .Y(_abc_15497_new_n938_));
NOR2X1 NOR2X1_81 ( .A(e_reg_3_), .B(_auto_iopadmap_cc_368_execute_22625_3_), .Y(_abc_15497_new_n958_));
NOR2X1 NOR2X1_82 ( .A(_abc_15497_new_n960_), .B(_abc_15497_new_n955_), .Y(_abc_15497_new_n961_));
NOR2X1 NOR2X1_83 ( .A(_abc_15497_new_n968_), .B(_abc_15497_new_n969_), .Y(_abc_15497_new_n970_));
NOR2X1 NOR2X1_84 ( .A(_auto_iopadmap_cc_368_execute_22625_4_), .B(_abc_15497_new_n883__bF_buf10), .Y(_abc_15497_new_n974_));
NOR2X1 NOR2X1_85 ( .A(e_reg_5_), .B(_auto_iopadmap_cc_368_execute_22625_5_), .Y(_abc_15497_new_n977_));
NOR2X1 NOR2X1_86 ( .A(_abc_15497_new_n979_), .B(_abc_15497_new_n976_), .Y(_abc_15497_new_n984_));
NOR2X1 NOR2X1_87 ( .A(_abc_15497_new_n978_), .B(_abc_15497_new_n984_), .Y(_abc_15497_new_n985_));
NOR2X1 NOR2X1_88 ( .A(_abc_15497_new_n986_), .B(_abc_15497_new_n985_), .Y(_abc_15497_new_n992_));
NOR2X1 NOR2X1_89 ( .A(_abc_15497_new_n991_), .B(_abc_15497_new_n992_), .Y(_abc_15497_new_n993_));
NOR2X1 NOR2X1_9 ( .A(c_reg_12_), .B(_auto_iopadmap_cc_368_execute_22625_76_), .Y(_abc_15497_new_n719_));
NOR2X1 NOR2X1_90 ( .A(e_reg_7_), .B(_auto_iopadmap_cc_368_execute_22625_7_), .Y(_abc_15497_new_n994_));
NOR2X1 NOR2X1_91 ( .A(_abc_15497_new_n998_), .B(_abc_15497_new_n993_), .Y(_abc_15497_new_n1001_));
NOR2X1 NOR2X1_92 ( .A(e_reg_8_), .B(_auto_iopadmap_cc_368_execute_22625_8_), .Y(_abc_15497_new_n1005_));
NOR2X1 NOR2X1_93 ( .A(_abc_15497_new_n1006_), .B(_abc_15497_new_n1007_), .Y(_abc_15497_new_n1008_));
NOR2X1 NOR2X1_94 ( .A(_abc_15497_new_n968_), .B(_abc_15497_new_n979_), .Y(_abc_15497_new_n1009_));
NOR2X1 NOR2X1_95 ( .A(_abc_15497_new_n986_), .B(_abc_15497_new_n997_), .Y(_abc_15497_new_n1010_));
NOR2X1 NOR2X1_96 ( .A(_abc_15497_new_n1011_), .B(_abc_15497_new_n969_), .Y(_abc_15497_new_n1012_));
NOR2X1 NOR2X1_97 ( .A(_abc_15497_new_n967_), .B(_abc_15497_new_n979_), .Y(_abc_15497_new_n1014_));
NOR2X1 NOR2X1_98 ( .A(_abc_15497_new_n1016_), .B(_abc_15497_new_n1012_), .Y(_abc_15497_new_n1017_));
NOR2X1 NOR2X1_99 ( .A(_abc_15497_new_n1005_), .B(_abc_15497_new_n1008_), .Y(_abc_15497_new_n1019_));
NOR3X1 NOR3X1_1 ( .A(_abc_15497_new_n2738_), .B(_abc_15497_new_n2768_), .C(_abc_15497_new_n2772_), .Y(_abc_15497_new_n2774_));
NOR3X1 NOR3X1_10 ( .A(_abc_15497_new_n3242_), .B(_abc_15497_new_n3243_), .C(_abc_15497_new_n3245_), .Y(_abc_15497_new_n3261_));
NOR3X1 NOR3X1_11 ( .A(_abc_15497_new_n2944_), .B(_abc_15497_new_n3268_), .C(_abc_15497_new_n3265_), .Y(_abc_15497_new_n3277_));
NOR3X1 NOR3X1_12 ( .A(_abc_15497_new_n3302_), .B(_abc_15497_new_n3303_), .C(_abc_15497_new_n3305_), .Y(_abc_15497_new_n3311_));
NOR3X1 NOR3X1_13 ( .A(_abc_15497_new_n2924__bF_buf1), .B(_abc_15497_new_n3326_), .C(_abc_15497_new_n3323_), .Y(_abc_15497_new_n3339_));
NOR3X1 NOR3X1_14 ( .A(_abc_15497_new_n3361_), .B(_abc_15497_new_n3362_), .C(_abc_15497_new_n3363_), .Y(_abc_15497_new_n3371_));
NOR3X1 NOR3X1_15 ( .A(_abc_15497_new_n3431_), .B(_abc_15497_new_n3432_), .C(_abc_15497_new_n3434_), .Y(_abc_15497_new_n3440_));
NOR3X1 NOR3X1_16 ( .A(_abc_15497_new_n2780__bF_buf0), .B(_abc_15497_new_n3515_), .C(_abc_15497_new_n3512_), .Y(_abc_15497_new_n3525_));
NOR3X1 NOR3X1_17 ( .A(_abc_15497_new_n3559_), .B(_abc_15497_new_n3560_), .C(_abc_15497_new_n3561_), .Y(_abc_15497_new_n3568_));
NOR3X1 NOR3X1_18 ( .A(_abc_15497_new_n2759__bF_buf2), .B(_abc_15497_new_n3581_), .C(_abc_15497_new_n3578_), .Y(_abc_15497_new_n3594_));
NOR3X1 NOR3X1_19 ( .A(_abc_15497_new_n3622_), .B(_abc_15497_new_n3623_), .C(_abc_15497_new_n3625_), .Y(_abc_15497_new_n3631_));
NOR3X1 NOR3X1_2 ( .A(_abc_15497_new_n2792_), .B(_abc_15497_new_n2793_), .C(_abc_15497_new_n2795_), .Y(_abc_15497_new_n2802_));
NOR3X1 NOR3X1_20 ( .A(_abc_15497_new_n2743__bF_buf4), .B(_abc_15497_new_n3646_), .C(_abc_15497_new_n3643_), .Y(_abc_15497_new_n3658_));
NOR3X1 NOR3X1_21 ( .A(_abc_15497_new_n3756_), .B(_abc_15497_new_n3757_), .C(_abc_15497_new_n3758_), .Y(_abc_15497_new_n3759_));
NOR3X1 NOR3X1_22 ( .A(_abc_15497_new_n4406_), .B(_abc_15497_new_n4433_), .C(_abc_15497_new_n4410_), .Y(_abc_15497_new_n4434_));
NOR3X1 NOR3X1_23 ( .A(w_mem_inst__abc_19396_new_n1615_), .B(w_mem_inst__abc_19396_new_n1599_), .C(w_mem_inst__abc_19396_new_n1608_), .Y(w_mem_inst__abc_19396_new_n1616_));
NOR3X1 NOR3X1_24 ( .A(w_mem_inst_w_ctr_reg_3_), .B(w_mem_inst_w_ctr_reg_2_), .C(w_mem_inst__abc_19396_new_n1605_), .Y(w_mem_inst__abc_19396_new_n1637_));
NOR3X1 NOR3X1_25 ( .A(w_mem_inst_w_ctr_reg_0_), .B(w_mem_inst__abc_19396_new_n1592_), .C(w_mem_inst__abc_19396_new_n1612_), .Y(w_mem_inst__abc_19396_new_n1638_));
NOR3X1 NOR3X1_26 ( .A(w_mem_inst__abc_19396_new_n1624_), .B(w_mem_inst__abc_19396_new_n1640_), .C(w_mem_inst__abc_19396_new_n1633_), .Y(w_mem_inst__abc_19396_new_n1641_));
NOR3X1 NOR3X1_27 ( .A(w_mem_inst__abc_19396_new_n1653_), .B(w_mem_inst__abc_19396_new_n1647_), .C(w_mem_inst__abc_19396_new_n1650_), .Y(w_mem_inst__abc_19396_new_n1654_));
NOR3X1 NOR3X1_28 ( .A(w_mem_inst__abc_19396_new_n1658_), .B(w_mem_inst__abc_19396_new_n1665_), .C(w_mem_inst__abc_19396_new_n1661_), .Y(w_mem_inst__abc_19396_new_n1666_));
NOR3X1 NOR3X1_29 ( .A(w_mem_inst__abc_19396_new_n1678_), .B(w_mem_inst__abc_19396_new_n1672_), .C(w_mem_inst__abc_19396_new_n1675_), .Y(w_mem_inst__abc_19396_new_n1679_));
NOR3X1 NOR3X1_3 ( .A(_abc_15497_new_n2827_), .B(_abc_15497_new_n2866_), .C(_abc_15497_new_n2862_), .Y(_abc_15497_new_n2867_));
NOR3X1 NOR3X1_30 ( .A(w_mem_inst__abc_19396_new_n1683_), .B(w_mem_inst__abc_19396_new_n1690_), .C(w_mem_inst__abc_19396_new_n1686_), .Y(w_mem_inst__abc_19396_new_n1691_));
NOR3X1 NOR3X1_31 ( .A(w_mem_inst__abc_19396_new_n1703_), .B(w_mem_inst__abc_19396_new_n1697_), .C(w_mem_inst__abc_19396_new_n1700_), .Y(w_mem_inst__abc_19396_new_n1704_));
NOR3X1 NOR3X1_32 ( .A(w_mem_inst__abc_19396_new_n1708_), .B(w_mem_inst__abc_19396_new_n1715_), .C(w_mem_inst__abc_19396_new_n1711_), .Y(w_mem_inst__abc_19396_new_n1716_));
NOR3X1 NOR3X1_33 ( .A(w_mem_inst__abc_19396_new_n1728_), .B(w_mem_inst__abc_19396_new_n1722_), .C(w_mem_inst__abc_19396_new_n1725_), .Y(w_mem_inst__abc_19396_new_n1729_));
NOR3X1 NOR3X1_34 ( .A(w_mem_inst__abc_19396_new_n1733_), .B(w_mem_inst__abc_19396_new_n1740_), .C(w_mem_inst__abc_19396_new_n1736_), .Y(w_mem_inst__abc_19396_new_n1741_));
NOR3X1 NOR3X1_35 ( .A(w_mem_inst__abc_19396_new_n1753_), .B(w_mem_inst__abc_19396_new_n1747_), .C(w_mem_inst__abc_19396_new_n1750_), .Y(w_mem_inst__abc_19396_new_n1754_));
NOR3X1 NOR3X1_36 ( .A(w_mem_inst__abc_19396_new_n1758_), .B(w_mem_inst__abc_19396_new_n1765_), .C(w_mem_inst__abc_19396_new_n1761_), .Y(w_mem_inst__abc_19396_new_n1766_));
NOR3X1 NOR3X1_37 ( .A(w_mem_inst__abc_19396_new_n1778_), .B(w_mem_inst__abc_19396_new_n1772_), .C(w_mem_inst__abc_19396_new_n1775_), .Y(w_mem_inst__abc_19396_new_n1779_));
NOR3X1 NOR3X1_38 ( .A(w_mem_inst__abc_19396_new_n1783_), .B(w_mem_inst__abc_19396_new_n1790_), .C(w_mem_inst__abc_19396_new_n1786_), .Y(w_mem_inst__abc_19396_new_n1791_));
NOR3X1 NOR3X1_39 ( .A(w_mem_inst__abc_19396_new_n1803_), .B(w_mem_inst__abc_19396_new_n1797_), .C(w_mem_inst__abc_19396_new_n1800_), .Y(w_mem_inst__abc_19396_new_n1804_));
NOR3X1 NOR3X1_4 ( .A(_abc_15497_new_n2885_), .B(_abc_15497_new_n2930_), .C(_abc_15497_new_n2933_), .Y(_abc_15497_new_n2940_));
NOR3X1 NOR3X1_40 ( .A(w_mem_inst__abc_19396_new_n1808_), .B(w_mem_inst__abc_19396_new_n1815_), .C(w_mem_inst__abc_19396_new_n1811_), .Y(w_mem_inst__abc_19396_new_n1816_));
NOR3X1 NOR3X1_41 ( .A(w_mem_inst__abc_19396_new_n1828_), .B(w_mem_inst__abc_19396_new_n1822_), .C(w_mem_inst__abc_19396_new_n1825_), .Y(w_mem_inst__abc_19396_new_n1829_));
NOR3X1 NOR3X1_42 ( .A(w_mem_inst__abc_19396_new_n1833_), .B(w_mem_inst__abc_19396_new_n1840_), .C(w_mem_inst__abc_19396_new_n1836_), .Y(w_mem_inst__abc_19396_new_n1841_));
NOR3X1 NOR3X1_43 ( .A(w_mem_inst__abc_19396_new_n1853_), .B(w_mem_inst__abc_19396_new_n1847_), .C(w_mem_inst__abc_19396_new_n1850_), .Y(w_mem_inst__abc_19396_new_n1854_));
NOR3X1 NOR3X1_44 ( .A(w_mem_inst__abc_19396_new_n1858_), .B(w_mem_inst__abc_19396_new_n1865_), .C(w_mem_inst__abc_19396_new_n1861_), .Y(w_mem_inst__abc_19396_new_n1866_));
NOR3X1 NOR3X1_45 ( .A(w_mem_inst__abc_19396_new_n1878_), .B(w_mem_inst__abc_19396_new_n1872_), .C(w_mem_inst__abc_19396_new_n1875_), .Y(w_mem_inst__abc_19396_new_n1879_));
NOR3X1 NOR3X1_46 ( .A(w_mem_inst__abc_19396_new_n1883_), .B(w_mem_inst__abc_19396_new_n1890_), .C(w_mem_inst__abc_19396_new_n1886_), .Y(w_mem_inst__abc_19396_new_n1891_));
NOR3X1 NOR3X1_47 ( .A(w_mem_inst__abc_19396_new_n1903_), .B(w_mem_inst__abc_19396_new_n1897_), .C(w_mem_inst__abc_19396_new_n1900_), .Y(w_mem_inst__abc_19396_new_n1904_));
NOR3X1 NOR3X1_48 ( .A(w_mem_inst__abc_19396_new_n1908_), .B(w_mem_inst__abc_19396_new_n1915_), .C(w_mem_inst__abc_19396_new_n1911_), .Y(w_mem_inst__abc_19396_new_n1916_));
NOR3X1 NOR3X1_49 ( .A(w_mem_inst__abc_19396_new_n1928_), .B(w_mem_inst__abc_19396_new_n1922_), .C(w_mem_inst__abc_19396_new_n1925_), .Y(w_mem_inst__abc_19396_new_n1929_));
NOR3X1 NOR3X1_5 ( .A(_abc_15497_new_n3018_), .B(_abc_15497_new_n3019_), .C(_abc_15497_new_n3021_), .Y(_abc_15497_new_n3028_));
NOR3X1 NOR3X1_50 ( .A(w_mem_inst__abc_19396_new_n1933_), .B(w_mem_inst__abc_19396_new_n1940_), .C(w_mem_inst__abc_19396_new_n1936_), .Y(w_mem_inst__abc_19396_new_n1941_));
NOR3X1 NOR3X1_51 ( .A(w_mem_inst__abc_19396_new_n1953_), .B(w_mem_inst__abc_19396_new_n1947_), .C(w_mem_inst__abc_19396_new_n1950_), .Y(w_mem_inst__abc_19396_new_n1954_));
NOR3X1 NOR3X1_52 ( .A(w_mem_inst__abc_19396_new_n1958_), .B(w_mem_inst__abc_19396_new_n1965_), .C(w_mem_inst__abc_19396_new_n1961_), .Y(w_mem_inst__abc_19396_new_n1966_));
NOR3X1 NOR3X1_53 ( .A(w_mem_inst__abc_19396_new_n1978_), .B(w_mem_inst__abc_19396_new_n1972_), .C(w_mem_inst__abc_19396_new_n1975_), .Y(w_mem_inst__abc_19396_new_n1979_));
NOR3X1 NOR3X1_54 ( .A(w_mem_inst__abc_19396_new_n1983_), .B(w_mem_inst__abc_19396_new_n1990_), .C(w_mem_inst__abc_19396_new_n1986_), .Y(w_mem_inst__abc_19396_new_n1991_));
NOR3X1 NOR3X1_55 ( .A(w_mem_inst__abc_19396_new_n2003_), .B(w_mem_inst__abc_19396_new_n1997_), .C(w_mem_inst__abc_19396_new_n2000_), .Y(w_mem_inst__abc_19396_new_n2004_));
NOR3X1 NOR3X1_56 ( .A(w_mem_inst__abc_19396_new_n2008_), .B(w_mem_inst__abc_19396_new_n2015_), .C(w_mem_inst__abc_19396_new_n2011_), .Y(w_mem_inst__abc_19396_new_n2016_));
NOR3X1 NOR3X1_57 ( .A(w_mem_inst__abc_19396_new_n2028_), .B(w_mem_inst__abc_19396_new_n2022_), .C(w_mem_inst__abc_19396_new_n2025_), .Y(w_mem_inst__abc_19396_new_n2029_));
NOR3X1 NOR3X1_58 ( .A(w_mem_inst__abc_19396_new_n2033_), .B(w_mem_inst__abc_19396_new_n2040_), .C(w_mem_inst__abc_19396_new_n2036_), .Y(w_mem_inst__abc_19396_new_n2041_));
NOR3X1 NOR3X1_59 ( .A(w_mem_inst__abc_19396_new_n2053_), .B(w_mem_inst__abc_19396_new_n2047_), .C(w_mem_inst__abc_19396_new_n2050_), .Y(w_mem_inst__abc_19396_new_n2054_));
NOR3X1 NOR3X1_6 ( .A(_abc_15497_new_n2944_), .B(_abc_15497_new_n3040_), .C(_abc_15497_new_n3035_), .Y(_abc_15497_new_n3050_));
NOR3X1 NOR3X1_60 ( .A(w_mem_inst__abc_19396_new_n2058_), .B(w_mem_inst__abc_19396_new_n2065_), .C(w_mem_inst__abc_19396_new_n2061_), .Y(w_mem_inst__abc_19396_new_n2066_));
NOR3X1 NOR3X1_61 ( .A(w_mem_inst__abc_19396_new_n2078_), .B(w_mem_inst__abc_19396_new_n2072_), .C(w_mem_inst__abc_19396_new_n2075_), .Y(w_mem_inst__abc_19396_new_n2079_));
NOR3X1 NOR3X1_62 ( .A(w_mem_inst__abc_19396_new_n2083_), .B(w_mem_inst__abc_19396_new_n2090_), .C(w_mem_inst__abc_19396_new_n2086_), .Y(w_mem_inst__abc_19396_new_n2091_));
NOR3X1 NOR3X1_63 ( .A(w_mem_inst__abc_19396_new_n2103_), .B(w_mem_inst__abc_19396_new_n2097_), .C(w_mem_inst__abc_19396_new_n2100_), .Y(w_mem_inst__abc_19396_new_n2104_));
NOR3X1 NOR3X1_64 ( .A(w_mem_inst__abc_19396_new_n2108_), .B(w_mem_inst__abc_19396_new_n2115_), .C(w_mem_inst__abc_19396_new_n2111_), .Y(w_mem_inst__abc_19396_new_n2116_));
NOR3X1 NOR3X1_65 ( .A(w_mem_inst__abc_19396_new_n2128_), .B(w_mem_inst__abc_19396_new_n2122_), .C(w_mem_inst__abc_19396_new_n2125_), .Y(w_mem_inst__abc_19396_new_n2129_));
NOR3X1 NOR3X1_66 ( .A(w_mem_inst__abc_19396_new_n2133_), .B(w_mem_inst__abc_19396_new_n2140_), .C(w_mem_inst__abc_19396_new_n2136_), .Y(w_mem_inst__abc_19396_new_n2141_));
NOR3X1 NOR3X1_67 ( .A(w_mem_inst__abc_19396_new_n2153_), .B(w_mem_inst__abc_19396_new_n2147_), .C(w_mem_inst__abc_19396_new_n2150_), .Y(w_mem_inst__abc_19396_new_n2154_));
NOR3X1 NOR3X1_68 ( .A(w_mem_inst__abc_19396_new_n2158_), .B(w_mem_inst__abc_19396_new_n2165_), .C(w_mem_inst__abc_19396_new_n2161_), .Y(w_mem_inst__abc_19396_new_n2166_));
NOR3X1 NOR3X1_69 ( .A(w_mem_inst__abc_19396_new_n2178_), .B(w_mem_inst__abc_19396_new_n2172_), .C(w_mem_inst__abc_19396_new_n2175_), .Y(w_mem_inst__abc_19396_new_n2179_));
NOR3X1 NOR3X1_7 ( .A(_abc_15497_new_n3076_), .B(_abc_15497_new_n3077_), .C(_abc_15497_new_n3079_), .Y(_abc_15497_new_n3086_));
NOR3X1 NOR3X1_70 ( .A(w_mem_inst__abc_19396_new_n2183_), .B(w_mem_inst__abc_19396_new_n2190_), .C(w_mem_inst__abc_19396_new_n2186_), .Y(w_mem_inst__abc_19396_new_n2191_));
NOR3X1 NOR3X1_71 ( .A(w_mem_inst__abc_19396_new_n2203_), .B(w_mem_inst__abc_19396_new_n2197_), .C(w_mem_inst__abc_19396_new_n2200_), .Y(w_mem_inst__abc_19396_new_n2204_));
NOR3X1 NOR3X1_72 ( .A(w_mem_inst__abc_19396_new_n2208_), .B(w_mem_inst__abc_19396_new_n2215_), .C(w_mem_inst__abc_19396_new_n2211_), .Y(w_mem_inst__abc_19396_new_n2216_));
NOR3X1 NOR3X1_73 ( .A(w_mem_inst__abc_19396_new_n2228_), .B(w_mem_inst__abc_19396_new_n2222_), .C(w_mem_inst__abc_19396_new_n2225_), .Y(w_mem_inst__abc_19396_new_n2229_));
NOR3X1 NOR3X1_74 ( .A(w_mem_inst__abc_19396_new_n2233_), .B(w_mem_inst__abc_19396_new_n2240_), .C(w_mem_inst__abc_19396_new_n2236_), .Y(w_mem_inst__abc_19396_new_n2241_));
NOR3X1 NOR3X1_75 ( .A(w_mem_inst__abc_19396_new_n2253_), .B(w_mem_inst__abc_19396_new_n2247_), .C(w_mem_inst__abc_19396_new_n2250_), .Y(w_mem_inst__abc_19396_new_n2254_));
NOR3X1 NOR3X1_76 ( .A(w_mem_inst__abc_19396_new_n2258_), .B(w_mem_inst__abc_19396_new_n2265_), .C(w_mem_inst__abc_19396_new_n2261_), .Y(w_mem_inst__abc_19396_new_n2266_));
NOR3X1 NOR3X1_77 ( .A(w_mem_inst__abc_19396_new_n2278_), .B(w_mem_inst__abc_19396_new_n2272_), .C(w_mem_inst__abc_19396_new_n2275_), .Y(w_mem_inst__abc_19396_new_n2279_));
NOR3X1 NOR3X1_78 ( .A(w_mem_inst__abc_19396_new_n2283_), .B(w_mem_inst__abc_19396_new_n2290_), .C(w_mem_inst__abc_19396_new_n2286_), .Y(w_mem_inst__abc_19396_new_n2291_));
NOR3X1 NOR3X1_79 ( .A(w_mem_inst__abc_19396_new_n2303_), .B(w_mem_inst__abc_19396_new_n2297_), .C(w_mem_inst__abc_19396_new_n2300_), .Y(w_mem_inst__abc_19396_new_n2304_));
NOR3X1 NOR3X1_8 ( .A(_abc_15497_new_n2739_), .B(_abc_15497_new_n3098_), .C(_abc_15497_new_n3093_), .Y(_abc_15497_new_n3106_));
NOR3X1 NOR3X1_80 ( .A(w_mem_inst__abc_19396_new_n2308_), .B(w_mem_inst__abc_19396_new_n2315_), .C(w_mem_inst__abc_19396_new_n2311_), .Y(w_mem_inst__abc_19396_new_n2316_));
NOR3X1 NOR3X1_81 ( .A(w_mem_inst__abc_19396_new_n2328_), .B(w_mem_inst__abc_19396_new_n2322_), .C(w_mem_inst__abc_19396_new_n2325_), .Y(w_mem_inst__abc_19396_new_n2329_));
NOR3X1 NOR3X1_82 ( .A(w_mem_inst__abc_19396_new_n2333_), .B(w_mem_inst__abc_19396_new_n2340_), .C(w_mem_inst__abc_19396_new_n2336_), .Y(w_mem_inst__abc_19396_new_n2341_));
NOR3X1 NOR3X1_83 ( .A(w_mem_inst__abc_19396_new_n2353_), .B(w_mem_inst__abc_19396_new_n2347_), .C(w_mem_inst__abc_19396_new_n2350_), .Y(w_mem_inst__abc_19396_new_n2354_));
NOR3X1 NOR3X1_84 ( .A(w_mem_inst__abc_19396_new_n2358_), .B(w_mem_inst__abc_19396_new_n2365_), .C(w_mem_inst__abc_19396_new_n2361_), .Y(w_mem_inst__abc_19396_new_n2366_));
NOR3X1 NOR3X1_85 ( .A(w_mem_inst__abc_19396_new_n2378_), .B(w_mem_inst__abc_19396_new_n2372_), .C(w_mem_inst__abc_19396_new_n2375_), .Y(w_mem_inst__abc_19396_new_n2379_));
NOR3X1 NOR3X1_86 ( .A(w_mem_inst__abc_19396_new_n2383_), .B(w_mem_inst__abc_19396_new_n2390_), .C(w_mem_inst__abc_19396_new_n2386_), .Y(w_mem_inst__abc_19396_new_n2391_));
NOR3X1 NOR3X1_87 ( .A(w_mem_inst__abc_19396_new_n2403_), .B(w_mem_inst__abc_19396_new_n2397_), .C(w_mem_inst__abc_19396_new_n2400_), .Y(w_mem_inst__abc_19396_new_n2404_));
NOR3X1 NOR3X1_88 ( .A(w_mem_inst__abc_19396_new_n2408_), .B(w_mem_inst__abc_19396_new_n2415_), .C(w_mem_inst__abc_19396_new_n2411_), .Y(w_mem_inst__abc_19396_new_n2416_));
NOR3X1 NOR3X1_9 ( .A(_abc_15497_new_n3131_), .B(_abc_15497_new_n3132_), .C(_abc_15497_new_n3134_), .Y(_abc_15497_new_n3141_));
OAI21X1 OAI21X1_1 ( .A(_abc_15497_new_n707_), .B(_abc_15497_new_n714_), .C(_abc_15497_new_n715_), .Y(_abc_15497_new_n716_));
OAI21X1 OAI21X1_10 ( .A(_abc_15497_new_n698_), .B(_abc_15497_new_n866_), .C(_abc_15497_new_n874_), .Y(_abc_15497_new_n877_));
OAI21X1 OAI21X1_100 ( .A(_abc_15497_new_n1270_), .B(_abc_15497_new_n1272_), .C(_abc_15497_new_n1282_), .Y(_abc_15497_new_n1283_));
OAI21X1 OAI21X1_1000 ( .A(w_mem_inst__abc_19396_new_n1873_), .B(w_mem_inst__abc_19396_new_n1604__bF_buf4), .C(w_mem_inst__abc_19396_new_n1874_), .Y(w_mem_inst__abc_19396_new_n1875_));
OAI21X1 OAI21X1_1001 ( .A(w_mem_inst__abc_19396_new_n1876_), .B(w_mem_inst__abc_19396_new_n1611__bF_buf4), .C(w_mem_inst__abc_19396_new_n1877_), .Y(w_mem_inst__abc_19396_new_n1878_));
OAI21X1 OAI21X1_1002 ( .A(w_mem_inst__abc_19396_new_n1896_), .B(w_mem_inst__abc_19396_new_n1598__bF_buf3), .C(w_mem_inst__abc_19396_new_n1586__bF_buf2), .Y(w_mem_inst__abc_19396_new_n1897_));
OAI21X1 OAI21X1_1003 ( .A(w_mem_inst__abc_19396_new_n1898_), .B(w_mem_inst__abc_19396_new_n1604__bF_buf3), .C(w_mem_inst__abc_19396_new_n1899_), .Y(w_mem_inst__abc_19396_new_n1900_));
OAI21X1 OAI21X1_1004 ( .A(w_mem_inst__abc_19396_new_n1901_), .B(w_mem_inst__abc_19396_new_n1611__bF_buf3), .C(w_mem_inst__abc_19396_new_n1902_), .Y(w_mem_inst__abc_19396_new_n1903_));
OAI21X1 OAI21X1_1005 ( .A(w_mem_inst__abc_19396_new_n1921_), .B(w_mem_inst__abc_19396_new_n1598__bF_buf2), .C(w_mem_inst__abc_19396_new_n1586__bF_buf1), .Y(w_mem_inst__abc_19396_new_n1922_));
OAI21X1 OAI21X1_1006 ( .A(w_mem_inst__abc_19396_new_n1923_), .B(w_mem_inst__abc_19396_new_n1604__bF_buf2), .C(w_mem_inst__abc_19396_new_n1924_), .Y(w_mem_inst__abc_19396_new_n1925_));
OAI21X1 OAI21X1_1007 ( .A(w_mem_inst__abc_19396_new_n1926_), .B(w_mem_inst__abc_19396_new_n1611__bF_buf2), .C(w_mem_inst__abc_19396_new_n1927_), .Y(w_mem_inst__abc_19396_new_n1928_));
OAI21X1 OAI21X1_1008 ( .A(w_mem_inst__abc_19396_new_n1946_), .B(w_mem_inst__abc_19396_new_n1598__bF_buf1), .C(w_mem_inst__abc_19396_new_n1586__bF_buf0), .Y(w_mem_inst__abc_19396_new_n1947_));
OAI21X1 OAI21X1_1009 ( .A(w_mem_inst__abc_19396_new_n1948_), .B(w_mem_inst__abc_19396_new_n1604__bF_buf1), .C(w_mem_inst__abc_19396_new_n1949_), .Y(w_mem_inst__abc_19396_new_n1950_));
OAI21X1 OAI21X1_101 ( .A(_abc_15497_new_n1281_), .B(_abc_15497_new_n1285_), .C(digest_update_bF_buf6), .Y(_abc_15497_new_n1287_));
OAI21X1 OAI21X1_1010 ( .A(w_mem_inst__abc_19396_new_n1951_), .B(w_mem_inst__abc_19396_new_n1611__bF_buf1), .C(w_mem_inst__abc_19396_new_n1952_), .Y(w_mem_inst__abc_19396_new_n1953_));
OAI21X1 OAI21X1_1011 ( .A(w_mem_inst__abc_19396_new_n1971_), .B(w_mem_inst__abc_19396_new_n1598__bF_buf0), .C(w_mem_inst__abc_19396_new_n1586__bF_buf4), .Y(w_mem_inst__abc_19396_new_n1972_));
OAI21X1 OAI21X1_1012 ( .A(w_mem_inst__abc_19396_new_n1973_), .B(w_mem_inst__abc_19396_new_n1604__bF_buf0), .C(w_mem_inst__abc_19396_new_n1974_), .Y(w_mem_inst__abc_19396_new_n1975_));
OAI21X1 OAI21X1_1013 ( .A(w_mem_inst__abc_19396_new_n1976_), .B(w_mem_inst__abc_19396_new_n1611__bF_buf0), .C(w_mem_inst__abc_19396_new_n1977_), .Y(w_mem_inst__abc_19396_new_n1978_));
OAI21X1 OAI21X1_1014 ( .A(w_mem_inst__abc_19396_new_n1996_), .B(w_mem_inst__abc_19396_new_n1598__bF_buf4), .C(w_mem_inst__abc_19396_new_n1586__bF_buf3), .Y(w_mem_inst__abc_19396_new_n1997_));
OAI21X1 OAI21X1_1015 ( .A(w_mem_inst__abc_19396_new_n1998_), .B(w_mem_inst__abc_19396_new_n1604__bF_buf4), .C(w_mem_inst__abc_19396_new_n1999_), .Y(w_mem_inst__abc_19396_new_n2000_));
OAI21X1 OAI21X1_1016 ( .A(w_mem_inst__abc_19396_new_n2001_), .B(w_mem_inst__abc_19396_new_n1611__bF_buf4), .C(w_mem_inst__abc_19396_new_n2002_), .Y(w_mem_inst__abc_19396_new_n2003_));
OAI21X1 OAI21X1_1017 ( .A(w_mem_inst__abc_19396_new_n2021_), .B(w_mem_inst__abc_19396_new_n1598__bF_buf3), .C(w_mem_inst__abc_19396_new_n1586__bF_buf2), .Y(w_mem_inst__abc_19396_new_n2022_));
OAI21X1 OAI21X1_1018 ( .A(w_mem_inst__abc_19396_new_n2023_), .B(w_mem_inst__abc_19396_new_n1604__bF_buf3), .C(w_mem_inst__abc_19396_new_n2024_), .Y(w_mem_inst__abc_19396_new_n2025_));
OAI21X1 OAI21X1_1019 ( .A(w_mem_inst__abc_19396_new_n2026_), .B(w_mem_inst__abc_19396_new_n1611__bF_buf3), .C(w_mem_inst__abc_19396_new_n2027_), .Y(w_mem_inst__abc_19396_new_n2028_));
OAI21X1 OAI21X1_102 ( .A(_auto_iopadmap_cc_368_execute_22625_30_), .B(_abc_15497_new_n883__bF_buf10), .C(_abc_15497_new_n870__bF_buf11), .Y(_abc_15497_new_n1288_));
OAI21X1 OAI21X1_1020 ( .A(w_mem_inst__abc_19396_new_n2046_), .B(w_mem_inst__abc_19396_new_n1598__bF_buf2), .C(w_mem_inst__abc_19396_new_n1586__bF_buf1), .Y(w_mem_inst__abc_19396_new_n2047_));
OAI21X1 OAI21X1_1021 ( .A(w_mem_inst__abc_19396_new_n2048_), .B(w_mem_inst__abc_19396_new_n1604__bF_buf2), .C(w_mem_inst__abc_19396_new_n2049_), .Y(w_mem_inst__abc_19396_new_n2050_));
OAI21X1 OAI21X1_1022 ( .A(w_mem_inst__abc_19396_new_n2051_), .B(w_mem_inst__abc_19396_new_n1611__bF_buf2), .C(w_mem_inst__abc_19396_new_n2052_), .Y(w_mem_inst__abc_19396_new_n2053_));
OAI21X1 OAI21X1_1023 ( .A(w_mem_inst__abc_19396_new_n2071_), .B(w_mem_inst__abc_19396_new_n1598__bF_buf1), .C(w_mem_inst__abc_19396_new_n1586__bF_buf0), .Y(w_mem_inst__abc_19396_new_n2072_));
OAI21X1 OAI21X1_1024 ( .A(w_mem_inst__abc_19396_new_n2073_), .B(w_mem_inst__abc_19396_new_n1604__bF_buf1), .C(w_mem_inst__abc_19396_new_n2074_), .Y(w_mem_inst__abc_19396_new_n2075_));
OAI21X1 OAI21X1_1025 ( .A(w_mem_inst__abc_19396_new_n2076_), .B(w_mem_inst__abc_19396_new_n1611__bF_buf1), .C(w_mem_inst__abc_19396_new_n2077_), .Y(w_mem_inst__abc_19396_new_n2078_));
OAI21X1 OAI21X1_1026 ( .A(w_mem_inst__abc_19396_new_n2096_), .B(w_mem_inst__abc_19396_new_n1598__bF_buf0), .C(w_mem_inst__abc_19396_new_n1586__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2097_));
OAI21X1 OAI21X1_1027 ( .A(w_mem_inst__abc_19396_new_n2098_), .B(w_mem_inst__abc_19396_new_n1604__bF_buf0), .C(w_mem_inst__abc_19396_new_n2099_), .Y(w_mem_inst__abc_19396_new_n2100_));
OAI21X1 OAI21X1_1028 ( .A(w_mem_inst__abc_19396_new_n2101_), .B(w_mem_inst__abc_19396_new_n1611__bF_buf0), .C(w_mem_inst__abc_19396_new_n2102_), .Y(w_mem_inst__abc_19396_new_n2103_));
OAI21X1 OAI21X1_1029 ( .A(w_mem_inst__abc_19396_new_n2121_), .B(w_mem_inst__abc_19396_new_n1598__bF_buf4), .C(w_mem_inst__abc_19396_new_n1586__bF_buf3), .Y(w_mem_inst__abc_19396_new_n2122_));
OAI21X1 OAI21X1_103 ( .A(_abc_15497_new_n1286_), .B(_abc_15497_new_n1287_), .C(_abc_15497_new_n1288_), .Y(_0H4_reg_31_0__30_));
OAI21X1 OAI21X1_1030 ( .A(w_mem_inst__abc_19396_new_n2123_), .B(w_mem_inst__abc_19396_new_n1604__bF_buf4), .C(w_mem_inst__abc_19396_new_n2124_), .Y(w_mem_inst__abc_19396_new_n2125_));
OAI21X1 OAI21X1_1031 ( .A(w_mem_inst__abc_19396_new_n2126_), .B(w_mem_inst__abc_19396_new_n1611__bF_buf4), .C(w_mem_inst__abc_19396_new_n2127_), .Y(w_mem_inst__abc_19396_new_n2128_));
OAI21X1 OAI21X1_1032 ( .A(w_mem_inst__abc_19396_new_n2146_), .B(w_mem_inst__abc_19396_new_n1598__bF_buf3), .C(w_mem_inst__abc_19396_new_n1586__bF_buf2), .Y(w_mem_inst__abc_19396_new_n2147_));
OAI21X1 OAI21X1_1033 ( .A(w_mem_inst__abc_19396_new_n2148_), .B(w_mem_inst__abc_19396_new_n1604__bF_buf3), .C(w_mem_inst__abc_19396_new_n2149_), .Y(w_mem_inst__abc_19396_new_n2150_));
OAI21X1 OAI21X1_1034 ( .A(w_mem_inst__abc_19396_new_n2151_), .B(w_mem_inst__abc_19396_new_n1611__bF_buf3), .C(w_mem_inst__abc_19396_new_n2152_), .Y(w_mem_inst__abc_19396_new_n2153_));
OAI21X1 OAI21X1_1035 ( .A(w_mem_inst__abc_19396_new_n2171_), .B(w_mem_inst__abc_19396_new_n1598__bF_buf2), .C(w_mem_inst__abc_19396_new_n1586__bF_buf1), .Y(w_mem_inst__abc_19396_new_n2172_));
OAI21X1 OAI21X1_1036 ( .A(w_mem_inst__abc_19396_new_n2173_), .B(w_mem_inst__abc_19396_new_n1604__bF_buf2), .C(w_mem_inst__abc_19396_new_n2174_), .Y(w_mem_inst__abc_19396_new_n2175_));
OAI21X1 OAI21X1_1037 ( .A(w_mem_inst__abc_19396_new_n2176_), .B(w_mem_inst__abc_19396_new_n1611__bF_buf2), .C(w_mem_inst__abc_19396_new_n2177_), .Y(w_mem_inst__abc_19396_new_n2178_));
OAI21X1 OAI21X1_1038 ( .A(w_mem_inst__abc_19396_new_n2196_), .B(w_mem_inst__abc_19396_new_n1598__bF_buf1), .C(w_mem_inst__abc_19396_new_n1586__bF_buf0), .Y(w_mem_inst__abc_19396_new_n2197_));
OAI21X1 OAI21X1_1039 ( .A(w_mem_inst__abc_19396_new_n2198_), .B(w_mem_inst__abc_19396_new_n1604__bF_buf1), .C(w_mem_inst__abc_19396_new_n2199_), .Y(w_mem_inst__abc_19396_new_n2200_));
OAI21X1 OAI21X1_104 ( .A(_abc_15497_new_n1281_), .B(_abc_15497_new_n1285_), .C(_abc_15497_new_n1290_), .Y(_abc_15497_new_n1291_));
OAI21X1 OAI21X1_1040 ( .A(w_mem_inst__abc_19396_new_n2201_), .B(w_mem_inst__abc_19396_new_n1611__bF_buf1), .C(w_mem_inst__abc_19396_new_n2202_), .Y(w_mem_inst__abc_19396_new_n2203_));
OAI21X1 OAI21X1_1041 ( .A(w_mem_inst__abc_19396_new_n2221_), .B(w_mem_inst__abc_19396_new_n1598__bF_buf0), .C(w_mem_inst__abc_19396_new_n1586__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2222_));
OAI21X1 OAI21X1_1042 ( .A(w_mem_inst__abc_19396_new_n2223_), .B(w_mem_inst__abc_19396_new_n1604__bF_buf0), .C(w_mem_inst__abc_19396_new_n2224_), .Y(w_mem_inst__abc_19396_new_n2225_));
OAI21X1 OAI21X1_1043 ( .A(w_mem_inst__abc_19396_new_n2226_), .B(w_mem_inst__abc_19396_new_n1611__bF_buf0), .C(w_mem_inst__abc_19396_new_n2227_), .Y(w_mem_inst__abc_19396_new_n2228_));
OAI21X1 OAI21X1_1044 ( .A(w_mem_inst__abc_19396_new_n2246_), .B(w_mem_inst__abc_19396_new_n1598__bF_buf4), .C(w_mem_inst__abc_19396_new_n1586__bF_buf3), .Y(w_mem_inst__abc_19396_new_n2247_));
OAI21X1 OAI21X1_1045 ( .A(w_mem_inst__abc_19396_new_n2248_), .B(w_mem_inst__abc_19396_new_n1604__bF_buf4), .C(w_mem_inst__abc_19396_new_n2249_), .Y(w_mem_inst__abc_19396_new_n2250_));
OAI21X1 OAI21X1_1046 ( .A(w_mem_inst__abc_19396_new_n2251_), .B(w_mem_inst__abc_19396_new_n1611__bF_buf4), .C(w_mem_inst__abc_19396_new_n2252_), .Y(w_mem_inst__abc_19396_new_n2253_));
OAI21X1 OAI21X1_1047 ( .A(w_mem_inst__abc_19396_new_n2271_), .B(w_mem_inst__abc_19396_new_n1598__bF_buf3), .C(w_mem_inst__abc_19396_new_n1586__bF_buf2), .Y(w_mem_inst__abc_19396_new_n2272_));
OAI21X1 OAI21X1_1048 ( .A(w_mem_inst__abc_19396_new_n2273_), .B(w_mem_inst__abc_19396_new_n1604__bF_buf3), .C(w_mem_inst__abc_19396_new_n2274_), .Y(w_mem_inst__abc_19396_new_n2275_));
OAI21X1 OAI21X1_1049 ( .A(w_mem_inst__abc_19396_new_n2276_), .B(w_mem_inst__abc_19396_new_n1611__bF_buf3), .C(w_mem_inst__abc_19396_new_n2277_), .Y(w_mem_inst__abc_19396_new_n2278_));
OAI21X1 OAI21X1_105 ( .A(_abc_15497_new_n1293_), .B(_abc_15497_new_n1294_), .C(digest_update_bF_buf5), .Y(_abc_15497_new_n1295_));
OAI21X1 OAI21X1_1050 ( .A(w_mem_inst__abc_19396_new_n2296_), .B(w_mem_inst__abc_19396_new_n1598__bF_buf2), .C(w_mem_inst__abc_19396_new_n1586__bF_buf1), .Y(w_mem_inst__abc_19396_new_n2297_));
OAI21X1 OAI21X1_1051 ( .A(w_mem_inst__abc_19396_new_n2298_), .B(w_mem_inst__abc_19396_new_n1604__bF_buf2), .C(w_mem_inst__abc_19396_new_n2299_), .Y(w_mem_inst__abc_19396_new_n2300_));
OAI21X1 OAI21X1_1052 ( .A(w_mem_inst__abc_19396_new_n2301_), .B(w_mem_inst__abc_19396_new_n1611__bF_buf2), .C(w_mem_inst__abc_19396_new_n2302_), .Y(w_mem_inst__abc_19396_new_n2303_));
OAI21X1 OAI21X1_1053 ( .A(w_mem_inst__abc_19396_new_n2321_), .B(w_mem_inst__abc_19396_new_n1598__bF_buf1), .C(w_mem_inst__abc_19396_new_n1586__bF_buf0), .Y(w_mem_inst__abc_19396_new_n2322_));
OAI21X1 OAI21X1_1054 ( .A(w_mem_inst__abc_19396_new_n2323_), .B(w_mem_inst__abc_19396_new_n1604__bF_buf1), .C(w_mem_inst__abc_19396_new_n2324_), .Y(w_mem_inst__abc_19396_new_n2325_));
OAI21X1 OAI21X1_1055 ( .A(w_mem_inst__abc_19396_new_n2326_), .B(w_mem_inst__abc_19396_new_n1611__bF_buf1), .C(w_mem_inst__abc_19396_new_n2327_), .Y(w_mem_inst__abc_19396_new_n2328_));
OAI21X1 OAI21X1_1056 ( .A(w_mem_inst__abc_19396_new_n2346_), .B(w_mem_inst__abc_19396_new_n1598__bF_buf0), .C(w_mem_inst__abc_19396_new_n1586__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2347_));
OAI21X1 OAI21X1_1057 ( .A(w_mem_inst__abc_19396_new_n2348_), .B(w_mem_inst__abc_19396_new_n1604__bF_buf0), .C(w_mem_inst__abc_19396_new_n2349_), .Y(w_mem_inst__abc_19396_new_n2350_));
OAI21X1 OAI21X1_1058 ( .A(w_mem_inst__abc_19396_new_n2351_), .B(w_mem_inst__abc_19396_new_n1611__bF_buf0), .C(w_mem_inst__abc_19396_new_n2352_), .Y(w_mem_inst__abc_19396_new_n2353_));
OAI21X1 OAI21X1_1059 ( .A(w_mem_inst__abc_19396_new_n2371_), .B(w_mem_inst__abc_19396_new_n1598__bF_buf4), .C(w_mem_inst__abc_19396_new_n1586__bF_buf3), .Y(w_mem_inst__abc_19396_new_n2372_));
OAI21X1 OAI21X1_106 ( .A(_auto_iopadmap_cc_368_execute_22625_31_), .B(_abc_15497_new_n883__bF_buf9), .C(_abc_15497_new_n870__bF_buf10), .Y(_abc_15497_new_n1296_));
OAI21X1 OAI21X1_1060 ( .A(w_mem_inst__abc_19396_new_n2373_), .B(w_mem_inst__abc_19396_new_n1604__bF_buf4), .C(w_mem_inst__abc_19396_new_n2374_), .Y(w_mem_inst__abc_19396_new_n2375_));
OAI21X1 OAI21X1_1061 ( .A(w_mem_inst__abc_19396_new_n2376_), .B(w_mem_inst__abc_19396_new_n1611__bF_buf4), .C(w_mem_inst__abc_19396_new_n2377_), .Y(w_mem_inst__abc_19396_new_n2378_));
OAI21X1 OAI21X1_1062 ( .A(w_mem_inst__abc_19396_new_n2396_), .B(w_mem_inst__abc_19396_new_n1598__bF_buf3), .C(w_mem_inst__abc_19396_new_n1586__bF_buf2), .Y(w_mem_inst__abc_19396_new_n2397_));
OAI21X1 OAI21X1_1063 ( .A(w_mem_inst__abc_19396_new_n2398_), .B(w_mem_inst__abc_19396_new_n1604__bF_buf3), .C(w_mem_inst__abc_19396_new_n2399_), .Y(w_mem_inst__abc_19396_new_n2400_));
OAI21X1 OAI21X1_1064 ( .A(w_mem_inst__abc_19396_new_n2401_), .B(w_mem_inst__abc_19396_new_n1611__bF_buf3), .C(w_mem_inst__abc_19396_new_n2402_), .Y(w_mem_inst__abc_19396_new_n2403_));
OAI21X1 OAI21X1_1065 ( .A(w_mem_inst__abc_19396_new_n2419_), .B(w_mem_inst__abc_19396_new_n1586__bF_buf1), .C(w_mem_inst__abc_19396_new_n2420__bF_buf60), .Y(w_mem_inst__abc_19396_new_n2421_));
OAI21X1 OAI21X1_1066 ( .A(w_mem_inst_w_ctr_reg_5_), .B(w_mem_inst__abc_19396_new_n1585_), .C(round_ctr_inc_bF_buf1), .Y(w_mem_inst__abc_19396_new_n2422_));
OAI21X1 OAI21X1_1067 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf59), .B(w_mem_inst__abc_19396_new_n2423_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf96), .Y(w_mem_inst__abc_19396_new_n2424_));
OAI21X1 OAI21X1_1068 ( .A(w_mem_inst_w_mem_14__0_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf95), .C(w_mem_inst__abc_19396_new_n2424_), .Y(w_mem_inst__abc_19396_new_n2425_));
OAI21X1 OAI21X1_1069 ( .A(w_mem_inst__abc_19396_new_n2418_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf60), .C(w_mem_inst__abc_19396_new_n2425_), .Y(w_mem_inst__0w_mem_13__31_0__0_));
OAI21X1 OAI21X1_107 ( .A(_auto_iopadmap_cc_368_execute_22625_32_), .B(d_reg_0_), .C(digest_update_bF_buf4), .Y(_abc_15497_new_n1301_));
OAI21X1 OAI21X1_1070 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf58), .B(w_mem_inst__abc_19396_new_n2428_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf94), .Y(w_mem_inst__abc_19396_new_n2429_));
OAI21X1 OAI21X1_1071 ( .A(w_mem_inst_w_mem_14__1_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf93), .C(w_mem_inst__abc_19396_new_n2429_), .Y(w_mem_inst__abc_19396_new_n2430_));
OAI21X1 OAI21X1_1072 ( .A(w_mem_inst__abc_19396_new_n2427_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf59), .C(w_mem_inst__abc_19396_new_n2430_), .Y(w_mem_inst__0w_mem_13__31_0__1_));
OAI21X1 OAI21X1_1073 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf57), .B(w_mem_inst__abc_19396_new_n2433_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf92), .Y(w_mem_inst__abc_19396_new_n2434_));
OAI21X1 OAI21X1_1074 ( .A(w_mem_inst_w_mem_14__2_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf91), .C(w_mem_inst__abc_19396_new_n2434_), .Y(w_mem_inst__abc_19396_new_n2435_));
OAI21X1 OAI21X1_1075 ( .A(w_mem_inst__abc_19396_new_n2432_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf58), .C(w_mem_inst__abc_19396_new_n2435_), .Y(w_mem_inst__0w_mem_13__31_0__2_));
OAI21X1 OAI21X1_1076 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf56), .B(w_mem_inst__abc_19396_new_n2438_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf90), .Y(w_mem_inst__abc_19396_new_n2439_));
OAI21X1 OAI21X1_1077 ( .A(w_mem_inst_w_mem_14__3_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf89), .C(w_mem_inst__abc_19396_new_n2439_), .Y(w_mem_inst__abc_19396_new_n2440_));
OAI21X1 OAI21X1_1078 ( .A(w_mem_inst__abc_19396_new_n2437_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf57), .C(w_mem_inst__abc_19396_new_n2440_), .Y(w_mem_inst__0w_mem_13__31_0__3_));
OAI21X1 OAI21X1_1079 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf55), .B(w_mem_inst__abc_19396_new_n2443_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf88), .Y(w_mem_inst__abc_19396_new_n2444_));
OAI21X1 OAI21X1_108 ( .A(_abc_15497_new_n1307_), .B(_abc_15497_new_n1308_), .C(_abc_15497_new_n1309_), .Y(_abc_15497_new_n1310_));
OAI21X1 OAI21X1_1080 ( .A(w_mem_inst_w_mem_14__4_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf87), .C(w_mem_inst__abc_19396_new_n2444_), .Y(w_mem_inst__abc_19396_new_n2445_));
OAI21X1 OAI21X1_1081 ( .A(w_mem_inst__abc_19396_new_n2442_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf56), .C(w_mem_inst__abc_19396_new_n2445_), .Y(w_mem_inst__0w_mem_13__31_0__4_));
OAI21X1 OAI21X1_1082 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf54), .B(w_mem_inst__abc_19396_new_n2448_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf86), .Y(w_mem_inst__abc_19396_new_n2449_));
OAI21X1 OAI21X1_1083 ( .A(w_mem_inst_w_mem_14__5_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf85), .C(w_mem_inst__abc_19396_new_n2449_), .Y(w_mem_inst__abc_19396_new_n2450_));
OAI21X1 OAI21X1_1084 ( .A(w_mem_inst__abc_19396_new_n2447_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf55), .C(w_mem_inst__abc_19396_new_n2450_), .Y(w_mem_inst__0w_mem_13__31_0__5_));
OAI21X1 OAI21X1_1085 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf53), .B(w_mem_inst__abc_19396_new_n2453_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf84), .Y(w_mem_inst__abc_19396_new_n2454_));
OAI21X1 OAI21X1_1086 ( .A(w_mem_inst_w_mem_14__6_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf83), .C(w_mem_inst__abc_19396_new_n2454_), .Y(w_mem_inst__abc_19396_new_n2455_));
OAI21X1 OAI21X1_1087 ( .A(w_mem_inst__abc_19396_new_n2452_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf54), .C(w_mem_inst__abc_19396_new_n2455_), .Y(w_mem_inst__0w_mem_13__31_0__6_));
OAI21X1 OAI21X1_1088 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf52), .B(w_mem_inst__abc_19396_new_n2458_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf82), .Y(w_mem_inst__abc_19396_new_n2459_));
OAI21X1 OAI21X1_1089 ( .A(w_mem_inst_w_mem_14__7_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf81), .C(w_mem_inst__abc_19396_new_n2459_), .Y(w_mem_inst__abc_19396_new_n2460_));
OAI21X1 OAI21X1_109 ( .A(_abc_15497_new_n1322_), .B(_abc_15497_new_n1318_), .C(digest_update_bF_buf1), .Y(_abc_15497_new_n1324_));
OAI21X1 OAI21X1_1090 ( .A(w_mem_inst__abc_19396_new_n2457_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf53), .C(w_mem_inst__abc_19396_new_n2460_), .Y(w_mem_inst__0w_mem_13__31_0__7_));
OAI21X1 OAI21X1_1091 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf51), .B(w_mem_inst__abc_19396_new_n2463_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf80), .Y(w_mem_inst__abc_19396_new_n2464_));
OAI21X1 OAI21X1_1092 ( .A(w_mem_inst_w_mem_14__8_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf79), .C(w_mem_inst__abc_19396_new_n2464_), .Y(w_mem_inst__abc_19396_new_n2465_));
OAI21X1 OAI21X1_1093 ( .A(w_mem_inst__abc_19396_new_n2462_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf52), .C(w_mem_inst__abc_19396_new_n2465_), .Y(w_mem_inst__0w_mem_13__31_0__8_));
OAI21X1 OAI21X1_1094 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf50), .B(w_mem_inst__abc_19396_new_n2468_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf78), .Y(w_mem_inst__abc_19396_new_n2469_));
OAI21X1 OAI21X1_1095 ( .A(w_mem_inst_w_mem_14__9_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf77), .C(w_mem_inst__abc_19396_new_n2469_), .Y(w_mem_inst__abc_19396_new_n2470_));
OAI21X1 OAI21X1_1096 ( .A(w_mem_inst__abc_19396_new_n2467_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf51), .C(w_mem_inst__abc_19396_new_n2470_), .Y(w_mem_inst__0w_mem_13__31_0__9_));
OAI21X1 OAI21X1_1097 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf49), .B(w_mem_inst__abc_19396_new_n2473_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf76), .Y(w_mem_inst__abc_19396_new_n2474_));
OAI21X1 OAI21X1_1098 ( .A(w_mem_inst_w_mem_14__10_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf75), .C(w_mem_inst__abc_19396_new_n2474_), .Y(w_mem_inst__abc_19396_new_n2475_));
OAI21X1 OAI21X1_1099 ( .A(w_mem_inst__abc_19396_new_n2472_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf50), .C(w_mem_inst__abc_19396_new_n2475_), .Y(w_mem_inst__0w_mem_13__31_0__10_));
OAI21X1 OAI21X1_11 ( .A(_auto_iopadmap_cc_368_execute_22625_91_), .B(_abc_15497_new_n883__bF_buf13), .C(_abc_15497_new_n870__bF_buf10), .Y(_abc_15497_new_n884_));
OAI21X1 OAI21X1_110 ( .A(_abc_15497_new_n1319_), .B(_abc_15497_new_n1318_), .C(_abc_15497_new_n1327_), .Y(_abc_15497_new_n1328_));
OAI21X1 OAI21X1_1100 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf48), .B(w_mem_inst__abc_19396_new_n2478_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf74), .Y(w_mem_inst__abc_19396_new_n2479_));
OAI21X1 OAI21X1_1101 ( .A(w_mem_inst_w_mem_14__11_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf73), .C(w_mem_inst__abc_19396_new_n2479_), .Y(w_mem_inst__abc_19396_new_n2480_));
OAI21X1 OAI21X1_1102 ( .A(w_mem_inst__abc_19396_new_n2477_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf49), .C(w_mem_inst__abc_19396_new_n2480_), .Y(w_mem_inst__0w_mem_13__31_0__11_));
OAI21X1 OAI21X1_1103 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf47), .B(w_mem_inst__abc_19396_new_n2483_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf72), .Y(w_mem_inst__abc_19396_new_n2484_));
OAI21X1 OAI21X1_1104 ( .A(w_mem_inst_w_mem_14__12_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf71), .C(w_mem_inst__abc_19396_new_n2484_), .Y(w_mem_inst__abc_19396_new_n2485_));
OAI21X1 OAI21X1_1105 ( .A(w_mem_inst__abc_19396_new_n2482_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf48), .C(w_mem_inst__abc_19396_new_n2485_), .Y(w_mem_inst__0w_mem_13__31_0__12_));
OAI21X1 OAI21X1_1106 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf46), .B(w_mem_inst__abc_19396_new_n2488_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf70), .Y(w_mem_inst__abc_19396_new_n2489_));
OAI21X1 OAI21X1_1107 ( .A(w_mem_inst_w_mem_14__13_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf69), .C(w_mem_inst__abc_19396_new_n2489_), .Y(w_mem_inst__abc_19396_new_n2490_));
OAI21X1 OAI21X1_1108 ( .A(w_mem_inst__abc_19396_new_n2487_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf47), .C(w_mem_inst__abc_19396_new_n2490_), .Y(w_mem_inst__0w_mem_13__31_0__13_));
OAI21X1 OAI21X1_1109 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf45), .B(w_mem_inst__abc_19396_new_n2493_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf68), .Y(w_mem_inst__abc_19396_new_n2494_));
OAI21X1 OAI21X1_111 ( .A(_abc_15497_new_n1332_), .B(_abc_15497_new_n1333_), .C(_abc_15497_new_n1334_), .Y(_abc_15497_new_n1335_));
OAI21X1 OAI21X1_1110 ( .A(w_mem_inst_w_mem_14__14_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf67), .C(w_mem_inst__abc_19396_new_n2494_), .Y(w_mem_inst__abc_19396_new_n2495_));
OAI21X1 OAI21X1_1111 ( .A(w_mem_inst__abc_19396_new_n2492_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf46), .C(w_mem_inst__abc_19396_new_n2495_), .Y(w_mem_inst__0w_mem_13__31_0__14_));
OAI21X1 OAI21X1_1112 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf44), .B(w_mem_inst__abc_19396_new_n2498_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf66), .Y(w_mem_inst__abc_19396_new_n2499_));
OAI21X1 OAI21X1_1113 ( .A(w_mem_inst_w_mem_14__15_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf65), .C(w_mem_inst__abc_19396_new_n2499_), .Y(w_mem_inst__abc_19396_new_n2500_));
OAI21X1 OAI21X1_1114 ( .A(w_mem_inst__abc_19396_new_n2497_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf45), .C(w_mem_inst__abc_19396_new_n2500_), .Y(w_mem_inst__0w_mem_13__31_0__15_));
OAI21X1 OAI21X1_1115 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf43), .B(w_mem_inst__abc_19396_new_n2503_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf64), .Y(w_mem_inst__abc_19396_new_n2504_));
OAI21X1 OAI21X1_1116 ( .A(w_mem_inst_w_mem_14__16_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf63), .C(w_mem_inst__abc_19396_new_n2504_), .Y(w_mem_inst__abc_19396_new_n2505_));
OAI21X1 OAI21X1_1117 ( .A(w_mem_inst__abc_19396_new_n2502_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf44), .C(w_mem_inst__abc_19396_new_n2505_), .Y(w_mem_inst__0w_mem_13__31_0__16_));
OAI21X1 OAI21X1_1118 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf42), .B(w_mem_inst__abc_19396_new_n2508_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf62), .Y(w_mem_inst__abc_19396_new_n2509_));
OAI21X1 OAI21X1_1119 ( .A(w_mem_inst_w_mem_14__17_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf61), .C(w_mem_inst__abc_19396_new_n2509_), .Y(w_mem_inst__abc_19396_new_n2510_));
OAI21X1 OAI21X1_112 ( .A(_auto_iopadmap_cc_368_execute_22625_37_), .B(_abc_15497_new_n883__bF_buf5), .C(_abc_15497_new_n870__bF_buf9), .Y(_abc_15497_new_n1340_));
OAI21X1 OAI21X1_1120 ( .A(w_mem_inst__abc_19396_new_n2507_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf43), .C(w_mem_inst__abc_19396_new_n2510_), .Y(w_mem_inst__0w_mem_13__31_0__17_));
OAI21X1 OAI21X1_1121 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf41), .B(w_mem_inst__abc_19396_new_n2513_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf60), .Y(w_mem_inst__abc_19396_new_n2514_));
OAI21X1 OAI21X1_1122 ( .A(w_mem_inst_w_mem_14__18_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf59), .C(w_mem_inst__abc_19396_new_n2514_), .Y(w_mem_inst__abc_19396_new_n2515_));
OAI21X1 OAI21X1_1123 ( .A(w_mem_inst__abc_19396_new_n2512_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf42), .C(w_mem_inst__abc_19396_new_n2515_), .Y(w_mem_inst__0w_mem_13__31_0__18_));
OAI21X1 OAI21X1_1124 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf40), .B(w_mem_inst__abc_19396_new_n2518_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf58), .Y(w_mem_inst__abc_19396_new_n2519_));
OAI21X1 OAI21X1_1125 ( .A(w_mem_inst_w_mem_14__19_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf57), .C(w_mem_inst__abc_19396_new_n2519_), .Y(w_mem_inst__abc_19396_new_n2520_));
OAI21X1 OAI21X1_1126 ( .A(w_mem_inst__abc_19396_new_n2517_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf41), .C(w_mem_inst__abc_19396_new_n2520_), .Y(w_mem_inst__0w_mem_13__31_0__19_));
OAI21X1 OAI21X1_1127 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf39), .B(w_mem_inst__abc_19396_new_n2523_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf56), .Y(w_mem_inst__abc_19396_new_n2524_));
OAI21X1 OAI21X1_1128 ( .A(w_mem_inst_w_mem_14__20_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf55), .C(w_mem_inst__abc_19396_new_n2524_), .Y(w_mem_inst__abc_19396_new_n2525_));
OAI21X1 OAI21X1_1129 ( .A(w_mem_inst__abc_19396_new_n2522_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf40), .C(w_mem_inst__abc_19396_new_n2525_), .Y(w_mem_inst__0w_mem_13__31_0__20_));
OAI21X1 OAI21X1_113 ( .A(_abc_15497_new_n1337_), .B(_abc_15497_new_n1339_), .C(_abc_15497_new_n1340_), .Y(_0H3_reg_31_0__5_));
OAI21X1 OAI21X1_1130 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf38), .B(w_mem_inst__abc_19396_new_n2528_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf54), .Y(w_mem_inst__abc_19396_new_n2529_));
OAI21X1 OAI21X1_1131 ( .A(w_mem_inst_w_mem_14__21_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf53), .C(w_mem_inst__abc_19396_new_n2529_), .Y(w_mem_inst__abc_19396_new_n2530_));
OAI21X1 OAI21X1_1132 ( .A(w_mem_inst__abc_19396_new_n2527_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf39), .C(w_mem_inst__abc_19396_new_n2530_), .Y(w_mem_inst__0w_mem_13__31_0__21_));
OAI21X1 OAI21X1_1133 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf37), .B(w_mem_inst__abc_19396_new_n2533_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf52), .Y(w_mem_inst__abc_19396_new_n2534_));
OAI21X1 OAI21X1_1134 ( .A(w_mem_inst_w_mem_14__22_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf51), .C(w_mem_inst__abc_19396_new_n2534_), .Y(w_mem_inst__abc_19396_new_n2535_));
OAI21X1 OAI21X1_1135 ( .A(w_mem_inst__abc_19396_new_n2532_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf38), .C(w_mem_inst__abc_19396_new_n2535_), .Y(w_mem_inst__0w_mem_13__31_0__22_));
OAI21X1 OAI21X1_1136 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf36), .B(w_mem_inst__abc_19396_new_n2538_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf50), .Y(w_mem_inst__abc_19396_new_n2539_));
OAI21X1 OAI21X1_1137 ( .A(w_mem_inst_w_mem_14__23_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf49), .C(w_mem_inst__abc_19396_new_n2539_), .Y(w_mem_inst__abc_19396_new_n2540_));
OAI21X1 OAI21X1_1138 ( .A(w_mem_inst__abc_19396_new_n2537_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf37), .C(w_mem_inst__abc_19396_new_n2540_), .Y(w_mem_inst__0w_mem_13__31_0__23_));
OAI21X1 OAI21X1_1139 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf35), .B(w_mem_inst__abc_19396_new_n2543_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf48), .Y(w_mem_inst__abc_19396_new_n2544_));
OAI21X1 OAI21X1_114 ( .A(_abc_15497_new_n1342_), .B(_abc_15497_new_n1343_), .C(_abc_15497_new_n1338_), .Y(_abc_15497_new_n1344_));
OAI21X1 OAI21X1_1140 ( .A(w_mem_inst_w_mem_14__24_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf47), .C(w_mem_inst__abc_19396_new_n2544_), .Y(w_mem_inst__abc_19396_new_n2545_));
OAI21X1 OAI21X1_1141 ( .A(w_mem_inst__abc_19396_new_n2542_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf36), .C(w_mem_inst__abc_19396_new_n2545_), .Y(w_mem_inst__0w_mem_13__31_0__24_));
OAI21X1 OAI21X1_1142 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf34), .B(w_mem_inst__abc_19396_new_n2548_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf46), .Y(w_mem_inst__abc_19396_new_n2549_));
OAI21X1 OAI21X1_1143 ( .A(w_mem_inst_w_mem_14__25_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf45), .C(w_mem_inst__abc_19396_new_n2549_), .Y(w_mem_inst__abc_19396_new_n2550_));
OAI21X1 OAI21X1_1144 ( .A(w_mem_inst__abc_19396_new_n2547_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf35), .C(w_mem_inst__abc_19396_new_n2550_), .Y(w_mem_inst__0w_mem_13__31_0__25_));
OAI21X1 OAI21X1_1145 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf33), .B(w_mem_inst__abc_19396_new_n2553_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf44), .Y(w_mem_inst__abc_19396_new_n2554_));
OAI21X1 OAI21X1_1146 ( .A(w_mem_inst_w_mem_14__26_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf43), .C(w_mem_inst__abc_19396_new_n2554_), .Y(w_mem_inst__abc_19396_new_n2555_));
OAI21X1 OAI21X1_1147 ( .A(w_mem_inst__abc_19396_new_n2552_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf34), .C(w_mem_inst__abc_19396_new_n2555_), .Y(w_mem_inst__0w_mem_13__31_0__26_));
OAI21X1 OAI21X1_1148 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf32), .B(w_mem_inst__abc_19396_new_n2558_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf42), .Y(w_mem_inst__abc_19396_new_n2559_));
OAI21X1 OAI21X1_1149 ( .A(w_mem_inst_w_mem_14__27_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf41), .C(w_mem_inst__abc_19396_new_n2559_), .Y(w_mem_inst__abc_19396_new_n2560_));
OAI21X1 OAI21X1_115 ( .A(_auto_iopadmap_cc_368_execute_22625_38_), .B(_abc_15497_new_n883__bF_buf4), .C(_abc_15497_new_n870__bF_buf8), .Y(_abc_15497_new_n1349_));
OAI21X1 OAI21X1_1150 ( .A(w_mem_inst__abc_19396_new_n2557_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf33), .C(w_mem_inst__abc_19396_new_n2560_), .Y(w_mem_inst__0w_mem_13__31_0__27_));
OAI21X1 OAI21X1_1151 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf31), .B(w_mem_inst__abc_19396_new_n2563_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf40), .Y(w_mem_inst__abc_19396_new_n2564_));
OAI21X1 OAI21X1_1152 ( .A(w_mem_inst_w_mem_14__28_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf39), .C(w_mem_inst__abc_19396_new_n2564_), .Y(w_mem_inst__abc_19396_new_n2565_));
OAI21X1 OAI21X1_1153 ( .A(w_mem_inst__abc_19396_new_n2562_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf32), .C(w_mem_inst__abc_19396_new_n2565_), .Y(w_mem_inst__0w_mem_13__31_0__28_));
OAI21X1 OAI21X1_1154 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf30), .B(w_mem_inst__abc_19396_new_n2568_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf38), .Y(w_mem_inst__abc_19396_new_n2569_));
OAI21X1 OAI21X1_1155 ( .A(w_mem_inst_w_mem_14__29_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf37), .C(w_mem_inst__abc_19396_new_n2569_), .Y(w_mem_inst__abc_19396_new_n2570_));
OAI21X1 OAI21X1_1156 ( .A(w_mem_inst__abc_19396_new_n2567_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf31), .C(w_mem_inst__abc_19396_new_n2570_), .Y(w_mem_inst__0w_mem_13__31_0__29_));
OAI21X1 OAI21X1_1157 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf29), .B(w_mem_inst__abc_19396_new_n2573_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf36), .Y(w_mem_inst__abc_19396_new_n2574_));
OAI21X1 OAI21X1_1158 ( .A(w_mem_inst_w_mem_14__30_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf35), .C(w_mem_inst__abc_19396_new_n2574_), .Y(w_mem_inst__abc_19396_new_n2575_));
OAI21X1 OAI21X1_1159 ( .A(w_mem_inst__abc_19396_new_n2572_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf30), .C(w_mem_inst__abc_19396_new_n2575_), .Y(w_mem_inst__0w_mem_13__31_0__30_));
OAI21X1 OAI21X1_116 ( .A(_abc_15497_new_n1346_), .B(_abc_15497_new_n1348_), .C(_abc_15497_new_n1349_), .Y(_0H3_reg_31_0__6_));
OAI21X1 OAI21X1_1160 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf28), .B(w_mem_inst__abc_19396_new_n2578_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf34), .Y(w_mem_inst__abc_19396_new_n2579_));
OAI21X1 OAI21X1_1161 ( .A(w_mem_inst_w_mem_14__31_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf33), .C(w_mem_inst__abc_19396_new_n2579_), .Y(w_mem_inst__abc_19396_new_n2580_));
OAI21X1 OAI21X1_1162 ( .A(w_mem_inst__abc_19396_new_n2577_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf29), .C(w_mem_inst__abc_19396_new_n2580_), .Y(w_mem_inst__0w_mem_13__31_0__31_));
OAI21X1 OAI21X1_1163 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf27), .B(w_mem_inst__abc_19396_new_n2648_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf31), .Y(w_mem_inst__abc_19396_new_n2649_));
OAI21X1 OAI21X1_1164 ( .A(w_mem_inst_w_mem_15__0_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf30), .C(w_mem_inst__abc_19396_new_n2649_), .Y(w_mem_inst__abc_19396_new_n2650_));
OAI21X1 OAI21X1_1165 ( .A(w_mem_inst__abc_19396_new_n2647_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf28), .C(w_mem_inst__abc_19396_new_n2650_), .Y(w_mem_inst__0w_mem_14__31_0__0_));
OAI21X1 OAI21X1_1166 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf26), .B(w_mem_inst__abc_19396_new_n2653_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf29), .Y(w_mem_inst__abc_19396_new_n2654_));
OAI21X1 OAI21X1_1167 ( .A(w_mem_inst_w_mem_15__1_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf28), .C(w_mem_inst__abc_19396_new_n2654_), .Y(w_mem_inst__abc_19396_new_n2655_));
OAI21X1 OAI21X1_1168 ( .A(w_mem_inst__abc_19396_new_n2652_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf27), .C(w_mem_inst__abc_19396_new_n2655_), .Y(w_mem_inst__0w_mem_14__31_0__1_));
OAI21X1 OAI21X1_1169 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf25), .B(w_mem_inst__abc_19396_new_n2658_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf27), .Y(w_mem_inst__abc_19396_new_n2659_));
OAI21X1 OAI21X1_117 ( .A(_abc_15497_new_n1356_), .B(_abc_15497_new_n1357_), .C(_abc_15497_new_n1347_), .Y(_abc_15497_new_n1358_));
OAI21X1 OAI21X1_1170 ( .A(w_mem_inst_w_mem_15__2_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf26), .C(w_mem_inst__abc_19396_new_n2659_), .Y(w_mem_inst__abc_19396_new_n2660_));
OAI21X1 OAI21X1_1171 ( .A(w_mem_inst__abc_19396_new_n2657_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf26), .C(w_mem_inst__abc_19396_new_n2660_), .Y(w_mem_inst__0w_mem_14__31_0__2_));
OAI21X1 OAI21X1_1172 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf24), .B(w_mem_inst__abc_19396_new_n2663_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf25), .Y(w_mem_inst__abc_19396_new_n2664_));
OAI21X1 OAI21X1_1173 ( .A(w_mem_inst_w_mem_15__3_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf24), .C(w_mem_inst__abc_19396_new_n2664_), .Y(w_mem_inst__abc_19396_new_n2665_));
OAI21X1 OAI21X1_1174 ( .A(w_mem_inst__abc_19396_new_n2662_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf25), .C(w_mem_inst__abc_19396_new_n2665_), .Y(w_mem_inst__0w_mem_14__31_0__3_));
OAI21X1 OAI21X1_1175 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf23), .B(w_mem_inst__abc_19396_new_n2668_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf23), .Y(w_mem_inst__abc_19396_new_n2669_));
OAI21X1 OAI21X1_1176 ( .A(w_mem_inst_w_mem_15__4_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf22), .C(w_mem_inst__abc_19396_new_n2669_), .Y(w_mem_inst__abc_19396_new_n2670_));
OAI21X1 OAI21X1_1177 ( .A(w_mem_inst__abc_19396_new_n2667_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf24), .C(w_mem_inst__abc_19396_new_n2670_), .Y(w_mem_inst__0w_mem_14__31_0__4_));
OAI21X1 OAI21X1_1178 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf22), .B(w_mem_inst__abc_19396_new_n2673_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf21), .Y(w_mem_inst__abc_19396_new_n2674_));
OAI21X1 OAI21X1_1179 ( .A(w_mem_inst_w_mem_15__5_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf20), .C(w_mem_inst__abc_19396_new_n2674_), .Y(w_mem_inst__abc_19396_new_n2675_));
OAI21X1 OAI21X1_118 ( .A(_abc_15497_new_n1367_), .B(_abc_15497_new_n1362_), .C(digest_update_bF_buf6), .Y(_abc_15497_new_n1369_));
OAI21X1 OAI21X1_1180 ( .A(w_mem_inst__abc_19396_new_n2672_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf23), .C(w_mem_inst__abc_19396_new_n2675_), .Y(w_mem_inst__0w_mem_14__31_0__5_));
OAI21X1 OAI21X1_1181 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf21), .B(w_mem_inst__abc_19396_new_n2678_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf19), .Y(w_mem_inst__abc_19396_new_n2679_));
OAI21X1 OAI21X1_1182 ( .A(w_mem_inst_w_mem_15__6_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf18), .C(w_mem_inst__abc_19396_new_n2679_), .Y(w_mem_inst__abc_19396_new_n2680_));
OAI21X1 OAI21X1_1183 ( .A(w_mem_inst__abc_19396_new_n2677_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf22), .C(w_mem_inst__abc_19396_new_n2680_), .Y(w_mem_inst__0w_mem_14__31_0__6_));
OAI21X1 OAI21X1_1184 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf20), .B(w_mem_inst__abc_19396_new_n2683_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf17), .Y(w_mem_inst__abc_19396_new_n2684_));
OAI21X1 OAI21X1_1185 ( .A(w_mem_inst_w_mem_15__7_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf16), .C(w_mem_inst__abc_19396_new_n2684_), .Y(w_mem_inst__abc_19396_new_n2685_));
OAI21X1 OAI21X1_1186 ( .A(w_mem_inst__abc_19396_new_n2682_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf21), .C(w_mem_inst__abc_19396_new_n2685_), .Y(w_mem_inst__0w_mem_14__31_0__7_));
OAI21X1 OAI21X1_1187 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf19), .B(w_mem_inst__abc_19396_new_n2688_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf15), .Y(w_mem_inst__abc_19396_new_n2689_));
OAI21X1 OAI21X1_1188 ( .A(w_mem_inst_w_mem_15__8_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf14), .C(w_mem_inst__abc_19396_new_n2689_), .Y(w_mem_inst__abc_19396_new_n2690_));
OAI21X1 OAI21X1_1189 ( .A(w_mem_inst__abc_19396_new_n2687_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf20), .C(w_mem_inst__abc_19396_new_n2690_), .Y(w_mem_inst__0w_mem_14__31_0__8_));
OAI21X1 OAI21X1_119 ( .A(_abc_15497_new_n1361_), .B(_abc_15497_new_n1364_), .C(_abc_15497_new_n1377_), .Y(_abc_15497_new_n1378_));
OAI21X1 OAI21X1_1190 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf18), .B(w_mem_inst__abc_19396_new_n2693_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf13), .Y(w_mem_inst__abc_19396_new_n2694_));
OAI21X1 OAI21X1_1191 ( .A(w_mem_inst_w_mem_15__9_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf12), .C(w_mem_inst__abc_19396_new_n2694_), .Y(w_mem_inst__abc_19396_new_n2695_));
OAI21X1 OAI21X1_1192 ( .A(w_mem_inst__abc_19396_new_n2692_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf19), .C(w_mem_inst__abc_19396_new_n2695_), .Y(w_mem_inst__0w_mem_14__31_0__9_));
OAI21X1 OAI21X1_1193 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf17), .B(w_mem_inst__abc_19396_new_n2698_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf11), .Y(w_mem_inst__abc_19396_new_n2699_));
OAI21X1 OAI21X1_1194 ( .A(w_mem_inst_w_mem_15__10_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf10), .C(w_mem_inst__abc_19396_new_n2699_), .Y(w_mem_inst__abc_19396_new_n2700_));
OAI21X1 OAI21X1_1195 ( .A(w_mem_inst__abc_19396_new_n2697_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf18), .C(w_mem_inst__abc_19396_new_n2700_), .Y(w_mem_inst__0w_mem_14__31_0__10_));
OAI21X1 OAI21X1_1196 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf16), .B(w_mem_inst__abc_19396_new_n2703_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf9), .Y(w_mem_inst__abc_19396_new_n2704_));
OAI21X1 OAI21X1_1197 ( .A(w_mem_inst_w_mem_15__11_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf8), .C(w_mem_inst__abc_19396_new_n2704_), .Y(w_mem_inst__abc_19396_new_n2705_));
OAI21X1 OAI21X1_1198 ( .A(w_mem_inst__abc_19396_new_n2702_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf17), .C(w_mem_inst__abc_19396_new_n2705_), .Y(w_mem_inst__0w_mem_14__31_0__11_));
OAI21X1 OAI21X1_1199 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf15), .B(w_mem_inst__abc_19396_new_n2708_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf7), .Y(w_mem_inst__abc_19396_new_n2709_));
OAI21X1 OAI21X1_12 ( .A(_abc_15497_new_n870__bF_buf9), .B(_abc_15497_new_n882_), .C(_abc_15497_new_n884_), .Y(_0H2_reg_31_0__27_));
OAI21X1 OAI21X1_120 ( .A(_abc_15497_new_n1365_), .B(_abc_15497_new_n1372_), .C(_abc_15497_new_n1376_), .Y(_abc_15497_new_n1379_));
OAI21X1 OAI21X1_1200 ( .A(w_mem_inst_w_mem_15__12_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf6), .C(w_mem_inst__abc_19396_new_n2709_), .Y(w_mem_inst__abc_19396_new_n2710_));
OAI21X1 OAI21X1_1201 ( .A(w_mem_inst__abc_19396_new_n2707_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf16), .C(w_mem_inst__abc_19396_new_n2710_), .Y(w_mem_inst__0w_mem_14__31_0__12_));
OAI21X1 OAI21X1_1202 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf14), .B(w_mem_inst__abc_19396_new_n2713_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf5), .Y(w_mem_inst__abc_19396_new_n2714_));
OAI21X1 OAI21X1_1203 ( .A(w_mem_inst_w_mem_15__13_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf4), .C(w_mem_inst__abc_19396_new_n2714_), .Y(w_mem_inst__abc_19396_new_n2715_));
OAI21X1 OAI21X1_1204 ( .A(w_mem_inst__abc_19396_new_n2712_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf15), .C(w_mem_inst__abc_19396_new_n2715_), .Y(w_mem_inst__0w_mem_14__31_0__13_));
OAI21X1 OAI21X1_1205 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf13), .B(w_mem_inst__abc_19396_new_n2718_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf3), .Y(w_mem_inst__abc_19396_new_n2719_));
OAI21X1 OAI21X1_1206 ( .A(w_mem_inst_w_mem_15__14_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf2), .C(w_mem_inst__abc_19396_new_n2719_), .Y(w_mem_inst__abc_19396_new_n2720_));
OAI21X1 OAI21X1_1207 ( .A(w_mem_inst__abc_19396_new_n2717_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf14), .C(w_mem_inst__abc_19396_new_n2720_), .Y(w_mem_inst__0w_mem_14__31_0__14_));
OAI21X1 OAI21X1_1208 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf12), .B(w_mem_inst__abc_19396_new_n2723_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf1), .Y(w_mem_inst__abc_19396_new_n2724_));
OAI21X1 OAI21X1_1209 ( .A(w_mem_inst_w_mem_15__15_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf0), .C(w_mem_inst__abc_19396_new_n2724_), .Y(w_mem_inst__abc_19396_new_n2725_));
OAI21X1 OAI21X1_121 ( .A(_abc_15497_new_n1372_), .B(_abc_15497_new_n1378_), .C(_abc_15497_new_n1379_), .Y(_abc_15497_new_n1380_));
OAI21X1 OAI21X1_1210 ( .A(w_mem_inst__abc_19396_new_n2722_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf13), .C(w_mem_inst__abc_19396_new_n2725_), .Y(w_mem_inst__0w_mem_14__31_0__15_));
OAI21X1 OAI21X1_1211 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf11), .B(w_mem_inst__abc_19396_new_n2728_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf96), .Y(w_mem_inst__abc_19396_new_n2729_));
OAI21X1 OAI21X1_1212 ( .A(w_mem_inst_w_mem_15__16_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf95), .C(w_mem_inst__abc_19396_new_n2729_), .Y(w_mem_inst__abc_19396_new_n2730_));
OAI21X1 OAI21X1_1213 ( .A(w_mem_inst__abc_19396_new_n2727_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf12), .C(w_mem_inst__abc_19396_new_n2730_), .Y(w_mem_inst__0w_mem_14__31_0__16_));
OAI21X1 OAI21X1_1214 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf10), .B(w_mem_inst__abc_19396_new_n2733_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf94), .Y(w_mem_inst__abc_19396_new_n2734_));
OAI21X1 OAI21X1_1215 ( .A(w_mem_inst_w_mem_15__17_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf93), .C(w_mem_inst__abc_19396_new_n2734_), .Y(w_mem_inst__abc_19396_new_n2735_));
OAI21X1 OAI21X1_1216 ( .A(w_mem_inst__abc_19396_new_n2732_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf11), .C(w_mem_inst__abc_19396_new_n2735_), .Y(w_mem_inst__0w_mem_14__31_0__17_));
OAI21X1 OAI21X1_1217 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf9), .B(w_mem_inst__abc_19396_new_n2738_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf92), .Y(w_mem_inst__abc_19396_new_n2739_));
OAI21X1 OAI21X1_1218 ( .A(w_mem_inst_w_mem_15__18_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf91), .C(w_mem_inst__abc_19396_new_n2739_), .Y(w_mem_inst__abc_19396_new_n2740_));
OAI21X1 OAI21X1_1219 ( .A(w_mem_inst__abc_19396_new_n2737_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf10), .C(w_mem_inst__abc_19396_new_n2740_), .Y(w_mem_inst__0w_mem_14__31_0__18_));
OAI21X1 OAI21X1_122 ( .A(_abc_15497_new_n1383_), .B(_abc_15497_new_n1362_), .C(_abc_15497_new_n1384_), .Y(_abc_15497_new_n1385_));
OAI21X1 OAI21X1_1220 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf8), .B(w_mem_inst__abc_19396_new_n2743_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf90), .Y(w_mem_inst__abc_19396_new_n2744_));
OAI21X1 OAI21X1_1221 ( .A(w_mem_inst_w_mem_15__19_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf89), .C(w_mem_inst__abc_19396_new_n2744_), .Y(w_mem_inst__abc_19396_new_n2745_));
OAI21X1 OAI21X1_1222 ( .A(w_mem_inst__abc_19396_new_n2742_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf9), .C(w_mem_inst__abc_19396_new_n2745_), .Y(w_mem_inst__0w_mem_14__31_0__19_));
OAI21X1 OAI21X1_1223 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf7), .B(w_mem_inst__abc_19396_new_n2748_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf88), .Y(w_mem_inst__abc_19396_new_n2749_));
OAI21X1 OAI21X1_1224 ( .A(w_mem_inst_w_mem_15__20_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf87), .C(w_mem_inst__abc_19396_new_n2749_), .Y(w_mem_inst__abc_19396_new_n2750_));
OAI21X1 OAI21X1_1225 ( .A(w_mem_inst__abc_19396_new_n2747_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf8), .C(w_mem_inst__abc_19396_new_n2750_), .Y(w_mem_inst__0w_mem_14__31_0__20_));
OAI21X1 OAI21X1_1226 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf6), .B(w_mem_inst__abc_19396_new_n2753_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf86), .Y(w_mem_inst__abc_19396_new_n2754_));
OAI21X1 OAI21X1_1227 ( .A(w_mem_inst_w_mem_15__21_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf85), .C(w_mem_inst__abc_19396_new_n2754_), .Y(w_mem_inst__abc_19396_new_n2755_));
OAI21X1 OAI21X1_1228 ( .A(w_mem_inst__abc_19396_new_n2752_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf7), .C(w_mem_inst__abc_19396_new_n2755_), .Y(w_mem_inst__0w_mem_14__31_0__21_));
OAI21X1 OAI21X1_1229 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf5), .B(w_mem_inst__abc_19396_new_n2758_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf84), .Y(w_mem_inst__abc_19396_new_n2759_));
OAI21X1 OAI21X1_123 ( .A(_abc_15497_new_n1385_), .B(_abc_15497_new_n1389_), .C(_abc_15497_new_n1391_), .Y(_abc_15497_new_n1392_));
OAI21X1 OAI21X1_1230 ( .A(w_mem_inst_w_mem_15__22_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf83), .C(w_mem_inst__abc_19396_new_n2759_), .Y(w_mem_inst__abc_19396_new_n2760_));
OAI21X1 OAI21X1_1231 ( .A(w_mem_inst__abc_19396_new_n2757_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf6), .C(w_mem_inst__abc_19396_new_n2760_), .Y(w_mem_inst__0w_mem_14__31_0__22_));
OAI21X1 OAI21X1_1232 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf4), .B(w_mem_inst__abc_19396_new_n2763_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf82), .Y(w_mem_inst__abc_19396_new_n2764_));
OAI21X1 OAI21X1_1233 ( .A(w_mem_inst_w_mem_15__23_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf81), .C(w_mem_inst__abc_19396_new_n2764_), .Y(w_mem_inst__abc_19396_new_n2765_));
OAI21X1 OAI21X1_1234 ( .A(w_mem_inst__abc_19396_new_n2762_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf5), .C(w_mem_inst__abc_19396_new_n2765_), .Y(w_mem_inst__0w_mem_14__31_0__23_));
OAI21X1 OAI21X1_1235 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf3), .B(w_mem_inst__abc_19396_new_n2768_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf80), .Y(w_mem_inst__abc_19396_new_n2769_));
OAI21X1 OAI21X1_1236 ( .A(w_mem_inst_w_mem_15__24_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf79), .C(w_mem_inst__abc_19396_new_n2769_), .Y(w_mem_inst__abc_19396_new_n2770_));
OAI21X1 OAI21X1_1237 ( .A(w_mem_inst__abc_19396_new_n2767_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf4), .C(w_mem_inst__abc_19396_new_n2770_), .Y(w_mem_inst__0w_mem_14__31_0__24_));
OAI21X1 OAI21X1_1238 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf2), .B(w_mem_inst__abc_19396_new_n2773_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf78), .Y(w_mem_inst__abc_19396_new_n2774_));
OAI21X1 OAI21X1_1239 ( .A(w_mem_inst_w_mem_15__25_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf77), .C(w_mem_inst__abc_19396_new_n2774_), .Y(w_mem_inst__abc_19396_new_n2775_));
OAI21X1 OAI21X1_124 ( .A(_auto_iopadmap_cc_368_execute_22625_42_), .B(_abc_15497_new_n883__bF_buf3), .C(_abc_15497_new_n870__bF_buf4), .Y(_abc_15497_new_n1393_));
OAI21X1 OAI21X1_1240 ( .A(w_mem_inst__abc_19396_new_n2772_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf3), .C(w_mem_inst__abc_19396_new_n2775_), .Y(w_mem_inst__0w_mem_14__31_0__25_));
OAI21X1 OAI21X1_1241 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf1), .B(w_mem_inst__abc_19396_new_n2778_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf76), .Y(w_mem_inst__abc_19396_new_n2779_));
OAI21X1 OAI21X1_1242 ( .A(w_mem_inst_w_mem_15__26_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf75), .C(w_mem_inst__abc_19396_new_n2779_), .Y(w_mem_inst__abc_19396_new_n2780_));
OAI21X1 OAI21X1_1243 ( .A(w_mem_inst__abc_19396_new_n2777_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf2), .C(w_mem_inst__abc_19396_new_n2780_), .Y(w_mem_inst__0w_mem_14__31_0__26_));
OAI21X1 OAI21X1_1244 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf0), .B(w_mem_inst__abc_19396_new_n2783_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf74), .Y(w_mem_inst__abc_19396_new_n2784_));
OAI21X1 OAI21X1_1245 ( .A(w_mem_inst_w_mem_15__27_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf73), .C(w_mem_inst__abc_19396_new_n2784_), .Y(w_mem_inst__abc_19396_new_n2785_));
OAI21X1 OAI21X1_1246 ( .A(w_mem_inst__abc_19396_new_n2782_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf1), .C(w_mem_inst__abc_19396_new_n2785_), .Y(w_mem_inst__0w_mem_14__31_0__27_));
OAI21X1 OAI21X1_1247 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf60), .B(w_mem_inst__abc_19396_new_n2788_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf72), .Y(w_mem_inst__abc_19396_new_n2789_));
OAI21X1 OAI21X1_1248 ( .A(w_mem_inst_w_mem_15__28_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf71), .C(w_mem_inst__abc_19396_new_n2789_), .Y(w_mem_inst__abc_19396_new_n2790_));
OAI21X1 OAI21X1_1249 ( .A(w_mem_inst__abc_19396_new_n2787_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf0), .C(w_mem_inst__abc_19396_new_n2790_), .Y(w_mem_inst__0w_mem_14__31_0__28_));
OAI21X1 OAI21X1_125 ( .A(_abc_15497_new_n1401_), .B(_abc_15497_new_n1396_), .C(digest_update_bF_buf5), .Y(_abc_15497_new_n1403_));
OAI21X1 OAI21X1_1250 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf59), .B(w_mem_inst__abc_19396_new_n2793_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf70), .Y(w_mem_inst__abc_19396_new_n2794_));
OAI21X1 OAI21X1_1251 ( .A(w_mem_inst_w_mem_15__29_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf69), .C(w_mem_inst__abc_19396_new_n2794_), .Y(w_mem_inst__abc_19396_new_n2795_));
OAI21X1 OAI21X1_1252 ( .A(w_mem_inst__abc_19396_new_n2792_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf60), .C(w_mem_inst__abc_19396_new_n2795_), .Y(w_mem_inst__0w_mem_14__31_0__29_));
OAI21X1 OAI21X1_1253 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf58), .B(w_mem_inst__abc_19396_new_n2798_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf68), .Y(w_mem_inst__abc_19396_new_n2799_));
OAI21X1 OAI21X1_1254 ( .A(w_mem_inst_w_mem_15__30_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf67), .C(w_mem_inst__abc_19396_new_n2799_), .Y(w_mem_inst__abc_19396_new_n2800_));
OAI21X1 OAI21X1_1255 ( .A(w_mem_inst__abc_19396_new_n2797_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf59), .C(w_mem_inst__abc_19396_new_n2800_), .Y(w_mem_inst__0w_mem_14__31_0__30_));
OAI21X1 OAI21X1_1256 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf57), .B(w_mem_inst__abc_19396_new_n2803_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf66), .Y(w_mem_inst__abc_19396_new_n2804_));
OAI21X1 OAI21X1_1257 ( .A(w_mem_inst_w_mem_15__31_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf65), .C(w_mem_inst__abc_19396_new_n2804_), .Y(w_mem_inst__abc_19396_new_n2805_));
OAI21X1 OAI21X1_1258 ( .A(w_mem_inst__abc_19396_new_n2802_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf58), .C(w_mem_inst__abc_19396_new_n2805_), .Y(w_mem_inst__0w_mem_14__31_0__31_));
OAI21X1 OAI21X1_1259 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf56), .B(w_mem_inst__abc_19396_new_n2808_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf64), .Y(w_mem_inst__abc_19396_new_n2809_));
OAI21X1 OAI21X1_126 ( .A(_abc_15497_new_n1405_), .B(_abc_15497_new_n1384_), .C(_abc_15497_new_n1408_), .Y(_abc_15497_new_n1409_));
OAI21X1 OAI21X1_1260 ( .A(w_mem_inst_w_mem_11__0_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf63), .C(w_mem_inst__abc_19396_new_n2809_), .Y(w_mem_inst__abc_19396_new_n2810_));
OAI21X1 OAI21X1_1261 ( .A(w_mem_inst__abc_19396_new_n2807_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf57), .C(w_mem_inst__abc_19396_new_n2810_), .Y(w_mem_inst__0w_mem_10__31_0__0_));
OAI21X1 OAI21X1_1262 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf55), .B(w_mem_inst__abc_19396_new_n2813_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf62), .Y(w_mem_inst__abc_19396_new_n2814_));
OAI21X1 OAI21X1_1263 ( .A(w_mem_inst_w_mem_11__1_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf61), .C(w_mem_inst__abc_19396_new_n2814_), .Y(w_mem_inst__abc_19396_new_n2815_));
OAI21X1 OAI21X1_1264 ( .A(w_mem_inst__abc_19396_new_n2812_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf56), .C(w_mem_inst__abc_19396_new_n2815_), .Y(w_mem_inst__0w_mem_10__31_0__1_));
OAI21X1 OAI21X1_1265 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf54), .B(w_mem_inst__abc_19396_new_n2818_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf60), .Y(w_mem_inst__abc_19396_new_n2819_));
OAI21X1 OAI21X1_1266 ( .A(w_mem_inst_w_mem_11__2_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf59), .C(w_mem_inst__abc_19396_new_n2819_), .Y(w_mem_inst__abc_19396_new_n2820_));
OAI21X1 OAI21X1_1267 ( .A(w_mem_inst__abc_19396_new_n2817_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf55), .C(w_mem_inst__abc_19396_new_n2820_), .Y(w_mem_inst__0w_mem_10__31_0__2_));
OAI21X1 OAI21X1_1268 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf53), .B(w_mem_inst__abc_19396_new_n2823_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf58), .Y(w_mem_inst__abc_19396_new_n2824_));
OAI21X1 OAI21X1_1269 ( .A(w_mem_inst_w_mem_11__3_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf57), .C(w_mem_inst__abc_19396_new_n2824_), .Y(w_mem_inst__abc_19396_new_n2825_));
OAI21X1 OAI21X1_127 ( .A(_abc_15497_new_n1407_), .B(_abc_15497_new_n1362_), .C(_abc_15497_new_n1410_), .Y(_abc_15497_new_n1411_));
OAI21X1 OAI21X1_1270 ( .A(w_mem_inst__abc_19396_new_n2822_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf54), .C(w_mem_inst__abc_19396_new_n2825_), .Y(w_mem_inst__0w_mem_10__31_0__3_));
OAI21X1 OAI21X1_1271 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf52), .B(w_mem_inst__abc_19396_new_n2828_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf56), .Y(w_mem_inst__abc_19396_new_n2829_));
OAI21X1 OAI21X1_1272 ( .A(w_mem_inst_w_mem_11__4_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf55), .C(w_mem_inst__abc_19396_new_n2829_), .Y(w_mem_inst__abc_19396_new_n2830_));
OAI21X1 OAI21X1_1273 ( .A(w_mem_inst__abc_19396_new_n2827_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf53), .C(w_mem_inst__abc_19396_new_n2830_), .Y(w_mem_inst__0w_mem_10__31_0__4_));
OAI21X1 OAI21X1_1274 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf51), .B(w_mem_inst__abc_19396_new_n2833_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf54), .Y(w_mem_inst__abc_19396_new_n2834_));
OAI21X1 OAI21X1_1275 ( .A(w_mem_inst_w_mem_11__5_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf53), .C(w_mem_inst__abc_19396_new_n2834_), .Y(w_mem_inst__abc_19396_new_n2835_));
OAI21X1 OAI21X1_1276 ( .A(w_mem_inst__abc_19396_new_n2832_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf52), .C(w_mem_inst__abc_19396_new_n2835_), .Y(w_mem_inst__0w_mem_10__31_0__5_));
OAI21X1 OAI21X1_1277 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf50), .B(w_mem_inst__abc_19396_new_n2838_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf52), .Y(w_mem_inst__abc_19396_new_n2839_));
OAI21X1 OAI21X1_1278 ( .A(w_mem_inst_w_mem_11__6_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf51), .C(w_mem_inst__abc_19396_new_n2839_), .Y(w_mem_inst__abc_19396_new_n2840_));
OAI21X1 OAI21X1_1279 ( .A(w_mem_inst__abc_19396_new_n2837_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf51), .C(w_mem_inst__abc_19396_new_n2840_), .Y(w_mem_inst__0w_mem_10__31_0__6_));
OAI21X1 OAI21X1_128 ( .A(_auto_iopadmap_cc_368_execute_22625_44_), .B(_abc_15497_new_n883__bF_buf2), .C(_abc_15497_new_n870__bF_buf3), .Y(_abc_15497_new_n1420_));
OAI21X1 OAI21X1_1280 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf49), .B(w_mem_inst__abc_19396_new_n2843_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf50), .Y(w_mem_inst__abc_19396_new_n2844_));
OAI21X1 OAI21X1_1281 ( .A(w_mem_inst_w_mem_11__7_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf49), .C(w_mem_inst__abc_19396_new_n2844_), .Y(w_mem_inst__abc_19396_new_n2845_));
OAI21X1 OAI21X1_1282 ( .A(w_mem_inst__abc_19396_new_n2842_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf50), .C(w_mem_inst__abc_19396_new_n2845_), .Y(w_mem_inst__0w_mem_10__31_0__7_));
OAI21X1 OAI21X1_1283 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf48), .B(w_mem_inst__abc_19396_new_n2848_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf48), .Y(w_mem_inst__abc_19396_new_n2849_));
OAI21X1 OAI21X1_1284 ( .A(w_mem_inst_w_mem_11__8_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf47), .C(w_mem_inst__abc_19396_new_n2849_), .Y(w_mem_inst__abc_19396_new_n2850_));
OAI21X1 OAI21X1_1285 ( .A(w_mem_inst__abc_19396_new_n2847_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf49), .C(w_mem_inst__abc_19396_new_n2850_), .Y(w_mem_inst__0w_mem_10__31_0__8_));
OAI21X1 OAI21X1_1286 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf47), .B(w_mem_inst__abc_19396_new_n2853_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf46), .Y(w_mem_inst__abc_19396_new_n2854_));
OAI21X1 OAI21X1_1287 ( .A(w_mem_inst_w_mem_11__9_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf45), .C(w_mem_inst__abc_19396_new_n2854_), .Y(w_mem_inst__abc_19396_new_n2855_));
OAI21X1 OAI21X1_1288 ( .A(w_mem_inst__abc_19396_new_n2852_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf48), .C(w_mem_inst__abc_19396_new_n2855_), .Y(w_mem_inst__0w_mem_10__31_0__9_));
OAI21X1 OAI21X1_1289 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf46), .B(w_mem_inst__abc_19396_new_n2858_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf44), .Y(w_mem_inst__abc_19396_new_n2859_));
OAI21X1 OAI21X1_129 ( .A(_abc_15497_new_n1417_), .B(_abc_15497_new_n1419_), .C(_abc_15497_new_n1420_), .Y(_0H3_reg_31_0__12_));
OAI21X1 OAI21X1_1290 ( .A(w_mem_inst_w_mem_11__10_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf43), .C(w_mem_inst__abc_19396_new_n2859_), .Y(w_mem_inst__abc_19396_new_n2860_));
OAI21X1 OAI21X1_1291 ( .A(w_mem_inst__abc_19396_new_n2857_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf47), .C(w_mem_inst__abc_19396_new_n2860_), .Y(w_mem_inst__0w_mem_10__31_0__10_));
OAI21X1 OAI21X1_1292 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf45), .B(w_mem_inst__abc_19396_new_n2863_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf42), .Y(w_mem_inst__abc_19396_new_n2864_));
OAI21X1 OAI21X1_1293 ( .A(w_mem_inst_w_mem_11__11_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf41), .C(w_mem_inst__abc_19396_new_n2864_), .Y(w_mem_inst__abc_19396_new_n2865_));
OAI21X1 OAI21X1_1294 ( .A(w_mem_inst__abc_19396_new_n2862_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf46), .C(w_mem_inst__abc_19396_new_n2865_), .Y(w_mem_inst__0w_mem_10__31_0__11_));
OAI21X1 OAI21X1_1295 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf44), .B(w_mem_inst__abc_19396_new_n2868_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf40), .Y(w_mem_inst__abc_19396_new_n2869_));
OAI21X1 OAI21X1_1296 ( .A(w_mem_inst_w_mem_11__12_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf39), .C(w_mem_inst__abc_19396_new_n2869_), .Y(w_mem_inst__abc_19396_new_n2870_));
OAI21X1 OAI21X1_1297 ( .A(w_mem_inst__abc_19396_new_n2867_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf45), .C(w_mem_inst__abc_19396_new_n2870_), .Y(w_mem_inst__0w_mem_10__31_0__12_));
OAI21X1 OAI21X1_1298 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf43), .B(w_mem_inst__abc_19396_new_n2873_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf38), .Y(w_mem_inst__abc_19396_new_n2874_));
OAI21X1 OAI21X1_1299 ( .A(w_mem_inst_w_mem_11__13_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf37), .C(w_mem_inst__abc_19396_new_n2874_), .Y(w_mem_inst__abc_19396_new_n2875_));
OAI21X1 OAI21X1_13 ( .A(_abc_15497_new_n878_), .B(_abc_15497_new_n889_), .C(_abc_15497_new_n879_), .Y(_abc_15497_new_n890_));
OAI21X1 OAI21X1_130 ( .A(_abc_15497_new_n1415_), .B(_abc_15497_new_n1423_), .C(_abc_15497_new_n1427_), .Y(_abc_15497_new_n1429_));
OAI21X1 OAI21X1_1300 ( .A(w_mem_inst__abc_19396_new_n2872_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf44), .C(w_mem_inst__abc_19396_new_n2875_), .Y(w_mem_inst__0w_mem_10__31_0__13_));
OAI21X1 OAI21X1_1301 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf42), .B(w_mem_inst__abc_19396_new_n2878_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf36), .Y(w_mem_inst__abc_19396_new_n2879_));
OAI21X1 OAI21X1_1302 ( .A(w_mem_inst_w_mem_11__14_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf35), .C(w_mem_inst__abc_19396_new_n2879_), .Y(w_mem_inst__abc_19396_new_n2880_));
OAI21X1 OAI21X1_1303 ( .A(w_mem_inst__abc_19396_new_n2877_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf43), .C(w_mem_inst__abc_19396_new_n2880_), .Y(w_mem_inst__0w_mem_10__31_0__14_));
OAI21X1 OAI21X1_1304 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf41), .B(w_mem_inst__abc_19396_new_n2883_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf34), .Y(w_mem_inst__abc_19396_new_n2884_));
OAI21X1 OAI21X1_1305 ( .A(w_mem_inst_w_mem_11__15_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf33), .C(w_mem_inst__abc_19396_new_n2884_), .Y(w_mem_inst__abc_19396_new_n2885_));
OAI21X1 OAI21X1_1306 ( .A(w_mem_inst__abc_19396_new_n2882_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf42), .C(w_mem_inst__abc_19396_new_n2885_), .Y(w_mem_inst__0w_mem_10__31_0__15_));
OAI21X1 OAI21X1_1307 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf40), .B(w_mem_inst__abc_19396_new_n2888_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf32), .Y(w_mem_inst__abc_19396_new_n2889_));
OAI21X1 OAI21X1_1308 ( .A(w_mem_inst_w_mem_11__16_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf31), .C(w_mem_inst__abc_19396_new_n2889_), .Y(w_mem_inst__abc_19396_new_n2890_));
OAI21X1 OAI21X1_1309 ( .A(w_mem_inst__abc_19396_new_n2887_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf41), .C(w_mem_inst__abc_19396_new_n2890_), .Y(w_mem_inst__0w_mem_10__31_0__16_));
OAI21X1 OAI21X1_131 ( .A(_abc_15497_new_n1423_), .B(_abc_15497_new_n1428_), .C(_abc_15497_new_n1429_), .Y(_abc_15497_new_n1430_));
OAI21X1 OAI21X1_1310 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf39), .B(w_mem_inst__abc_19396_new_n2893_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf30), .Y(w_mem_inst__abc_19396_new_n2894_));
OAI21X1 OAI21X1_1311 ( .A(w_mem_inst_w_mem_11__17_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf29), .C(w_mem_inst__abc_19396_new_n2894_), .Y(w_mem_inst__abc_19396_new_n2895_));
OAI21X1 OAI21X1_1312 ( .A(w_mem_inst__abc_19396_new_n2892_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf40), .C(w_mem_inst__abc_19396_new_n2895_), .Y(w_mem_inst__0w_mem_10__31_0__17_));
OAI21X1 OAI21X1_1313 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf38), .B(w_mem_inst__abc_19396_new_n2898_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf28), .Y(w_mem_inst__abc_19396_new_n2899_));
OAI21X1 OAI21X1_1314 ( .A(w_mem_inst_w_mem_11__18_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf27), .C(w_mem_inst__abc_19396_new_n2899_), .Y(w_mem_inst__abc_19396_new_n2900_));
OAI21X1 OAI21X1_1315 ( .A(w_mem_inst__abc_19396_new_n2897_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf39), .C(w_mem_inst__abc_19396_new_n2900_), .Y(w_mem_inst__0w_mem_10__31_0__18_));
OAI21X1 OAI21X1_1316 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf37), .B(w_mem_inst__abc_19396_new_n2903_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf26), .Y(w_mem_inst__abc_19396_new_n2904_));
OAI21X1 OAI21X1_1317 ( .A(w_mem_inst_w_mem_11__19_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf25), .C(w_mem_inst__abc_19396_new_n2904_), .Y(w_mem_inst__abc_19396_new_n2905_));
OAI21X1 OAI21X1_1318 ( .A(w_mem_inst__abc_19396_new_n2902_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf38), .C(w_mem_inst__abc_19396_new_n2905_), .Y(w_mem_inst__0w_mem_10__31_0__19_));
OAI21X1 OAI21X1_1319 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf36), .B(w_mem_inst__abc_19396_new_n2908_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf24), .Y(w_mem_inst__abc_19396_new_n2909_));
OAI21X1 OAI21X1_132 ( .A(_abc_15497_new_n1439_), .B(_abc_15497_new_n1434_), .C(digest_update_bF_buf3), .Y(_abc_15497_new_n1441_));
OAI21X1 OAI21X1_1320 ( .A(w_mem_inst_w_mem_11__20_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf23), .C(w_mem_inst__abc_19396_new_n2909_), .Y(w_mem_inst__abc_19396_new_n2910_));
OAI21X1 OAI21X1_1321 ( .A(w_mem_inst__abc_19396_new_n2907_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf37), .C(w_mem_inst__abc_19396_new_n2910_), .Y(w_mem_inst__0w_mem_10__31_0__20_));
OAI21X1 OAI21X1_1322 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf35), .B(w_mem_inst__abc_19396_new_n2913_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf22), .Y(w_mem_inst__abc_19396_new_n2914_));
OAI21X1 OAI21X1_1323 ( .A(w_mem_inst_w_mem_11__21_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf21), .C(w_mem_inst__abc_19396_new_n2914_), .Y(w_mem_inst__abc_19396_new_n2915_));
OAI21X1 OAI21X1_1324 ( .A(w_mem_inst__abc_19396_new_n2912_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf36), .C(w_mem_inst__abc_19396_new_n2915_), .Y(w_mem_inst__0w_mem_10__31_0__21_));
OAI21X1 OAI21X1_1325 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf34), .B(w_mem_inst__abc_19396_new_n2918_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf20), .Y(w_mem_inst__abc_19396_new_n2919_));
OAI21X1 OAI21X1_1326 ( .A(w_mem_inst_w_mem_11__22_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf19), .C(w_mem_inst__abc_19396_new_n2919_), .Y(w_mem_inst__abc_19396_new_n2920_));
OAI21X1 OAI21X1_1327 ( .A(w_mem_inst__abc_19396_new_n2917_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf35), .C(w_mem_inst__abc_19396_new_n2920_), .Y(w_mem_inst__0w_mem_10__31_0__22_));
OAI21X1 OAI21X1_1328 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf33), .B(w_mem_inst__abc_19396_new_n2923_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf18), .Y(w_mem_inst__abc_19396_new_n2924_));
OAI21X1 OAI21X1_1329 ( .A(w_mem_inst_w_mem_11__23_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf17), .C(w_mem_inst__abc_19396_new_n2924_), .Y(w_mem_inst__abc_19396_new_n2925_));
OAI21X1 OAI21X1_133 ( .A(_auto_iopadmap_cc_368_execute_22625_46_), .B(_abc_15497_new_n883__bF_buf1), .C(_abc_15497_new_n870__bF_buf1), .Y(_abc_15497_new_n1442_));
OAI21X1 OAI21X1_1330 ( .A(w_mem_inst__abc_19396_new_n2922_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf34), .C(w_mem_inst__abc_19396_new_n2925_), .Y(w_mem_inst__0w_mem_10__31_0__23_));
OAI21X1 OAI21X1_1331 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf32), .B(w_mem_inst__abc_19396_new_n2928_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf16), .Y(w_mem_inst__abc_19396_new_n2929_));
OAI21X1 OAI21X1_1332 ( .A(w_mem_inst_w_mem_11__24_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf15), .C(w_mem_inst__abc_19396_new_n2929_), .Y(w_mem_inst__abc_19396_new_n2930_));
OAI21X1 OAI21X1_1333 ( .A(w_mem_inst__abc_19396_new_n2927_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf33), .C(w_mem_inst__abc_19396_new_n2930_), .Y(w_mem_inst__0w_mem_10__31_0__24_));
OAI21X1 OAI21X1_1334 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf31), .B(w_mem_inst__abc_19396_new_n2933_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf14), .Y(w_mem_inst__abc_19396_new_n2934_));
OAI21X1 OAI21X1_1335 ( .A(w_mem_inst_w_mem_11__25_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf13), .C(w_mem_inst__abc_19396_new_n2934_), .Y(w_mem_inst__abc_19396_new_n2935_));
OAI21X1 OAI21X1_1336 ( .A(w_mem_inst__abc_19396_new_n2932_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf32), .C(w_mem_inst__abc_19396_new_n2935_), .Y(w_mem_inst__0w_mem_10__31_0__25_));
OAI21X1 OAI21X1_1337 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf30), .B(w_mem_inst__abc_19396_new_n2938_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf12), .Y(w_mem_inst__abc_19396_new_n2939_));
OAI21X1 OAI21X1_1338 ( .A(w_mem_inst_w_mem_11__26_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf11), .C(w_mem_inst__abc_19396_new_n2939_), .Y(w_mem_inst__abc_19396_new_n2940_));
OAI21X1 OAI21X1_1339 ( .A(w_mem_inst__abc_19396_new_n2937_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf31), .C(w_mem_inst__abc_19396_new_n2940_), .Y(w_mem_inst__0w_mem_10__31_0__26_));
OAI21X1 OAI21X1_134 ( .A(_abc_15497_new_n1440_), .B(_abc_15497_new_n1441_), .C(_abc_15497_new_n1442_), .Y(_0H3_reg_31_0__14_));
OAI21X1 OAI21X1_1340 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf29), .B(w_mem_inst__abc_19396_new_n2943_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf10), .Y(w_mem_inst__abc_19396_new_n2944_));
OAI21X1 OAI21X1_1341 ( .A(w_mem_inst_w_mem_11__27_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf9), .C(w_mem_inst__abc_19396_new_n2944_), .Y(w_mem_inst__abc_19396_new_n2945_));
OAI21X1 OAI21X1_1342 ( .A(w_mem_inst__abc_19396_new_n2942_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf30), .C(w_mem_inst__abc_19396_new_n2945_), .Y(w_mem_inst__0w_mem_10__31_0__27_));
OAI21X1 OAI21X1_1343 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf28), .B(w_mem_inst__abc_19396_new_n2948_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf8), .Y(w_mem_inst__abc_19396_new_n2949_));
OAI21X1 OAI21X1_1344 ( .A(w_mem_inst_w_mem_11__28_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf7), .C(w_mem_inst__abc_19396_new_n2949_), .Y(w_mem_inst__abc_19396_new_n2950_));
OAI21X1 OAI21X1_1345 ( .A(w_mem_inst__abc_19396_new_n2947_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf29), .C(w_mem_inst__abc_19396_new_n2950_), .Y(w_mem_inst__0w_mem_10__31_0__28_));
OAI21X1 OAI21X1_1346 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf27), .B(w_mem_inst__abc_19396_new_n2953_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf6), .Y(w_mem_inst__abc_19396_new_n2954_));
OAI21X1 OAI21X1_1347 ( .A(w_mem_inst_w_mem_11__29_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf5), .C(w_mem_inst__abc_19396_new_n2954_), .Y(w_mem_inst__abc_19396_new_n2955_));
OAI21X1 OAI21X1_1348 ( .A(w_mem_inst__abc_19396_new_n2952_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf28), .C(w_mem_inst__abc_19396_new_n2955_), .Y(w_mem_inst__0w_mem_10__31_0__29_));
OAI21X1 OAI21X1_1349 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf26), .B(w_mem_inst__abc_19396_new_n2958_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf4), .Y(w_mem_inst__abc_19396_new_n2959_));
OAI21X1 OAI21X1_135 ( .A(_abc_15497_new_n1435_), .B(_abc_15497_new_n1434_), .C(_abc_15497_new_n1436_), .Y(_abc_15497_new_n1445_));
OAI21X1 OAI21X1_1350 ( .A(w_mem_inst_w_mem_11__30_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf3), .C(w_mem_inst__abc_19396_new_n2959_), .Y(w_mem_inst__abc_19396_new_n2960_));
OAI21X1 OAI21X1_1351 ( .A(w_mem_inst__abc_19396_new_n2957_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf27), .C(w_mem_inst__abc_19396_new_n2960_), .Y(w_mem_inst__0w_mem_10__31_0__30_));
OAI21X1 OAI21X1_1352 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf25), .B(w_mem_inst__abc_19396_new_n2963_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf2), .Y(w_mem_inst__abc_19396_new_n2964_));
OAI21X1 OAI21X1_1353 ( .A(w_mem_inst_w_mem_11__31_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf1), .C(w_mem_inst__abc_19396_new_n2964_), .Y(w_mem_inst__abc_19396_new_n2965_));
OAI21X1 OAI21X1_1354 ( .A(w_mem_inst__abc_19396_new_n2962_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf26), .C(w_mem_inst__abc_19396_new_n2965_), .Y(w_mem_inst__0w_mem_10__31_0__31_));
OAI21X1 OAI21X1_1355 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf24), .B(w_mem_inst__abc_19396_new_n2968_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf0), .Y(w_mem_inst__abc_19396_new_n2969_));
OAI21X1 OAI21X1_1356 ( .A(w_mem_inst_w_mem_13__0_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf96), .C(w_mem_inst__abc_19396_new_n2969_), .Y(w_mem_inst__abc_19396_new_n2970_));
OAI21X1 OAI21X1_1357 ( .A(w_mem_inst__abc_19396_new_n2967_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf25), .C(w_mem_inst__abc_19396_new_n2970_), .Y(w_mem_inst__0w_mem_12__31_0__0_));
OAI21X1 OAI21X1_1358 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf23), .B(w_mem_inst__abc_19396_new_n2973_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf95), .Y(w_mem_inst__abc_19396_new_n2974_));
OAI21X1 OAI21X1_1359 ( .A(w_mem_inst_w_mem_13__1_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf94), .C(w_mem_inst__abc_19396_new_n2974_), .Y(w_mem_inst__abc_19396_new_n2975_));
OAI21X1 OAI21X1_136 ( .A(_abc_15497_new_n1453_), .B(_abc_15497_new_n1432_), .C(_abc_15497_new_n1454_), .Y(_abc_15497_new_n1455_));
OAI21X1 OAI21X1_1360 ( .A(w_mem_inst__abc_19396_new_n2972_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf24), .C(w_mem_inst__abc_19396_new_n2975_), .Y(w_mem_inst__0w_mem_12__31_0__1_));
OAI21X1 OAI21X1_1361 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf22), .B(w_mem_inst__abc_19396_new_n2978_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf93), .Y(w_mem_inst__abc_19396_new_n2979_));
OAI21X1 OAI21X1_1362 ( .A(w_mem_inst_w_mem_13__2_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf92), .C(w_mem_inst__abc_19396_new_n2979_), .Y(w_mem_inst__abc_19396_new_n2980_));
OAI21X1 OAI21X1_1363 ( .A(w_mem_inst__abc_19396_new_n2977_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf23), .C(w_mem_inst__abc_19396_new_n2980_), .Y(w_mem_inst__0w_mem_12__31_0__2_));
OAI21X1 OAI21X1_1364 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf21), .B(w_mem_inst__abc_19396_new_n2983_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf91), .Y(w_mem_inst__abc_19396_new_n2984_));
OAI21X1 OAI21X1_1365 ( .A(w_mem_inst_w_mem_13__3_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf90), .C(w_mem_inst__abc_19396_new_n2984_), .Y(w_mem_inst__abc_19396_new_n2985_));
OAI21X1 OAI21X1_1366 ( .A(w_mem_inst__abc_19396_new_n2982_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf22), .C(w_mem_inst__abc_19396_new_n2985_), .Y(w_mem_inst__0w_mem_12__31_0__3_));
OAI21X1 OAI21X1_1367 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf20), .B(w_mem_inst__abc_19396_new_n2988_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf89), .Y(w_mem_inst__abc_19396_new_n2989_));
OAI21X1 OAI21X1_1368 ( .A(w_mem_inst_w_mem_13__4_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf88), .C(w_mem_inst__abc_19396_new_n2989_), .Y(w_mem_inst__abc_19396_new_n2990_));
OAI21X1 OAI21X1_1369 ( .A(w_mem_inst__abc_19396_new_n2987_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf21), .C(w_mem_inst__abc_19396_new_n2990_), .Y(w_mem_inst__0w_mem_12__31_0__4_));
OAI21X1 OAI21X1_137 ( .A(_abc_15497_new_n1459_), .B(_abc_15497_new_n1362_), .C(_abc_15497_new_n1458_), .Y(_abc_15497_new_n1460_));
OAI21X1 OAI21X1_1370 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf19), .B(w_mem_inst__abc_19396_new_n2993_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf87), .Y(w_mem_inst__abc_19396_new_n2994_));
OAI21X1 OAI21X1_1371 ( .A(w_mem_inst_w_mem_13__5_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf86), .C(w_mem_inst__abc_19396_new_n2994_), .Y(w_mem_inst__abc_19396_new_n2995_));
OAI21X1 OAI21X1_1372 ( .A(w_mem_inst__abc_19396_new_n2992_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf20), .C(w_mem_inst__abc_19396_new_n2995_), .Y(w_mem_inst__0w_mem_12__31_0__5_));
OAI21X1 OAI21X1_1373 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf18), .B(w_mem_inst__abc_19396_new_n2998_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf85), .Y(w_mem_inst__abc_19396_new_n2999_));
OAI21X1 OAI21X1_1374 ( .A(w_mem_inst_w_mem_13__6_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf84), .C(w_mem_inst__abc_19396_new_n2999_), .Y(w_mem_inst__abc_19396_new_n3000_));
OAI21X1 OAI21X1_1375 ( .A(w_mem_inst__abc_19396_new_n2997_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf19), .C(w_mem_inst__abc_19396_new_n3000_), .Y(w_mem_inst__0w_mem_12__31_0__6_));
OAI21X1 OAI21X1_1376 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf17), .B(w_mem_inst__abc_19396_new_n3003_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf83), .Y(w_mem_inst__abc_19396_new_n3004_));
OAI21X1 OAI21X1_1377 ( .A(w_mem_inst_w_mem_13__7_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf82), .C(w_mem_inst__abc_19396_new_n3004_), .Y(w_mem_inst__abc_19396_new_n3005_));
OAI21X1 OAI21X1_1378 ( .A(w_mem_inst__abc_19396_new_n3002_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf18), .C(w_mem_inst__abc_19396_new_n3005_), .Y(w_mem_inst__0w_mem_12__31_0__7_));
OAI21X1 OAI21X1_1379 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf16), .B(w_mem_inst__abc_19396_new_n3008_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf81), .Y(w_mem_inst__abc_19396_new_n3009_));
OAI21X1 OAI21X1_138 ( .A(_abc_15497_new_n1473_), .B(_abc_15497_new_n1472_), .C(digest_update_bF_buf2), .Y(_abc_15497_new_n1474_));
OAI21X1 OAI21X1_1380 ( .A(w_mem_inst_w_mem_13__8_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf80), .C(w_mem_inst__abc_19396_new_n3009_), .Y(w_mem_inst__abc_19396_new_n3010_));
OAI21X1 OAI21X1_1381 ( .A(w_mem_inst__abc_19396_new_n3007_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf17), .C(w_mem_inst__abc_19396_new_n3010_), .Y(w_mem_inst__0w_mem_12__31_0__8_));
OAI21X1 OAI21X1_1382 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf15), .B(w_mem_inst__abc_19396_new_n3013_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf79), .Y(w_mem_inst__abc_19396_new_n3014_));
OAI21X1 OAI21X1_1383 ( .A(w_mem_inst_w_mem_13__9_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf78), .C(w_mem_inst__abc_19396_new_n3014_), .Y(w_mem_inst__abc_19396_new_n3015_));
OAI21X1 OAI21X1_1384 ( .A(w_mem_inst__abc_19396_new_n3012_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf16), .C(w_mem_inst__abc_19396_new_n3015_), .Y(w_mem_inst__0w_mem_12__31_0__9_));
OAI21X1 OAI21X1_1385 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf14), .B(w_mem_inst__abc_19396_new_n3018_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf77), .Y(w_mem_inst__abc_19396_new_n3019_));
OAI21X1 OAI21X1_1386 ( .A(w_mem_inst_w_mem_13__10_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf76), .C(w_mem_inst__abc_19396_new_n3019_), .Y(w_mem_inst__abc_19396_new_n3020_));
OAI21X1 OAI21X1_1387 ( .A(w_mem_inst__abc_19396_new_n3017_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf15), .C(w_mem_inst__abc_19396_new_n3020_), .Y(w_mem_inst__0w_mem_12__31_0__10_));
OAI21X1 OAI21X1_1388 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf13), .B(w_mem_inst__abc_19396_new_n3023_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf75), .Y(w_mem_inst__abc_19396_new_n3024_));
OAI21X1 OAI21X1_1389 ( .A(w_mem_inst_w_mem_13__11_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf74), .C(w_mem_inst__abc_19396_new_n3024_), .Y(w_mem_inst__abc_19396_new_n3025_));
OAI21X1 OAI21X1_139 ( .A(_auto_iopadmap_cc_368_execute_22625_49_), .B(_abc_15497_new_n883__bF_buf0), .C(_abc_15497_new_n870__bF_buf10), .Y(_abc_15497_new_n1475_));
OAI21X1 OAI21X1_1390 ( .A(w_mem_inst__abc_19396_new_n3022_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf14), .C(w_mem_inst__abc_19396_new_n3025_), .Y(w_mem_inst__0w_mem_12__31_0__11_));
OAI21X1 OAI21X1_1391 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf12), .B(w_mem_inst__abc_19396_new_n3028_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf73), .Y(w_mem_inst__abc_19396_new_n3029_));
OAI21X1 OAI21X1_1392 ( .A(w_mem_inst_w_mem_13__12_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf72), .C(w_mem_inst__abc_19396_new_n3029_), .Y(w_mem_inst__abc_19396_new_n3030_));
OAI21X1 OAI21X1_1393 ( .A(w_mem_inst__abc_19396_new_n3027_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf13), .C(w_mem_inst__abc_19396_new_n3030_), .Y(w_mem_inst__0w_mem_12__31_0__12_));
OAI21X1 OAI21X1_1394 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf11), .B(w_mem_inst__abc_19396_new_n3033_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf71), .Y(w_mem_inst__abc_19396_new_n3034_));
OAI21X1 OAI21X1_1395 ( .A(w_mem_inst_w_mem_13__13_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf70), .C(w_mem_inst__abc_19396_new_n3034_), .Y(w_mem_inst__abc_19396_new_n3035_));
OAI21X1 OAI21X1_1396 ( .A(w_mem_inst__abc_19396_new_n3032_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf12), .C(w_mem_inst__abc_19396_new_n3035_), .Y(w_mem_inst__0w_mem_12__31_0__13_));
OAI21X1 OAI21X1_1397 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf10), .B(w_mem_inst__abc_19396_new_n3038_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf69), .Y(w_mem_inst__abc_19396_new_n3039_));
OAI21X1 OAI21X1_1398 ( .A(w_mem_inst_w_mem_13__14_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf68), .C(w_mem_inst__abc_19396_new_n3039_), .Y(w_mem_inst__abc_19396_new_n3040_));
OAI21X1 OAI21X1_1399 ( .A(w_mem_inst__abc_19396_new_n3037_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf11), .C(w_mem_inst__abc_19396_new_n3040_), .Y(w_mem_inst__0w_mem_12__31_0__14_));
OAI21X1 OAI21X1_14 ( .A(_abc_15497_new_n887_), .B(_abc_15497_new_n848_), .C(_abc_15497_new_n891_), .Y(_abc_15497_new_n892_));
OAI21X1 OAI21X1_140 ( .A(_abc_15497_new_n1489_), .B(_abc_15497_new_n1482_), .C(digest_update_bF_buf1), .Y(_abc_15497_new_n1490_));
OAI21X1 OAI21X1_1400 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf9), .B(w_mem_inst__abc_19396_new_n3043_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf67), .Y(w_mem_inst__abc_19396_new_n3044_));
OAI21X1 OAI21X1_1401 ( .A(w_mem_inst_w_mem_13__15_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf66), .C(w_mem_inst__abc_19396_new_n3044_), .Y(w_mem_inst__abc_19396_new_n3045_));
OAI21X1 OAI21X1_1402 ( .A(w_mem_inst__abc_19396_new_n3042_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf10), .C(w_mem_inst__abc_19396_new_n3045_), .Y(w_mem_inst__0w_mem_12__31_0__15_));
OAI21X1 OAI21X1_1403 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf8), .B(w_mem_inst__abc_19396_new_n3048_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf65), .Y(w_mem_inst__abc_19396_new_n3049_));
OAI21X1 OAI21X1_1404 ( .A(w_mem_inst_w_mem_13__16_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf64), .C(w_mem_inst__abc_19396_new_n3049_), .Y(w_mem_inst__abc_19396_new_n3050_));
OAI21X1 OAI21X1_1405 ( .A(w_mem_inst__abc_19396_new_n3047_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf9), .C(w_mem_inst__abc_19396_new_n3050_), .Y(w_mem_inst__0w_mem_12__31_0__16_));
OAI21X1 OAI21X1_1406 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf7), .B(w_mem_inst__abc_19396_new_n3053_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf63), .Y(w_mem_inst__abc_19396_new_n3054_));
OAI21X1 OAI21X1_1407 ( .A(w_mem_inst_w_mem_13__17_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf62), .C(w_mem_inst__abc_19396_new_n3054_), .Y(w_mem_inst__abc_19396_new_n3055_));
OAI21X1 OAI21X1_1408 ( .A(w_mem_inst__abc_19396_new_n3052_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf8), .C(w_mem_inst__abc_19396_new_n3055_), .Y(w_mem_inst__0w_mem_12__31_0__17_));
OAI21X1 OAI21X1_1409 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf6), .B(w_mem_inst__abc_19396_new_n3058_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf61), .Y(w_mem_inst__abc_19396_new_n3059_));
OAI21X1 OAI21X1_141 ( .A(_abc_15497_new_n1498_), .B(_abc_15497_new_n1493_), .C(digest_update_bF_buf0), .Y(_abc_15497_new_n1500_));
OAI21X1 OAI21X1_1410 ( .A(w_mem_inst_w_mem_13__18_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf60), .C(w_mem_inst__abc_19396_new_n3059_), .Y(w_mem_inst__abc_19396_new_n3060_));
OAI21X1 OAI21X1_1411 ( .A(w_mem_inst__abc_19396_new_n3057_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf7), .C(w_mem_inst__abc_19396_new_n3060_), .Y(w_mem_inst__0w_mem_12__31_0__18_));
OAI21X1 OAI21X1_1412 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf5), .B(w_mem_inst__abc_19396_new_n3063_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf59), .Y(w_mem_inst__abc_19396_new_n3064_));
OAI21X1 OAI21X1_1413 ( .A(w_mem_inst_w_mem_13__19_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf58), .C(w_mem_inst__abc_19396_new_n3064_), .Y(w_mem_inst__abc_19396_new_n3065_));
OAI21X1 OAI21X1_1414 ( .A(w_mem_inst__abc_19396_new_n3062_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf6), .C(w_mem_inst__abc_19396_new_n3065_), .Y(w_mem_inst__0w_mem_12__31_0__19_));
OAI21X1 OAI21X1_1415 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf4), .B(w_mem_inst__abc_19396_new_n3068_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf57), .Y(w_mem_inst__abc_19396_new_n3069_));
OAI21X1 OAI21X1_1416 ( .A(w_mem_inst_w_mem_13__20_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf56), .C(w_mem_inst__abc_19396_new_n3069_), .Y(w_mem_inst__abc_19396_new_n3070_));
OAI21X1 OAI21X1_1417 ( .A(w_mem_inst__abc_19396_new_n3067_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf5), .C(w_mem_inst__abc_19396_new_n3070_), .Y(w_mem_inst__0w_mem_12__31_0__20_));
OAI21X1 OAI21X1_1418 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf3), .B(w_mem_inst__abc_19396_new_n3073_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf55), .Y(w_mem_inst__abc_19396_new_n3074_));
OAI21X1 OAI21X1_1419 ( .A(w_mem_inst_w_mem_13__21_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf54), .C(w_mem_inst__abc_19396_new_n3074_), .Y(w_mem_inst__abc_19396_new_n3075_));
OAI21X1 OAI21X1_142 ( .A(_abc_15497_new_n1478_), .B(_abc_15497_new_n1503_), .C(_abc_15497_new_n1505_), .Y(_abc_15497_new_n1506_));
OAI21X1 OAI21X1_1420 ( .A(w_mem_inst__abc_19396_new_n3072_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf4), .C(w_mem_inst__abc_19396_new_n3075_), .Y(w_mem_inst__0w_mem_12__31_0__21_));
OAI21X1 OAI21X1_1421 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf2), .B(w_mem_inst__abc_19396_new_n3078_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf53), .Y(w_mem_inst__abc_19396_new_n3079_));
OAI21X1 OAI21X1_1422 ( .A(w_mem_inst_w_mem_13__22_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf52), .C(w_mem_inst__abc_19396_new_n3079_), .Y(w_mem_inst__abc_19396_new_n3080_));
OAI21X1 OAI21X1_1423 ( .A(w_mem_inst__abc_19396_new_n3077_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf3), .C(w_mem_inst__abc_19396_new_n3080_), .Y(w_mem_inst__0w_mem_12__31_0__22_));
OAI21X1 OAI21X1_1424 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf1), .B(w_mem_inst__abc_19396_new_n3083_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf51), .Y(w_mem_inst__abc_19396_new_n3084_));
OAI21X1 OAI21X1_1425 ( .A(w_mem_inst_w_mem_13__23_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf50), .C(w_mem_inst__abc_19396_new_n3084_), .Y(w_mem_inst__abc_19396_new_n3085_));
OAI21X1 OAI21X1_1426 ( .A(w_mem_inst__abc_19396_new_n3082_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf2), .C(w_mem_inst__abc_19396_new_n3085_), .Y(w_mem_inst__0w_mem_12__31_0__23_));
OAI21X1 OAI21X1_1427 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf0), .B(w_mem_inst__abc_19396_new_n3088_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf49), .Y(w_mem_inst__abc_19396_new_n3089_));
OAI21X1 OAI21X1_1428 ( .A(w_mem_inst_w_mem_13__24_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf48), .C(w_mem_inst__abc_19396_new_n3089_), .Y(w_mem_inst__abc_19396_new_n3090_));
OAI21X1 OAI21X1_1429 ( .A(w_mem_inst__abc_19396_new_n3087_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf1), .C(w_mem_inst__abc_19396_new_n3090_), .Y(w_mem_inst__0w_mem_12__31_0__24_));
OAI21X1 OAI21X1_143 ( .A(_abc_15497_new_n1515_), .B(_abc_15497_new_n1507_), .C(digest_update_bF_buf8), .Y(_abc_15497_new_n1516_));
OAI21X1 OAI21X1_1430 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf60), .B(w_mem_inst__abc_19396_new_n3093_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf47), .Y(w_mem_inst__abc_19396_new_n3094_));
OAI21X1 OAI21X1_1431 ( .A(w_mem_inst_w_mem_13__25_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf46), .C(w_mem_inst__abc_19396_new_n3094_), .Y(w_mem_inst__abc_19396_new_n3095_));
OAI21X1 OAI21X1_1432 ( .A(w_mem_inst__abc_19396_new_n3092_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf0), .C(w_mem_inst__abc_19396_new_n3095_), .Y(w_mem_inst__0w_mem_12__31_0__25_));
OAI21X1 OAI21X1_1433 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf59), .B(w_mem_inst__abc_19396_new_n3098_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf45), .Y(w_mem_inst__abc_19396_new_n3099_));
OAI21X1 OAI21X1_1434 ( .A(w_mem_inst_w_mem_13__26_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf44), .C(w_mem_inst__abc_19396_new_n3099_), .Y(w_mem_inst__abc_19396_new_n3100_));
OAI21X1 OAI21X1_1435 ( .A(w_mem_inst__abc_19396_new_n3097_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf60), .C(w_mem_inst__abc_19396_new_n3100_), .Y(w_mem_inst__0w_mem_12__31_0__26_));
OAI21X1 OAI21X1_1436 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf58), .B(w_mem_inst__abc_19396_new_n3103_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf43), .Y(w_mem_inst__abc_19396_new_n3104_));
OAI21X1 OAI21X1_1437 ( .A(w_mem_inst_w_mem_13__27_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf42), .C(w_mem_inst__abc_19396_new_n3104_), .Y(w_mem_inst__abc_19396_new_n3105_));
OAI21X1 OAI21X1_1438 ( .A(w_mem_inst__abc_19396_new_n3102_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf59), .C(w_mem_inst__abc_19396_new_n3105_), .Y(w_mem_inst__0w_mem_12__31_0__27_));
OAI21X1 OAI21X1_1439 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf57), .B(w_mem_inst__abc_19396_new_n3108_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf41), .Y(w_mem_inst__abc_19396_new_n3109_));
OAI21X1 OAI21X1_144 ( .A(_auto_iopadmap_cc_368_execute_22625_52_), .B(_abc_15497_new_n883__bF_buf13), .C(_abc_15497_new_n870__bF_buf9), .Y(_abc_15497_new_n1517_));
OAI21X1 OAI21X1_1440 ( .A(w_mem_inst_w_mem_13__28_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf40), .C(w_mem_inst__abc_19396_new_n3109_), .Y(w_mem_inst__abc_19396_new_n3110_));
OAI21X1 OAI21X1_1441 ( .A(w_mem_inst__abc_19396_new_n3107_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf58), .C(w_mem_inst__abc_19396_new_n3110_), .Y(w_mem_inst__0w_mem_12__31_0__28_));
OAI21X1 OAI21X1_1442 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf56), .B(w_mem_inst__abc_19396_new_n3113_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf39), .Y(w_mem_inst__abc_19396_new_n3114_));
OAI21X1 OAI21X1_1443 ( .A(w_mem_inst_w_mem_13__29_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf38), .C(w_mem_inst__abc_19396_new_n3114_), .Y(w_mem_inst__abc_19396_new_n3115_));
OAI21X1 OAI21X1_1444 ( .A(w_mem_inst__abc_19396_new_n3112_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf57), .C(w_mem_inst__abc_19396_new_n3115_), .Y(w_mem_inst__0w_mem_12__31_0__29_));
OAI21X1 OAI21X1_1445 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf55), .B(w_mem_inst__abc_19396_new_n3118_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf37), .Y(w_mem_inst__abc_19396_new_n3119_));
OAI21X1 OAI21X1_1446 ( .A(w_mem_inst_w_mem_13__30_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf36), .C(w_mem_inst__abc_19396_new_n3119_), .Y(w_mem_inst__abc_19396_new_n3120_));
OAI21X1 OAI21X1_1447 ( .A(w_mem_inst__abc_19396_new_n3117_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf56), .C(w_mem_inst__abc_19396_new_n3120_), .Y(w_mem_inst__0w_mem_12__31_0__30_));
OAI21X1 OAI21X1_1448 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf54), .B(w_mem_inst__abc_19396_new_n3123_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf35), .Y(w_mem_inst__abc_19396_new_n3124_));
OAI21X1 OAI21X1_1449 ( .A(w_mem_inst_w_mem_13__31_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf34), .C(w_mem_inst__abc_19396_new_n3124_), .Y(w_mem_inst__abc_19396_new_n3125_));
OAI21X1 OAI21X1_145 ( .A(_abc_15497_new_n1516_), .B(_abc_15497_new_n1514_), .C(_abc_15497_new_n1517_), .Y(_0H3_reg_31_0__20_));
OAI21X1 OAI21X1_1450 ( .A(w_mem_inst__abc_19396_new_n3122_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf55), .C(w_mem_inst__abc_19396_new_n3125_), .Y(w_mem_inst__0w_mem_12__31_0__31_));
OAI21X1 OAI21X1_1451 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf53), .B(w_mem_inst__abc_19396_new_n3128_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf33), .Y(w_mem_inst__abc_19396_new_n3129_));
OAI21X1 OAI21X1_1452 ( .A(w_mem_inst_w_mem_12__0_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf32), .C(w_mem_inst__abc_19396_new_n3129_), .Y(w_mem_inst__abc_19396_new_n3130_));
OAI21X1 OAI21X1_1453 ( .A(w_mem_inst__abc_19396_new_n3127_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf54), .C(w_mem_inst__abc_19396_new_n3130_), .Y(w_mem_inst__0w_mem_11__31_0__0_));
OAI21X1 OAI21X1_1454 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf52), .B(w_mem_inst__abc_19396_new_n3133_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf31), .Y(w_mem_inst__abc_19396_new_n3134_));
OAI21X1 OAI21X1_1455 ( .A(w_mem_inst_w_mem_12__1_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf30), .C(w_mem_inst__abc_19396_new_n3134_), .Y(w_mem_inst__abc_19396_new_n3135_));
OAI21X1 OAI21X1_1456 ( .A(w_mem_inst__abc_19396_new_n3132_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf53), .C(w_mem_inst__abc_19396_new_n3135_), .Y(w_mem_inst__0w_mem_11__31_0__1_));
OAI21X1 OAI21X1_1457 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf51), .B(w_mem_inst__abc_19396_new_n3138_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf29), .Y(w_mem_inst__abc_19396_new_n3139_));
OAI21X1 OAI21X1_1458 ( .A(w_mem_inst_w_mem_12__2_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf28), .C(w_mem_inst__abc_19396_new_n3139_), .Y(w_mem_inst__abc_19396_new_n3140_));
OAI21X1 OAI21X1_1459 ( .A(w_mem_inst__abc_19396_new_n3137_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf52), .C(w_mem_inst__abc_19396_new_n3140_), .Y(w_mem_inst__0w_mem_11__31_0__2_));
OAI21X1 OAI21X1_146 ( .A(_abc_15497_new_n1509_), .B(_abc_15497_new_n1507_), .C(_abc_15497_new_n1519_), .Y(_abc_15497_new_n1520_));
OAI21X1 OAI21X1_1460 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf50), .B(w_mem_inst__abc_19396_new_n3143_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf27), .Y(w_mem_inst__abc_19396_new_n3144_));
OAI21X1 OAI21X1_1461 ( .A(w_mem_inst_w_mem_12__3_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf26), .C(w_mem_inst__abc_19396_new_n3144_), .Y(w_mem_inst__abc_19396_new_n3145_));
OAI21X1 OAI21X1_1462 ( .A(w_mem_inst__abc_19396_new_n3142_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf51), .C(w_mem_inst__abc_19396_new_n3145_), .Y(w_mem_inst__0w_mem_11__31_0__3_));
OAI21X1 OAI21X1_1463 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf49), .B(w_mem_inst__abc_19396_new_n3148_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf25), .Y(w_mem_inst__abc_19396_new_n3149_));
OAI21X1 OAI21X1_1464 ( .A(w_mem_inst_w_mem_12__4_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf24), .C(w_mem_inst__abc_19396_new_n3149_), .Y(w_mem_inst__abc_19396_new_n3150_));
OAI21X1 OAI21X1_1465 ( .A(w_mem_inst__abc_19396_new_n3147_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf50), .C(w_mem_inst__abc_19396_new_n3150_), .Y(w_mem_inst__0w_mem_11__31_0__4_));
OAI21X1 OAI21X1_1466 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf48), .B(w_mem_inst__abc_19396_new_n3153_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf23), .Y(w_mem_inst__abc_19396_new_n3154_));
OAI21X1 OAI21X1_1467 ( .A(w_mem_inst_w_mem_12__5_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf22), .C(w_mem_inst__abc_19396_new_n3154_), .Y(w_mem_inst__abc_19396_new_n3155_));
OAI21X1 OAI21X1_1468 ( .A(w_mem_inst__abc_19396_new_n3152_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf49), .C(w_mem_inst__abc_19396_new_n3155_), .Y(w_mem_inst__0w_mem_11__31_0__5_));
OAI21X1 OAI21X1_1469 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf47), .B(w_mem_inst__abc_19396_new_n3158_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf21), .Y(w_mem_inst__abc_19396_new_n3159_));
OAI21X1 OAI21X1_147 ( .A(_auto_iopadmap_cc_368_execute_22625_53_), .B(_abc_15497_new_n883__bF_buf12), .C(_abc_15497_new_n870__bF_buf8), .Y(_abc_15497_new_n1526_));
OAI21X1 OAI21X1_1470 ( .A(w_mem_inst_w_mem_12__6_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf20), .C(w_mem_inst__abc_19396_new_n3159_), .Y(w_mem_inst__abc_19396_new_n3160_));
OAI21X1 OAI21X1_1471 ( .A(w_mem_inst__abc_19396_new_n3157_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf48), .C(w_mem_inst__abc_19396_new_n3160_), .Y(w_mem_inst__0w_mem_11__31_0__6_));
OAI21X1 OAI21X1_1472 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf46), .B(w_mem_inst__abc_19396_new_n3163_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf19), .Y(w_mem_inst__abc_19396_new_n3164_));
OAI21X1 OAI21X1_1473 ( .A(w_mem_inst_w_mem_12__7_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf18), .C(w_mem_inst__abc_19396_new_n3164_), .Y(w_mem_inst__abc_19396_new_n3165_));
OAI21X1 OAI21X1_1474 ( .A(w_mem_inst__abc_19396_new_n3162_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf47), .C(w_mem_inst__abc_19396_new_n3165_), .Y(w_mem_inst__0w_mem_11__31_0__7_));
OAI21X1 OAI21X1_1475 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf45), .B(w_mem_inst__abc_19396_new_n3168_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf17), .Y(w_mem_inst__abc_19396_new_n3169_));
OAI21X1 OAI21X1_1476 ( .A(w_mem_inst_w_mem_12__8_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf16), .C(w_mem_inst__abc_19396_new_n3169_), .Y(w_mem_inst__abc_19396_new_n3170_));
OAI21X1 OAI21X1_1477 ( .A(w_mem_inst__abc_19396_new_n3167_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf46), .C(w_mem_inst__abc_19396_new_n3170_), .Y(w_mem_inst__0w_mem_11__31_0__8_));
OAI21X1 OAI21X1_1478 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf44), .B(w_mem_inst__abc_19396_new_n3173_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf15), .Y(w_mem_inst__abc_19396_new_n3174_));
OAI21X1 OAI21X1_1479 ( .A(w_mem_inst_w_mem_12__9_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf14), .C(w_mem_inst__abc_19396_new_n3174_), .Y(w_mem_inst__abc_19396_new_n3175_));
OAI21X1 OAI21X1_148 ( .A(_abc_15497_new_n870__bF_buf7), .B(_abc_15497_new_n1525_), .C(_abc_15497_new_n1526_), .Y(_0H3_reg_31_0__21_));
OAI21X1 OAI21X1_1480 ( .A(w_mem_inst__abc_19396_new_n3172_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf45), .C(w_mem_inst__abc_19396_new_n3175_), .Y(w_mem_inst__0w_mem_11__31_0__9_));
OAI21X1 OAI21X1_1481 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf43), .B(w_mem_inst__abc_19396_new_n3178_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf13), .Y(w_mem_inst__abc_19396_new_n3179_));
OAI21X1 OAI21X1_1482 ( .A(w_mem_inst_w_mem_12__10_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf12), .C(w_mem_inst__abc_19396_new_n3179_), .Y(w_mem_inst__abc_19396_new_n3180_));
OAI21X1 OAI21X1_1483 ( .A(w_mem_inst__abc_19396_new_n3177_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf44), .C(w_mem_inst__abc_19396_new_n3180_), .Y(w_mem_inst__0w_mem_11__31_0__10_));
OAI21X1 OAI21X1_1484 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf42), .B(w_mem_inst__abc_19396_new_n3183_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf11), .Y(w_mem_inst__abc_19396_new_n3184_));
OAI21X1 OAI21X1_1485 ( .A(w_mem_inst_w_mem_12__11_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf10), .C(w_mem_inst__abc_19396_new_n3184_), .Y(w_mem_inst__abc_19396_new_n3185_));
OAI21X1 OAI21X1_1486 ( .A(w_mem_inst__abc_19396_new_n3182_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf43), .C(w_mem_inst__abc_19396_new_n3185_), .Y(w_mem_inst__0w_mem_11__31_0__11_));
OAI21X1 OAI21X1_1487 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf41), .B(w_mem_inst__abc_19396_new_n3188_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf9), .Y(w_mem_inst__abc_19396_new_n3189_));
OAI21X1 OAI21X1_1488 ( .A(w_mem_inst_w_mem_12__12_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf8), .C(w_mem_inst__abc_19396_new_n3189_), .Y(w_mem_inst__abc_19396_new_n3190_));
OAI21X1 OAI21X1_1489 ( .A(w_mem_inst__abc_19396_new_n3187_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf42), .C(w_mem_inst__abc_19396_new_n3190_), .Y(w_mem_inst__0w_mem_11__31_0__12_));
OAI21X1 OAI21X1_149 ( .A(_abc_15497_new_n1521_), .B(_abc_15497_new_n1519_), .C(_abc_15497_new_n1523_), .Y(_abc_15497_new_n1534_));
OAI21X1 OAI21X1_1490 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf40), .B(w_mem_inst__abc_19396_new_n3193_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf7), .Y(w_mem_inst__abc_19396_new_n3194_));
OAI21X1 OAI21X1_1491 ( .A(w_mem_inst_w_mem_12__13_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf6), .C(w_mem_inst__abc_19396_new_n3194_), .Y(w_mem_inst__abc_19396_new_n3195_));
OAI21X1 OAI21X1_1492 ( .A(w_mem_inst__abc_19396_new_n3192_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf41), .C(w_mem_inst__abc_19396_new_n3195_), .Y(w_mem_inst__0w_mem_11__31_0__13_));
OAI21X1 OAI21X1_1493 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf39), .B(w_mem_inst__abc_19396_new_n3198_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf5), .Y(w_mem_inst__abc_19396_new_n3199_));
OAI21X1 OAI21X1_1494 ( .A(w_mem_inst_w_mem_12__14_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf4), .C(w_mem_inst__abc_19396_new_n3199_), .Y(w_mem_inst__abc_19396_new_n3200_));
OAI21X1 OAI21X1_1495 ( .A(w_mem_inst__abc_19396_new_n3197_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf40), .C(w_mem_inst__abc_19396_new_n3200_), .Y(w_mem_inst__0w_mem_11__31_0__14_));
OAI21X1 OAI21X1_1496 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf38), .B(w_mem_inst__abc_19396_new_n3203_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf3), .Y(w_mem_inst__abc_19396_new_n3204_));
OAI21X1 OAI21X1_1497 ( .A(w_mem_inst_w_mem_12__15_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf2), .C(w_mem_inst__abc_19396_new_n3204_), .Y(w_mem_inst__abc_19396_new_n3205_));
OAI21X1 OAI21X1_1498 ( .A(w_mem_inst__abc_19396_new_n3202_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf39), .C(w_mem_inst__abc_19396_new_n3205_), .Y(w_mem_inst__0w_mem_11__31_0__15_));
OAI21X1 OAI21X1_1499 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf37), .B(w_mem_inst__abc_19396_new_n3208_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf1), .Y(w_mem_inst__abc_19396_new_n3209_));
OAI21X1 OAI21X1_15 ( .A(_abc_15497_new_n892_), .B(_abc_15497_new_n896_), .C(_abc_15497_new_n897_), .Y(_abc_15497_new_n898_));
OAI21X1 OAI21X1_150 ( .A(_abc_15497_new_n1533_), .B(_abc_15497_new_n1536_), .C(digest_update_bF_buf7), .Y(_abc_15497_new_n1538_));
OAI21X1 OAI21X1_1500 ( .A(w_mem_inst_w_mem_12__16_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf0), .C(w_mem_inst__abc_19396_new_n3209_), .Y(w_mem_inst__abc_19396_new_n3210_));
OAI21X1 OAI21X1_1501 ( .A(w_mem_inst__abc_19396_new_n3207_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf38), .C(w_mem_inst__abc_19396_new_n3210_), .Y(w_mem_inst__0w_mem_11__31_0__16_));
OAI21X1 OAI21X1_1502 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf36), .B(w_mem_inst__abc_19396_new_n3213_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf96), .Y(w_mem_inst__abc_19396_new_n3214_));
OAI21X1 OAI21X1_1503 ( .A(w_mem_inst_w_mem_12__17_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf95), .C(w_mem_inst__abc_19396_new_n3214_), .Y(w_mem_inst__abc_19396_new_n3215_));
OAI21X1 OAI21X1_1504 ( .A(w_mem_inst__abc_19396_new_n3212_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf37), .C(w_mem_inst__abc_19396_new_n3215_), .Y(w_mem_inst__0w_mem_11__31_0__17_));
OAI21X1 OAI21X1_1505 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf35), .B(w_mem_inst__abc_19396_new_n3218_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf94), .Y(w_mem_inst__abc_19396_new_n3219_));
OAI21X1 OAI21X1_1506 ( .A(w_mem_inst_w_mem_12__18_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf93), .C(w_mem_inst__abc_19396_new_n3219_), .Y(w_mem_inst__abc_19396_new_n3220_));
OAI21X1 OAI21X1_1507 ( .A(w_mem_inst__abc_19396_new_n3217_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf36), .C(w_mem_inst__abc_19396_new_n3220_), .Y(w_mem_inst__0w_mem_11__31_0__18_));
OAI21X1 OAI21X1_1508 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf34), .B(w_mem_inst__abc_19396_new_n3223_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf92), .Y(w_mem_inst__abc_19396_new_n3224_));
OAI21X1 OAI21X1_1509 ( .A(w_mem_inst_w_mem_12__19_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf91), .C(w_mem_inst__abc_19396_new_n3224_), .Y(w_mem_inst__abc_19396_new_n3225_));
OAI21X1 OAI21X1_151 ( .A(_abc_15497_new_n1546_), .B(_abc_15497_new_n1542_), .C(digest_update_bF_buf6), .Y(_abc_15497_new_n1548_));
OAI21X1 OAI21X1_1510 ( .A(w_mem_inst__abc_19396_new_n3222_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf35), .C(w_mem_inst__abc_19396_new_n3225_), .Y(w_mem_inst__0w_mem_11__31_0__19_));
OAI21X1 OAI21X1_1511 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf33), .B(w_mem_inst__abc_19396_new_n3228_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf90), .Y(w_mem_inst__abc_19396_new_n3229_));
OAI21X1 OAI21X1_1512 ( .A(w_mem_inst_w_mem_12__20_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf89), .C(w_mem_inst__abc_19396_new_n3229_), .Y(w_mem_inst__abc_19396_new_n3230_));
OAI21X1 OAI21X1_1513 ( .A(w_mem_inst__abc_19396_new_n3227_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf34), .C(w_mem_inst__abc_19396_new_n3230_), .Y(w_mem_inst__0w_mem_11__31_0__20_));
OAI21X1 OAI21X1_1514 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf32), .B(w_mem_inst__abc_19396_new_n3233_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf88), .Y(w_mem_inst__abc_19396_new_n3234_));
OAI21X1 OAI21X1_1515 ( .A(w_mem_inst_w_mem_12__21_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf87), .C(w_mem_inst__abc_19396_new_n3234_), .Y(w_mem_inst__abc_19396_new_n3235_));
OAI21X1 OAI21X1_1516 ( .A(w_mem_inst__abc_19396_new_n3232_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf33), .C(w_mem_inst__abc_19396_new_n3235_), .Y(w_mem_inst__0w_mem_11__31_0__21_));
OAI21X1 OAI21X1_1517 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf31), .B(w_mem_inst__abc_19396_new_n3238_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf86), .Y(w_mem_inst__abc_19396_new_n3239_));
OAI21X1 OAI21X1_1518 ( .A(w_mem_inst_w_mem_12__22_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf85), .C(w_mem_inst__abc_19396_new_n3239_), .Y(w_mem_inst__abc_19396_new_n3240_));
OAI21X1 OAI21X1_1519 ( .A(w_mem_inst__abc_19396_new_n3237_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf32), .C(w_mem_inst__abc_19396_new_n3240_), .Y(w_mem_inst__0w_mem_11__31_0__22_));
OAI21X1 OAI21X1_152 ( .A(_abc_15497_new_n1528_), .B(_abc_15497_new_n1530_), .C(_abc_15497_new_n1545_), .Y(_abc_15497_new_n1552_));
OAI21X1 OAI21X1_1520 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf30), .B(w_mem_inst__abc_19396_new_n3243_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf84), .Y(w_mem_inst__abc_19396_new_n3244_));
OAI21X1 OAI21X1_1521 ( .A(w_mem_inst_w_mem_12__23_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf83), .C(w_mem_inst__abc_19396_new_n3244_), .Y(w_mem_inst__abc_19396_new_n3245_));
OAI21X1 OAI21X1_1522 ( .A(w_mem_inst__abc_19396_new_n3242_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf31), .C(w_mem_inst__abc_19396_new_n3245_), .Y(w_mem_inst__0w_mem_11__31_0__23_));
OAI21X1 OAI21X1_1523 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf29), .B(w_mem_inst__abc_19396_new_n3248_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf82), .Y(w_mem_inst__abc_19396_new_n3249_));
OAI21X1 OAI21X1_1524 ( .A(w_mem_inst_w_mem_12__24_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf81), .C(w_mem_inst__abc_19396_new_n3249_), .Y(w_mem_inst__abc_19396_new_n3250_));
OAI21X1 OAI21X1_1525 ( .A(w_mem_inst__abc_19396_new_n3247_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf30), .C(w_mem_inst__abc_19396_new_n3250_), .Y(w_mem_inst__0w_mem_11__31_0__24_));
OAI21X1 OAI21X1_1526 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf28), .B(w_mem_inst__abc_19396_new_n3253_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf80), .Y(w_mem_inst__abc_19396_new_n3254_));
OAI21X1 OAI21X1_1527 ( .A(w_mem_inst_w_mem_12__25_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf79), .C(w_mem_inst__abc_19396_new_n3254_), .Y(w_mem_inst__abc_19396_new_n3255_));
OAI21X1 OAI21X1_1528 ( .A(w_mem_inst__abc_19396_new_n3252_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf29), .C(w_mem_inst__abc_19396_new_n3255_), .Y(w_mem_inst__0w_mem_11__31_0__25_));
OAI21X1 OAI21X1_1529 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf27), .B(w_mem_inst__abc_19396_new_n3258_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf78), .Y(w_mem_inst__abc_19396_new_n3259_));
OAI21X1 OAI21X1_153 ( .A(_abc_15497_new_n1555_), .B(_abc_15497_new_n1551_), .C(_abc_15497_new_n1554_), .Y(_abc_15497_new_n1556_));
OAI21X1 OAI21X1_1530 ( .A(w_mem_inst_w_mem_12__26_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf77), .C(w_mem_inst__abc_19396_new_n3259_), .Y(w_mem_inst__abc_19396_new_n3260_));
OAI21X1 OAI21X1_1531 ( .A(w_mem_inst__abc_19396_new_n3257_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf28), .C(w_mem_inst__abc_19396_new_n3260_), .Y(w_mem_inst__0w_mem_11__31_0__26_));
OAI21X1 OAI21X1_1532 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf26), .B(w_mem_inst__abc_19396_new_n3263_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf76), .Y(w_mem_inst__abc_19396_new_n3264_));
OAI21X1 OAI21X1_1533 ( .A(w_mem_inst_w_mem_12__27_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf75), .C(w_mem_inst__abc_19396_new_n3264_), .Y(w_mem_inst__abc_19396_new_n3265_));
OAI21X1 OAI21X1_1534 ( .A(w_mem_inst__abc_19396_new_n3262_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf27), .C(w_mem_inst__abc_19396_new_n3265_), .Y(w_mem_inst__0w_mem_11__31_0__27_));
OAI21X1 OAI21X1_1535 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf25), .B(w_mem_inst__abc_19396_new_n3268_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf74), .Y(w_mem_inst__abc_19396_new_n3269_));
OAI21X1 OAI21X1_1536 ( .A(w_mem_inst_w_mem_12__28_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf73), .C(w_mem_inst__abc_19396_new_n3269_), .Y(w_mem_inst__abc_19396_new_n3270_));
OAI21X1 OAI21X1_1537 ( .A(w_mem_inst__abc_19396_new_n3267_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf26), .C(w_mem_inst__abc_19396_new_n3270_), .Y(w_mem_inst__0w_mem_11__31_0__28_));
OAI21X1 OAI21X1_1538 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf24), .B(w_mem_inst__abc_19396_new_n3273_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf72), .Y(w_mem_inst__abc_19396_new_n3274_));
OAI21X1 OAI21X1_1539 ( .A(w_mem_inst_w_mem_12__29_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf71), .C(w_mem_inst__abc_19396_new_n3274_), .Y(w_mem_inst__abc_19396_new_n3275_));
OAI21X1 OAI21X1_154 ( .A(_abc_15497_new_n1566_), .B(_abc_15497_new_n1559_), .C(digest_update_bF_buf5), .Y(_abc_15497_new_n1567_));
OAI21X1 OAI21X1_1540 ( .A(w_mem_inst__abc_19396_new_n3272_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf25), .C(w_mem_inst__abc_19396_new_n3275_), .Y(w_mem_inst__0w_mem_11__31_0__29_));
OAI21X1 OAI21X1_1541 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf23), .B(w_mem_inst__abc_19396_new_n3278_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf70), .Y(w_mem_inst__abc_19396_new_n3279_));
OAI21X1 OAI21X1_1542 ( .A(w_mem_inst_w_mem_12__30_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf69), .C(w_mem_inst__abc_19396_new_n3279_), .Y(w_mem_inst__abc_19396_new_n3280_));
OAI21X1 OAI21X1_1543 ( .A(w_mem_inst__abc_19396_new_n3277_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf24), .C(w_mem_inst__abc_19396_new_n3280_), .Y(w_mem_inst__0w_mem_11__31_0__30_));
OAI21X1 OAI21X1_1544 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf22), .B(w_mem_inst__abc_19396_new_n3283_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf68), .Y(w_mem_inst__abc_19396_new_n3284_));
OAI21X1 OAI21X1_1545 ( .A(w_mem_inst_w_mem_12__31_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf67), .C(w_mem_inst__abc_19396_new_n3284_), .Y(w_mem_inst__abc_19396_new_n3285_));
OAI21X1 OAI21X1_1546 ( .A(w_mem_inst__abc_19396_new_n3282_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf23), .C(w_mem_inst__abc_19396_new_n3285_), .Y(w_mem_inst__0w_mem_11__31_0__31_));
OAI21X1 OAI21X1_1547 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf21), .B(w_mem_inst__abc_19396_new_n3287_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf66), .Y(w_mem_inst__abc_19396_new_n3288_));
OAI21X1 OAI21X1_1548 ( .A(w_mem_inst_w_mem_8__0_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf65), .C(w_mem_inst__abc_19396_new_n3288_), .Y(w_mem_inst__abc_19396_new_n3289_));
OAI21X1 OAI21X1_1549 ( .A(w_mem_inst__abc_19396_new_n1609_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf22), .C(w_mem_inst__abc_19396_new_n3289_), .Y(w_mem_inst__0w_mem_7__31_0__0_));
OAI21X1 OAI21X1_155 ( .A(_abc_15497_new_n1550_), .B(_abc_15497_new_n1562_), .C(_abc_15497_new_n1575_), .Y(_abc_15497_new_n1576_));
OAI21X1 OAI21X1_1550 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf20), .B(w_mem_inst__abc_19396_new_n3291_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf64), .Y(w_mem_inst__abc_19396_new_n3292_));
OAI21X1 OAI21X1_1551 ( .A(w_mem_inst_w_mem_8__1_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf63), .C(w_mem_inst__abc_19396_new_n3292_), .Y(w_mem_inst__abc_19396_new_n3293_));
OAI21X1 OAI21X1_1552 ( .A(w_mem_inst__abc_19396_new_n1651_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf21), .C(w_mem_inst__abc_19396_new_n3293_), .Y(w_mem_inst__0w_mem_7__31_0__1_));
OAI21X1 OAI21X1_1553 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf19), .B(w_mem_inst__abc_19396_new_n3295_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf62), .Y(w_mem_inst__abc_19396_new_n3296_));
OAI21X1 OAI21X1_1554 ( .A(w_mem_inst_w_mem_8__2_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf61), .C(w_mem_inst__abc_19396_new_n3296_), .Y(w_mem_inst__abc_19396_new_n3297_));
OAI21X1 OAI21X1_1555 ( .A(w_mem_inst__abc_19396_new_n1676_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf20), .C(w_mem_inst__abc_19396_new_n3297_), .Y(w_mem_inst__0w_mem_7__31_0__2_));
OAI21X1 OAI21X1_1556 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf18), .B(w_mem_inst__abc_19396_new_n3299_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf60), .Y(w_mem_inst__abc_19396_new_n3300_));
OAI21X1 OAI21X1_1557 ( .A(w_mem_inst_w_mem_8__3_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf59), .C(w_mem_inst__abc_19396_new_n3300_), .Y(w_mem_inst__abc_19396_new_n3301_));
OAI21X1 OAI21X1_1558 ( .A(w_mem_inst__abc_19396_new_n1701_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf19), .C(w_mem_inst__abc_19396_new_n3301_), .Y(w_mem_inst__0w_mem_7__31_0__3_));
OAI21X1 OAI21X1_1559 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf17), .B(w_mem_inst__abc_19396_new_n3303_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf58), .Y(w_mem_inst__abc_19396_new_n3304_));
OAI21X1 OAI21X1_156 ( .A(_abc_15497_new_n1563_), .B(_abc_15497_new_n1570_), .C(_abc_15497_new_n1574_), .Y(_abc_15497_new_n1577_));
OAI21X1 OAI21X1_1560 ( .A(w_mem_inst_w_mem_8__4_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf57), .C(w_mem_inst__abc_19396_new_n3304_), .Y(w_mem_inst__abc_19396_new_n3305_));
OAI21X1 OAI21X1_1561 ( .A(w_mem_inst__abc_19396_new_n1726_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf18), .C(w_mem_inst__abc_19396_new_n3305_), .Y(w_mem_inst__0w_mem_7__31_0__4_));
OAI21X1 OAI21X1_1562 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf16), .B(w_mem_inst__abc_19396_new_n3307_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf56), .Y(w_mem_inst__abc_19396_new_n3308_));
OAI21X1 OAI21X1_1563 ( .A(w_mem_inst_w_mem_8__5_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf55), .C(w_mem_inst__abc_19396_new_n3308_), .Y(w_mem_inst__abc_19396_new_n3309_));
OAI21X1 OAI21X1_1564 ( .A(w_mem_inst__abc_19396_new_n1751_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf17), .C(w_mem_inst__abc_19396_new_n3309_), .Y(w_mem_inst__0w_mem_7__31_0__5_));
OAI21X1 OAI21X1_1565 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf15), .B(w_mem_inst__abc_19396_new_n3311_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf54), .Y(w_mem_inst__abc_19396_new_n3312_));
OAI21X1 OAI21X1_1566 ( .A(w_mem_inst_w_mem_8__6_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf53), .C(w_mem_inst__abc_19396_new_n3312_), .Y(w_mem_inst__abc_19396_new_n3313_));
OAI21X1 OAI21X1_1567 ( .A(w_mem_inst__abc_19396_new_n1776_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf16), .C(w_mem_inst__abc_19396_new_n3313_), .Y(w_mem_inst__0w_mem_7__31_0__6_));
OAI21X1 OAI21X1_1568 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf14), .B(w_mem_inst__abc_19396_new_n3315_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf52), .Y(w_mem_inst__abc_19396_new_n3316_));
OAI21X1 OAI21X1_1569 ( .A(w_mem_inst_w_mem_8__7_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf51), .C(w_mem_inst__abc_19396_new_n3316_), .Y(w_mem_inst__abc_19396_new_n3317_));
OAI21X1 OAI21X1_157 ( .A(_abc_15497_new_n1570_), .B(_abc_15497_new_n1576_), .C(_abc_15497_new_n1577_), .Y(_abc_15497_new_n1578_));
OAI21X1 OAI21X1_1570 ( .A(w_mem_inst__abc_19396_new_n1801_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf15), .C(w_mem_inst__abc_19396_new_n3317_), .Y(w_mem_inst__0w_mem_7__31_0__7_));
OAI21X1 OAI21X1_1571 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf13), .B(w_mem_inst__abc_19396_new_n3319_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf50), .Y(w_mem_inst__abc_19396_new_n3320_));
OAI21X1 OAI21X1_1572 ( .A(w_mem_inst_w_mem_8__8_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf49), .C(w_mem_inst__abc_19396_new_n3320_), .Y(w_mem_inst__abc_19396_new_n3321_));
OAI21X1 OAI21X1_1573 ( .A(w_mem_inst__abc_19396_new_n1826_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf14), .C(w_mem_inst__abc_19396_new_n3321_), .Y(w_mem_inst__0w_mem_7__31_0__8_));
OAI21X1 OAI21X1_1574 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf12), .B(w_mem_inst__abc_19396_new_n3323_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf48), .Y(w_mem_inst__abc_19396_new_n3324_));
OAI21X1 OAI21X1_1575 ( .A(w_mem_inst_w_mem_8__9_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf47), .C(w_mem_inst__abc_19396_new_n3324_), .Y(w_mem_inst__abc_19396_new_n3325_));
OAI21X1 OAI21X1_1576 ( .A(w_mem_inst__abc_19396_new_n1851_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf13), .C(w_mem_inst__abc_19396_new_n3325_), .Y(w_mem_inst__0w_mem_7__31_0__9_));
OAI21X1 OAI21X1_1577 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf11), .B(w_mem_inst__abc_19396_new_n3327_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf46), .Y(w_mem_inst__abc_19396_new_n3328_));
OAI21X1 OAI21X1_1578 ( .A(w_mem_inst_w_mem_8__10_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf45), .C(w_mem_inst__abc_19396_new_n3328_), .Y(w_mem_inst__abc_19396_new_n3329_));
OAI21X1 OAI21X1_1579 ( .A(w_mem_inst__abc_19396_new_n1876_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf12), .C(w_mem_inst__abc_19396_new_n3329_), .Y(w_mem_inst__0w_mem_7__31_0__10_));
OAI21X1 OAI21X1_158 ( .A(_abc_15497_new_n1589_), .B(_abc_15497_new_n1584_), .C(digest_update_bF_buf4), .Y(_abc_15497_new_n1591_));
OAI21X1 OAI21X1_1580 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf10), .B(w_mem_inst__abc_19396_new_n3331_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf44), .Y(w_mem_inst__abc_19396_new_n3332_));
OAI21X1 OAI21X1_1581 ( .A(w_mem_inst_w_mem_8__11_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf43), .C(w_mem_inst__abc_19396_new_n3332_), .Y(w_mem_inst__abc_19396_new_n3333_));
OAI21X1 OAI21X1_1582 ( .A(w_mem_inst__abc_19396_new_n1901_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf11), .C(w_mem_inst__abc_19396_new_n3333_), .Y(w_mem_inst__0w_mem_7__31_0__11_));
OAI21X1 OAI21X1_1583 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf9), .B(w_mem_inst__abc_19396_new_n3335_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf42), .Y(w_mem_inst__abc_19396_new_n3336_));
OAI21X1 OAI21X1_1584 ( .A(w_mem_inst_w_mem_8__12_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf41), .C(w_mem_inst__abc_19396_new_n3336_), .Y(w_mem_inst__abc_19396_new_n3337_));
OAI21X1 OAI21X1_1585 ( .A(w_mem_inst__abc_19396_new_n1926_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf10), .C(w_mem_inst__abc_19396_new_n3337_), .Y(w_mem_inst__0w_mem_7__31_0__12_));
OAI21X1 OAI21X1_1586 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf8), .B(w_mem_inst__abc_19396_new_n3339_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf40), .Y(w_mem_inst__abc_19396_new_n3340_));
OAI21X1 OAI21X1_1587 ( .A(w_mem_inst_w_mem_8__13_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf39), .C(w_mem_inst__abc_19396_new_n3340_), .Y(w_mem_inst__abc_19396_new_n3341_));
OAI21X1 OAI21X1_1588 ( .A(w_mem_inst__abc_19396_new_n1951_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf9), .C(w_mem_inst__abc_19396_new_n3341_), .Y(w_mem_inst__0w_mem_7__31_0__13_));
OAI21X1 OAI21X1_1589 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf7), .B(w_mem_inst__abc_19396_new_n3343_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf38), .Y(w_mem_inst__abc_19396_new_n3344_));
OAI21X1 OAI21X1_159 ( .A(_abc_15497_new_n1580_), .B(_abc_15497_new_n1586_), .C(_abc_15497_new_n1599_), .Y(_abc_15497_new_n1600_));
OAI21X1 OAI21X1_1590 ( .A(w_mem_inst_w_mem_8__14_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf37), .C(w_mem_inst__abc_19396_new_n3344_), .Y(w_mem_inst__abc_19396_new_n3345_));
OAI21X1 OAI21X1_1591 ( .A(w_mem_inst__abc_19396_new_n1976_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf8), .C(w_mem_inst__abc_19396_new_n3345_), .Y(w_mem_inst__0w_mem_7__31_0__14_));
OAI21X1 OAI21X1_1592 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf6), .B(w_mem_inst__abc_19396_new_n3347_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf36), .Y(w_mem_inst__abc_19396_new_n3348_));
OAI21X1 OAI21X1_1593 ( .A(w_mem_inst_w_mem_8__15_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf35), .C(w_mem_inst__abc_19396_new_n3348_), .Y(w_mem_inst__abc_19396_new_n3349_));
OAI21X1 OAI21X1_1594 ( .A(w_mem_inst__abc_19396_new_n2001_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf7), .C(w_mem_inst__abc_19396_new_n3349_), .Y(w_mem_inst__0w_mem_7__31_0__15_));
OAI21X1 OAI21X1_1595 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf5), .B(w_mem_inst__abc_19396_new_n3351_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf34), .Y(w_mem_inst__abc_19396_new_n3352_));
OAI21X1 OAI21X1_1596 ( .A(w_mem_inst_w_mem_8__16_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf33), .C(w_mem_inst__abc_19396_new_n3352_), .Y(w_mem_inst__abc_19396_new_n3353_));
OAI21X1 OAI21X1_1597 ( .A(w_mem_inst__abc_19396_new_n2026_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf6), .C(w_mem_inst__abc_19396_new_n3353_), .Y(w_mem_inst__0w_mem_7__31_0__16_));
OAI21X1 OAI21X1_1598 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf4), .B(w_mem_inst__abc_19396_new_n3355_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf32), .Y(w_mem_inst__abc_19396_new_n3356_));
OAI21X1 OAI21X1_1599 ( .A(w_mem_inst_w_mem_8__17_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf31), .C(w_mem_inst__abc_19396_new_n3356_), .Y(w_mem_inst__abc_19396_new_n3357_));
OAI21X1 OAI21X1_16 ( .A(_auto_iopadmap_cc_368_execute_22625_92_), .B(_abc_15497_new_n883__bF_buf12), .C(_abc_15497_new_n870__bF_buf7), .Y(_abc_15497_new_n899_));
OAI21X1 OAI21X1_160 ( .A(_abc_15497_new_n1587_), .B(_abc_15497_new_n1594_), .C(_abc_15497_new_n1598_), .Y(_abc_15497_new_n1601_));
OAI21X1 OAI21X1_1600 ( .A(w_mem_inst__abc_19396_new_n2051_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf5), .C(w_mem_inst__abc_19396_new_n3357_), .Y(w_mem_inst__0w_mem_7__31_0__17_));
OAI21X1 OAI21X1_1601 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf3), .B(w_mem_inst__abc_19396_new_n3359_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf30), .Y(w_mem_inst__abc_19396_new_n3360_));
OAI21X1 OAI21X1_1602 ( .A(w_mem_inst_w_mem_8__18_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf29), .C(w_mem_inst__abc_19396_new_n3360_), .Y(w_mem_inst__abc_19396_new_n3361_));
OAI21X1 OAI21X1_1603 ( .A(w_mem_inst__abc_19396_new_n2076_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf4), .C(w_mem_inst__abc_19396_new_n3361_), .Y(w_mem_inst__0w_mem_7__31_0__18_));
OAI21X1 OAI21X1_1604 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf2), .B(w_mem_inst__abc_19396_new_n3363_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf28), .Y(w_mem_inst__abc_19396_new_n3364_));
OAI21X1 OAI21X1_1605 ( .A(w_mem_inst_w_mem_8__19_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf27), .C(w_mem_inst__abc_19396_new_n3364_), .Y(w_mem_inst__abc_19396_new_n3365_));
OAI21X1 OAI21X1_1606 ( .A(w_mem_inst__abc_19396_new_n2101_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf3), .C(w_mem_inst__abc_19396_new_n3365_), .Y(w_mem_inst__0w_mem_7__31_0__19_));
OAI21X1 OAI21X1_1607 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf1), .B(w_mem_inst__abc_19396_new_n3367_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf26), .Y(w_mem_inst__abc_19396_new_n3368_));
OAI21X1 OAI21X1_1608 ( .A(w_mem_inst_w_mem_8__20_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf25), .C(w_mem_inst__abc_19396_new_n3368_), .Y(w_mem_inst__abc_19396_new_n3369_));
OAI21X1 OAI21X1_1609 ( .A(w_mem_inst__abc_19396_new_n2126_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf2), .C(w_mem_inst__abc_19396_new_n3369_), .Y(w_mem_inst__0w_mem_7__31_0__20_));
OAI21X1 OAI21X1_161 ( .A(_abc_15497_new_n1594_), .B(_abc_15497_new_n1600_), .C(_abc_15497_new_n1601_), .Y(_abc_15497_new_n1602_));
OAI21X1 OAI21X1_1610 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf0), .B(w_mem_inst__abc_19396_new_n3371_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf24), .Y(w_mem_inst__abc_19396_new_n3372_));
OAI21X1 OAI21X1_1611 ( .A(w_mem_inst_w_mem_8__21_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf23), .C(w_mem_inst__abc_19396_new_n3372_), .Y(w_mem_inst__abc_19396_new_n3373_));
OAI21X1 OAI21X1_1612 ( .A(w_mem_inst__abc_19396_new_n2151_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf1), .C(w_mem_inst__abc_19396_new_n3373_), .Y(w_mem_inst__0w_mem_7__31_0__21_));
OAI21X1 OAI21X1_1613 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf60), .B(w_mem_inst__abc_19396_new_n3375_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf22), .Y(w_mem_inst__abc_19396_new_n3376_));
OAI21X1 OAI21X1_1614 ( .A(w_mem_inst_w_mem_8__22_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf21), .C(w_mem_inst__abc_19396_new_n3376_), .Y(w_mem_inst__abc_19396_new_n3377_));
OAI21X1 OAI21X1_1615 ( .A(w_mem_inst__abc_19396_new_n2176_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf0), .C(w_mem_inst__abc_19396_new_n3377_), .Y(w_mem_inst__0w_mem_7__31_0__22_));
OAI21X1 OAI21X1_1616 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf59), .B(w_mem_inst__abc_19396_new_n3379_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf20), .Y(w_mem_inst__abc_19396_new_n3380_));
OAI21X1 OAI21X1_1617 ( .A(w_mem_inst_w_mem_8__23_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf19), .C(w_mem_inst__abc_19396_new_n3380_), .Y(w_mem_inst__abc_19396_new_n3381_));
OAI21X1 OAI21X1_1618 ( .A(w_mem_inst__abc_19396_new_n2201_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf60), .C(w_mem_inst__abc_19396_new_n3381_), .Y(w_mem_inst__0w_mem_7__31_0__23_));
OAI21X1 OAI21X1_1619 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf58), .B(w_mem_inst__abc_19396_new_n3383_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf18), .Y(w_mem_inst__abc_19396_new_n3384_));
OAI21X1 OAI21X1_162 ( .A(_abc_15497_new_n1582_), .B(_abc_15497_new_n1606_), .C(_abc_15497_new_n1607_), .Y(_abc_15497_new_n1608_));
OAI21X1 OAI21X1_1620 ( .A(w_mem_inst_w_mem_8__24_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf17), .C(w_mem_inst__abc_19396_new_n3384_), .Y(w_mem_inst__abc_19396_new_n3385_));
OAI21X1 OAI21X1_1621 ( .A(w_mem_inst__abc_19396_new_n2226_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf59), .C(w_mem_inst__abc_19396_new_n3385_), .Y(w_mem_inst__0w_mem_7__31_0__24_));
OAI21X1 OAI21X1_1622 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf57), .B(w_mem_inst__abc_19396_new_n3387_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf16), .Y(w_mem_inst__abc_19396_new_n3388_));
OAI21X1 OAI21X1_1623 ( .A(w_mem_inst_w_mem_8__25_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf15), .C(w_mem_inst__abc_19396_new_n3388_), .Y(w_mem_inst__abc_19396_new_n3389_));
OAI21X1 OAI21X1_1624 ( .A(w_mem_inst__abc_19396_new_n2251_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf58), .C(w_mem_inst__abc_19396_new_n3389_), .Y(w_mem_inst__0w_mem_7__31_0__25_));
OAI21X1 OAI21X1_1625 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf56), .B(w_mem_inst__abc_19396_new_n3391_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf14), .Y(w_mem_inst__abc_19396_new_n3392_));
OAI21X1 OAI21X1_1626 ( .A(w_mem_inst_w_mem_8__26_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf13), .C(w_mem_inst__abc_19396_new_n3392_), .Y(w_mem_inst__abc_19396_new_n3393_));
OAI21X1 OAI21X1_1627 ( .A(w_mem_inst__abc_19396_new_n2276_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf57), .C(w_mem_inst__abc_19396_new_n3393_), .Y(w_mem_inst__0w_mem_7__31_0__26_));
OAI21X1 OAI21X1_1628 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf55), .B(w_mem_inst__abc_19396_new_n3395_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf12), .Y(w_mem_inst__abc_19396_new_n3396_));
OAI21X1 OAI21X1_1629 ( .A(w_mem_inst_w_mem_8__27_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf11), .C(w_mem_inst__abc_19396_new_n3396_), .Y(w_mem_inst__abc_19396_new_n3397_));
OAI21X1 OAI21X1_163 ( .A(_abc_15497_new_n1605_), .B(_abc_15497_new_n1559_), .C(_abc_15497_new_n1609_), .Y(_abc_15497_new_n1610_));
OAI21X1 OAI21X1_1630 ( .A(w_mem_inst__abc_19396_new_n2301_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf56), .C(w_mem_inst__abc_19396_new_n3397_), .Y(w_mem_inst__0w_mem_7__31_0__27_));
OAI21X1 OAI21X1_1631 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf54), .B(w_mem_inst__abc_19396_new_n3399_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf10), .Y(w_mem_inst__abc_19396_new_n3400_));
OAI21X1 OAI21X1_1632 ( .A(w_mem_inst_w_mem_8__28_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf9), .C(w_mem_inst__abc_19396_new_n3400_), .Y(w_mem_inst__abc_19396_new_n3401_));
OAI21X1 OAI21X1_1633 ( .A(w_mem_inst__abc_19396_new_n2326_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf55), .C(w_mem_inst__abc_19396_new_n3401_), .Y(w_mem_inst__0w_mem_7__31_0__28_));
OAI21X1 OAI21X1_1634 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf53), .B(w_mem_inst__abc_19396_new_n3403_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf8), .Y(w_mem_inst__abc_19396_new_n3404_));
OAI21X1 OAI21X1_1635 ( .A(w_mem_inst_w_mem_8__29_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf7), .C(w_mem_inst__abc_19396_new_n3404_), .Y(w_mem_inst__abc_19396_new_n3405_));
OAI21X1 OAI21X1_1636 ( .A(w_mem_inst__abc_19396_new_n2351_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf54), .C(w_mem_inst__abc_19396_new_n3405_), .Y(w_mem_inst__0w_mem_7__31_0__29_));
OAI21X1 OAI21X1_1637 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf52), .B(w_mem_inst__abc_19396_new_n3407_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf6), .Y(w_mem_inst__abc_19396_new_n3408_));
OAI21X1 OAI21X1_1638 ( .A(w_mem_inst_w_mem_8__30_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf5), .C(w_mem_inst__abc_19396_new_n3408_), .Y(w_mem_inst__abc_19396_new_n3409_));
OAI21X1 OAI21X1_1639 ( .A(w_mem_inst__abc_19396_new_n2376_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf53), .C(w_mem_inst__abc_19396_new_n3409_), .Y(w_mem_inst__0w_mem_7__31_0__30_));
OAI21X1 OAI21X1_164 ( .A(_auto_iopadmap_cc_368_execute_22625_60_), .B(_abc_15497_new_n883__bF_buf11), .C(_abc_15497_new_n870__bF_buf4), .Y(_abc_15497_new_n1615_));
OAI21X1 OAI21X1_1640 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf51), .B(w_mem_inst__abc_19396_new_n3411_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf4), .Y(w_mem_inst__abc_19396_new_n3412_));
OAI21X1 OAI21X1_1641 ( .A(w_mem_inst_w_mem_8__31_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf3), .C(w_mem_inst__abc_19396_new_n3412_), .Y(w_mem_inst__abc_19396_new_n3413_));
OAI21X1 OAI21X1_1642 ( .A(w_mem_inst__abc_19396_new_n2401_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf52), .C(w_mem_inst__abc_19396_new_n3413_), .Y(w_mem_inst__0w_mem_7__31_0__31_));
OAI21X1 OAI21X1_1643 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf50), .B(w_mem_inst__abc_19396_new_n3416_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf2), .Y(w_mem_inst__abc_19396_new_n3417_));
OAI21X1 OAI21X1_1644 ( .A(w_mem_inst_w_mem_10__0_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf1), .C(w_mem_inst__abc_19396_new_n3417_), .Y(w_mem_inst__abc_19396_new_n3418_));
OAI21X1 OAI21X1_1645 ( .A(w_mem_inst__abc_19396_new_n3415_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf51), .C(w_mem_inst__abc_19396_new_n3418_), .Y(w_mem_inst__0w_mem_9__31_0__0_));
OAI21X1 OAI21X1_1646 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf49), .B(w_mem_inst__abc_19396_new_n3421_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf0), .Y(w_mem_inst__abc_19396_new_n3422_));
OAI21X1 OAI21X1_1647 ( .A(w_mem_inst_w_mem_10__1_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf96), .C(w_mem_inst__abc_19396_new_n3422_), .Y(w_mem_inst__abc_19396_new_n3423_));
OAI21X1 OAI21X1_1648 ( .A(w_mem_inst__abc_19396_new_n3420_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf50), .C(w_mem_inst__abc_19396_new_n3423_), .Y(w_mem_inst__0w_mem_9__31_0__1_));
OAI21X1 OAI21X1_1649 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf48), .B(w_mem_inst__abc_19396_new_n3426_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf95), .Y(w_mem_inst__abc_19396_new_n3427_));
OAI21X1 OAI21X1_165 ( .A(_abc_15497_new_n1612_), .B(_abc_15497_new_n1614_), .C(_abc_15497_new_n1615_), .Y(_0H3_reg_31_0__28_));
OAI21X1 OAI21X1_1650 ( .A(w_mem_inst_w_mem_10__2_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf94), .C(w_mem_inst__abc_19396_new_n3427_), .Y(w_mem_inst__abc_19396_new_n3428_));
OAI21X1 OAI21X1_1651 ( .A(w_mem_inst__abc_19396_new_n3425_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf49), .C(w_mem_inst__abc_19396_new_n3428_), .Y(w_mem_inst__0w_mem_9__31_0__2_));
OAI21X1 OAI21X1_1652 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf47), .B(w_mem_inst__abc_19396_new_n3431_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf93), .Y(w_mem_inst__abc_19396_new_n3432_));
OAI21X1 OAI21X1_1653 ( .A(w_mem_inst_w_mem_10__3_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf92), .C(w_mem_inst__abc_19396_new_n3432_), .Y(w_mem_inst__abc_19396_new_n3433_));
OAI21X1 OAI21X1_1654 ( .A(w_mem_inst__abc_19396_new_n3430_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf48), .C(w_mem_inst__abc_19396_new_n3433_), .Y(w_mem_inst__0w_mem_9__31_0__3_));
OAI21X1 OAI21X1_1655 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf46), .B(w_mem_inst__abc_19396_new_n3436_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf91), .Y(w_mem_inst__abc_19396_new_n3437_));
OAI21X1 OAI21X1_1656 ( .A(w_mem_inst_w_mem_10__4_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf90), .C(w_mem_inst__abc_19396_new_n3437_), .Y(w_mem_inst__abc_19396_new_n3438_));
OAI21X1 OAI21X1_1657 ( .A(w_mem_inst__abc_19396_new_n3435_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf47), .C(w_mem_inst__abc_19396_new_n3438_), .Y(w_mem_inst__0w_mem_9__31_0__4_));
OAI21X1 OAI21X1_1658 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf45), .B(w_mem_inst__abc_19396_new_n3441_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf89), .Y(w_mem_inst__abc_19396_new_n3442_));
OAI21X1 OAI21X1_1659 ( .A(w_mem_inst_w_mem_10__5_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf88), .C(w_mem_inst__abc_19396_new_n3442_), .Y(w_mem_inst__abc_19396_new_n3443_));
OAI21X1 OAI21X1_166 ( .A(_abc_15497_new_n871__bF_buf1), .B(_abc_15497_new_n872__bF_buf1), .C(_auto_iopadmap_cc_368_execute_22625_61_), .Y(_abc_15497_new_n1617_));
OAI21X1 OAI21X1_1660 ( .A(w_mem_inst__abc_19396_new_n3440_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf46), .C(w_mem_inst__abc_19396_new_n3443_), .Y(w_mem_inst__0w_mem_9__31_0__5_));
OAI21X1 OAI21X1_1661 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf44), .B(w_mem_inst__abc_19396_new_n3446_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf87), .Y(w_mem_inst__abc_19396_new_n3447_));
OAI21X1 OAI21X1_1662 ( .A(w_mem_inst_w_mem_10__6_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf86), .C(w_mem_inst__abc_19396_new_n3447_), .Y(w_mem_inst__abc_19396_new_n3448_));
OAI21X1 OAI21X1_1663 ( .A(w_mem_inst__abc_19396_new_n3445_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf45), .C(w_mem_inst__abc_19396_new_n3448_), .Y(w_mem_inst__0w_mem_9__31_0__6_));
OAI21X1 OAI21X1_1664 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf43), .B(w_mem_inst__abc_19396_new_n3451_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf85), .Y(w_mem_inst__abc_19396_new_n3452_));
OAI21X1 OAI21X1_1665 ( .A(w_mem_inst_w_mem_10__7_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf84), .C(w_mem_inst__abc_19396_new_n3452_), .Y(w_mem_inst__abc_19396_new_n3453_));
OAI21X1 OAI21X1_1666 ( .A(w_mem_inst__abc_19396_new_n3450_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf44), .C(w_mem_inst__abc_19396_new_n3453_), .Y(w_mem_inst__0w_mem_9__31_0__7_));
OAI21X1 OAI21X1_1667 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf42), .B(w_mem_inst__abc_19396_new_n3456_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf83), .Y(w_mem_inst__abc_19396_new_n3457_));
OAI21X1 OAI21X1_1668 ( .A(w_mem_inst_w_mem_10__8_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf82), .C(w_mem_inst__abc_19396_new_n3457_), .Y(w_mem_inst__abc_19396_new_n3458_));
OAI21X1 OAI21X1_1669 ( .A(w_mem_inst__abc_19396_new_n3455_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf43), .C(w_mem_inst__abc_19396_new_n3458_), .Y(w_mem_inst__0w_mem_9__31_0__8_));
OAI21X1 OAI21X1_167 ( .A(_abc_15497_new_n1624_), .B(_abc_15497_new_n1619_), .C(digest_update_bF_buf2), .Y(_abc_15497_new_n1625_));
OAI21X1 OAI21X1_1670 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf41), .B(w_mem_inst__abc_19396_new_n3461_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf81), .Y(w_mem_inst__abc_19396_new_n3462_));
OAI21X1 OAI21X1_1671 ( .A(w_mem_inst_w_mem_10__9_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf80), .C(w_mem_inst__abc_19396_new_n3462_), .Y(w_mem_inst__abc_19396_new_n3463_));
OAI21X1 OAI21X1_1672 ( .A(w_mem_inst__abc_19396_new_n3460_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf42), .C(w_mem_inst__abc_19396_new_n3463_), .Y(w_mem_inst__0w_mem_9__31_0__9_));
OAI21X1 OAI21X1_1673 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf40), .B(w_mem_inst__abc_19396_new_n3466_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf79), .Y(w_mem_inst__abc_19396_new_n3467_));
OAI21X1 OAI21X1_1674 ( .A(w_mem_inst_w_mem_10__10_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf78), .C(w_mem_inst__abc_19396_new_n3467_), .Y(w_mem_inst__abc_19396_new_n3468_));
OAI21X1 OAI21X1_1675 ( .A(w_mem_inst__abc_19396_new_n3465_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf41), .C(w_mem_inst__abc_19396_new_n3468_), .Y(w_mem_inst__0w_mem_9__31_0__10_));
OAI21X1 OAI21X1_1676 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf39), .B(w_mem_inst__abc_19396_new_n3471_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf77), .Y(w_mem_inst__abc_19396_new_n3472_));
OAI21X1 OAI21X1_1677 ( .A(w_mem_inst_w_mem_10__11_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf76), .C(w_mem_inst__abc_19396_new_n3472_), .Y(w_mem_inst__abc_19396_new_n3473_));
OAI21X1 OAI21X1_1678 ( .A(w_mem_inst__abc_19396_new_n3470_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf40), .C(w_mem_inst__abc_19396_new_n3473_), .Y(w_mem_inst__0w_mem_9__31_0__11_));
OAI21X1 OAI21X1_1679 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf38), .B(w_mem_inst__abc_19396_new_n3476_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf75), .Y(w_mem_inst__abc_19396_new_n3477_));
OAI21X1 OAI21X1_168 ( .A(_abc_15497_new_n1618_), .B(_abc_15497_new_n1620_), .C(_abc_15497_new_n1631_), .Y(_abc_15497_new_n1632_));
OAI21X1 OAI21X1_1680 ( .A(w_mem_inst_w_mem_10__12_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf74), .C(w_mem_inst__abc_19396_new_n3477_), .Y(w_mem_inst__abc_19396_new_n3478_));
OAI21X1 OAI21X1_1681 ( .A(w_mem_inst__abc_19396_new_n3475_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf39), .C(w_mem_inst__abc_19396_new_n3478_), .Y(w_mem_inst__0w_mem_9__31_0__12_));
OAI21X1 OAI21X1_1682 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf37), .B(w_mem_inst__abc_19396_new_n3481_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf73), .Y(w_mem_inst__abc_19396_new_n3482_));
OAI21X1 OAI21X1_1683 ( .A(w_mem_inst_w_mem_10__13_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf72), .C(w_mem_inst__abc_19396_new_n3482_), .Y(w_mem_inst__abc_19396_new_n3483_));
OAI21X1 OAI21X1_1684 ( .A(w_mem_inst__abc_19396_new_n3480_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf38), .C(w_mem_inst__abc_19396_new_n3483_), .Y(w_mem_inst__0w_mem_9__31_0__13_));
OAI21X1 OAI21X1_1685 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf36), .B(w_mem_inst__abc_19396_new_n3486_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf71), .Y(w_mem_inst__abc_19396_new_n3487_));
OAI21X1 OAI21X1_1686 ( .A(w_mem_inst_w_mem_10__14_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf70), .C(w_mem_inst__abc_19396_new_n3487_), .Y(w_mem_inst__abc_19396_new_n3488_));
OAI21X1 OAI21X1_1687 ( .A(w_mem_inst__abc_19396_new_n3485_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf37), .C(w_mem_inst__abc_19396_new_n3488_), .Y(w_mem_inst__0w_mem_9__31_0__14_));
OAI21X1 OAI21X1_1688 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf35), .B(w_mem_inst__abc_19396_new_n3491_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf69), .Y(w_mem_inst__abc_19396_new_n3492_));
OAI21X1 OAI21X1_1689 ( .A(w_mem_inst_w_mem_10__15_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf68), .C(w_mem_inst__abc_19396_new_n3492_), .Y(w_mem_inst__abc_19396_new_n3493_));
OAI21X1 OAI21X1_169 ( .A(_abc_15497_new_n1630_), .B(_abc_15497_new_n1634_), .C(_abc_15497_new_n1638_), .Y(_abc_15497_new_n1639_));
OAI21X1 OAI21X1_1690 ( .A(w_mem_inst__abc_19396_new_n3490_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf36), .C(w_mem_inst__abc_19396_new_n3493_), .Y(w_mem_inst__0w_mem_9__31_0__15_));
OAI21X1 OAI21X1_1691 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf34), .B(w_mem_inst__abc_19396_new_n3496_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf67), .Y(w_mem_inst__abc_19396_new_n3497_));
OAI21X1 OAI21X1_1692 ( .A(w_mem_inst_w_mem_10__16_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf66), .C(w_mem_inst__abc_19396_new_n3497_), .Y(w_mem_inst__abc_19396_new_n3498_));
OAI21X1 OAI21X1_1693 ( .A(w_mem_inst__abc_19396_new_n3495_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf35), .C(w_mem_inst__abc_19396_new_n3498_), .Y(w_mem_inst__0w_mem_9__31_0__16_));
OAI21X1 OAI21X1_1694 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf33), .B(w_mem_inst__abc_19396_new_n3501_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf65), .Y(w_mem_inst__abc_19396_new_n3502_));
OAI21X1 OAI21X1_1695 ( .A(w_mem_inst_w_mem_10__17_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf64), .C(w_mem_inst__abc_19396_new_n3502_), .Y(w_mem_inst__abc_19396_new_n3503_));
OAI21X1 OAI21X1_1696 ( .A(w_mem_inst__abc_19396_new_n3500_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf34), .C(w_mem_inst__abc_19396_new_n3503_), .Y(w_mem_inst__0w_mem_9__31_0__17_));
OAI21X1 OAI21X1_1697 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf32), .B(w_mem_inst__abc_19396_new_n3506_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf63), .Y(w_mem_inst__abc_19396_new_n3507_));
OAI21X1 OAI21X1_1698 ( .A(w_mem_inst_w_mem_10__18_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf62), .C(w_mem_inst__abc_19396_new_n3507_), .Y(w_mem_inst__abc_19396_new_n3508_));
OAI21X1 OAI21X1_1699 ( .A(w_mem_inst__abc_19396_new_n3505_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf33), .C(w_mem_inst__abc_19396_new_n3508_), .Y(w_mem_inst__0w_mem_9__31_0__18_));
OAI21X1 OAI21X1_17 ( .A(_abc_15497_new_n907_), .B(_abc_15497_new_n902_), .C(digest_update_bF_buf6), .Y(_abc_15497_new_n909_));
OAI21X1 OAI21X1_170 ( .A(_abc_15497_new_n1640_), .B(_abc_15497_new_n1639_), .C(digest_update_bF_buf1), .Y(_abc_15497_new_n1642_));
OAI21X1 OAI21X1_1700 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf31), .B(w_mem_inst__abc_19396_new_n3511_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf61), .Y(w_mem_inst__abc_19396_new_n3512_));
OAI21X1 OAI21X1_1701 ( .A(w_mem_inst_w_mem_10__19_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf60), .C(w_mem_inst__abc_19396_new_n3512_), .Y(w_mem_inst__abc_19396_new_n3513_));
OAI21X1 OAI21X1_1702 ( .A(w_mem_inst__abc_19396_new_n3510_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf32), .C(w_mem_inst__abc_19396_new_n3513_), .Y(w_mem_inst__0w_mem_9__31_0__19_));
OAI21X1 OAI21X1_1703 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf30), .B(w_mem_inst__abc_19396_new_n3516_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf59), .Y(w_mem_inst__abc_19396_new_n3517_));
OAI21X1 OAI21X1_1704 ( .A(w_mem_inst_w_mem_10__20_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf58), .C(w_mem_inst__abc_19396_new_n3517_), .Y(w_mem_inst__abc_19396_new_n3518_));
OAI21X1 OAI21X1_1705 ( .A(w_mem_inst__abc_19396_new_n3515_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf31), .C(w_mem_inst__abc_19396_new_n3518_), .Y(w_mem_inst__0w_mem_9__31_0__20_));
OAI21X1 OAI21X1_1706 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf29), .B(w_mem_inst__abc_19396_new_n3521_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf57), .Y(w_mem_inst__abc_19396_new_n3522_));
OAI21X1 OAI21X1_1707 ( .A(w_mem_inst_w_mem_10__21_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf56), .C(w_mem_inst__abc_19396_new_n3522_), .Y(w_mem_inst__abc_19396_new_n3523_));
OAI21X1 OAI21X1_1708 ( .A(w_mem_inst__abc_19396_new_n3520_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf30), .C(w_mem_inst__abc_19396_new_n3523_), .Y(w_mem_inst__0w_mem_9__31_0__21_));
OAI21X1 OAI21X1_1709 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf28), .B(w_mem_inst__abc_19396_new_n3526_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf55), .Y(w_mem_inst__abc_19396_new_n3527_));
OAI21X1 OAI21X1_171 ( .A(next), .B(init), .C(_auto_iopadmap_cc_368_execute_22788), .Y(_abc_15497_new_n1644_));
OAI21X1 OAI21X1_1710 ( .A(w_mem_inst_w_mem_10__22_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf54), .C(w_mem_inst__abc_19396_new_n3527_), .Y(w_mem_inst__abc_19396_new_n3528_));
OAI21X1 OAI21X1_1711 ( .A(w_mem_inst__abc_19396_new_n3525_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf29), .C(w_mem_inst__abc_19396_new_n3528_), .Y(w_mem_inst__0w_mem_9__31_0__22_));
OAI21X1 OAI21X1_1712 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf27), .B(w_mem_inst__abc_19396_new_n3531_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf53), .Y(w_mem_inst__abc_19396_new_n3532_));
OAI21X1 OAI21X1_1713 ( .A(w_mem_inst_w_mem_10__23_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf52), .C(w_mem_inst__abc_19396_new_n3532_), .Y(w_mem_inst__abc_19396_new_n3533_));
OAI21X1 OAI21X1_1714 ( .A(w_mem_inst__abc_19396_new_n3530_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf28), .C(w_mem_inst__abc_19396_new_n3533_), .Y(w_mem_inst__0w_mem_9__31_0__23_));
OAI21X1 OAI21X1_1715 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf26), .B(w_mem_inst__abc_19396_new_n3536_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf51), .Y(w_mem_inst__abc_19396_new_n3537_));
OAI21X1 OAI21X1_1716 ( .A(w_mem_inst_w_mem_10__24_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf50), .C(w_mem_inst__abc_19396_new_n3537_), .Y(w_mem_inst__abc_19396_new_n3538_));
OAI21X1 OAI21X1_1717 ( .A(w_mem_inst__abc_19396_new_n3535_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf27), .C(w_mem_inst__abc_19396_new_n3538_), .Y(w_mem_inst__0w_mem_9__31_0__24_));
OAI21X1 OAI21X1_1718 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf25), .B(w_mem_inst__abc_19396_new_n3541_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf49), .Y(w_mem_inst__abc_19396_new_n3542_));
OAI21X1 OAI21X1_1719 ( .A(w_mem_inst_w_mem_10__25_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf48), .C(w_mem_inst__abc_19396_new_n3542_), .Y(w_mem_inst__abc_19396_new_n3543_));
OAI21X1 OAI21X1_172 ( .A(_abc_15497_new_n871__bF_buf0), .B(_abc_15497_new_n1647_), .C(_abc_15497_new_n1646_), .Y(_abc_15497_new_n1648_));
OAI21X1 OAI21X1_1720 ( .A(w_mem_inst__abc_19396_new_n3540_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf26), .C(w_mem_inst__abc_19396_new_n3543_), .Y(w_mem_inst__0w_mem_9__31_0__25_));
OAI21X1 OAI21X1_1721 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf24), .B(w_mem_inst__abc_19396_new_n3546_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf47), .Y(w_mem_inst__abc_19396_new_n3547_));
OAI21X1 OAI21X1_1722 ( .A(w_mem_inst_w_mem_10__26_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf46), .C(w_mem_inst__abc_19396_new_n3547_), .Y(w_mem_inst__abc_19396_new_n3548_));
OAI21X1 OAI21X1_1723 ( .A(w_mem_inst__abc_19396_new_n3545_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf25), .C(w_mem_inst__abc_19396_new_n3548_), .Y(w_mem_inst__0w_mem_9__31_0__26_));
OAI21X1 OAI21X1_1724 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf23), .B(w_mem_inst__abc_19396_new_n3551_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf45), .Y(w_mem_inst__abc_19396_new_n3552_));
OAI21X1 OAI21X1_1725 ( .A(w_mem_inst_w_mem_10__27_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf44), .C(w_mem_inst__abc_19396_new_n3552_), .Y(w_mem_inst__abc_19396_new_n3553_));
OAI21X1 OAI21X1_1726 ( .A(w_mem_inst__abc_19396_new_n3550_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf24), .C(w_mem_inst__abc_19396_new_n3553_), .Y(w_mem_inst__0w_mem_9__31_0__27_));
OAI21X1 OAI21X1_1727 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf22), .B(w_mem_inst__abc_19396_new_n3556_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf43), .Y(w_mem_inst__abc_19396_new_n3557_));
OAI21X1 OAI21X1_1728 ( .A(w_mem_inst_w_mem_10__28_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf42), .C(w_mem_inst__abc_19396_new_n3557_), .Y(w_mem_inst__abc_19396_new_n3558_));
OAI21X1 OAI21X1_1729 ( .A(w_mem_inst__abc_19396_new_n3555_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf23), .C(w_mem_inst__abc_19396_new_n3558_), .Y(w_mem_inst__0w_mem_9__31_0__28_));
OAI21X1 OAI21X1_173 ( .A(_abc_15497_new_n937_), .B(_abc_15497_new_n1648__bF_buf8), .C(_abc_15497_new_n1651_), .Y(_0e_reg_31_0__0_));
OAI21X1 OAI21X1_1730 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf21), .B(w_mem_inst__abc_19396_new_n3561_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf41), .Y(w_mem_inst__abc_19396_new_n3562_));
OAI21X1 OAI21X1_1731 ( .A(w_mem_inst_w_mem_10__29_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf40), .C(w_mem_inst__abc_19396_new_n3562_), .Y(w_mem_inst__abc_19396_new_n3563_));
OAI21X1 OAI21X1_1732 ( .A(w_mem_inst__abc_19396_new_n3560_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf22), .C(w_mem_inst__abc_19396_new_n3563_), .Y(w_mem_inst__0w_mem_9__31_0__29_));
OAI21X1 OAI21X1_1733 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf20), .B(w_mem_inst__abc_19396_new_n3566_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf39), .Y(w_mem_inst__abc_19396_new_n3567_));
OAI21X1 OAI21X1_1734 ( .A(w_mem_inst_w_mem_10__30_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf38), .C(w_mem_inst__abc_19396_new_n3567_), .Y(w_mem_inst__abc_19396_new_n3568_));
OAI21X1 OAI21X1_1735 ( .A(w_mem_inst__abc_19396_new_n3565_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf21), .C(w_mem_inst__abc_19396_new_n3568_), .Y(w_mem_inst__0w_mem_9__31_0__30_));
OAI21X1 OAI21X1_1736 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf19), .B(w_mem_inst__abc_19396_new_n3571_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf37), .Y(w_mem_inst__abc_19396_new_n3572_));
OAI21X1 OAI21X1_1737 ( .A(w_mem_inst_w_mem_10__31_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf36), .C(w_mem_inst__abc_19396_new_n3572_), .Y(w_mem_inst__abc_19396_new_n3573_));
OAI21X1 OAI21X1_1738 ( .A(w_mem_inst__abc_19396_new_n3570_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf20), .C(w_mem_inst__abc_19396_new_n3573_), .Y(w_mem_inst__0w_mem_9__31_0__31_));
OAI21X1 OAI21X1_1739 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf18), .B(w_mem_inst__abc_19396_new_n3575_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf35), .Y(w_mem_inst__abc_19396_new_n3576_));
OAI21X1 OAI21X1_174 ( .A(_abc_15497_new_n947_), .B(_abc_15497_new_n1648__bF_buf7), .C(_abc_15497_new_n1654_), .Y(_0e_reg_31_0__1_));
OAI21X1 OAI21X1_1740 ( .A(w_mem_inst_w_mem_9__0_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf34), .C(w_mem_inst__abc_19396_new_n3576_), .Y(w_mem_inst__abc_19396_new_n3577_));
OAI21X1 OAI21X1_1741 ( .A(w_mem_inst__abc_19396_new_n1600_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf19), .C(w_mem_inst__abc_19396_new_n3577_), .Y(w_mem_inst__0w_mem_8__31_0__0_));
OAI21X1 OAI21X1_1742 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf17), .B(w_mem_inst__abc_19396_new_n3579_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf33), .Y(w_mem_inst__abc_19396_new_n3580_));
OAI21X1 OAI21X1_1743 ( .A(w_mem_inst_w_mem_9__1_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf32), .C(w_mem_inst__abc_19396_new_n3580_), .Y(w_mem_inst__abc_19396_new_n3581_));
OAI21X1 OAI21X1_1744 ( .A(w_mem_inst__abc_19396_new_n1648_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf18), .C(w_mem_inst__abc_19396_new_n3581_), .Y(w_mem_inst__0w_mem_8__31_0__1_));
OAI21X1 OAI21X1_1745 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf16), .B(w_mem_inst__abc_19396_new_n3583_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf31), .Y(w_mem_inst__abc_19396_new_n3584_));
OAI21X1 OAI21X1_1746 ( .A(w_mem_inst_w_mem_9__2_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf30), .C(w_mem_inst__abc_19396_new_n3584_), .Y(w_mem_inst__abc_19396_new_n3585_));
OAI21X1 OAI21X1_1747 ( .A(w_mem_inst__abc_19396_new_n1673_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf17), .C(w_mem_inst__abc_19396_new_n3585_), .Y(w_mem_inst__0w_mem_8__31_0__2_));
OAI21X1 OAI21X1_1748 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf15), .B(w_mem_inst__abc_19396_new_n3587_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf29), .Y(w_mem_inst__abc_19396_new_n3588_));
OAI21X1 OAI21X1_1749 ( .A(w_mem_inst_w_mem_9__3_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf28), .C(w_mem_inst__abc_19396_new_n3588_), .Y(w_mem_inst__abc_19396_new_n3589_));
OAI21X1 OAI21X1_175 ( .A(_abc_15497_new_n956_), .B(_abc_15497_new_n1648__bF_buf6), .C(_abc_15497_new_n1657_), .Y(_0e_reg_31_0__2_));
OAI21X1 OAI21X1_1750 ( .A(w_mem_inst__abc_19396_new_n1698_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf16), .C(w_mem_inst__abc_19396_new_n3589_), .Y(w_mem_inst__0w_mem_8__31_0__3_));
OAI21X1 OAI21X1_1751 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf14), .B(w_mem_inst__abc_19396_new_n3591_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf27), .Y(w_mem_inst__abc_19396_new_n3592_));
OAI21X1 OAI21X1_1752 ( .A(w_mem_inst_w_mem_9__4_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf26), .C(w_mem_inst__abc_19396_new_n3592_), .Y(w_mem_inst__abc_19396_new_n3593_));
OAI21X1 OAI21X1_1753 ( .A(w_mem_inst__abc_19396_new_n1723_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf15), .C(w_mem_inst__abc_19396_new_n3593_), .Y(w_mem_inst__0w_mem_8__31_0__4_));
OAI21X1 OAI21X1_1754 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf13), .B(w_mem_inst__abc_19396_new_n3595_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf25), .Y(w_mem_inst__abc_19396_new_n3596_));
OAI21X1 OAI21X1_1755 ( .A(w_mem_inst_w_mem_9__5_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf24), .C(w_mem_inst__abc_19396_new_n3596_), .Y(w_mem_inst__abc_19396_new_n3597_));
OAI21X1 OAI21X1_1756 ( .A(w_mem_inst__abc_19396_new_n1748_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf14), .C(w_mem_inst__abc_19396_new_n3597_), .Y(w_mem_inst__0w_mem_8__31_0__5_));
OAI21X1 OAI21X1_1757 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf12), .B(w_mem_inst__abc_19396_new_n3599_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf23), .Y(w_mem_inst__abc_19396_new_n3600_));
OAI21X1 OAI21X1_1758 ( .A(w_mem_inst_w_mem_9__6_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf22), .C(w_mem_inst__abc_19396_new_n3600_), .Y(w_mem_inst__abc_19396_new_n3601_));
OAI21X1 OAI21X1_1759 ( .A(w_mem_inst__abc_19396_new_n1773_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf13), .C(w_mem_inst__abc_19396_new_n3601_), .Y(w_mem_inst__0w_mem_8__31_0__6_));
OAI21X1 OAI21X1_176 ( .A(_abc_15497_new_n960_), .B(_abc_15497_new_n1648__bF_buf5), .C(_abc_15497_new_n1660_), .Y(_0e_reg_31_0__3_));
OAI21X1 OAI21X1_1760 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf11), .B(w_mem_inst__abc_19396_new_n3603_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf21), .Y(w_mem_inst__abc_19396_new_n3604_));
OAI21X1 OAI21X1_1761 ( .A(w_mem_inst_w_mem_9__7_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf20), .C(w_mem_inst__abc_19396_new_n3604_), .Y(w_mem_inst__abc_19396_new_n3605_));
OAI21X1 OAI21X1_1762 ( .A(w_mem_inst__abc_19396_new_n1798_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf12), .C(w_mem_inst__abc_19396_new_n3605_), .Y(w_mem_inst__0w_mem_8__31_0__7_));
OAI21X1 OAI21X1_1763 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf10), .B(w_mem_inst__abc_19396_new_n3607_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf19), .Y(w_mem_inst__abc_19396_new_n3608_));
OAI21X1 OAI21X1_1764 ( .A(w_mem_inst_w_mem_9__8_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf18), .C(w_mem_inst__abc_19396_new_n3608_), .Y(w_mem_inst__abc_19396_new_n3609_));
OAI21X1 OAI21X1_1765 ( .A(w_mem_inst__abc_19396_new_n1823_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf11), .C(w_mem_inst__abc_19396_new_n3609_), .Y(w_mem_inst__0w_mem_8__31_0__8_));
OAI21X1 OAI21X1_1766 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf9), .B(w_mem_inst__abc_19396_new_n3611_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf17), .Y(w_mem_inst__abc_19396_new_n3612_));
OAI21X1 OAI21X1_1767 ( .A(w_mem_inst_w_mem_9__9_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf16), .C(w_mem_inst__abc_19396_new_n3612_), .Y(w_mem_inst__abc_19396_new_n3613_));
OAI21X1 OAI21X1_1768 ( .A(w_mem_inst__abc_19396_new_n1848_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf10), .C(w_mem_inst__abc_19396_new_n3613_), .Y(w_mem_inst__0w_mem_8__31_0__9_));
OAI21X1 OAI21X1_1769 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf8), .B(w_mem_inst__abc_19396_new_n3615_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf15), .Y(w_mem_inst__abc_19396_new_n3616_));
OAI21X1 OAI21X1_177 ( .A(_auto_iopadmap_cc_368_execute_22625_4_), .B(_abc_15497_new_n883__bF_buf6), .C(round_ctr_rst_bF_buf8), .Y(_abc_15497_new_n1662_));
OAI21X1 OAI21X1_1770 ( .A(w_mem_inst_w_mem_9__10_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf14), .C(w_mem_inst__abc_19396_new_n3616_), .Y(w_mem_inst__abc_19396_new_n3617_));
OAI21X1 OAI21X1_1771 ( .A(w_mem_inst__abc_19396_new_n1873_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf9), .C(w_mem_inst__abc_19396_new_n3617_), .Y(w_mem_inst__0w_mem_8__31_0__10_));
OAI21X1 OAI21X1_1772 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf7), .B(w_mem_inst__abc_19396_new_n3619_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf13), .Y(w_mem_inst__abc_19396_new_n3620_));
OAI21X1 OAI21X1_1773 ( .A(w_mem_inst_w_mem_9__11_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf12), .C(w_mem_inst__abc_19396_new_n3620_), .Y(w_mem_inst__abc_19396_new_n3621_));
OAI21X1 OAI21X1_1774 ( .A(w_mem_inst__abc_19396_new_n1898_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf8), .C(w_mem_inst__abc_19396_new_n3621_), .Y(w_mem_inst__0w_mem_8__31_0__11_));
OAI21X1 OAI21X1_1775 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf6), .B(w_mem_inst__abc_19396_new_n3623_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf11), .Y(w_mem_inst__abc_19396_new_n3624_));
OAI21X1 OAI21X1_1776 ( .A(w_mem_inst_w_mem_9__12_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf10), .C(w_mem_inst__abc_19396_new_n3624_), .Y(w_mem_inst__abc_19396_new_n3625_));
OAI21X1 OAI21X1_1777 ( .A(w_mem_inst__abc_19396_new_n1923_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf7), .C(w_mem_inst__abc_19396_new_n3625_), .Y(w_mem_inst__0w_mem_8__31_0__12_));
OAI21X1 OAI21X1_1778 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf5), .B(w_mem_inst__abc_19396_new_n3627_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf9), .Y(w_mem_inst__abc_19396_new_n3628_));
OAI21X1 OAI21X1_1779 ( .A(w_mem_inst_w_mem_9__13_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf8), .C(w_mem_inst__abc_19396_new_n3628_), .Y(w_mem_inst__abc_19396_new_n3629_));
OAI21X1 OAI21X1_178 ( .A(round_ctr_inc_bF_buf6), .B(_abc_15497_new_n1662_), .C(_abc_15497_new_n1664_), .Y(_0e_reg_31_0__4_));
OAI21X1 OAI21X1_1780 ( .A(w_mem_inst__abc_19396_new_n1948_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf6), .C(w_mem_inst__abc_19396_new_n3629_), .Y(w_mem_inst__0w_mem_8__31_0__13_));
OAI21X1 OAI21X1_1781 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf4), .B(w_mem_inst__abc_19396_new_n3631_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf7), .Y(w_mem_inst__abc_19396_new_n3632_));
OAI21X1 OAI21X1_1782 ( .A(w_mem_inst_w_mem_9__14_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf6), .C(w_mem_inst__abc_19396_new_n3632_), .Y(w_mem_inst__abc_19396_new_n3633_));
OAI21X1 OAI21X1_1783 ( .A(w_mem_inst__abc_19396_new_n1973_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf5), .C(w_mem_inst__abc_19396_new_n3633_), .Y(w_mem_inst__0w_mem_8__31_0__14_));
OAI21X1 OAI21X1_1784 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf3), .B(w_mem_inst__abc_19396_new_n3635_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf5), .Y(w_mem_inst__abc_19396_new_n3636_));
OAI21X1 OAI21X1_1785 ( .A(w_mem_inst_w_mem_9__15_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf4), .C(w_mem_inst__abc_19396_new_n3636_), .Y(w_mem_inst__abc_19396_new_n3637_));
OAI21X1 OAI21X1_1786 ( .A(w_mem_inst__abc_19396_new_n1998_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf4), .C(w_mem_inst__abc_19396_new_n3637_), .Y(w_mem_inst__0w_mem_8__31_0__15_));
OAI21X1 OAI21X1_1787 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf2), .B(w_mem_inst__abc_19396_new_n3639_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf3), .Y(w_mem_inst__abc_19396_new_n3640_));
OAI21X1 OAI21X1_1788 ( .A(w_mem_inst_w_mem_9__16_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf2), .C(w_mem_inst__abc_19396_new_n3640_), .Y(w_mem_inst__abc_19396_new_n3641_));
OAI21X1 OAI21X1_1789 ( .A(w_mem_inst__abc_19396_new_n2023_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf3), .C(w_mem_inst__abc_19396_new_n3641_), .Y(w_mem_inst__0w_mem_8__31_0__16_));
OAI21X1 OAI21X1_179 ( .A(_auto_iopadmap_cc_368_execute_22625_5_), .B(_abc_15497_new_n883__bF_buf5), .C(round_ctr_rst_bF_buf7), .Y(_abc_15497_new_n1666_));
OAI21X1 OAI21X1_1790 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf1), .B(w_mem_inst__abc_19396_new_n3643_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf1), .Y(w_mem_inst__abc_19396_new_n3644_));
OAI21X1 OAI21X1_1791 ( .A(w_mem_inst_w_mem_9__17_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf0), .C(w_mem_inst__abc_19396_new_n3644_), .Y(w_mem_inst__abc_19396_new_n3645_));
OAI21X1 OAI21X1_1792 ( .A(w_mem_inst__abc_19396_new_n2048_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf2), .C(w_mem_inst__abc_19396_new_n3645_), .Y(w_mem_inst__0w_mem_8__31_0__17_));
OAI21X1 OAI21X1_1793 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf0), .B(w_mem_inst__abc_19396_new_n3647_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf96), .Y(w_mem_inst__abc_19396_new_n3648_));
OAI21X1 OAI21X1_1794 ( .A(w_mem_inst_w_mem_9__18_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf95), .C(w_mem_inst__abc_19396_new_n3648_), .Y(w_mem_inst__abc_19396_new_n3649_));
OAI21X1 OAI21X1_1795 ( .A(w_mem_inst__abc_19396_new_n2073_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf1), .C(w_mem_inst__abc_19396_new_n3649_), .Y(w_mem_inst__0w_mem_8__31_0__18_));
OAI21X1 OAI21X1_1796 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf60), .B(w_mem_inst__abc_19396_new_n3651_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf94), .Y(w_mem_inst__abc_19396_new_n3652_));
OAI21X1 OAI21X1_1797 ( .A(w_mem_inst_w_mem_9__19_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf93), .C(w_mem_inst__abc_19396_new_n3652_), .Y(w_mem_inst__abc_19396_new_n3653_));
OAI21X1 OAI21X1_1798 ( .A(w_mem_inst__abc_19396_new_n2098_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf0), .C(w_mem_inst__abc_19396_new_n3653_), .Y(w_mem_inst__0w_mem_8__31_0__19_));
OAI21X1 OAI21X1_1799 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf59), .B(w_mem_inst__abc_19396_new_n3655_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf92), .Y(w_mem_inst__abc_19396_new_n3656_));
OAI21X1 OAI21X1_18 ( .A(_abc_15497_new_n894_), .B(_abc_15497_new_n903_), .C(_abc_15497_new_n915_), .Y(_abc_15497_new_n916_));
OAI21X1 OAI21X1_180 ( .A(round_ctr_inc_bF_buf4), .B(_abc_15497_new_n1666_), .C(_abc_15497_new_n1667_), .Y(_0e_reg_31_0__5_));
OAI21X1 OAI21X1_1800 ( .A(w_mem_inst_w_mem_9__20_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf91), .C(w_mem_inst__abc_19396_new_n3656_), .Y(w_mem_inst__abc_19396_new_n3657_));
OAI21X1 OAI21X1_1801 ( .A(w_mem_inst__abc_19396_new_n2123_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf60), .C(w_mem_inst__abc_19396_new_n3657_), .Y(w_mem_inst__0w_mem_8__31_0__20_));
OAI21X1 OAI21X1_1802 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf58), .B(w_mem_inst__abc_19396_new_n3659_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf90), .Y(w_mem_inst__abc_19396_new_n3660_));
OAI21X1 OAI21X1_1803 ( .A(w_mem_inst_w_mem_9__21_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf89), .C(w_mem_inst__abc_19396_new_n3660_), .Y(w_mem_inst__abc_19396_new_n3661_));
OAI21X1 OAI21X1_1804 ( .A(w_mem_inst__abc_19396_new_n2148_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf59), .C(w_mem_inst__abc_19396_new_n3661_), .Y(w_mem_inst__0w_mem_8__31_0__21_));
OAI21X1 OAI21X1_1805 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf57), .B(w_mem_inst__abc_19396_new_n3663_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf88), .Y(w_mem_inst__abc_19396_new_n3664_));
OAI21X1 OAI21X1_1806 ( .A(w_mem_inst_w_mem_9__22_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf87), .C(w_mem_inst__abc_19396_new_n3664_), .Y(w_mem_inst__abc_19396_new_n3665_));
OAI21X1 OAI21X1_1807 ( .A(w_mem_inst__abc_19396_new_n2173_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf58), .C(w_mem_inst__abc_19396_new_n3665_), .Y(w_mem_inst__0w_mem_8__31_0__22_));
OAI21X1 OAI21X1_1808 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf56), .B(w_mem_inst__abc_19396_new_n3667_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf86), .Y(w_mem_inst__abc_19396_new_n3668_));
OAI21X1 OAI21X1_1809 ( .A(w_mem_inst_w_mem_9__23_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf85), .C(w_mem_inst__abc_19396_new_n3668_), .Y(w_mem_inst__abc_19396_new_n3669_));
OAI21X1 OAI21X1_181 ( .A(_auto_iopadmap_cc_368_execute_22625_6_), .B(_abc_15497_new_n883__bF_buf4), .C(round_ctr_rst_bF_buf6), .Y(_abc_15497_new_n1669_));
OAI21X1 OAI21X1_1810 ( .A(w_mem_inst__abc_19396_new_n2198_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf57), .C(w_mem_inst__abc_19396_new_n3669_), .Y(w_mem_inst__0w_mem_8__31_0__23_));
OAI21X1 OAI21X1_1811 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf55), .B(w_mem_inst__abc_19396_new_n3671_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf84), .Y(w_mem_inst__abc_19396_new_n3672_));
OAI21X1 OAI21X1_1812 ( .A(w_mem_inst_w_mem_9__24_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf83), .C(w_mem_inst__abc_19396_new_n3672_), .Y(w_mem_inst__abc_19396_new_n3673_));
OAI21X1 OAI21X1_1813 ( .A(w_mem_inst__abc_19396_new_n2223_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf56), .C(w_mem_inst__abc_19396_new_n3673_), .Y(w_mem_inst__0w_mem_8__31_0__24_));
OAI21X1 OAI21X1_1814 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf54), .B(w_mem_inst__abc_19396_new_n3675_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf82), .Y(w_mem_inst__abc_19396_new_n3676_));
OAI21X1 OAI21X1_1815 ( .A(w_mem_inst_w_mem_9__25_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf81), .C(w_mem_inst__abc_19396_new_n3676_), .Y(w_mem_inst__abc_19396_new_n3677_));
OAI21X1 OAI21X1_1816 ( .A(w_mem_inst__abc_19396_new_n2248_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf55), .C(w_mem_inst__abc_19396_new_n3677_), .Y(w_mem_inst__0w_mem_8__31_0__25_));
OAI21X1 OAI21X1_1817 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf53), .B(w_mem_inst__abc_19396_new_n3679_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf80), .Y(w_mem_inst__abc_19396_new_n3680_));
OAI21X1 OAI21X1_1818 ( .A(w_mem_inst_w_mem_9__26_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf79), .C(w_mem_inst__abc_19396_new_n3680_), .Y(w_mem_inst__abc_19396_new_n3681_));
OAI21X1 OAI21X1_1819 ( .A(w_mem_inst__abc_19396_new_n2273_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf54), .C(w_mem_inst__abc_19396_new_n3681_), .Y(w_mem_inst__0w_mem_8__31_0__26_));
OAI21X1 OAI21X1_182 ( .A(round_ctr_inc_bF_buf2), .B(_abc_15497_new_n1669_), .C(_abc_15497_new_n1670_), .Y(_0e_reg_31_0__6_));
OAI21X1 OAI21X1_1820 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf52), .B(w_mem_inst__abc_19396_new_n3683_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf78), .Y(w_mem_inst__abc_19396_new_n3684_));
OAI21X1 OAI21X1_1821 ( .A(w_mem_inst_w_mem_9__27_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf77), .C(w_mem_inst__abc_19396_new_n3684_), .Y(w_mem_inst__abc_19396_new_n3685_));
OAI21X1 OAI21X1_1822 ( .A(w_mem_inst__abc_19396_new_n2298_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf53), .C(w_mem_inst__abc_19396_new_n3685_), .Y(w_mem_inst__0w_mem_8__31_0__27_));
OAI21X1 OAI21X1_1823 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf51), .B(w_mem_inst__abc_19396_new_n3687_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf76), .Y(w_mem_inst__abc_19396_new_n3688_));
OAI21X1 OAI21X1_1824 ( .A(w_mem_inst_w_mem_9__28_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf75), .C(w_mem_inst__abc_19396_new_n3688_), .Y(w_mem_inst__abc_19396_new_n3689_));
OAI21X1 OAI21X1_1825 ( .A(w_mem_inst__abc_19396_new_n2323_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf52), .C(w_mem_inst__abc_19396_new_n3689_), .Y(w_mem_inst__0w_mem_8__31_0__28_));
OAI21X1 OAI21X1_1826 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf50), .B(w_mem_inst__abc_19396_new_n3691_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf74), .Y(w_mem_inst__abc_19396_new_n3692_));
OAI21X1 OAI21X1_1827 ( .A(w_mem_inst_w_mem_9__29_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf73), .C(w_mem_inst__abc_19396_new_n3692_), .Y(w_mem_inst__abc_19396_new_n3693_));
OAI21X1 OAI21X1_1828 ( .A(w_mem_inst__abc_19396_new_n2348_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf51), .C(w_mem_inst__abc_19396_new_n3693_), .Y(w_mem_inst__0w_mem_8__31_0__29_));
OAI21X1 OAI21X1_1829 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf49), .B(w_mem_inst__abc_19396_new_n3695_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf72), .Y(w_mem_inst__abc_19396_new_n3696_));
OAI21X1 OAI21X1_183 ( .A(_auto_iopadmap_cc_368_execute_22625_7_), .B(_abc_15497_new_n883__bF_buf3), .C(round_ctr_rst_bF_buf5), .Y(_abc_15497_new_n1672_));
OAI21X1 OAI21X1_1830 ( .A(w_mem_inst_w_mem_9__30_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf71), .C(w_mem_inst__abc_19396_new_n3696_), .Y(w_mem_inst__abc_19396_new_n3697_));
OAI21X1 OAI21X1_1831 ( .A(w_mem_inst__abc_19396_new_n2373_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf50), .C(w_mem_inst__abc_19396_new_n3697_), .Y(w_mem_inst__0w_mem_8__31_0__30_));
OAI21X1 OAI21X1_1832 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf48), .B(w_mem_inst__abc_19396_new_n3699_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf70), .Y(w_mem_inst__abc_19396_new_n3700_));
OAI21X1 OAI21X1_1833 ( .A(w_mem_inst_w_mem_9__31_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf69), .C(w_mem_inst__abc_19396_new_n3700_), .Y(w_mem_inst__abc_19396_new_n3701_));
OAI21X1 OAI21X1_1834 ( .A(w_mem_inst__abc_19396_new_n2398_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf49), .C(w_mem_inst__abc_19396_new_n3701_), .Y(w_mem_inst__0w_mem_8__31_0__31_));
OAI21X1 OAI21X1_1835 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf47), .B(w_mem_inst__abc_19396_new_n3704_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf68), .Y(w_mem_inst__abc_19396_new_n3705_));
OAI21X1 OAI21X1_1836 ( .A(w_mem_inst_w_mem_5__0_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf67), .C(w_mem_inst__abc_19396_new_n3705_), .Y(w_mem_inst__abc_19396_new_n3706_));
OAI21X1 OAI21X1_1837 ( .A(w_mem_inst__abc_19396_new_n3703_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf48), .C(w_mem_inst__abc_19396_new_n3706_), .Y(w_mem_inst__0w_mem_4__31_0__0_));
OAI21X1 OAI21X1_1838 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf46), .B(w_mem_inst__abc_19396_new_n3709_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf66), .Y(w_mem_inst__abc_19396_new_n3710_));
OAI21X1 OAI21X1_1839 ( .A(w_mem_inst_w_mem_5__1_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf65), .C(w_mem_inst__abc_19396_new_n3710_), .Y(w_mem_inst__abc_19396_new_n3711_));
OAI21X1 OAI21X1_184 ( .A(round_ctr_inc_bF_buf0), .B(_abc_15497_new_n1672_), .C(_abc_15497_new_n1673_), .Y(_0e_reg_31_0__7_));
OAI21X1 OAI21X1_1840 ( .A(w_mem_inst__abc_19396_new_n3708_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf47), .C(w_mem_inst__abc_19396_new_n3711_), .Y(w_mem_inst__0w_mem_4__31_0__1_));
OAI21X1 OAI21X1_1841 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf45), .B(w_mem_inst__abc_19396_new_n3714_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf64), .Y(w_mem_inst__abc_19396_new_n3715_));
OAI21X1 OAI21X1_1842 ( .A(w_mem_inst_w_mem_5__2_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf63), .C(w_mem_inst__abc_19396_new_n3715_), .Y(w_mem_inst__abc_19396_new_n3716_));
OAI21X1 OAI21X1_1843 ( .A(w_mem_inst__abc_19396_new_n3713_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf46), .C(w_mem_inst__abc_19396_new_n3716_), .Y(w_mem_inst__0w_mem_4__31_0__2_));
OAI21X1 OAI21X1_1844 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf44), .B(w_mem_inst__abc_19396_new_n3719_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf62), .Y(w_mem_inst__abc_19396_new_n3720_));
OAI21X1 OAI21X1_1845 ( .A(w_mem_inst_w_mem_5__3_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf61), .C(w_mem_inst__abc_19396_new_n3720_), .Y(w_mem_inst__abc_19396_new_n3721_));
OAI21X1 OAI21X1_1846 ( .A(w_mem_inst__abc_19396_new_n3718_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf45), .C(w_mem_inst__abc_19396_new_n3721_), .Y(w_mem_inst__0w_mem_4__31_0__3_));
OAI21X1 OAI21X1_1847 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf43), .B(w_mem_inst__abc_19396_new_n3724_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf60), .Y(w_mem_inst__abc_19396_new_n3725_));
OAI21X1 OAI21X1_1848 ( .A(w_mem_inst_w_mem_5__4_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf59), .C(w_mem_inst__abc_19396_new_n3725_), .Y(w_mem_inst__abc_19396_new_n3726_));
OAI21X1 OAI21X1_1849 ( .A(w_mem_inst__abc_19396_new_n3723_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf44), .C(w_mem_inst__abc_19396_new_n3726_), .Y(w_mem_inst__0w_mem_4__31_0__4_));
OAI21X1 OAI21X1_185 ( .A(_abc_15497_new_n871__bF_buf4), .B(_abc_15497_new_n872__bF_buf0), .C(_abc_15497_new_n1007_), .Y(_abc_15497_new_n1675_));
OAI21X1 OAI21X1_1850 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf42), .B(w_mem_inst__abc_19396_new_n3729_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf58), .Y(w_mem_inst__abc_19396_new_n3730_));
OAI21X1 OAI21X1_1851 ( .A(w_mem_inst_w_mem_5__5_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf57), .C(w_mem_inst__abc_19396_new_n3730_), .Y(w_mem_inst__abc_19396_new_n3731_));
OAI21X1 OAI21X1_1852 ( .A(w_mem_inst__abc_19396_new_n3728_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf43), .C(w_mem_inst__abc_19396_new_n3731_), .Y(w_mem_inst__0w_mem_4__31_0__5_));
OAI21X1 OAI21X1_1853 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf41), .B(w_mem_inst__abc_19396_new_n3734_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf56), .Y(w_mem_inst__abc_19396_new_n3735_));
OAI21X1 OAI21X1_1854 ( .A(w_mem_inst_w_mem_5__6_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf55), .C(w_mem_inst__abc_19396_new_n3735_), .Y(w_mem_inst__abc_19396_new_n3736_));
OAI21X1 OAI21X1_1855 ( .A(w_mem_inst__abc_19396_new_n3733_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf42), .C(w_mem_inst__abc_19396_new_n3736_), .Y(w_mem_inst__0w_mem_4__31_0__6_));
OAI21X1 OAI21X1_1856 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf40), .B(w_mem_inst__abc_19396_new_n3739_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf54), .Y(w_mem_inst__abc_19396_new_n3740_));
OAI21X1 OAI21X1_1857 ( .A(w_mem_inst_w_mem_5__7_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf53), .C(w_mem_inst__abc_19396_new_n3740_), .Y(w_mem_inst__abc_19396_new_n3741_));
OAI21X1 OAI21X1_1858 ( .A(w_mem_inst__abc_19396_new_n3738_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf41), .C(w_mem_inst__abc_19396_new_n3741_), .Y(w_mem_inst__0w_mem_4__31_0__7_));
OAI21X1 OAI21X1_1859 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf39), .B(w_mem_inst__abc_19396_new_n3744_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf52), .Y(w_mem_inst__abc_19396_new_n3745_));
OAI21X1 OAI21X1_186 ( .A(_abc_15497_new_n1006_), .B(_abc_15497_new_n1648__bF_buf3), .C(_abc_15497_new_n1676_), .Y(_0e_reg_31_0__8_));
OAI21X1 OAI21X1_1860 ( .A(w_mem_inst_w_mem_5__8_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf51), .C(w_mem_inst__abc_19396_new_n3745_), .Y(w_mem_inst__abc_19396_new_n3746_));
OAI21X1 OAI21X1_1861 ( .A(w_mem_inst__abc_19396_new_n3743_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf40), .C(w_mem_inst__abc_19396_new_n3746_), .Y(w_mem_inst__0w_mem_4__31_0__8_));
OAI21X1 OAI21X1_1862 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf38), .B(w_mem_inst__abc_19396_new_n3749_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf50), .Y(w_mem_inst__abc_19396_new_n3750_));
OAI21X1 OAI21X1_1863 ( .A(w_mem_inst_w_mem_5__9_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf49), .C(w_mem_inst__abc_19396_new_n3750_), .Y(w_mem_inst__abc_19396_new_n3751_));
OAI21X1 OAI21X1_1864 ( .A(w_mem_inst__abc_19396_new_n3748_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf39), .C(w_mem_inst__abc_19396_new_n3751_), .Y(w_mem_inst__0w_mem_4__31_0__9_));
OAI21X1 OAI21X1_1865 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf37), .B(w_mem_inst__abc_19396_new_n3754_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf48), .Y(w_mem_inst__abc_19396_new_n3755_));
OAI21X1 OAI21X1_1866 ( .A(w_mem_inst_w_mem_5__10_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf47), .C(w_mem_inst__abc_19396_new_n3755_), .Y(w_mem_inst__abc_19396_new_n3756_));
OAI21X1 OAI21X1_1867 ( .A(w_mem_inst__abc_19396_new_n3753_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf38), .C(w_mem_inst__abc_19396_new_n3756_), .Y(w_mem_inst__0w_mem_4__31_0__10_));
OAI21X1 OAI21X1_1868 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf36), .B(w_mem_inst__abc_19396_new_n3759_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf46), .Y(w_mem_inst__abc_19396_new_n3760_));
OAI21X1 OAI21X1_1869 ( .A(w_mem_inst_w_mem_5__11_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf45), .C(w_mem_inst__abc_19396_new_n3760_), .Y(w_mem_inst__abc_19396_new_n3761_));
OAI21X1 OAI21X1_187 ( .A(_abc_15497_new_n1034_), .B(_abc_15497_new_n1648__bF_buf2), .C(_abc_15497_new_n1679_), .Y(_0e_reg_31_0__9_));
OAI21X1 OAI21X1_1870 ( .A(w_mem_inst__abc_19396_new_n3758_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf37), .C(w_mem_inst__abc_19396_new_n3761_), .Y(w_mem_inst__0w_mem_4__31_0__11_));
OAI21X1 OAI21X1_1871 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf35), .B(w_mem_inst__abc_19396_new_n3764_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf44), .Y(w_mem_inst__abc_19396_new_n3765_));
OAI21X1 OAI21X1_1872 ( .A(w_mem_inst_w_mem_5__12_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf43), .C(w_mem_inst__abc_19396_new_n3765_), .Y(w_mem_inst__abc_19396_new_n3766_));
OAI21X1 OAI21X1_1873 ( .A(w_mem_inst__abc_19396_new_n3763_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf36), .C(w_mem_inst__abc_19396_new_n3766_), .Y(w_mem_inst__0w_mem_4__31_0__12_));
OAI21X1 OAI21X1_1874 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf34), .B(w_mem_inst__abc_19396_new_n3769_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf42), .Y(w_mem_inst__abc_19396_new_n3770_));
OAI21X1 OAI21X1_1875 ( .A(w_mem_inst_w_mem_5__13_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf41), .C(w_mem_inst__abc_19396_new_n3770_), .Y(w_mem_inst__abc_19396_new_n3771_));
OAI21X1 OAI21X1_1876 ( .A(w_mem_inst__abc_19396_new_n3768_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf35), .C(w_mem_inst__abc_19396_new_n3771_), .Y(w_mem_inst__0w_mem_4__31_0__13_));
OAI21X1 OAI21X1_1877 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf33), .B(w_mem_inst__abc_19396_new_n3774_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf40), .Y(w_mem_inst__abc_19396_new_n3775_));
OAI21X1 OAI21X1_1878 ( .A(w_mem_inst_w_mem_5__14_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf39), .C(w_mem_inst__abc_19396_new_n3775_), .Y(w_mem_inst__abc_19396_new_n3776_));
OAI21X1 OAI21X1_1879 ( .A(w_mem_inst__abc_19396_new_n3773_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf34), .C(w_mem_inst__abc_19396_new_n3776_), .Y(w_mem_inst__0w_mem_4__31_0__14_));
OAI21X1 OAI21X1_188 ( .A(_abc_15497_new_n1049_), .B(_abc_15497_new_n1648__bF_buf1), .C(_abc_15497_new_n1682_), .Y(_0e_reg_31_0__10_));
OAI21X1 OAI21X1_1880 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf32), .B(w_mem_inst__abc_19396_new_n3779_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf38), .Y(w_mem_inst__abc_19396_new_n3780_));
OAI21X1 OAI21X1_1881 ( .A(w_mem_inst_w_mem_5__15_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf37), .C(w_mem_inst__abc_19396_new_n3780_), .Y(w_mem_inst__abc_19396_new_n3781_));
OAI21X1 OAI21X1_1882 ( .A(w_mem_inst__abc_19396_new_n3778_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf33), .C(w_mem_inst__abc_19396_new_n3781_), .Y(w_mem_inst__0w_mem_4__31_0__15_));
OAI21X1 OAI21X1_1883 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf31), .B(w_mem_inst__abc_19396_new_n3784_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf36), .Y(w_mem_inst__abc_19396_new_n3785_));
OAI21X1 OAI21X1_1884 ( .A(w_mem_inst_w_mem_5__16_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf35), .C(w_mem_inst__abc_19396_new_n3785_), .Y(w_mem_inst__abc_19396_new_n3786_));
OAI21X1 OAI21X1_1885 ( .A(w_mem_inst__abc_19396_new_n3783_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf32), .C(w_mem_inst__abc_19396_new_n3786_), .Y(w_mem_inst__0w_mem_4__31_0__16_));
OAI21X1 OAI21X1_1886 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf30), .B(w_mem_inst__abc_19396_new_n3789_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf34), .Y(w_mem_inst__abc_19396_new_n3790_));
OAI21X1 OAI21X1_1887 ( .A(w_mem_inst_w_mem_5__17_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf33), .C(w_mem_inst__abc_19396_new_n3790_), .Y(w_mem_inst__abc_19396_new_n3791_));
OAI21X1 OAI21X1_1888 ( .A(w_mem_inst__abc_19396_new_n3788_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf31), .C(w_mem_inst__abc_19396_new_n3791_), .Y(w_mem_inst__0w_mem_4__31_0__17_));
OAI21X1 OAI21X1_1889 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf29), .B(w_mem_inst__abc_19396_new_n3794_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf32), .Y(w_mem_inst__abc_19396_new_n3795_));
OAI21X1 OAI21X1_189 ( .A(_abc_15497_new_n1684_), .B(_abc_15497_new_n1648__bF_buf0), .C(_abc_15497_new_n1686_), .Y(_0e_reg_31_0__11_));
OAI21X1 OAI21X1_1890 ( .A(w_mem_inst_w_mem_5__18_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf31), .C(w_mem_inst__abc_19396_new_n3795_), .Y(w_mem_inst__abc_19396_new_n3796_));
OAI21X1 OAI21X1_1891 ( .A(w_mem_inst__abc_19396_new_n3793_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf30), .C(w_mem_inst__abc_19396_new_n3796_), .Y(w_mem_inst__0w_mem_4__31_0__18_));
OAI21X1 OAI21X1_1892 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf28), .B(w_mem_inst__abc_19396_new_n3799_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf30), .Y(w_mem_inst__abc_19396_new_n3800_));
OAI21X1 OAI21X1_1893 ( .A(w_mem_inst_w_mem_5__19_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf29), .C(w_mem_inst__abc_19396_new_n3800_), .Y(w_mem_inst__abc_19396_new_n3801_));
OAI21X1 OAI21X1_1894 ( .A(w_mem_inst__abc_19396_new_n3798_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf29), .C(w_mem_inst__abc_19396_new_n3801_), .Y(w_mem_inst__0w_mem_4__31_0__19_));
OAI21X1 OAI21X1_1895 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf27), .B(w_mem_inst__abc_19396_new_n3804_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf28), .Y(w_mem_inst__abc_19396_new_n3805_));
OAI21X1 OAI21X1_1896 ( .A(w_mem_inst_w_mem_5__20_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf27), .C(w_mem_inst__abc_19396_new_n3805_), .Y(w_mem_inst__abc_19396_new_n3806_));
OAI21X1 OAI21X1_1897 ( .A(w_mem_inst__abc_19396_new_n3803_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf28), .C(w_mem_inst__abc_19396_new_n3806_), .Y(w_mem_inst__0w_mem_4__31_0__20_));
OAI21X1 OAI21X1_1898 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf26), .B(w_mem_inst__abc_19396_new_n3809_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf26), .Y(w_mem_inst__abc_19396_new_n3810_));
OAI21X1 OAI21X1_1899 ( .A(w_mem_inst_w_mem_5__21_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf25), .C(w_mem_inst__abc_19396_new_n3810_), .Y(w_mem_inst__abc_19396_new_n3811_));
OAI21X1 OAI21X1_19 ( .A(_abc_15497_new_n903_), .B(_abc_15497_new_n902_), .C(_abc_15497_new_n915_), .Y(_abc_15497_new_n922_));
OAI21X1 OAI21X1_190 ( .A(_abc_15497_new_n1064_), .B(_abc_15497_new_n1648__bF_buf8), .C(_abc_15497_new_n1689_), .Y(_0e_reg_31_0__12_));
OAI21X1 OAI21X1_1900 ( .A(w_mem_inst__abc_19396_new_n3808_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf27), .C(w_mem_inst__abc_19396_new_n3811_), .Y(w_mem_inst__0w_mem_4__31_0__21_));
OAI21X1 OAI21X1_1901 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf25), .B(w_mem_inst__abc_19396_new_n3814_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf24), .Y(w_mem_inst__abc_19396_new_n3815_));
OAI21X1 OAI21X1_1902 ( .A(w_mem_inst_w_mem_5__22_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf23), .C(w_mem_inst__abc_19396_new_n3815_), .Y(w_mem_inst__abc_19396_new_n3816_));
OAI21X1 OAI21X1_1903 ( .A(w_mem_inst__abc_19396_new_n3813_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf26), .C(w_mem_inst__abc_19396_new_n3816_), .Y(w_mem_inst__0w_mem_4__31_0__22_));
OAI21X1 OAI21X1_1904 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf24), .B(w_mem_inst__abc_19396_new_n3819_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf22), .Y(w_mem_inst__abc_19396_new_n3820_));
OAI21X1 OAI21X1_1905 ( .A(w_mem_inst_w_mem_5__23_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf21), .C(w_mem_inst__abc_19396_new_n3820_), .Y(w_mem_inst__abc_19396_new_n3821_));
OAI21X1 OAI21X1_1906 ( .A(w_mem_inst__abc_19396_new_n3818_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf25), .C(w_mem_inst__abc_19396_new_n3821_), .Y(w_mem_inst__0w_mem_4__31_0__23_));
OAI21X1 OAI21X1_1907 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf23), .B(w_mem_inst__abc_19396_new_n3824_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf20), .Y(w_mem_inst__abc_19396_new_n3825_));
OAI21X1 OAI21X1_1908 ( .A(w_mem_inst_w_mem_5__24_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf19), .C(w_mem_inst__abc_19396_new_n3825_), .Y(w_mem_inst__abc_19396_new_n3826_));
OAI21X1 OAI21X1_1909 ( .A(w_mem_inst__abc_19396_new_n3823_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf24), .C(w_mem_inst__abc_19396_new_n3826_), .Y(w_mem_inst__0w_mem_4__31_0__24_));
OAI21X1 OAI21X1_191 ( .A(_auto_iopadmap_cc_368_execute_22625_13_), .B(_abc_15497_new_n883__bF_buf12), .C(round_ctr_rst_bF_buf4), .Y(_abc_15497_new_n1691_));
OAI21X1 OAI21X1_1910 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf22), .B(w_mem_inst__abc_19396_new_n3829_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf18), .Y(w_mem_inst__abc_19396_new_n3830_));
OAI21X1 OAI21X1_1911 ( .A(w_mem_inst_w_mem_5__25_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf17), .C(w_mem_inst__abc_19396_new_n3830_), .Y(w_mem_inst__abc_19396_new_n3831_));
OAI21X1 OAI21X1_1912 ( .A(w_mem_inst__abc_19396_new_n3828_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf23), .C(w_mem_inst__abc_19396_new_n3831_), .Y(w_mem_inst__0w_mem_4__31_0__25_));
OAI21X1 OAI21X1_1913 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf21), .B(w_mem_inst__abc_19396_new_n3834_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf16), .Y(w_mem_inst__abc_19396_new_n3835_));
OAI21X1 OAI21X1_1914 ( .A(w_mem_inst_w_mem_5__26_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf15), .C(w_mem_inst__abc_19396_new_n3835_), .Y(w_mem_inst__abc_19396_new_n3836_));
OAI21X1 OAI21X1_1915 ( .A(w_mem_inst__abc_19396_new_n3833_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf22), .C(w_mem_inst__abc_19396_new_n3836_), .Y(w_mem_inst__0w_mem_4__31_0__26_));
OAI21X1 OAI21X1_1916 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf20), .B(w_mem_inst__abc_19396_new_n3839_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf14), .Y(w_mem_inst__abc_19396_new_n3840_));
OAI21X1 OAI21X1_1917 ( .A(w_mem_inst_w_mem_5__27_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf13), .C(w_mem_inst__abc_19396_new_n3840_), .Y(w_mem_inst__abc_19396_new_n3841_));
OAI21X1 OAI21X1_1918 ( .A(w_mem_inst__abc_19396_new_n3838_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf21), .C(w_mem_inst__abc_19396_new_n3841_), .Y(w_mem_inst__0w_mem_4__31_0__27_));
OAI21X1 OAI21X1_1919 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf19), .B(w_mem_inst__abc_19396_new_n3844_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf12), .Y(w_mem_inst__abc_19396_new_n3845_));
OAI21X1 OAI21X1_192 ( .A(round_ctr_inc_bF_buf7), .B(_abc_15497_new_n1691_), .C(_abc_15497_new_n1692_), .Y(_0e_reg_31_0__13_));
OAI21X1 OAI21X1_1920 ( .A(w_mem_inst_w_mem_5__28_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf11), .C(w_mem_inst__abc_19396_new_n3845_), .Y(w_mem_inst__abc_19396_new_n3846_));
OAI21X1 OAI21X1_1921 ( .A(w_mem_inst__abc_19396_new_n3843_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf20), .C(w_mem_inst__abc_19396_new_n3846_), .Y(w_mem_inst__0w_mem_4__31_0__28_));
OAI21X1 OAI21X1_1922 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf18), .B(w_mem_inst__abc_19396_new_n3849_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf10), .Y(w_mem_inst__abc_19396_new_n3850_));
OAI21X1 OAI21X1_1923 ( .A(w_mem_inst_w_mem_5__29_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf9), .C(w_mem_inst__abc_19396_new_n3850_), .Y(w_mem_inst__abc_19396_new_n3851_));
OAI21X1 OAI21X1_1924 ( .A(w_mem_inst__abc_19396_new_n3848_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf19), .C(w_mem_inst__abc_19396_new_n3851_), .Y(w_mem_inst__0w_mem_4__31_0__29_));
OAI21X1 OAI21X1_1925 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf17), .B(w_mem_inst__abc_19396_new_n3854_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf8), .Y(w_mem_inst__abc_19396_new_n3855_));
OAI21X1 OAI21X1_1926 ( .A(w_mem_inst_w_mem_5__30_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf7), .C(w_mem_inst__abc_19396_new_n3855_), .Y(w_mem_inst__abc_19396_new_n3856_));
OAI21X1 OAI21X1_1927 ( .A(w_mem_inst__abc_19396_new_n3853_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf18), .C(w_mem_inst__abc_19396_new_n3856_), .Y(w_mem_inst__0w_mem_4__31_0__30_));
OAI21X1 OAI21X1_1928 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf16), .B(w_mem_inst__abc_19396_new_n3859_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf6), .Y(w_mem_inst__abc_19396_new_n3860_));
OAI21X1 OAI21X1_1929 ( .A(w_mem_inst_w_mem_5__31_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf5), .C(w_mem_inst__abc_19396_new_n3860_), .Y(w_mem_inst__abc_19396_new_n3861_));
OAI21X1 OAI21X1_193 ( .A(_abc_15497_new_n871__bF_buf3), .B(_abc_15497_new_n872__bF_buf4), .C(_abc_15497_new_n1081_), .Y(_abc_15497_new_n1694_));
OAI21X1 OAI21X1_1930 ( .A(w_mem_inst__abc_19396_new_n3858_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf17), .C(w_mem_inst__abc_19396_new_n3861_), .Y(w_mem_inst__0w_mem_4__31_0__31_));
OAI21X1 OAI21X1_1931 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf15), .B(w_mem_inst__abc_19396_new_n3864_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf4), .Y(w_mem_inst__abc_19396_new_n3865_));
OAI21X1 OAI21X1_1932 ( .A(w_mem_inst_w_mem_7__0_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf3), .C(w_mem_inst__abc_19396_new_n3865_), .Y(w_mem_inst__abc_19396_new_n3866_));
OAI21X1 OAI21X1_1933 ( .A(w_mem_inst__abc_19396_new_n3863_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf16), .C(w_mem_inst__abc_19396_new_n3866_), .Y(w_mem_inst__0w_mem_6__31_0__0_));
OAI21X1 OAI21X1_1934 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf14), .B(w_mem_inst__abc_19396_new_n3869_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf2), .Y(w_mem_inst__abc_19396_new_n3870_));
OAI21X1 OAI21X1_1935 ( .A(w_mem_inst_w_mem_7__1_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf1), .C(w_mem_inst__abc_19396_new_n3870_), .Y(w_mem_inst__abc_19396_new_n3871_));
OAI21X1 OAI21X1_1936 ( .A(w_mem_inst__abc_19396_new_n3868_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf15), .C(w_mem_inst__abc_19396_new_n3871_), .Y(w_mem_inst__0w_mem_6__31_0__1_));
OAI21X1 OAI21X1_1937 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf13), .B(w_mem_inst__abc_19396_new_n3874_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf0), .Y(w_mem_inst__abc_19396_new_n3875_));
OAI21X1 OAI21X1_1938 ( .A(w_mem_inst_w_mem_7__2_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf96), .C(w_mem_inst__abc_19396_new_n3875_), .Y(w_mem_inst__abc_19396_new_n3876_));
OAI21X1 OAI21X1_1939 ( .A(w_mem_inst__abc_19396_new_n3873_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf14), .C(w_mem_inst__abc_19396_new_n3876_), .Y(w_mem_inst__0w_mem_6__31_0__2_));
OAI21X1 OAI21X1_194 ( .A(_abc_15497_new_n1080_), .B(_abc_15497_new_n1648__bF_buf7), .C(_abc_15497_new_n1695_), .Y(_0e_reg_31_0__14_));
OAI21X1 OAI21X1_1940 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf12), .B(w_mem_inst__abc_19396_new_n3879_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf95), .Y(w_mem_inst__abc_19396_new_n3880_));
OAI21X1 OAI21X1_1941 ( .A(w_mem_inst_w_mem_7__3_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf94), .C(w_mem_inst__abc_19396_new_n3880_), .Y(w_mem_inst__abc_19396_new_n3881_));
OAI21X1 OAI21X1_1942 ( .A(w_mem_inst__abc_19396_new_n3878_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf13), .C(w_mem_inst__abc_19396_new_n3881_), .Y(w_mem_inst__0w_mem_6__31_0__3_));
OAI21X1 OAI21X1_1943 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf11), .B(w_mem_inst__abc_19396_new_n3884_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf93), .Y(w_mem_inst__abc_19396_new_n3885_));
OAI21X1 OAI21X1_1944 ( .A(w_mem_inst_w_mem_7__4_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf92), .C(w_mem_inst__abc_19396_new_n3885_), .Y(w_mem_inst__abc_19396_new_n3886_));
OAI21X1 OAI21X1_1945 ( .A(w_mem_inst__abc_19396_new_n3883_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf12), .C(w_mem_inst__abc_19396_new_n3886_), .Y(w_mem_inst__0w_mem_6__31_0__4_));
OAI21X1 OAI21X1_1946 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf10), .B(w_mem_inst__abc_19396_new_n3889_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf91), .Y(w_mem_inst__abc_19396_new_n3890_));
OAI21X1 OAI21X1_1947 ( .A(w_mem_inst_w_mem_7__5_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf90), .C(w_mem_inst__abc_19396_new_n3890_), .Y(w_mem_inst__abc_19396_new_n3891_));
OAI21X1 OAI21X1_1948 ( .A(w_mem_inst__abc_19396_new_n3888_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf11), .C(w_mem_inst__abc_19396_new_n3891_), .Y(w_mem_inst__0w_mem_6__31_0__5_));
OAI21X1 OAI21X1_1949 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf9), .B(w_mem_inst__abc_19396_new_n3894_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf89), .Y(w_mem_inst__abc_19396_new_n3895_));
OAI21X1 OAI21X1_195 ( .A(_auto_iopadmap_cc_368_execute_22625_15_), .B(_abc_15497_new_n883__bF_buf11), .C(round_ctr_rst_bF_buf3), .Y(_abc_15497_new_n1697_));
OAI21X1 OAI21X1_1950 ( .A(w_mem_inst_w_mem_7__6_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf88), .C(w_mem_inst__abc_19396_new_n3895_), .Y(w_mem_inst__abc_19396_new_n3896_));
OAI21X1 OAI21X1_1951 ( .A(w_mem_inst__abc_19396_new_n3893_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf10), .C(w_mem_inst__abc_19396_new_n3896_), .Y(w_mem_inst__0w_mem_6__31_0__6_));
OAI21X1 OAI21X1_1952 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf8), .B(w_mem_inst__abc_19396_new_n3899_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf87), .Y(w_mem_inst__abc_19396_new_n3900_));
OAI21X1 OAI21X1_1953 ( .A(w_mem_inst_w_mem_7__7_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf86), .C(w_mem_inst__abc_19396_new_n3900_), .Y(w_mem_inst__abc_19396_new_n3901_));
OAI21X1 OAI21X1_1954 ( .A(w_mem_inst__abc_19396_new_n3898_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf9), .C(w_mem_inst__abc_19396_new_n3901_), .Y(w_mem_inst__0w_mem_6__31_0__7_));
OAI21X1 OAI21X1_1955 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf7), .B(w_mem_inst__abc_19396_new_n3904_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf85), .Y(w_mem_inst__abc_19396_new_n3905_));
OAI21X1 OAI21X1_1956 ( .A(w_mem_inst_w_mem_7__8_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf84), .C(w_mem_inst__abc_19396_new_n3905_), .Y(w_mem_inst__abc_19396_new_n3906_));
OAI21X1 OAI21X1_1957 ( .A(w_mem_inst__abc_19396_new_n3903_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf8), .C(w_mem_inst__abc_19396_new_n3906_), .Y(w_mem_inst__0w_mem_6__31_0__8_));
OAI21X1 OAI21X1_1958 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf6), .B(w_mem_inst__abc_19396_new_n3909_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf83), .Y(w_mem_inst__abc_19396_new_n3910_));
OAI21X1 OAI21X1_1959 ( .A(w_mem_inst_w_mem_7__9_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf82), .C(w_mem_inst__abc_19396_new_n3910_), .Y(w_mem_inst__abc_19396_new_n3911_));
OAI21X1 OAI21X1_196 ( .A(round_ctr_inc_bF_buf4), .B(_abc_15497_new_n1697_), .C(_abc_15497_new_n1698_), .Y(_0e_reg_31_0__15_));
OAI21X1 OAI21X1_1960 ( .A(w_mem_inst__abc_19396_new_n3908_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf7), .C(w_mem_inst__abc_19396_new_n3911_), .Y(w_mem_inst__0w_mem_6__31_0__9_));
OAI21X1 OAI21X1_1961 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf5), .B(w_mem_inst__abc_19396_new_n3914_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf81), .Y(w_mem_inst__abc_19396_new_n3915_));
OAI21X1 OAI21X1_1962 ( .A(w_mem_inst_w_mem_7__10_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf80), .C(w_mem_inst__abc_19396_new_n3915_), .Y(w_mem_inst__abc_19396_new_n3916_));
OAI21X1 OAI21X1_1963 ( .A(w_mem_inst__abc_19396_new_n3913_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf6), .C(w_mem_inst__abc_19396_new_n3916_), .Y(w_mem_inst__0w_mem_6__31_0__10_));
OAI21X1 OAI21X1_1964 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf4), .B(w_mem_inst__abc_19396_new_n3919_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf79), .Y(w_mem_inst__abc_19396_new_n3920_));
OAI21X1 OAI21X1_1965 ( .A(w_mem_inst_w_mem_7__11_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf78), .C(w_mem_inst__abc_19396_new_n3920_), .Y(w_mem_inst__abc_19396_new_n3921_));
OAI21X1 OAI21X1_1966 ( .A(w_mem_inst__abc_19396_new_n3918_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf5), .C(w_mem_inst__abc_19396_new_n3921_), .Y(w_mem_inst__0w_mem_6__31_0__11_));
OAI21X1 OAI21X1_1967 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf3), .B(w_mem_inst__abc_19396_new_n3924_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf77), .Y(w_mem_inst__abc_19396_new_n3925_));
OAI21X1 OAI21X1_1968 ( .A(w_mem_inst_w_mem_7__12_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf76), .C(w_mem_inst__abc_19396_new_n3925_), .Y(w_mem_inst__abc_19396_new_n3926_));
OAI21X1 OAI21X1_1969 ( .A(w_mem_inst__abc_19396_new_n3923_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf4), .C(w_mem_inst__abc_19396_new_n3926_), .Y(w_mem_inst__0w_mem_6__31_0__12_));
OAI21X1 OAI21X1_197 ( .A(_abc_15497_new_n1112_), .B(_abc_15497_new_n1648__bF_buf6), .C(_abc_15497_new_n1701_), .Y(_0e_reg_31_0__16_));
OAI21X1 OAI21X1_1970 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf2), .B(w_mem_inst__abc_19396_new_n3929_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf75), .Y(w_mem_inst__abc_19396_new_n3930_));
OAI21X1 OAI21X1_1971 ( .A(w_mem_inst_w_mem_7__13_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf74), .C(w_mem_inst__abc_19396_new_n3930_), .Y(w_mem_inst__abc_19396_new_n3931_));
OAI21X1 OAI21X1_1972 ( .A(w_mem_inst__abc_19396_new_n3928_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf3), .C(w_mem_inst__abc_19396_new_n3931_), .Y(w_mem_inst__0w_mem_6__31_0__13_));
OAI21X1 OAI21X1_1973 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf1), .B(w_mem_inst__abc_19396_new_n3934_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf73), .Y(w_mem_inst__abc_19396_new_n3935_));
OAI21X1 OAI21X1_1974 ( .A(w_mem_inst_w_mem_7__14_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf72), .C(w_mem_inst__abc_19396_new_n3935_), .Y(w_mem_inst__abc_19396_new_n3936_));
OAI21X1 OAI21X1_1975 ( .A(w_mem_inst__abc_19396_new_n3933_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf2), .C(w_mem_inst__abc_19396_new_n3936_), .Y(w_mem_inst__0w_mem_6__31_0__14_));
OAI21X1 OAI21X1_1976 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf0), .B(w_mem_inst__abc_19396_new_n3939_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf71), .Y(w_mem_inst__abc_19396_new_n3940_));
OAI21X1 OAI21X1_1977 ( .A(w_mem_inst_w_mem_7__15_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf70), .C(w_mem_inst__abc_19396_new_n3940_), .Y(w_mem_inst__abc_19396_new_n3941_));
OAI21X1 OAI21X1_1978 ( .A(w_mem_inst__abc_19396_new_n3938_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf1), .C(w_mem_inst__abc_19396_new_n3941_), .Y(w_mem_inst__0w_mem_6__31_0__15_));
OAI21X1 OAI21X1_1979 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf60), .B(w_mem_inst__abc_19396_new_n3944_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf69), .Y(w_mem_inst__abc_19396_new_n3945_));
OAI21X1 OAI21X1_198 ( .A(_abc_15497_new_n871__bF_buf2), .B(_abc_15497_new_n872__bF_buf3), .C(_abc_15497_new_n1122_), .Y(_abc_15497_new_n1703_));
OAI21X1 OAI21X1_1980 ( .A(w_mem_inst_w_mem_7__16_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf68), .C(w_mem_inst__abc_19396_new_n3945_), .Y(w_mem_inst__abc_19396_new_n3946_));
OAI21X1 OAI21X1_1981 ( .A(w_mem_inst__abc_19396_new_n3943_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf0), .C(w_mem_inst__abc_19396_new_n3946_), .Y(w_mem_inst__0w_mem_6__31_0__16_));
OAI21X1 OAI21X1_1982 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf59), .B(w_mem_inst__abc_19396_new_n3949_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf67), .Y(w_mem_inst__abc_19396_new_n3950_));
OAI21X1 OAI21X1_1983 ( .A(w_mem_inst_w_mem_7__17_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf66), .C(w_mem_inst__abc_19396_new_n3950_), .Y(w_mem_inst__abc_19396_new_n3951_));
OAI21X1 OAI21X1_1984 ( .A(w_mem_inst__abc_19396_new_n3948_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf60), .C(w_mem_inst__abc_19396_new_n3951_), .Y(w_mem_inst__0w_mem_6__31_0__17_));
OAI21X1 OAI21X1_1985 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf58), .B(w_mem_inst__abc_19396_new_n3954_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf65), .Y(w_mem_inst__abc_19396_new_n3955_));
OAI21X1 OAI21X1_1986 ( .A(w_mem_inst_w_mem_7__18_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf64), .C(w_mem_inst__abc_19396_new_n3955_), .Y(w_mem_inst__abc_19396_new_n3956_));
OAI21X1 OAI21X1_1987 ( .A(w_mem_inst__abc_19396_new_n3953_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf59), .C(w_mem_inst__abc_19396_new_n3956_), .Y(w_mem_inst__0w_mem_6__31_0__18_));
OAI21X1 OAI21X1_1988 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf57), .B(w_mem_inst__abc_19396_new_n3959_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf63), .Y(w_mem_inst__abc_19396_new_n3960_));
OAI21X1 OAI21X1_1989 ( .A(w_mem_inst_w_mem_7__19_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf62), .C(w_mem_inst__abc_19396_new_n3960_), .Y(w_mem_inst__abc_19396_new_n3961_));
OAI21X1 OAI21X1_199 ( .A(_abc_15497_new_n1121_), .B(_abc_15497_new_n1648__bF_buf5), .C(_abc_15497_new_n1704_), .Y(_0e_reg_31_0__17_));
OAI21X1 OAI21X1_1990 ( .A(w_mem_inst__abc_19396_new_n3958_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf58), .C(w_mem_inst__abc_19396_new_n3961_), .Y(w_mem_inst__0w_mem_6__31_0__19_));
OAI21X1 OAI21X1_1991 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf56), .B(w_mem_inst__abc_19396_new_n3964_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf61), .Y(w_mem_inst__abc_19396_new_n3965_));
OAI21X1 OAI21X1_1992 ( .A(w_mem_inst_w_mem_7__20_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf60), .C(w_mem_inst__abc_19396_new_n3965_), .Y(w_mem_inst__abc_19396_new_n3966_));
OAI21X1 OAI21X1_1993 ( .A(w_mem_inst__abc_19396_new_n3963_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf57), .C(w_mem_inst__abc_19396_new_n3966_), .Y(w_mem_inst__0w_mem_6__31_0__20_));
OAI21X1 OAI21X1_1994 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf55), .B(w_mem_inst__abc_19396_new_n3969_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf59), .Y(w_mem_inst__abc_19396_new_n3970_));
OAI21X1 OAI21X1_1995 ( .A(w_mem_inst_w_mem_7__21_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf58), .C(w_mem_inst__abc_19396_new_n3970_), .Y(w_mem_inst__abc_19396_new_n3971_));
OAI21X1 OAI21X1_1996 ( .A(w_mem_inst__abc_19396_new_n3968_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf56), .C(w_mem_inst__abc_19396_new_n3971_), .Y(w_mem_inst__0w_mem_6__31_0__21_));
OAI21X1 OAI21X1_1997 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf54), .B(w_mem_inst__abc_19396_new_n3974_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf57), .Y(w_mem_inst__abc_19396_new_n3975_));
OAI21X1 OAI21X1_1998 ( .A(w_mem_inst_w_mem_7__22_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf56), .C(w_mem_inst__abc_19396_new_n3975_), .Y(w_mem_inst__abc_19396_new_n3976_));
OAI21X1 OAI21X1_1999 ( .A(w_mem_inst__abc_19396_new_n3973_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf55), .C(w_mem_inst__abc_19396_new_n3976_), .Y(w_mem_inst__0w_mem_6__31_0__22_));
OAI21X1 OAI21X1_2 ( .A(_abc_15497_new_n766_), .B(_abc_15497_new_n777_), .C(_abc_15497_new_n765_), .Y(_abc_15497_new_n778_));
OAI21X1 OAI21X1_20 ( .A(_abc_15497_new_n921_), .B(_abc_15497_new_n922_), .C(digest_update_bF_buf5), .Y(_abc_15497_new_n923_));
OAI21X1 OAI21X1_200 ( .A(_abc_15497_new_n1130_), .B(_abc_15497_new_n1648__bF_buf4), .C(_abc_15497_new_n1707_), .Y(_0e_reg_31_0__18_));
OAI21X1 OAI21X1_2000 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf53), .B(w_mem_inst__abc_19396_new_n3979_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf55), .Y(w_mem_inst__abc_19396_new_n3980_));
OAI21X1 OAI21X1_2001 ( .A(w_mem_inst_w_mem_7__23_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf54), .C(w_mem_inst__abc_19396_new_n3980_), .Y(w_mem_inst__abc_19396_new_n3981_));
OAI21X1 OAI21X1_2002 ( .A(w_mem_inst__abc_19396_new_n3978_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf54), .C(w_mem_inst__abc_19396_new_n3981_), .Y(w_mem_inst__0w_mem_6__31_0__23_));
OAI21X1 OAI21X1_2003 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf52), .B(w_mem_inst__abc_19396_new_n3984_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf53), .Y(w_mem_inst__abc_19396_new_n3985_));
OAI21X1 OAI21X1_2004 ( .A(w_mem_inst_w_mem_7__24_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf52), .C(w_mem_inst__abc_19396_new_n3985_), .Y(w_mem_inst__abc_19396_new_n3986_));
OAI21X1 OAI21X1_2005 ( .A(w_mem_inst__abc_19396_new_n3983_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf53), .C(w_mem_inst__abc_19396_new_n3986_), .Y(w_mem_inst__0w_mem_6__31_0__24_));
OAI21X1 OAI21X1_2006 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf51), .B(w_mem_inst__abc_19396_new_n3989_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf51), .Y(w_mem_inst__abc_19396_new_n3990_));
OAI21X1 OAI21X1_2007 ( .A(w_mem_inst_w_mem_7__25_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf50), .C(w_mem_inst__abc_19396_new_n3990_), .Y(w_mem_inst__abc_19396_new_n3991_));
OAI21X1 OAI21X1_2008 ( .A(w_mem_inst__abc_19396_new_n3988_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf52), .C(w_mem_inst__abc_19396_new_n3991_), .Y(w_mem_inst__0w_mem_6__31_0__25_));
OAI21X1 OAI21X1_2009 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf50), .B(w_mem_inst__abc_19396_new_n3994_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf49), .Y(w_mem_inst__abc_19396_new_n3995_));
OAI21X1 OAI21X1_201 ( .A(_abc_15497_new_n1146_), .B(_abc_15497_new_n1648__bF_buf3), .C(_abc_15497_new_n1710_), .Y(_0e_reg_31_0__19_));
OAI21X1 OAI21X1_2010 ( .A(w_mem_inst_w_mem_7__26_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf48), .C(w_mem_inst__abc_19396_new_n3995_), .Y(w_mem_inst__abc_19396_new_n3996_));
OAI21X1 OAI21X1_2011 ( .A(w_mem_inst__abc_19396_new_n3993_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf51), .C(w_mem_inst__abc_19396_new_n3996_), .Y(w_mem_inst__0w_mem_6__31_0__26_));
OAI21X1 OAI21X1_2012 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf49), .B(w_mem_inst__abc_19396_new_n3999_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf47), .Y(w_mem_inst__abc_19396_new_n4000_));
OAI21X1 OAI21X1_2013 ( .A(w_mem_inst_w_mem_7__27_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf46), .C(w_mem_inst__abc_19396_new_n4000_), .Y(w_mem_inst__abc_19396_new_n4001_));
OAI21X1 OAI21X1_2014 ( .A(w_mem_inst__abc_19396_new_n3998_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf50), .C(w_mem_inst__abc_19396_new_n4001_), .Y(w_mem_inst__0w_mem_6__31_0__27_));
OAI21X1 OAI21X1_2015 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf48), .B(w_mem_inst__abc_19396_new_n4004_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf45), .Y(w_mem_inst__abc_19396_new_n4005_));
OAI21X1 OAI21X1_2016 ( .A(w_mem_inst_w_mem_7__28_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf44), .C(w_mem_inst__abc_19396_new_n4005_), .Y(w_mem_inst__abc_19396_new_n4006_));
OAI21X1 OAI21X1_2017 ( .A(w_mem_inst__abc_19396_new_n4003_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf49), .C(w_mem_inst__abc_19396_new_n4006_), .Y(w_mem_inst__0w_mem_6__31_0__28_));
OAI21X1 OAI21X1_2018 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf47), .B(w_mem_inst__abc_19396_new_n4009_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf43), .Y(w_mem_inst__abc_19396_new_n4010_));
OAI21X1 OAI21X1_2019 ( .A(w_mem_inst_w_mem_7__29_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf42), .C(w_mem_inst__abc_19396_new_n4010_), .Y(w_mem_inst__abc_19396_new_n4011_));
OAI21X1 OAI21X1_202 ( .A(_abc_15497_new_n871__bF_buf1), .B(_abc_15497_new_n872__bF_buf2), .C(_abc_15497_new_n1163_), .Y(_abc_15497_new_n1712_));
OAI21X1 OAI21X1_2020 ( .A(w_mem_inst__abc_19396_new_n4008_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf48), .C(w_mem_inst__abc_19396_new_n4011_), .Y(w_mem_inst__0w_mem_6__31_0__29_));
OAI21X1 OAI21X1_2021 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf46), .B(w_mem_inst__abc_19396_new_n4014_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf41), .Y(w_mem_inst__abc_19396_new_n4015_));
OAI21X1 OAI21X1_2022 ( .A(w_mem_inst_w_mem_7__30_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf40), .C(w_mem_inst__abc_19396_new_n4015_), .Y(w_mem_inst__abc_19396_new_n4016_));
OAI21X1 OAI21X1_2023 ( .A(w_mem_inst__abc_19396_new_n4013_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf47), .C(w_mem_inst__abc_19396_new_n4016_), .Y(w_mem_inst__0w_mem_6__31_0__30_));
OAI21X1 OAI21X1_2024 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf45), .B(w_mem_inst__abc_19396_new_n4019_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf39), .Y(w_mem_inst__abc_19396_new_n4020_));
OAI21X1 OAI21X1_2025 ( .A(w_mem_inst_w_mem_7__31_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf38), .C(w_mem_inst__abc_19396_new_n4020_), .Y(w_mem_inst__abc_19396_new_n4021_));
OAI21X1 OAI21X1_2026 ( .A(w_mem_inst__abc_19396_new_n4018_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf46), .C(w_mem_inst__abc_19396_new_n4021_), .Y(w_mem_inst__0w_mem_6__31_0__31_));
OAI21X1 OAI21X1_2027 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf44), .B(w_mem_inst__abc_19396_new_n4023_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf37), .Y(w_mem_inst__abc_19396_new_n4024_));
OAI21X1 OAI21X1_2028 ( .A(w_mem_inst_w_mem_6__0_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf36), .C(w_mem_inst__abc_19396_new_n4024_), .Y(w_mem_inst__abc_19396_new_n4025_));
OAI21X1 OAI21X1_2029 ( .A(w_mem_inst__abc_19396_new_n1591_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf45), .C(w_mem_inst__abc_19396_new_n4025_), .Y(w_mem_inst__0w_mem_5__31_0__0_));
OAI21X1 OAI21X1_203 ( .A(_abc_15497_new_n1162_), .B(_abc_15497_new_n1648__bF_buf2), .C(_abc_15497_new_n1713_), .Y(_0e_reg_31_0__20_));
OAI21X1 OAI21X1_2030 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf43), .B(w_mem_inst__abc_19396_new_n4027_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf35), .Y(w_mem_inst__abc_19396_new_n4028_));
OAI21X1 OAI21X1_2031 ( .A(w_mem_inst_w_mem_6__1_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf34), .C(w_mem_inst__abc_19396_new_n4028_), .Y(w_mem_inst__abc_19396_new_n4029_));
OAI21X1 OAI21X1_2032 ( .A(w_mem_inst__abc_19396_new_n1646_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf44), .C(w_mem_inst__abc_19396_new_n4029_), .Y(w_mem_inst__0w_mem_5__31_0__1_));
OAI21X1 OAI21X1_2033 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf42), .B(w_mem_inst__abc_19396_new_n4031_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf33), .Y(w_mem_inst__abc_19396_new_n4032_));
OAI21X1 OAI21X1_2034 ( .A(w_mem_inst_w_mem_6__2_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf32), .C(w_mem_inst__abc_19396_new_n4032_), .Y(w_mem_inst__abc_19396_new_n4033_));
OAI21X1 OAI21X1_2035 ( .A(w_mem_inst__abc_19396_new_n1671_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf43), .C(w_mem_inst__abc_19396_new_n4033_), .Y(w_mem_inst__0w_mem_5__31_0__2_));
OAI21X1 OAI21X1_2036 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf41), .B(w_mem_inst__abc_19396_new_n4035_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf31), .Y(w_mem_inst__abc_19396_new_n4036_));
OAI21X1 OAI21X1_2037 ( .A(w_mem_inst_w_mem_6__3_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf30), .C(w_mem_inst__abc_19396_new_n4036_), .Y(w_mem_inst__abc_19396_new_n4037_));
OAI21X1 OAI21X1_2038 ( .A(w_mem_inst__abc_19396_new_n1696_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf42), .C(w_mem_inst__abc_19396_new_n4037_), .Y(w_mem_inst__0w_mem_5__31_0__3_));
OAI21X1 OAI21X1_2039 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf40), .B(w_mem_inst__abc_19396_new_n4039_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf29), .Y(w_mem_inst__abc_19396_new_n4040_));
OAI21X1 OAI21X1_204 ( .A(_abc_15497_new_n1173_), .B(_abc_15497_new_n1648__bF_buf1), .C(_abc_15497_new_n1716_), .Y(_0e_reg_31_0__21_));
OAI21X1 OAI21X1_2040 ( .A(w_mem_inst_w_mem_6__4_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf28), .C(w_mem_inst__abc_19396_new_n4040_), .Y(w_mem_inst__abc_19396_new_n4041_));
OAI21X1 OAI21X1_2041 ( .A(w_mem_inst__abc_19396_new_n1721_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf41), .C(w_mem_inst__abc_19396_new_n4041_), .Y(w_mem_inst__0w_mem_5__31_0__4_));
OAI21X1 OAI21X1_2042 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf39), .B(w_mem_inst__abc_19396_new_n4043_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf27), .Y(w_mem_inst__abc_19396_new_n4044_));
OAI21X1 OAI21X1_2043 ( .A(w_mem_inst_w_mem_6__5_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf26), .C(w_mem_inst__abc_19396_new_n4044_), .Y(w_mem_inst__abc_19396_new_n4045_));
OAI21X1 OAI21X1_2044 ( .A(w_mem_inst__abc_19396_new_n1746_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf40), .C(w_mem_inst__abc_19396_new_n4045_), .Y(w_mem_inst__0w_mem_5__31_0__5_));
OAI21X1 OAI21X1_2045 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf38), .B(w_mem_inst__abc_19396_new_n4047_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf25), .Y(w_mem_inst__abc_19396_new_n4048_));
OAI21X1 OAI21X1_2046 ( .A(w_mem_inst_w_mem_6__6_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf24), .C(w_mem_inst__abc_19396_new_n4048_), .Y(w_mem_inst__abc_19396_new_n4049_));
OAI21X1 OAI21X1_2047 ( .A(w_mem_inst__abc_19396_new_n1771_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf39), .C(w_mem_inst__abc_19396_new_n4049_), .Y(w_mem_inst__0w_mem_5__31_0__6_));
OAI21X1 OAI21X1_2048 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf37), .B(w_mem_inst__abc_19396_new_n4051_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf23), .Y(w_mem_inst__abc_19396_new_n4052_));
OAI21X1 OAI21X1_2049 ( .A(w_mem_inst_w_mem_6__7_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf22), .C(w_mem_inst__abc_19396_new_n4052_), .Y(w_mem_inst__abc_19396_new_n4053_));
OAI21X1 OAI21X1_205 ( .A(_auto_iopadmap_cc_368_execute_22625_22_), .B(_abc_15497_new_n883__bF_buf6), .C(round_ctr_rst_bF_buf2), .Y(_abc_15497_new_n1718_));
OAI21X1 OAI21X1_2050 ( .A(w_mem_inst__abc_19396_new_n1796_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf38), .C(w_mem_inst__abc_19396_new_n4053_), .Y(w_mem_inst__0w_mem_5__31_0__7_));
OAI21X1 OAI21X1_2051 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf36), .B(w_mem_inst__abc_19396_new_n4055_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf21), .Y(w_mem_inst__abc_19396_new_n4056_));
OAI21X1 OAI21X1_2052 ( .A(w_mem_inst_w_mem_6__8_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf20), .C(w_mem_inst__abc_19396_new_n4056_), .Y(w_mem_inst__abc_19396_new_n4057_));
OAI21X1 OAI21X1_2053 ( .A(w_mem_inst__abc_19396_new_n1821_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf37), .C(w_mem_inst__abc_19396_new_n4057_), .Y(w_mem_inst__0w_mem_5__31_0__8_));
OAI21X1 OAI21X1_2054 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf35), .B(w_mem_inst__abc_19396_new_n4059_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf19), .Y(w_mem_inst__abc_19396_new_n4060_));
OAI21X1 OAI21X1_2055 ( .A(w_mem_inst_w_mem_6__9_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf18), .C(w_mem_inst__abc_19396_new_n4060_), .Y(w_mem_inst__abc_19396_new_n4061_));
OAI21X1 OAI21X1_2056 ( .A(w_mem_inst__abc_19396_new_n1846_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf36), .C(w_mem_inst__abc_19396_new_n4061_), .Y(w_mem_inst__0w_mem_5__31_0__9_));
OAI21X1 OAI21X1_2057 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf34), .B(w_mem_inst__abc_19396_new_n4063_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf17), .Y(w_mem_inst__abc_19396_new_n4064_));
OAI21X1 OAI21X1_2058 ( .A(w_mem_inst_w_mem_6__10_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf16), .C(w_mem_inst__abc_19396_new_n4064_), .Y(w_mem_inst__abc_19396_new_n4065_));
OAI21X1 OAI21X1_2059 ( .A(w_mem_inst__abc_19396_new_n1871_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf35), .C(w_mem_inst__abc_19396_new_n4065_), .Y(w_mem_inst__0w_mem_5__31_0__10_));
OAI21X1 OAI21X1_206 ( .A(round_ctr_inc_bF_buf10), .B(_abc_15497_new_n1718_), .C(_abc_15497_new_n1719_), .Y(_0e_reg_31_0__22_));
OAI21X1 OAI21X1_2060 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf33), .B(w_mem_inst__abc_19396_new_n4067_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf15), .Y(w_mem_inst__abc_19396_new_n4068_));
OAI21X1 OAI21X1_2061 ( .A(w_mem_inst_w_mem_6__11_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf14), .C(w_mem_inst__abc_19396_new_n4068_), .Y(w_mem_inst__abc_19396_new_n4069_));
OAI21X1 OAI21X1_2062 ( .A(w_mem_inst__abc_19396_new_n1896_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf34), .C(w_mem_inst__abc_19396_new_n4069_), .Y(w_mem_inst__0w_mem_5__31_0__11_));
OAI21X1 OAI21X1_2063 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf32), .B(w_mem_inst__abc_19396_new_n4071_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf13), .Y(w_mem_inst__abc_19396_new_n4072_));
OAI21X1 OAI21X1_2064 ( .A(w_mem_inst_w_mem_6__12_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf12), .C(w_mem_inst__abc_19396_new_n4072_), .Y(w_mem_inst__abc_19396_new_n4073_));
OAI21X1 OAI21X1_2065 ( .A(w_mem_inst__abc_19396_new_n1921_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf33), .C(w_mem_inst__abc_19396_new_n4073_), .Y(w_mem_inst__0w_mem_5__31_0__12_));
OAI21X1 OAI21X1_2066 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf31), .B(w_mem_inst__abc_19396_new_n4075_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf11), .Y(w_mem_inst__abc_19396_new_n4076_));
OAI21X1 OAI21X1_2067 ( .A(w_mem_inst_w_mem_6__13_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf10), .C(w_mem_inst__abc_19396_new_n4076_), .Y(w_mem_inst__abc_19396_new_n4077_));
OAI21X1 OAI21X1_2068 ( .A(w_mem_inst__abc_19396_new_n1946_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf32), .C(w_mem_inst__abc_19396_new_n4077_), .Y(w_mem_inst__0w_mem_5__31_0__13_));
OAI21X1 OAI21X1_2069 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf30), .B(w_mem_inst__abc_19396_new_n4079_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf9), .Y(w_mem_inst__abc_19396_new_n4080_));
OAI21X1 OAI21X1_207 ( .A(_auto_iopadmap_cc_368_execute_22625_23_), .B(_abc_15497_new_n883__bF_buf5), .C(round_ctr_rst_bF_buf1), .Y(_abc_15497_new_n1721_));
OAI21X1 OAI21X1_2070 ( .A(w_mem_inst_w_mem_6__14_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf8), .C(w_mem_inst__abc_19396_new_n4080_), .Y(w_mem_inst__abc_19396_new_n4081_));
OAI21X1 OAI21X1_2071 ( .A(w_mem_inst__abc_19396_new_n1971_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf31), .C(w_mem_inst__abc_19396_new_n4081_), .Y(w_mem_inst__0w_mem_5__31_0__14_));
OAI21X1 OAI21X1_2072 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf29), .B(w_mem_inst__abc_19396_new_n4083_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf7), .Y(w_mem_inst__abc_19396_new_n4084_));
OAI21X1 OAI21X1_2073 ( .A(w_mem_inst_w_mem_6__15_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf6), .C(w_mem_inst__abc_19396_new_n4084_), .Y(w_mem_inst__abc_19396_new_n4085_));
OAI21X1 OAI21X1_2074 ( .A(w_mem_inst__abc_19396_new_n1996_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf30), .C(w_mem_inst__abc_19396_new_n4085_), .Y(w_mem_inst__0w_mem_5__31_0__15_));
OAI21X1 OAI21X1_2075 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf28), .B(w_mem_inst__abc_19396_new_n4087_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf5), .Y(w_mem_inst__abc_19396_new_n4088_));
OAI21X1 OAI21X1_2076 ( .A(w_mem_inst_w_mem_6__16_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf4), .C(w_mem_inst__abc_19396_new_n4088_), .Y(w_mem_inst__abc_19396_new_n4089_));
OAI21X1 OAI21X1_2077 ( .A(w_mem_inst__abc_19396_new_n2021_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf29), .C(w_mem_inst__abc_19396_new_n4089_), .Y(w_mem_inst__0w_mem_5__31_0__16_));
OAI21X1 OAI21X1_2078 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf27), .B(w_mem_inst__abc_19396_new_n4091_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf3), .Y(w_mem_inst__abc_19396_new_n4092_));
OAI21X1 OAI21X1_2079 ( .A(w_mem_inst_w_mem_6__17_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf2), .C(w_mem_inst__abc_19396_new_n4092_), .Y(w_mem_inst__abc_19396_new_n4093_));
OAI21X1 OAI21X1_208 ( .A(round_ctr_inc_bF_buf8), .B(_abc_15497_new_n1721_), .C(_abc_15497_new_n1722_), .Y(_0e_reg_31_0__23_));
OAI21X1 OAI21X1_2080 ( .A(w_mem_inst__abc_19396_new_n2046_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf28), .C(w_mem_inst__abc_19396_new_n4093_), .Y(w_mem_inst__0w_mem_5__31_0__17_));
OAI21X1 OAI21X1_2081 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf26), .B(w_mem_inst__abc_19396_new_n4095_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf1), .Y(w_mem_inst__abc_19396_new_n4096_));
OAI21X1 OAI21X1_2082 ( .A(w_mem_inst_w_mem_6__18_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf0), .C(w_mem_inst__abc_19396_new_n4096_), .Y(w_mem_inst__abc_19396_new_n4097_));
OAI21X1 OAI21X1_2083 ( .A(w_mem_inst__abc_19396_new_n2071_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf27), .C(w_mem_inst__abc_19396_new_n4097_), .Y(w_mem_inst__0w_mem_5__31_0__18_));
OAI21X1 OAI21X1_2084 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf25), .B(w_mem_inst__abc_19396_new_n4099_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf96), .Y(w_mem_inst__abc_19396_new_n4100_));
OAI21X1 OAI21X1_2085 ( .A(w_mem_inst_w_mem_6__19_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf95), .C(w_mem_inst__abc_19396_new_n4100_), .Y(w_mem_inst__abc_19396_new_n4101_));
OAI21X1 OAI21X1_2086 ( .A(w_mem_inst__abc_19396_new_n2096_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf26), .C(w_mem_inst__abc_19396_new_n4101_), .Y(w_mem_inst__0w_mem_5__31_0__19_));
OAI21X1 OAI21X1_2087 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf24), .B(w_mem_inst__abc_19396_new_n4103_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf94), .Y(w_mem_inst__abc_19396_new_n4104_));
OAI21X1 OAI21X1_2088 ( .A(w_mem_inst_w_mem_6__20_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf93), .C(w_mem_inst__abc_19396_new_n4104_), .Y(w_mem_inst__abc_19396_new_n4105_));
OAI21X1 OAI21X1_2089 ( .A(w_mem_inst__abc_19396_new_n2121_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf25), .C(w_mem_inst__abc_19396_new_n4105_), .Y(w_mem_inst__0w_mem_5__31_0__20_));
OAI21X1 OAI21X1_209 ( .A(_abc_15497_new_n871__bF_buf0), .B(_abc_15497_new_n872__bF_buf1), .C(_abc_15497_new_n1214_), .Y(_abc_15497_new_n1724_));
OAI21X1 OAI21X1_2090 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf23), .B(w_mem_inst__abc_19396_new_n4107_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf92), .Y(w_mem_inst__abc_19396_new_n4108_));
OAI21X1 OAI21X1_2091 ( .A(w_mem_inst_w_mem_6__21_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf91), .C(w_mem_inst__abc_19396_new_n4108_), .Y(w_mem_inst__abc_19396_new_n4109_));
OAI21X1 OAI21X1_2092 ( .A(w_mem_inst__abc_19396_new_n2146_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf24), .C(w_mem_inst__abc_19396_new_n4109_), .Y(w_mem_inst__0w_mem_5__31_0__21_));
OAI21X1 OAI21X1_2093 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf22), .B(w_mem_inst__abc_19396_new_n4111_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf90), .Y(w_mem_inst__abc_19396_new_n4112_));
OAI21X1 OAI21X1_2094 ( .A(w_mem_inst_w_mem_6__22_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf89), .C(w_mem_inst__abc_19396_new_n4112_), .Y(w_mem_inst__abc_19396_new_n4113_));
OAI21X1 OAI21X1_2095 ( .A(w_mem_inst__abc_19396_new_n2171_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf23), .C(w_mem_inst__abc_19396_new_n4113_), .Y(w_mem_inst__0w_mem_5__31_0__22_));
OAI21X1 OAI21X1_2096 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf21), .B(w_mem_inst__abc_19396_new_n4115_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf88), .Y(w_mem_inst__abc_19396_new_n4116_));
OAI21X1 OAI21X1_2097 ( .A(w_mem_inst_w_mem_6__23_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf87), .C(w_mem_inst__abc_19396_new_n4116_), .Y(w_mem_inst__abc_19396_new_n4117_));
OAI21X1 OAI21X1_2098 ( .A(w_mem_inst__abc_19396_new_n2196_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf22), .C(w_mem_inst__abc_19396_new_n4117_), .Y(w_mem_inst__0w_mem_5__31_0__23_));
OAI21X1 OAI21X1_2099 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf20), .B(w_mem_inst__abc_19396_new_n4119_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf86), .Y(w_mem_inst__abc_19396_new_n4120_));
OAI21X1 OAI21X1_21 ( .A(_abc_15497_new_n916_), .B(_abc_15497_new_n927_), .C(_abc_15497_new_n921_), .Y(_abc_15497_new_n928_));
OAI21X1 OAI21X1_210 ( .A(_abc_15497_new_n1213_), .B(_abc_15497_new_n1648__bF_buf0), .C(_abc_15497_new_n1725_), .Y(_0e_reg_31_0__24_));
OAI21X1 OAI21X1_2100 ( .A(w_mem_inst_w_mem_6__24_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf85), .C(w_mem_inst__abc_19396_new_n4120_), .Y(w_mem_inst__abc_19396_new_n4121_));
OAI21X1 OAI21X1_2101 ( .A(w_mem_inst__abc_19396_new_n2221_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf21), .C(w_mem_inst__abc_19396_new_n4121_), .Y(w_mem_inst__0w_mem_5__31_0__24_));
OAI21X1 OAI21X1_2102 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf19), .B(w_mem_inst__abc_19396_new_n4123_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf84), .Y(w_mem_inst__abc_19396_new_n4124_));
OAI21X1 OAI21X1_2103 ( .A(w_mem_inst_w_mem_6__25_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf83), .C(w_mem_inst__abc_19396_new_n4124_), .Y(w_mem_inst__abc_19396_new_n4125_));
OAI21X1 OAI21X1_2104 ( .A(w_mem_inst__abc_19396_new_n2246_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf20), .C(w_mem_inst__abc_19396_new_n4125_), .Y(w_mem_inst__0w_mem_5__31_0__25_));
OAI21X1 OAI21X1_2105 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf18), .B(w_mem_inst__abc_19396_new_n4127_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf82), .Y(w_mem_inst__abc_19396_new_n4128_));
OAI21X1 OAI21X1_2106 ( .A(w_mem_inst_w_mem_6__26_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf81), .C(w_mem_inst__abc_19396_new_n4128_), .Y(w_mem_inst__abc_19396_new_n4129_));
OAI21X1 OAI21X1_2107 ( .A(w_mem_inst__abc_19396_new_n2271_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf19), .C(w_mem_inst__abc_19396_new_n4129_), .Y(w_mem_inst__0w_mem_5__31_0__26_));
OAI21X1 OAI21X1_2108 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf17), .B(w_mem_inst__abc_19396_new_n4131_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf80), .Y(w_mem_inst__abc_19396_new_n4132_));
OAI21X1 OAI21X1_2109 ( .A(w_mem_inst_w_mem_6__27_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf79), .C(w_mem_inst__abc_19396_new_n4132_), .Y(w_mem_inst__abc_19396_new_n4133_));
OAI21X1 OAI21X1_211 ( .A(_auto_iopadmap_cc_368_execute_22625_25_), .B(_abc_15497_new_n883__bF_buf4), .C(round_ctr_rst_bF_buf0), .Y(_abc_15497_new_n1727_));
OAI21X1 OAI21X1_2110 ( .A(w_mem_inst__abc_19396_new_n2296_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf18), .C(w_mem_inst__abc_19396_new_n4133_), .Y(w_mem_inst__0w_mem_5__31_0__27_));
OAI21X1 OAI21X1_2111 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf16), .B(w_mem_inst__abc_19396_new_n4135_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf78), .Y(w_mem_inst__abc_19396_new_n4136_));
OAI21X1 OAI21X1_2112 ( .A(w_mem_inst_w_mem_6__28_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf77), .C(w_mem_inst__abc_19396_new_n4136_), .Y(w_mem_inst__abc_19396_new_n4137_));
OAI21X1 OAI21X1_2113 ( .A(w_mem_inst__abc_19396_new_n2321_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf17), .C(w_mem_inst__abc_19396_new_n4137_), .Y(w_mem_inst__0w_mem_5__31_0__28_));
OAI21X1 OAI21X1_2114 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf15), .B(w_mem_inst__abc_19396_new_n4139_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf76), .Y(w_mem_inst__abc_19396_new_n4140_));
OAI21X1 OAI21X1_2115 ( .A(w_mem_inst_w_mem_6__29_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf75), .C(w_mem_inst__abc_19396_new_n4140_), .Y(w_mem_inst__abc_19396_new_n4141_));
OAI21X1 OAI21X1_2116 ( .A(w_mem_inst__abc_19396_new_n2346_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf16), .C(w_mem_inst__abc_19396_new_n4141_), .Y(w_mem_inst__0w_mem_5__31_0__29_));
OAI21X1 OAI21X1_2117 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf14), .B(w_mem_inst__abc_19396_new_n4143_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf74), .Y(w_mem_inst__abc_19396_new_n4144_));
OAI21X1 OAI21X1_2118 ( .A(w_mem_inst_w_mem_6__30_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf73), .C(w_mem_inst__abc_19396_new_n4144_), .Y(w_mem_inst__abc_19396_new_n4145_));
OAI21X1 OAI21X1_2119 ( .A(w_mem_inst__abc_19396_new_n2371_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf15), .C(w_mem_inst__abc_19396_new_n4145_), .Y(w_mem_inst__0w_mem_5__31_0__30_));
OAI21X1 OAI21X1_212 ( .A(round_ctr_inc_bF_buf5), .B(_abc_15497_new_n1727_), .C(_abc_15497_new_n1728_), .Y(_0e_reg_31_0__25_));
OAI21X1 OAI21X1_2120 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf13), .B(w_mem_inst__abc_19396_new_n4147_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf72), .Y(w_mem_inst__abc_19396_new_n4148_));
OAI21X1 OAI21X1_2121 ( .A(w_mem_inst_w_mem_6__31_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf71), .C(w_mem_inst__abc_19396_new_n4148_), .Y(w_mem_inst__abc_19396_new_n4149_));
OAI21X1 OAI21X1_2122 ( .A(w_mem_inst__abc_19396_new_n2396_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf14), .C(w_mem_inst__abc_19396_new_n4149_), .Y(w_mem_inst__0w_mem_5__31_0__31_));
OAI21X1 OAI21X1_2123 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf12), .B(w_mem_inst__abc_19396_new_n4152_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf70), .Y(w_mem_inst__abc_19396_new_n4153_));
OAI21X1 OAI21X1_2124 ( .A(w_mem_inst_w_mem_2__0_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf69), .C(w_mem_inst__abc_19396_new_n4153_), .Y(w_mem_inst__abc_19396_new_n4154_));
OAI21X1 OAI21X1_2125 ( .A(w_mem_inst__abc_19396_new_n4151_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf13), .C(w_mem_inst__abc_19396_new_n4154_), .Y(w_mem_inst__0w_mem_1__31_0__0_));
OAI21X1 OAI21X1_2126 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf11), .B(w_mem_inst__abc_19396_new_n4157_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf68), .Y(w_mem_inst__abc_19396_new_n4158_));
OAI21X1 OAI21X1_2127 ( .A(w_mem_inst_w_mem_2__1_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf67), .C(w_mem_inst__abc_19396_new_n4158_), .Y(w_mem_inst__abc_19396_new_n4159_));
OAI21X1 OAI21X1_2128 ( .A(w_mem_inst__abc_19396_new_n4156_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf12), .C(w_mem_inst__abc_19396_new_n4159_), .Y(w_mem_inst__0w_mem_1__31_0__1_));
OAI21X1 OAI21X1_2129 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf10), .B(w_mem_inst__abc_19396_new_n4162_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf66), .Y(w_mem_inst__abc_19396_new_n4163_));
OAI21X1 OAI21X1_213 ( .A(_abc_15497_new_n1239_), .B(_abc_15497_new_n1648__bF_buf8), .C(_abc_15497_new_n1731_), .Y(_0e_reg_31_0__26_));
OAI21X1 OAI21X1_2130 ( .A(w_mem_inst_w_mem_2__2_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf65), .C(w_mem_inst__abc_19396_new_n4163_), .Y(w_mem_inst__abc_19396_new_n4164_));
OAI21X1 OAI21X1_2131 ( .A(w_mem_inst__abc_19396_new_n4161_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf11), .C(w_mem_inst__abc_19396_new_n4164_), .Y(w_mem_inst__0w_mem_1__31_0__2_));
OAI21X1 OAI21X1_2132 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf9), .B(w_mem_inst__abc_19396_new_n4167_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf64), .Y(w_mem_inst__abc_19396_new_n4168_));
OAI21X1 OAI21X1_2133 ( .A(w_mem_inst_w_mem_2__3_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf63), .C(w_mem_inst__abc_19396_new_n4168_), .Y(w_mem_inst__abc_19396_new_n4169_));
OAI21X1 OAI21X1_2134 ( .A(w_mem_inst__abc_19396_new_n4166_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf10), .C(w_mem_inst__abc_19396_new_n4169_), .Y(w_mem_inst__0w_mem_1__31_0__3_));
OAI21X1 OAI21X1_2135 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf8), .B(w_mem_inst__abc_19396_new_n4172_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf62), .Y(w_mem_inst__abc_19396_new_n4173_));
OAI21X1 OAI21X1_2136 ( .A(w_mem_inst_w_mem_2__4_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf61), .C(w_mem_inst__abc_19396_new_n4173_), .Y(w_mem_inst__abc_19396_new_n4174_));
OAI21X1 OAI21X1_2137 ( .A(w_mem_inst__abc_19396_new_n4171_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf9), .C(w_mem_inst__abc_19396_new_n4174_), .Y(w_mem_inst__0w_mem_1__31_0__4_));
OAI21X1 OAI21X1_2138 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf7), .B(w_mem_inst__abc_19396_new_n4177_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf60), .Y(w_mem_inst__abc_19396_new_n4178_));
OAI21X1 OAI21X1_2139 ( .A(w_mem_inst_w_mem_2__5_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf59), .C(w_mem_inst__abc_19396_new_n4178_), .Y(w_mem_inst__abc_19396_new_n4179_));
OAI21X1 OAI21X1_214 ( .A(_abc_15497_new_n1250_), .B(_abc_15497_new_n1648__bF_buf7), .C(_abc_15497_new_n1734_), .Y(_0e_reg_31_0__27_));
OAI21X1 OAI21X1_2140 ( .A(w_mem_inst__abc_19396_new_n4176_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf8), .C(w_mem_inst__abc_19396_new_n4179_), .Y(w_mem_inst__0w_mem_1__31_0__5_));
OAI21X1 OAI21X1_2141 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf6), .B(w_mem_inst__abc_19396_new_n4182_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf58), .Y(w_mem_inst__abc_19396_new_n4183_));
OAI21X1 OAI21X1_2142 ( .A(w_mem_inst_w_mem_2__6_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf57), .C(w_mem_inst__abc_19396_new_n4183_), .Y(w_mem_inst__abc_19396_new_n4184_));
OAI21X1 OAI21X1_2143 ( .A(w_mem_inst__abc_19396_new_n4181_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf7), .C(w_mem_inst__abc_19396_new_n4184_), .Y(w_mem_inst__0w_mem_1__31_0__6_));
OAI21X1 OAI21X1_2144 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf5), .B(w_mem_inst__abc_19396_new_n4187_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf56), .Y(w_mem_inst__abc_19396_new_n4188_));
OAI21X1 OAI21X1_2145 ( .A(w_mem_inst_w_mem_2__7_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf55), .C(w_mem_inst__abc_19396_new_n4188_), .Y(w_mem_inst__abc_19396_new_n4189_));
OAI21X1 OAI21X1_2146 ( .A(w_mem_inst__abc_19396_new_n4186_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf6), .C(w_mem_inst__abc_19396_new_n4189_), .Y(w_mem_inst__0w_mem_1__31_0__7_));
OAI21X1 OAI21X1_2147 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf4), .B(w_mem_inst__abc_19396_new_n4192_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf54), .Y(w_mem_inst__abc_19396_new_n4193_));
OAI21X1 OAI21X1_2148 ( .A(w_mem_inst_w_mem_2__8_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf53), .C(w_mem_inst__abc_19396_new_n4193_), .Y(w_mem_inst__abc_19396_new_n4194_));
OAI21X1 OAI21X1_2149 ( .A(w_mem_inst__abc_19396_new_n4191_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf5), .C(w_mem_inst__abc_19396_new_n4194_), .Y(w_mem_inst__0w_mem_1__31_0__8_));
OAI21X1 OAI21X1_215 ( .A(_abc_15497_new_n1736_), .B(_abc_15497_new_n1648__bF_buf6), .C(_abc_15497_new_n1738_), .Y(_0e_reg_31_0__28_));
OAI21X1 OAI21X1_2150 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf3), .B(w_mem_inst__abc_19396_new_n4197_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf52), .Y(w_mem_inst__abc_19396_new_n4198_));
OAI21X1 OAI21X1_2151 ( .A(w_mem_inst_w_mem_2__9_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf51), .C(w_mem_inst__abc_19396_new_n4198_), .Y(w_mem_inst__abc_19396_new_n4199_));
OAI21X1 OAI21X1_2152 ( .A(w_mem_inst__abc_19396_new_n4196_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf4), .C(w_mem_inst__abc_19396_new_n4199_), .Y(w_mem_inst__0w_mem_1__31_0__9_));
OAI21X1 OAI21X1_2153 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf2), .B(w_mem_inst__abc_19396_new_n4202_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf50), .Y(w_mem_inst__abc_19396_new_n4203_));
OAI21X1 OAI21X1_2154 ( .A(w_mem_inst_w_mem_2__10_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf49), .C(w_mem_inst__abc_19396_new_n4203_), .Y(w_mem_inst__abc_19396_new_n4204_));
OAI21X1 OAI21X1_2155 ( .A(w_mem_inst__abc_19396_new_n4201_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf3), .C(w_mem_inst__abc_19396_new_n4204_), .Y(w_mem_inst__0w_mem_1__31_0__10_));
OAI21X1 OAI21X1_2156 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf1), .B(w_mem_inst__abc_19396_new_n4207_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf48), .Y(w_mem_inst__abc_19396_new_n4208_));
OAI21X1 OAI21X1_2157 ( .A(w_mem_inst_w_mem_2__11_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf47), .C(w_mem_inst__abc_19396_new_n4208_), .Y(w_mem_inst__abc_19396_new_n4209_));
OAI21X1 OAI21X1_2158 ( .A(w_mem_inst__abc_19396_new_n4206_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf2), .C(w_mem_inst__abc_19396_new_n4209_), .Y(w_mem_inst__0w_mem_1__31_0__11_));
OAI21X1 OAI21X1_2159 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf0), .B(w_mem_inst__abc_19396_new_n4212_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf46), .Y(w_mem_inst__abc_19396_new_n4213_));
OAI21X1 OAI21X1_216 ( .A(_abc_15497_new_n1273_), .B(_abc_15497_new_n1648__bF_buf5), .C(_abc_15497_new_n1741_), .Y(_0e_reg_31_0__29_));
OAI21X1 OAI21X1_2160 ( .A(w_mem_inst_w_mem_2__12_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf45), .C(w_mem_inst__abc_19396_new_n4213_), .Y(w_mem_inst__abc_19396_new_n4214_));
OAI21X1 OAI21X1_2161 ( .A(w_mem_inst__abc_19396_new_n4211_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf1), .C(w_mem_inst__abc_19396_new_n4214_), .Y(w_mem_inst__0w_mem_1__31_0__12_));
OAI21X1 OAI21X1_2162 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf60), .B(w_mem_inst__abc_19396_new_n4217_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf44), .Y(w_mem_inst__abc_19396_new_n4218_));
OAI21X1 OAI21X1_2163 ( .A(w_mem_inst_w_mem_2__13_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf43), .C(w_mem_inst__abc_19396_new_n4218_), .Y(w_mem_inst__abc_19396_new_n4219_));
OAI21X1 OAI21X1_2164 ( .A(w_mem_inst__abc_19396_new_n4216_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf0), .C(w_mem_inst__abc_19396_new_n4219_), .Y(w_mem_inst__0w_mem_1__31_0__13_));
OAI21X1 OAI21X1_2165 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf59), .B(w_mem_inst__abc_19396_new_n4222_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf42), .Y(w_mem_inst__abc_19396_new_n4223_));
OAI21X1 OAI21X1_2166 ( .A(w_mem_inst_w_mem_2__14_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf41), .C(w_mem_inst__abc_19396_new_n4223_), .Y(w_mem_inst__abc_19396_new_n4224_));
OAI21X1 OAI21X1_2167 ( .A(w_mem_inst__abc_19396_new_n4221_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf60), .C(w_mem_inst__abc_19396_new_n4224_), .Y(w_mem_inst__0w_mem_1__31_0__14_));
OAI21X1 OAI21X1_2168 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf58), .B(w_mem_inst__abc_19396_new_n4227_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf40), .Y(w_mem_inst__abc_19396_new_n4228_));
OAI21X1 OAI21X1_2169 ( .A(w_mem_inst_w_mem_2__15_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf39), .C(w_mem_inst__abc_19396_new_n4228_), .Y(w_mem_inst__abc_19396_new_n4229_));
OAI21X1 OAI21X1_217 ( .A(_auto_iopadmap_cc_368_execute_22625_30_), .B(_abc_15497_new_n883__bF_buf13), .C(round_ctr_rst_bF_buf8), .Y(_abc_15497_new_n1743_));
OAI21X1 OAI21X1_2170 ( .A(w_mem_inst__abc_19396_new_n4226_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf59), .C(w_mem_inst__abc_19396_new_n4229_), .Y(w_mem_inst__0w_mem_1__31_0__15_));
OAI21X1 OAI21X1_2171 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf57), .B(w_mem_inst__abc_19396_new_n4232_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf38), .Y(w_mem_inst__abc_19396_new_n4233_));
OAI21X1 OAI21X1_2172 ( .A(w_mem_inst_w_mem_2__16_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf37), .C(w_mem_inst__abc_19396_new_n4233_), .Y(w_mem_inst__abc_19396_new_n4234_));
OAI21X1 OAI21X1_2173 ( .A(w_mem_inst__abc_19396_new_n4231_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf58), .C(w_mem_inst__abc_19396_new_n4234_), .Y(w_mem_inst__0w_mem_1__31_0__16_));
OAI21X1 OAI21X1_2174 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf56), .B(w_mem_inst__abc_19396_new_n4237_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf36), .Y(w_mem_inst__abc_19396_new_n4238_));
OAI21X1 OAI21X1_2175 ( .A(w_mem_inst_w_mem_2__17_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf35), .C(w_mem_inst__abc_19396_new_n4238_), .Y(w_mem_inst__abc_19396_new_n4239_));
OAI21X1 OAI21X1_2176 ( .A(w_mem_inst__abc_19396_new_n4236_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf57), .C(w_mem_inst__abc_19396_new_n4239_), .Y(w_mem_inst__0w_mem_1__31_0__17_));
OAI21X1 OAI21X1_2177 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf55), .B(w_mem_inst__abc_19396_new_n4242_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf34), .Y(w_mem_inst__abc_19396_new_n4243_));
OAI21X1 OAI21X1_2178 ( .A(w_mem_inst_w_mem_2__18_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf33), .C(w_mem_inst__abc_19396_new_n4243_), .Y(w_mem_inst__abc_19396_new_n4244_));
OAI21X1 OAI21X1_2179 ( .A(w_mem_inst__abc_19396_new_n4241_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf56), .C(w_mem_inst__abc_19396_new_n4244_), .Y(w_mem_inst__0w_mem_1__31_0__18_));
OAI21X1 OAI21X1_218 ( .A(round_ctr_inc_bF_buf13), .B(_abc_15497_new_n1743_), .C(_abc_15497_new_n1744_), .Y(_0e_reg_31_0__30_));
OAI21X1 OAI21X1_2180 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf54), .B(w_mem_inst__abc_19396_new_n4247_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf32), .Y(w_mem_inst__abc_19396_new_n4248_));
OAI21X1 OAI21X1_2181 ( .A(w_mem_inst_w_mem_2__19_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf31), .C(w_mem_inst__abc_19396_new_n4248_), .Y(w_mem_inst__abc_19396_new_n4249_));
OAI21X1 OAI21X1_2182 ( .A(w_mem_inst__abc_19396_new_n4246_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf55), .C(w_mem_inst__abc_19396_new_n4249_), .Y(w_mem_inst__0w_mem_1__31_0__19_));
OAI21X1 OAI21X1_2183 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf53), .B(w_mem_inst__abc_19396_new_n4252_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf30), .Y(w_mem_inst__abc_19396_new_n4253_));
OAI21X1 OAI21X1_2184 ( .A(w_mem_inst_w_mem_2__20_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf29), .C(w_mem_inst__abc_19396_new_n4253_), .Y(w_mem_inst__abc_19396_new_n4254_));
OAI21X1 OAI21X1_2185 ( .A(w_mem_inst__abc_19396_new_n4251_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf54), .C(w_mem_inst__abc_19396_new_n4254_), .Y(w_mem_inst__0w_mem_1__31_0__20_));
OAI21X1 OAI21X1_2186 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf52), .B(w_mem_inst__abc_19396_new_n4257_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf28), .Y(w_mem_inst__abc_19396_new_n4258_));
OAI21X1 OAI21X1_2187 ( .A(w_mem_inst_w_mem_2__21_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf27), .C(w_mem_inst__abc_19396_new_n4258_), .Y(w_mem_inst__abc_19396_new_n4259_));
OAI21X1 OAI21X1_2188 ( .A(w_mem_inst__abc_19396_new_n4256_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf53), .C(w_mem_inst__abc_19396_new_n4259_), .Y(w_mem_inst__0w_mem_1__31_0__21_));
OAI21X1 OAI21X1_2189 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf51), .B(w_mem_inst__abc_19396_new_n4262_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf26), .Y(w_mem_inst__abc_19396_new_n4263_));
OAI21X1 OAI21X1_219 ( .A(_auto_iopadmap_cc_368_execute_22625_31_), .B(_abc_15497_new_n883__bF_buf12), .C(_abc_15497_new_n1650__bF_buf8), .Y(_abc_15497_new_n1746_));
OAI21X1 OAI21X1_2190 ( .A(w_mem_inst_w_mem_2__22_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf25), .C(w_mem_inst__abc_19396_new_n4263_), .Y(w_mem_inst__abc_19396_new_n4264_));
OAI21X1 OAI21X1_2191 ( .A(w_mem_inst__abc_19396_new_n4261_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf52), .C(w_mem_inst__abc_19396_new_n4264_), .Y(w_mem_inst__0w_mem_1__31_0__22_));
OAI21X1 OAI21X1_2192 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf50), .B(w_mem_inst__abc_19396_new_n4267_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf24), .Y(w_mem_inst__abc_19396_new_n4268_));
OAI21X1 OAI21X1_2193 ( .A(w_mem_inst_w_mem_2__23_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf23), .C(w_mem_inst__abc_19396_new_n4268_), .Y(w_mem_inst__abc_19396_new_n4269_));
OAI21X1 OAI21X1_2194 ( .A(w_mem_inst__abc_19396_new_n4266_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf51), .C(w_mem_inst__abc_19396_new_n4269_), .Y(w_mem_inst__0w_mem_1__31_0__23_));
OAI21X1 OAI21X1_2195 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf49), .B(w_mem_inst__abc_19396_new_n4272_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf22), .Y(w_mem_inst__abc_19396_new_n4273_));
OAI21X1 OAI21X1_2196 ( .A(w_mem_inst_w_mem_2__24_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf21), .C(w_mem_inst__abc_19396_new_n4273_), .Y(w_mem_inst__abc_19396_new_n4274_));
OAI21X1 OAI21X1_2197 ( .A(w_mem_inst__abc_19396_new_n4271_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf50), .C(w_mem_inst__abc_19396_new_n4274_), .Y(w_mem_inst__0w_mem_1__31_0__24_));
OAI21X1 OAI21X1_2198 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf48), .B(w_mem_inst__abc_19396_new_n4277_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf20), .Y(w_mem_inst__abc_19396_new_n4278_));
OAI21X1 OAI21X1_2199 ( .A(w_mem_inst_w_mem_2__25_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf19), .C(w_mem_inst__abc_19396_new_n4278_), .Y(w_mem_inst__abc_19396_new_n4279_));
OAI21X1 OAI21X1_22 ( .A(_abc_15497_new_n925_), .B(_abc_15497_new_n920_), .C(_abc_15497_new_n931_), .Y(_abc_15497_new_n932_));
OAI21X1 OAI21X1_220 ( .A(_abc_15497_new_n1751_), .B(_abc_15497_new_n1752_), .C(digest_update_bF_buf0), .Y(_abc_15497_new_n1753_));
OAI21X1 OAI21X1_2200 ( .A(w_mem_inst__abc_19396_new_n4276_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf49), .C(w_mem_inst__abc_19396_new_n4279_), .Y(w_mem_inst__0w_mem_1__31_0__25_));
OAI21X1 OAI21X1_2201 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf47), .B(w_mem_inst__abc_19396_new_n4282_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf18), .Y(w_mem_inst__abc_19396_new_n4283_));
OAI21X1 OAI21X1_2202 ( .A(w_mem_inst_w_mem_2__26_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf17), .C(w_mem_inst__abc_19396_new_n4283_), .Y(w_mem_inst__abc_19396_new_n4284_));
OAI21X1 OAI21X1_2203 ( .A(w_mem_inst__abc_19396_new_n4281_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf48), .C(w_mem_inst__abc_19396_new_n4284_), .Y(w_mem_inst__0w_mem_1__31_0__26_));
OAI21X1 OAI21X1_2204 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf46), .B(w_mem_inst__abc_19396_new_n4287_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf16), .Y(w_mem_inst__abc_19396_new_n4288_));
OAI21X1 OAI21X1_2205 ( .A(w_mem_inst_w_mem_2__27_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf15), .C(w_mem_inst__abc_19396_new_n4288_), .Y(w_mem_inst__abc_19396_new_n4289_));
OAI21X1 OAI21X1_2206 ( .A(w_mem_inst__abc_19396_new_n4286_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf47), .C(w_mem_inst__abc_19396_new_n4289_), .Y(w_mem_inst__0w_mem_1__31_0__27_));
OAI21X1 OAI21X1_2207 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf45), .B(w_mem_inst__abc_19396_new_n4292_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf14), .Y(w_mem_inst__abc_19396_new_n4293_));
OAI21X1 OAI21X1_2208 ( .A(w_mem_inst_w_mem_2__28_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf13), .C(w_mem_inst__abc_19396_new_n4293_), .Y(w_mem_inst__abc_19396_new_n4294_));
OAI21X1 OAI21X1_2209 ( .A(w_mem_inst__abc_19396_new_n4291_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf46), .C(w_mem_inst__abc_19396_new_n4294_), .Y(w_mem_inst__0w_mem_1__31_0__28_));
OAI21X1 OAI21X1_221 ( .A(_auto_iopadmap_cc_368_execute_22625_96_), .B(_abc_15497_new_n883__bF_buf11), .C(_abc_15497_new_n870__bF_buf1), .Y(_abc_15497_new_n1754_));
OAI21X1 OAI21X1_2210 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf44), .B(w_mem_inst__abc_19396_new_n4297_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf12), .Y(w_mem_inst__abc_19396_new_n4298_));
OAI21X1 OAI21X1_2211 ( .A(w_mem_inst_w_mem_2__29_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf11), .C(w_mem_inst__abc_19396_new_n4298_), .Y(w_mem_inst__abc_19396_new_n4299_));
OAI21X1 OAI21X1_2212 ( .A(w_mem_inst__abc_19396_new_n4296_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf45), .C(w_mem_inst__abc_19396_new_n4299_), .Y(w_mem_inst__0w_mem_1__31_0__29_));
OAI21X1 OAI21X1_2213 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf43), .B(w_mem_inst__abc_19396_new_n4302_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf10), .Y(w_mem_inst__abc_19396_new_n4303_));
OAI21X1 OAI21X1_2214 ( .A(w_mem_inst_w_mem_2__30_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf9), .C(w_mem_inst__abc_19396_new_n4303_), .Y(w_mem_inst__abc_19396_new_n4304_));
OAI21X1 OAI21X1_2215 ( .A(w_mem_inst__abc_19396_new_n4301_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf44), .C(w_mem_inst__abc_19396_new_n4304_), .Y(w_mem_inst__0w_mem_1__31_0__30_));
OAI21X1 OAI21X1_2216 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf42), .B(w_mem_inst__abc_19396_new_n4307_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf8), .Y(w_mem_inst__abc_19396_new_n4308_));
OAI21X1 OAI21X1_2217 ( .A(w_mem_inst_w_mem_2__31_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf7), .C(w_mem_inst__abc_19396_new_n4308_), .Y(w_mem_inst__abc_19396_new_n4309_));
OAI21X1 OAI21X1_2218 ( .A(w_mem_inst__abc_19396_new_n4306_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf43), .C(w_mem_inst__abc_19396_new_n4309_), .Y(w_mem_inst__0w_mem_1__31_0__31_));
OAI21X1 OAI21X1_2219 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf41), .B(w_mem_inst__abc_19396_new_n4312_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf6), .Y(w_mem_inst__abc_19396_new_n4313_));
OAI21X1 OAI21X1_222 ( .A(_abc_15497_new_n1750_), .B(_abc_15497_new_n1753_), .C(_abc_15497_new_n1754_), .Y(_0H1_reg_31_0__0_));
OAI21X1 OAI21X1_2220 ( .A(w_mem_inst_w_mem_4__0_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf5), .C(w_mem_inst__abc_19396_new_n4313_), .Y(w_mem_inst__abc_19396_new_n4314_));
OAI21X1 OAI21X1_2221 ( .A(w_mem_inst__abc_19396_new_n4311_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf42), .C(w_mem_inst__abc_19396_new_n4314_), .Y(w_mem_inst__0w_mem_3__31_0__0_));
OAI21X1 OAI21X1_2222 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf40), .B(w_mem_inst__abc_19396_new_n4317_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf4), .Y(w_mem_inst__abc_19396_new_n4318_));
OAI21X1 OAI21X1_2223 ( .A(w_mem_inst_w_mem_4__1_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf3), .C(w_mem_inst__abc_19396_new_n4318_), .Y(w_mem_inst__abc_19396_new_n4319_));
OAI21X1 OAI21X1_2224 ( .A(w_mem_inst__abc_19396_new_n4316_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf41), .C(w_mem_inst__abc_19396_new_n4319_), .Y(w_mem_inst__0w_mem_3__31_0__1_));
OAI21X1 OAI21X1_2225 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf39), .B(w_mem_inst__abc_19396_new_n4322_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf2), .Y(w_mem_inst__abc_19396_new_n4323_));
OAI21X1 OAI21X1_2226 ( .A(w_mem_inst_w_mem_4__2_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf1), .C(w_mem_inst__abc_19396_new_n4323_), .Y(w_mem_inst__abc_19396_new_n4324_));
OAI21X1 OAI21X1_2227 ( .A(w_mem_inst__abc_19396_new_n4321_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf40), .C(w_mem_inst__abc_19396_new_n4324_), .Y(w_mem_inst__0w_mem_3__31_0__2_));
OAI21X1 OAI21X1_2228 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf38), .B(w_mem_inst__abc_19396_new_n4327_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf0), .Y(w_mem_inst__abc_19396_new_n4328_));
OAI21X1 OAI21X1_2229 ( .A(w_mem_inst_w_mem_4__3_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf96), .C(w_mem_inst__abc_19396_new_n4328_), .Y(w_mem_inst__abc_19396_new_n4329_));
OAI21X1 OAI21X1_223 ( .A(_abc_15497_new_n1757_), .B(_abc_15497_new_n1758_), .C(_abc_15497_new_n1759_), .Y(_abc_15497_new_n1760_));
OAI21X1 OAI21X1_2230 ( .A(w_mem_inst__abc_19396_new_n4326_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf39), .C(w_mem_inst__abc_19396_new_n4329_), .Y(w_mem_inst__0w_mem_3__31_0__3_));
OAI21X1 OAI21X1_2231 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf37), .B(w_mem_inst__abc_19396_new_n4332_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf95), .Y(w_mem_inst__abc_19396_new_n4333_));
OAI21X1 OAI21X1_2232 ( .A(w_mem_inst_w_mem_4__4_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf94), .C(w_mem_inst__abc_19396_new_n4333_), .Y(w_mem_inst__abc_19396_new_n4334_));
OAI21X1 OAI21X1_2233 ( .A(w_mem_inst__abc_19396_new_n4331_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf38), .C(w_mem_inst__abc_19396_new_n4334_), .Y(w_mem_inst__0w_mem_3__31_0__4_));
OAI21X1 OAI21X1_2234 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf36), .B(w_mem_inst__abc_19396_new_n4337_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf93), .Y(w_mem_inst__abc_19396_new_n4338_));
OAI21X1 OAI21X1_2235 ( .A(w_mem_inst_w_mem_4__5_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf92), .C(w_mem_inst__abc_19396_new_n4338_), .Y(w_mem_inst__abc_19396_new_n4339_));
OAI21X1 OAI21X1_2236 ( .A(w_mem_inst__abc_19396_new_n4336_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf37), .C(w_mem_inst__abc_19396_new_n4339_), .Y(w_mem_inst__0w_mem_3__31_0__5_));
OAI21X1 OAI21X1_2237 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf35), .B(w_mem_inst__abc_19396_new_n4342_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf91), .Y(w_mem_inst__abc_19396_new_n4343_));
OAI21X1 OAI21X1_2238 ( .A(w_mem_inst_w_mem_4__6_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf90), .C(w_mem_inst__abc_19396_new_n4343_), .Y(w_mem_inst__abc_19396_new_n4344_));
OAI21X1 OAI21X1_2239 ( .A(w_mem_inst__abc_19396_new_n4341_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf36), .C(w_mem_inst__abc_19396_new_n4344_), .Y(w_mem_inst__0w_mem_3__31_0__6_));
OAI21X1 OAI21X1_224 ( .A(_abc_15497_new_n1756_), .B(_abc_15497_new_n873__bF_buf2), .C(_abc_15497_new_n1760_), .Y(_0H1_reg_31_0__1_));
OAI21X1 OAI21X1_2240 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf34), .B(w_mem_inst__abc_19396_new_n4347_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf89), .Y(w_mem_inst__abc_19396_new_n4348_));
OAI21X1 OAI21X1_2241 ( .A(w_mem_inst_w_mem_4__7_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf88), .C(w_mem_inst__abc_19396_new_n4348_), .Y(w_mem_inst__abc_19396_new_n4349_));
OAI21X1 OAI21X1_2242 ( .A(w_mem_inst__abc_19396_new_n4346_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf35), .C(w_mem_inst__abc_19396_new_n4349_), .Y(w_mem_inst__0w_mem_3__31_0__7_));
OAI21X1 OAI21X1_2243 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf33), .B(w_mem_inst__abc_19396_new_n4352_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf87), .Y(w_mem_inst__abc_19396_new_n4353_));
OAI21X1 OAI21X1_2244 ( .A(w_mem_inst_w_mem_4__8_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf86), .C(w_mem_inst__abc_19396_new_n4353_), .Y(w_mem_inst__abc_19396_new_n4354_));
OAI21X1 OAI21X1_2245 ( .A(w_mem_inst__abc_19396_new_n4351_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf34), .C(w_mem_inst__abc_19396_new_n4354_), .Y(w_mem_inst__0w_mem_3__31_0__8_));
OAI21X1 OAI21X1_2246 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf32), .B(w_mem_inst__abc_19396_new_n4357_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf85), .Y(w_mem_inst__abc_19396_new_n4358_));
OAI21X1 OAI21X1_2247 ( .A(w_mem_inst_w_mem_4__9_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf84), .C(w_mem_inst__abc_19396_new_n4358_), .Y(w_mem_inst__abc_19396_new_n4359_));
OAI21X1 OAI21X1_2248 ( .A(w_mem_inst__abc_19396_new_n4356_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf33), .C(w_mem_inst__abc_19396_new_n4359_), .Y(w_mem_inst__0w_mem_3__31_0__9_));
OAI21X1 OAI21X1_2249 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf31), .B(w_mem_inst__abc_19396_new_n4362_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf83), .Y(w_mem_inst__abc_19396_new_n4363_));
OAI21X1 OAI21X1_225 ( .A(_abc_15497_new_n1756_), .B(_abc_15497_new_n1763_), .C(_abc_15497_new_n1764_), .Y(_abc_15497_new_n1765_));
OAI21X1 OAI21X1_2250 ( .A(w_mem_inst_w_mem_4__10_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf82), .C(w_mem_inst__abc_19396_new_n4363_), .Y(w_mem_inst__abc_19396_new_n4364_));
OAI21X1 OAI21X1_2251 ( .A(w_mem_inst__abc_19396_new_n4361_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf32), .C(w_mem_inst__abc_19396_new_n4364_), .Y(w_mem_inst__0w_mem_3__31_0__10_));
OAI21X1 OAI21X1_2252 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf30), .B(w_mem_inst__abc_19396_new_n4367_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf81), .Y(w_mem_inst__abc_19396_new_n4368_));
OAI21X1 OAI21X1_2253 ( .A(w_mem_inst_w_mem_4__11_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf80), .C(w_mem_inst__abc_19396_new_n4368_), .Y(w_mem_inst__abc_19396_new_n4369_));
OAI21X1 OAI21X1_2254 ( .A(w_mem_inst__abc_19396_new_n4366_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf31), .C(w_mem_inst__abc_19396_new_n4369_), .Y(w_mem_inst__0w_mem_3__31_0__11_));
OAI21X1 OAI21X1_2255 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf29), .B(w_mem_inst__abc_19396_new_n4372_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf79), .Y(w_mem_inst__abc_19396_new_n4373_));
OAI21X1 OAI21X1_2256 ( .A(w_mem_inst_w_mem_4__12_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf78), .C(w_mem_inst__abc_19396_new_n4373_), .Y(w_mem_inst__abc_19396_new_n4374_));
OAI21X1 OAI21X1_2257 ( .A(w_mem_inst__abc_19396_new_n4371_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf30), .C(w_mem_inst__abc_19396_new_n4374_), .Y(w_mem_inst__0w_mem_3__31_0__12_));
OAI21X1 OAI21X1_2258 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf28), .B(w_mem_inst__abc_19396_new_n4377_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf77), .Y(w_mem_inst__abc_19396_new_n4378_));
OAI21X1 OAI21X1_2259 ( .A(w_mem_inst_w_mem_4__13_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf76), .C(w_mem_inst__abc_19396_new_n4378_), .Y(w_mem_inst__abc_19396_new_n4379_));
OAI21X1 OAI21X1_226 ( .A(_abc_15497_new_n1766_), .B(_abc_15497_new_n1765_), .C(digest_update_bF_buf8), .Y(_abc_15497_new_n1769_));
OAI21X1 OAI21X1_2260 ( .A(w_mem_inst__abc_19396_new_n4376_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf29), .C(w_mem_inst__abc_19396_new_n4379_), .Y(w_mem_inst__0w_mem_3__31_0__13_));
OAI21X1 OAI21X1_2261 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf27), .B(w_mem_inst__abc_19396_new_n4382_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf75), .Y(w_mem_inst__abc_19396_new_n4383_));
OAI21X1 OAI21X1_2262 ( .A(w_mem_inst_w_mem_4__14_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf74), .C(w_mem_inst__abc_19396_new_n4383_), .Y(w_mem_inst__abc_19396_new_n4384_));
OAI21X1 OAI21X1_2263 ( .A(w_mem_inst__abc_19396_new_n4381_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf28), .C(w_mem_inst__abc_19396_new_n4384_), .Y(w_mem_inst__0w_mem_3__31_0__14_));
OAI21X1 OAI21X1_2264 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf26), .B(w_mem_inst__abc_19396_new_n4387_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf73), .Y(w_mem_inst__abc_19396_new_n4388_));
OAI21X1 OAI21X1_2265 ( .A(w_mem_inst_w_mem_4__15_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf72), .C(w_mem_inst__abc_19396_new_n4388_), .Y(w_mem_inst__abc_19396_new_n4389_));
OAI21X1 OAI21X1_2266 ( .A(w_mem_inst__abc_19396_new_n4386_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf27), .C(w_mem_inst__abc_19396_new_n4389_), .Y(w_mem_inst__0w_mem_3__31_0__15_));
OAI21X1 OAI21X1_2267 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf25), .B(w_mem_inst__abc_19396_new_n4392_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf71), .Y(w_mem_inst__abc_19396_new_n4393_));
OAI21X1 OAI21X1_2268 ( .A(w_mem_inst_w_mem_4__16_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf70), .C(w_mem_inst__abc_19396_new_n4393_), .Y(w_mem_inst__abc_19396_new_n4394_));
OAI21X1 OAI21X1_2269 ( .A(w_mem_inst__abc_19396_new_n4391_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf26), .C(w_mem_inst__abc_19396_new_n4394_), .Y(w_mem_inst__0w_mem_3__31_0__16_));
OAI21X1 OAI21X1_227 ( .A(_abc_15497_new_n1762_), .B(_abc_15497_new_n1771_), .C(_abc_15497_new_n1767_), .Y(_abc_15497_new_n1772_));
OAI21X1 OAI21X1_2270 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf24), .B(w_mem_inst__abc_19396_new_n4397_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf69), .Y(w_mem_inst__abc_19396_new_n4398_));
OAI21X1 OAI21X1_2271 ( .A(w_mem_inst_w_mem_4__17_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf68), .C(w_mem_inst__abc_19396_new_n4398_), .Y(w_mem_inst__abc_19396_new_n4399_));
OAI21X1 OAI21X1_2272 ( .A(w_mem_inst__abc_19396_new_n4396_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf25), .C(w_mem_inst__abc_19396_new_n4399_), .Y(w_mem_inst__0w_mem_3__31_0__17_));
OAI21X1 OAI21X1_2273 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf23), .B(w_mem_inst__abc_19396_new_n4402_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf67), .Y(w_mem_inst__abc_19396_new_n4403_));
OAI21X1 OAI21X1_2274 ( .A(w_mem_inst_w_mem_4__18_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf66), .C(w_mem_inst__abc_19396_new_n4403_), .Y(w_mem_inst__abc_19396_new_n4404_));
OAI21X1 OAI21X1_2275 ( .A(w_mem_inst__abc_19396_new_n4401_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf24), .C(w_mem_inst__abc_19396_new_n4404_), .Y(w_mem_inst__0w_mem_3__31_0__18_));
OAI21X1 OAI21X1_2276 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf22), .B(w_mem_inst__abc_19396_new_n4407_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf65), .Y(w_mem_inst__abc_19396_new_n4408_));
OAI21X1 OAI21X1_2277 ( .A(w_mem_inst_w_mem_4__19_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf64), .C(w_mem_inst__abc_19396_new_n4408_), .Y(w_mem_inst__abc_19396_new_n4409_));
OAI21X1 OAI21X1_2278 ( .A(w_mem_inst__abc_19396_new_n4406_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf23), .C(w_mem_inst__abc_19396_new_n4409_), .Y(w_mem_inst__0w_mem_3__31_0__19_));
OAI21X1 OAI21X1_2279 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf21), .B(w_mem_inst__abc_19396_new_n4412_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf63), .Y(w_mem_inst__abc_19396_new_n4413_));
OAI21X1 OAI21X1_228 ( .A(_auto_iopadmap_cc_368_execute_22625_99_), .B(_abc_15497_new_n883__bF_buf10), .C(_abc_15497_new_n870__bF_buf11), .Y(_abc_15497_new_n1777_));
OAI21X1 OAI21X1_2280 ( .A(w_mem_inst_w_mem_4__20_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf62), .C(w_mem_inst__abc_19396_new_n4413_), .Y(w_mem_inst__abc_19396_new_n4414_));
OAI21X1 OAI21X1_2281 ( .A(w_mem_inst__abc_19396_new_n4411_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf22), .C(w_mem_inst__abc_19396_new_n4414_), .Y(w_mem_inst__0w_mem_3__31_0__20_));
OAI21X1 OAI21X1_2282 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf20), .B(w_mem_inst__abc_19396_new_n4417_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf61), .Y(w_mem_inst__abc_19396_new_n4418_));
OAI21X1 OAI21X1_2283 ( .A(w_mem_inst_w_mem_4__21_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf60), .C(w_mem_inst__abc_19396_new_n4418_), .Y(w_mem_inst__abc_19396_new_n4419_));
OAI21X1 OAI21X1_2284 ( .A(w_mem_inst__abc_19396_new_n4416_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf21), .C(w_mem_inst__abc_19396_new_n4419_), .Y(w_mem_inst__0w_mem_3__31_0__21_));
OAI21X1 OAI21X1_2285 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf19), .B(w_mem_inst__abc_19396_new_n4422_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf59), .Y(w_mem_inst__abc_19396_new_n4423_));
OAI21X1 OAI21X1_2286 ( .A(w_mem_inst_w_mem_4__22_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf58), .C(w_mem_inst__abc_19396_new_n4423_), .Y(w_mem_inst__abc_19396_new_n4424_));
OAI21X1 OAI21X1_2287 ( .A(w_mem_inst__abc_19396_new_n4421_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf20), .C(w_mem_inst__abc_19396_new_n4424_), .Y(w_mem_inst__0w_mem_3__31_0__22_));
OAI21X1 OAI21X1_2288 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf18), .B(w_mem_inst__abc_19396_new_n4427_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf57), .Y(w_mem_inst__abc_19396_new_n4428_));
OAI21X1 OAI21X1_2289 ( .A(w_mem_inst_w_mem_4__23_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf56), .C(w_mem_inst__abc_19396_new_n4428_), .Y(w_mem_inst__abc_19396_new_n4429_));
OAI21X1 OAI21X1_229 ( .A(_abc_15497_new_n870__bF_buf10), .B(_abc_15497_new_n1776_), .C(_abc_15497_new_n1777_), .Y(_0H1_reg_31_0__3_));
OAI21X1 OAI21X1_2290 ( .A(w_mem_inst__abc_19396_new_n4426_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf19), .C(w_mem_inst__abc_19396_new_n4429_), .Y(w_mem_inst__0w_mem_3__31_0__23_));
OAI21X1 OAI21X1_2291 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf17), .B(w_mem_inst__abc_19396_new_n4432_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf55), .Y(w_mem_inst__abc_19396_new_n4433_));
OAI21X1 OAI21X1_2292 ( .A(w_mem_inst_w_mem_4__24_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf54), .C(w_mem_inst__abc_19396_new_n4433_), .Y(w_mem_inst__abc_19396_new_n4434_));
OAI21X1 OAI21X1_2293 ( .A(w_mem_inst__abc_19396_new_n4431_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf18), .C(w_mem_inst__abc_19396_new_n4434_), .Y(w_mem_inst__0w_mem_3__31_0__24_));
OAI21X1 OAI21X1_2294 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf16), .B(w_mem_inst__abc_19396_new_n4437_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf53), .Y(w_mem_inst__abc_19396_new_n4438_));
OAI21X1 OAI21X1_2295 ( .A(w_mem_inst_w_mem_4__25_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf52), .C(w_mem_inst__abc_19396_new_n4438_), .Y(w_mem_inst__abc_19396_new_n4439_));
OAI21X1 OAI21X1_2296 ( .A(w_mem_inst__abc_19396_new_n4436_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf17), .C(w_mem_inst__abc_19396_new_n4439_), .Y(w_mem_inst__0w_mem_3__31_0__25_));
OAI21X1 OAI21X1_2297 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf15), .B(w_mem_inst__abc_19396_new_n4442_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf51), .Y(w_mem_inst__abc_19396_new_n4443_));
OAI21X1 OAI21X1_2298 ( .A(w_mem_inst_w_mem_4__26_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf50), .C(w_mem_inst__abc_19396_new_n4443_), .Y(w_mem_inst__abc_19396_new_n4444_));
OAI21X1 OAI21X1_2299 ( .A(w_mem_inst__abc_19396_new_n4441_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf16), .C(w_mem_inst__abc_19396_new_n4444_), .Y(w_mem_inst__0w_mem_3__31_0__26_));
OAI21X1 OAI21X1_23 ( .A(_auto_iopadmap_cc_368_execute_22625_95_), .B(_abc_15497_new_n883__bF_buf11), .C(_abc_15497_new_n870__bF_buf6), .Y(_abc_15497_new_n934_));
OAI21X1 OAI21X1_230 ( .A(_abc_15497_new_n1791_), .B(_abc_15497_new_n1793_), .C(_abc_15497_new_n1790_), .Y(_abc_15497_new_n1794_));
OAI21X1 OAI21X1_2300 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf14), .B(w_mem_inst__abc_19396_new_n4447_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf49), .Y(w_mem_inst__abc_19396_new_n4448_));
OAI21X1 OAI21X1_2301 ( .A(w_mem_inst_w_mem_4__27_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf48), .C(w_mem_inst__abc_19396_new_n4448_), .Y(w_mem_inst__abc_19396_new_n4449_));
OAI21X1 OAI21X1_2302 ( .A(w_mem_inst__abc_19396_new_n4446_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf15), .C(w_mem_inst__abc_19396_new_n4449_), .Y(w_mem_inst__0w_mem_3__31_0__27_));
OAI21X1 OAI21X1_2303 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf13), .B(w_mem_inst__abc_19396_new_n4452_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf47), .Y(w_mem_inst__abc_19396_new_n4453_));
OAI21X1 OAI21X1_2304 ( .A(w_mem_inst_w_mem_4__28_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf46), .C(w_mem_inst__abc_19396_new_n4453_), .Y(w_mem_inst__abc_19396_new_n4454_));
OAI21X1 OAI21X1_2305 ( .A(w_mem_inst__abc_19396_new_n4451_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf14), .C(w_mem_inst__abc_19396_new_n4454_), .Y(w_mem_inst__0w_mem_3__31_0__28_));
OAI21X1 OAI21X1_2306 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf12), .B(w_mem_inst__abc_19396_new_n4457_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf45), .Y(w_mem_inst__abc_19396_new_n4458_));
OAI21X1 OAI21X1_2307 ( .A(w_mem_inst_w_mem_4__29_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf44), .C(w_mem_inst__abc_19396_new_n4458_), .Y(w_mem_inst__abc_19396_new_n4459_));
OAI21X1 OAI21X1_2308 ( .A(w_mem_inst__abc_19396_new_n4456_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf13), .C(w_mem_inst__abc_19396_new_n4459_), .Y(w_mem_inst__0w_mem_3__31_0__29_));
OAI21X1 OAI21X1_2309 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf11), .B(w_mem_inst__abc_19396_new_n4462_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf43), .Y(w_mem_inst__abc_19396_new_n4463_));
OAI21X1 OAI21X1_231 ( .A(_abc_15497_new_n1789_), .B(_abc_15497_new_n1783_), .C(_abc_15497_new_n1795_), .Y(_abc_15497_new_n1796_));
OAI21X1 OAI21X1_2310 ( .A(w_mem_inst_w_mem_4__30_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf42), .C(w_mem_inst__abc_19396_new_n4463_), .Y(w_mem_inst__abc_19396_new_n4464_));
OAI21X1 OAI21X1_2311 ( .A(w_mem_inst__abc_19396_new_n4461_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf12), .C(w_mem_inst__abc_19396_new_n4464_), .Y(w_mem_inst__0w_mem_3__31_0__30_));
OAI21X1 OAI21X1_2312 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf10), .B(w_mem_inst__abc_19396_new_n4467_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf41), .Y(w_mem_inst__abc_19396_new_n4468_));
OAI21X1 OAI21X1_2313 ( .A(w_mem_inst_w_mem_4__31_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf40), .C(w_mem_inst__abc_19396_new_n4468_), .Y(w_mem_inst__abc_19396_new_n4469_));
OAI21X1 OAI21X1_2314 ( .A(w_mem_inst__abc_19396_new_n4466_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf11), .C(w_mem_inst__abc_19396_new_n4469_), .Y(w_mem_inst__0w_mem_3__31_0__31_));
OAI21X1 OAI21X1_2315 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf9), .B(w_mem_inst__abc_19396_new_n4472_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf39), .Y(w_mem_inst__abc_19396_new_n4473_));
OAI21X1 OAI21X1_2316 ( .A(w_mem_inst_w_mem_3__0_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf38), .C(w_mem_inst__abc_19396_new_n4473_), .Y(w_mem_inst__abc_19396_new_n4474_));
OAI21X1 OAI21X1_2317 ( .A(w_mem_inst__abc_19396_new_n4471_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf10), .C(w_mem_inst__abc_19396_new_n4474_), .Y(w_mem_inst__0w_mem_2__31_0__0_));
OAI21X1 OAI21X1_2318 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf8), .B(w_mem_inst__abc_19396_new_n4477_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf37), .Y(w_mem_inst__abc_19396_new_n4478_));
OAI21X1 OAI21X1_2319 ( .A(w_mem_inst_w_mem_3__1_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf36), .C(w_mem_inst__abc_19396_new_n4478_), .Y(w_mem_inst__abc_19396_new_n4479_));
OAI21X1 OAI21X1_232 ( .A(_abc_15497_new_n1787_), .B(_abc_15497_new_n1792_), .C(_abc_15497_new_n1796_), .Y(_abc_15497_new_n1800_));
OAI21X1 OAI21X1_2320 ( .A(w_mem_inst__abc_19396_new_n4476_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf9), .C(w_mem_inst__abc_19396_new_n4479_), .Y(w_mem_inst__0w_mem_2__31_0__1_));
OAI21X1 OAI21X1_2321 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf7), .B(w_mem_inst__abc_19396_new_n4482_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf35), .Y(w_mem_inst__abc_19396_new_n4483_));
OAI21X1 OAI21X1_2322 ( .A(w_mem_inst_w_mem_3__2_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf34), .C(w_mem_inst__abc_19396_new_n4483_), .Y(w_mem_inst__abc_19396_new_n4484_));
OAI21X1 OAI21X1_2323 ( .A(w_mem_inst__abc_19396_new_n4481_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf8), .C(w_mem_inst__abc_19396_new_n4484_), .Y(w_mem_inst__0w_mem_2__31_0__2_));
OAI21X1 OAI21X1_2324 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf6), .B(w_mem_inst__abc_19396_new_n4487_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf33), .Y(w_mem_inst__abc_19396_new_n4488_));
OAI21X1 OAI21X1_2325 ( .A(w_mem_inst_w_mem_3__3_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf32), .C(w_mem_inst__abc_19396_new_n4488_), .Y(w_mem_inst__abc_19396_new_n4489_));
OAI21X1 OAI21X1_2326 ( .A(w_mem_inst__abc_19396_new_n4486_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf7), .C(w_mem_inst__abc_19396_new_n4489_), .Y(w_mem_inst__0w_mem_2__31_0__3_));
OAI21X1 OAI21X1_2327 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf5), .B(w_mem_inst__abc_19396_new_n4492_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf31), .Y(w_mem_inst__abc_19396_new_n4493_));
OAI21X1 OAI21X1_2328 ( .A(w_mem_inst_w_mem_3__4_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf30), .C(w_mem_inst__abc_19396_new_n4493_), .Y(w_mem_inst__abc_19396_new_n4494_));
OAI21X1 OAI21X1_2329 ( .A(w_mem_inst__abc_19396_new_n4491_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf6), .C(w_mem_inst__abc_19396_new_n4494_), .Y(w_mem_inst__0w_mem_2__31_0__4_));
OAI21X1 OAI21X1_233 ( .A(_abc_15497_new_n1814_), .B(_abc_15497_new_n1813_), .C(digest_update_bF_buf6), .Y(_abc_15497_new_n1815_));
OAI21X1 OAI21X1_2330 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf4), .B(w_mem_inst__abc_19396_new_n4497_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf29), .Y(w_mem_inst__abc_19396_new_n4498_));
OAI21X1 OAI21X1_2331 ( .A(w_mem_inst_w_mem_3__5_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf28), .C(w_mem_inst__abc_19396_new_n4498_), .Y(w_mem_inst__abc_19396_new_n4499_));
OAI21X1 OAI21X1_2332 ( .A(w_mem_inst__abc_19396_new_n4496_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf5), .C(w_mem_inst__abc_19396_new_n4499_), .Y(w_mem_inst__0w_mem_2__31_0__5_));
OAI21X1 OAI21X1_2333 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf3), .B(w_mem_inst__abc_19396_new_n4502_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf27), .Y(w_mem_inst__abc_19396_new_n4503_));
OAI21X1 OAI21X1_2334 ( .A(w_mem_inst_w_mem_3__6_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf26), .C(w_mem_inst__abc_19396_new_n4503_), .Y(w_mem_inst__abc_19396_new_n4504_));
OAI21X1 OAI21X1_2335 ( .A(w_mem_inst__abc_19396_new_n4501_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf4), .C(w_mem_inst__abc_19396_new_n4504_), .Y(w_mem_inst__0w_mem_2__31_0__6_));
OAI21X1 OAI21X1_2336 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf2), .B(w_mem_inst__abc_19396_new_n4507_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf25), .Y(w_mem_inst__abc_19396_new_n4508_));
OAI21X1 OAI21X1_2337 ( .A(w_mem_inst_w_mem_3__7_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf24), .C(w_mem_inst__abc_19396_new_n4508_), .Y(w_mem_inst__abc_19396_new_n4509_));
OAI21X1 OAI21X1_2338 ( .A(w_mem_inst__abc_19396_new_n4506_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf3), .C(w_mem_inst__abc_19396_new_n4509_), .Y(w_mem_inst__0w_mem_2__31_0__7_));
OAI21X1 OAI21X1_2339 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf1), .B(w_mem_inst__abc_19396_new_n4512_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf23), .Y(w_mem_inst__abc_19396_new_n4513_));
OAI21X1 OAI21X1_234 ( .A(_auto_iopadmap_cc_368_execute_22625_103_), .B(_abc_15497_new_n883__bF_buf9), .C(_abc_15497_new_n870__bF_buf7), .Y(_abc_15497_new_n1816_));
OAI21X1 OAI21X1_2340 ( .A(w_mem_inst_w_mem_3__8_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf22), .C(w_mem_inst__abc_19396_new_n4513_), .Y(w_mem_inst__abc_19396_new_n4514_));
OAI21X1 OAI21X1_2341 ( .A(w_mem_inst__abc_19396_new_n4511_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf2), .C(w_mem_inst__abc_19396_new_n4514_), .Y(w_mem_inst__0w_mem_2__31_0__8_));
OAI21X1 OAI21X1_2342 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf0), .B(w_mem_inst__abc_19396_new_n4517_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf21), .Y(w_mem_inst__abc_19396_new_n4518_));
OAI21X1 OAI21X1_2343 ( .A(w_mem_inst_w_mem_3__9_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf20), .C(w_mem_inst__abc_19396_new_n4518_), .Y(w_mem_inst__abc_19396_new_n4519_));
OAI21X1 OAI21X1_2344 ( .A(w_mem_inst__abc_19396_new_n4516_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf1), .C(w_mem_inst__abc_19396_new_n4519_), .Y(w_mem_inst__0w_mem_2__31_0__9_));
OAI21X1 OAI21X1_2345 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf60), .B(w_mem_inst__abc_19396_new_n4522_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf19), .Y(w_mem_inst__abc_19396_new_n4523_));
OAI21X1 OAI21X1_2346 ( .A(w_mem_inst_w_mem_3__10_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf18), .C(w_mem_inst__abc_19396_new_n4523_), .Y(w_mem_inst__abc_19396_new_n4524_));
OAI21X1 OAI21X1_2347 ( .A(w_mem_inst__abc_19396_new_n4521_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf0), .C(w_mem_inst__abc_19396_new_n4524_), .Y(w_mem_inst__0w_mem_2__31_0__10_));
OAI21X1 OAI21X1_2348 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf59), .B(w_mem_inst__abc_19396_new_n4527_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf17), .Y(w_mem_inst__abc_19396_new_n4528_));
OAI21X1 OAI21X1_2349 ( .A(w_mem_inst_w_mem_3__11_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf16), .C(w_mem_inst__abc_19396_new_n4528_), .Y(w_mem_inst__abc_19396_new_n4529_));
OAI21X1 OAI21X1_235 ( .A(_auto_iopadmap_cc_368_execute_22625_103_), .B(b_reg_7_), .C(_abc_15497_new_n1823_), .Y(_abc_15497_new_n1824_));
OAI21X1 OAI21X1_2350 ( .A(w_mem_inst__abc_19396_new_n4526_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf60), .C(w_mem_inst__abc_19396_new_n4529_), .Y(w_mem_inst__0w_mem_2__31_0__11_));
OAI21X1 OAI21X1_2351 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf58), .B(w_mem_inst__abc_19396_new_n4532_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf15), .Y(w_mem_inst__abc_19396_new_n4533_));
OAI21X1 OAI21X1_2352 ( .A(w_mem_inst_w_mem_3__12_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf14), .C(w_mem_inst__abc_19396_new_n4533_), .Y(w_mem_inst__abc_19396_new_n4534_));
OAI21X1 OAI21X1_2353 ( .A(w_mem_inst__abc_19396_new_n4531_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf59), .C(w_mem_inst__abc_19396_new_n4534_), .Y(w_mem_inst__0w_mem_2__31_0__12_));
OAI21X1 OAI21X1_2354 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf57), .B(w_mem_inst__abc_19396_new_n4537_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf13), .Y(w_mem_inst__abc_19396_new_n4538_));
OAI21X1 OAI21X1_2355 ( .A(w_mem_inst_w_mem_3__13_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf12), .C(w_mem_inst__abc_19396_new_n4538_), .Y(w_mem_inst__abc_19396_new_n4539_));
OAI21X1 OAI21X1_2356 ( .A(w_mem_inst__abc_19396_new_n4536_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf58), .C(w_mem_inst__abc_19396_new_n4539_), .Y(w_mem_inst__0w_mem_2__31_0__13_));
OAI21X1 OAI21X1_2357 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf56), .B(w_mem_inst__abc_19396_new_n4542_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf11), .Y(w_mem_inst__abc_19396_new_n4543_));
OAI21X1 OAI21X1_2358 ( .A(w_mem_inst_w_mem_3__14_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf10), .C(w_mem_inst__abc_19396_new_n4543_), .Y(w_mem_inst__abc_19396_new_n4544_));
OAI21X1 OAI21X1_2359 ( .A(w_mem_inst__abc_19396_new_n4541_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf57), .C(w_mem_inst__abc_19396_new_n4544_), .Y(w_mem_inst__0w_mem_2__31_0__14_));
OAI21X1 OAI21X1_236 ( .A(_auto_iopadmap_cc_368_execute_22625_104_), .B(_abc_15497_new_n883__bF_buf8), .C(_abc_15497_new_n870__bF_buf6), .Y(_abc_15497_new_n1827_));
OAI21X1 OAI21X1_2360 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf55), .B(w_mem_inst__abc_19396_new_n4547_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf9), .Y(w_mem_inst__abc_19396_new_n4548_));
OAI21X1 OAI21X1_2361 ( .A(w_mem_inst_w_mem_3__15_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf8), .C(w_mem_inst__abc_19396_new_n4548_), .Y(w_mem_inst__abc_19396_new_n4549_));
OAI21X1 OAI21X1_2362 ( .A(w_mem_inst__abc_19396_new_n4546_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf56), .C(w_mem_inst__abc_19396_new_n4549_), .Y(w_mem_inst__0w_mem_2__31_0__15_));
OAI21X1 OAI21X1_2363 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf54), .B(w_mem_inst__abc_19396_new_n4552_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf7), .Y(w_mem_inst__abc_19396_new_n4553_));
OAI21X1 OAI21X1_2364 ( .A(w_mem_inst_w_mem_3__16_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf6), .C(w_mem_inst__abc_19396_new_n4553_), .Y(w_mem_inst__abc_19396_new_n4554_));
OAI21X1 OAI21X1_2365 ( .A(w_mem_inst__abc_19396_new_n4551_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf55), .C(w_mem_inst__abc_19396_new_n4554_), .Y(w_mem_inst__0w_mem_2__31_0__16_));
OAI21X1 OAI21X1_2366 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf53), .B(w_mem_inst__abc_19396_new_n4557_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf5), .Y(w_mem_inst__abc_19396_new_n4558_));
OAI21X1 OAI21X1_2367 ( .A(w_mem_inst_w_mem_3__17_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf4), .C(w_mem_inst__abc_19396_new_n4558_), .Y(w_mem_inst__abc_19396_new_n4559_));
OAI21X1 OAI21X1_2368 ( .A(w_mem_inst__abc_19396_new_n4556_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf54), .C(w_mem_inst__abc_19396_new_n4559_), .Y(w_mem_inst__0w_mem_2__31_0__17_));
OAI21X1 OAI21X1_2369 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf52), .B(w_mem_inst__abc_19396_new_n4562_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf3), .Y(w_mem_inst__abc_19396_new_n4563_));
OAI21X1 OAI21X1_237 ( .A(_abc_15497_new_n870__bF_buf5), .B(_abc_15497_new_n1826_), .C(_abc_15497_new_n1827_), .Y(_0H1_reg_31_0__8_));
OAI21X1 OAI21X1_2370 ( .A(w_mem_inst_w_mem_3__18_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf2), .C(w_mem_inst__abc_19396_new_n4563_), .Y(w_mem_inst__abc_19396_new_n4564_));
OAI21X1 OAI21X1_2371 ( .A(w_mem_inst__abc_19396_new_n4561_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf53), .C(w_mem_inst__abc_19396_new_n4564_), .Y(w_mem_inst__0w_mem_2__31_0__18_));
OAI21X1 OAI21X1_2372 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf51), .B(w_mem_inst__abc_19396_new_n4567_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf1), .Y(w_mem_inst__abc_19396_new_n4568_));
OAI21X1 OAI21X1_2373 ( .A(w_mem_inst_w_mem_3__19_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf0), .C(w_mem_inst__abc_19396_new_n4568_), .Y(w_mem_inst__abc_19396_new_n4569_));
OAI21X1 OAI21X1_2374 ( .A(w_mem_inst__abc_19396_new_n4566_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf52), .C(w_mem_inst__abc_19396_new_n4569_), .Y(w_mem_inst__0w_mem_2__31_0__19_));
OAI21X1 OAI21X1_2375 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf50), .B(w_mem_inst__abc_19396_new_n4572_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf96), .Y(w_mem_inst__abc_19396_new_n4573_));
OAI21X1 OAI21X1_2376 ( .A(w_mem_inst_w_mem_3__20_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf95), .C(w_mem_inst__abc_19396_new_n4573_), .Y(w_mem_inst__abc_19396_new_n4574_));
OAI21X1 OAI21X1_2377 ( .A(w_mem_inst__abc_19396_new_n4571_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf51), .C(w_mem_inst__abc_19396_new_n4574_), .Y(w_mem_inst__0w_mem_2__31_0__20_));
OAI21X1 OAI21X1_2378 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf49), .B(w_mem_inst__abc_19396_new_n4577_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf94), .Y(w_mem_inst__abc_19396_new_n4578_));
OAI21X1 OAI21X1_2379 ( .A(w_mem_inst_w_mem_3__21_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf93), .C(w_mem_inst__abc_19396_new_n4578_), .Y(w_mem_inst__abc_19396_new_n4579_));
OAI21X1 OAI21X1_238 ( .A(_auto_iopadmap_cc_368_execute_22625_105_), .B(_abc_15497_new_n883__bF_buf7), .C(_abc_15497_new_n870__bF_buf4), .Y(_abc_15497_new_n1834_));
OAI21X1 OAI21X1_2380 ( .A(w_mem_inst__abc_19396_new_n4576_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf50), .C(w_mem_inst__abc_19396_new_n4579_), .Y(w_mem_inst__0w_mem_2__31_0__21_));
OAI21X1 OAI21X1_2381 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf48), .B(w_mem_inst__abc_19396_new_n4582_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf92), .Y(w_mem_inst__abc_19396_new_n4583_));
OAI21X1 OAI21X1_2382 ( .A(w_mem_inst_w_mem_3__22_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf91), .C(w_mem_inst__abc_19396_new_n4583_), .Y(w_mem_inst__abc_19396_new_n4584_));
OAI21X1 OAI21X1_2383 ( .A(w_mem_inst__abc_19396_new_n4581_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf49), .C(w_mem_inst__abc_19396_new_n4584_), .Y(w_mem_inst__0w_mem_2__31_0__22_));
OAI21X1 OAI21X1_2384 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf47), .B(w_mem_inst__abc_19396_new_n4587_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf90), .Y(w_mem_inst__abc_19396_new_n4588_));
OAI21X1 OAI21X1_2385 ( .A(w_mem_inst_w_mem_3__23_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf89), .C(w_mem_inst__abc_19396_new_n4588_), .Y(w_mem_inst__abc_19396_new_n4589_));
OAI21X1 OAI21X1_2386 ( .A(w_mem_inst__abc_19396_new_n4586_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf48), .C(w_mem_inst__abc_19396_new_n4589_), .Y(w_mem_inst__0w_mem_2__31_0__23_));
OAI21X1 OAI21X1_2387 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf46), .B(w_mem_inst__abc_19396_new_n4592_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf88), .Y(w_mem_inst__abc_19396_new_n4593_));
OAI21X1 OAI21X1_2388 ( .A(w_mem_inst_w_mem_3__24_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf87), .C(w_mem_inst__abc_19396_new_n4593_), .Y(w_mem_inst__abc_19396_new_n4594_));
OAI21X1 OAI21X1_2389 ( .A(w_mem_inst__abc_19396_new_n4591_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf47), .C(w_mem_inst__abc_19396_new_n4594_), .Y(w_mem_inst__0w_mem_2__31_0__24_));
OAI21X1 OAI21X1_239 ( .A(_abc_15497_new_n870__bF_buf3), .B(_abc_15497_new_n1833_), .C(_abc_15497_new_n1834_), .Y(_0H1_reg_31_0__9_));
OAI21X1 OAI21X1_2390 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf45), .B(w_mem_inst__abc_19396_new_n4597_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf86), .Y(w_mem_inst__abc_19396_new_n4598_));
OAI21X1 OAI21X1_2391 ( .A(w_mem_inst_w_mem_3__25_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf85), .C(w_mem_inst__abc_19396_new_n4598_), .Y(w_mem_inst__abc_19396_new_n4599_));
OAI21X1 OAI21X1_2392 ( .A(w_mem_inst__abc_19396_new_n4596_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf46), .C(w_mem_inst__abc_19396_new_n4599_), .Y(w_mem_inst__0w_mem_2__31_0__25_));
OAI21X1 OAI21X1_2393 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf44), .B(w_mem_inst__abc_19396_new_n4602_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf84), .Y(w_mem_inst__abc_19396_new_n4603_));
OAI21X1 OAI21X1_2394 ( .A(w_mem_inst_w_mem_3__26_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf83), .C(w_mem_inst__abc_19396_new_n4603_), .Y(w_mem_inst__abc_19396_new_n4604_));
OAI21X1 OAI21X1_2395 ( .A(w_mem_inst__abc_19396_new_n4601_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf45), .C(w_mem_inst__abc_19396_new_n4604_), .Y(w_mem_inst__0w_mem_2__31_0__26_));
OAI21X1 OAI21X1_2396 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf43), .B(w_mem_inst__abc_19396_new_n4607_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf82), .Y(w_mem_inst__abc_19396_new_n4608_));
OAI21X1 OAI21X1_2397 ( .A(w_mem_inst_w_mem_3__27_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf81), .C(w_mem_inst__abc_19396_new_n4608_), .Y(w_mem_inst__abc_19396_new_n4609_));
OAI21X1 OAI21X1_2398 ( .A(w_mem_inst__abc_19396_new_n4606_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf44), .C(w_mem_inst__abc_19396_new_n4609_), .Y(w_mem_inst__0w_mem_2__31_0__27_));
OAI21X1 OAI21X1_2399 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf42), .B(w_mem_inst__abc_19396_new_n4612_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf80), .Y(w_mem_inst__abc_19396_new_n4613_));
OAI21X1 OAI21X1_24 ( .A(_abc_15497_new_n870__bF_buf5), .B(_abc_15497_new_n933_), .C(_abc_15497_new_n934_), .Y(_0H2_reg_31_0__31_));
OAI21X1 OAI21X1_240 ( .A(_abc_15497_new_n1837_), .B(_abc_15497_new_n1824_), .C(_abc_15497_new_n1838_), .Y(_abc_15497_new_n1839_));
OAI21X1 OAI21X1_2400 ( .A(w_mem_inst_w_mem_3__28_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf79), .C(w_mem_inst__abc_19396_new_n4613_), .Y(w_mem_inst__abc_19396_new_n4614_));
OAI21X1 OAI21X1_2401 ( .A(w_mem_inst__abc_19396_new_n4611_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf43), .C(w_mem_inst__abc_19396_new_n4614_), .Y(w_mem_inst__0w_mem_2__31_0__28_));
OAI21X1 OAI21X1_2402 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf41), .B(w_mem_inst__abc_19396_new_n4617_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf78), .Y(w_mem_inst__abc_19396_new_n4618_));
OAI21X1 OAI21X1_2403 ( .A(w_mem_inst_w_mem_3__29_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf77), .C(w_mem_inst__abc_19396_new_n4618_), .Y(w_mem_inst__abc_19396_new_n4619_));
OAI21X1 OAI21X1_2404 ( .A(w_mem_inst__abc_19396_new_n4616_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf42), .C(w_mem_inst__abc_19396_new_n4619_), .Y(w_mem_inst__0w_mem_2__31_0__29_));
OAI21X1 OAI21X1_2405 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf40), .B(w_mem_inst__abc_19396_new_n4622_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf76), .Y(w_mem_inst__abc_19396_new_n4623_));
OAI21X1 OAI21X1_2406 ( .A(w_mem_inst_w_mem_3__30_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf75), .C(w_mem_inst__abc_19396_new_n4623_), .Y(w_mem_inst__abc_19396_new_n4624_));
OAI21X1 OAI21X1_2407 ( .A(w_mem_inst__abc_19396_new_n4621_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf41), .C(w_mem_inst__abc_19396_new_n4624_), .Y(w_mem_inst__0w_mem_2__31_0__30_));
OAI21X1 OAI21X1_2408 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf39), .B(w_mem_inst__abc_19396_new_n4627_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf74), .Y(w_mem_inst__abc_19396_new_n4628_));
OAI21X1 OAI21X1_2409 ( .A(w_mem_inst_w_mem_3__31_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf73), .C(w_mem_inst__abc_19396_new_n4628_), .Y(w_mem_inst__abc_19396_new_n4629_));
OAI21X1 OAI21X1_241 ( .A(_abc_15497_new_n1836_), .B(_abc_15497_new_n1841_), .C(_abc_15497_new_n1845_), .Y(_abc_15497_new_n1848_));
OAI21X1 OAI21X1_2410 ( .A(w_mem_inst__abc_19396_new_n4626_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf40), .C(w_mem_inst__abc_19396_new_n4629_), .Y(w_mem_inst__0w_mem_2__31_0__31_));
OAI21X1 OAI21X1_2411 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf38), .B(w_mem_inst__abc_19396_new_n4632_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf72), .Y(w_mem_inst__abc_19396_new_n4633_));
OAI21X1 OAI21X1_2412 ( .A(w_mem_inst_w_mem_1__0_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf71), .C(w_mem_inst__abc_19396_new_n4633_), .Y(w_mem_inst__abc_19396_new_n4634_));
OAI21X1 OAI21X1_2413 ( .A(w_mem_inst__abc_19396_new_n4631_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf39), .C(w_mem_inst__abc_19396_new_n4634_), .Y(w_mem_inst__0w_mem_0__31_0__0_));
OAI21X1 OAI21X1_2414 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf37), .B(w_mem_inst__abc_19396_new_n4637_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf70), .Y(w_mem_inst__abc_19396_new_n4638_));
OAI21X1 OAI21X1_2415 ( .A(w_mem_inst_w_mem_1__1_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf69), .C(w_mem_inst__abc_19396_new_n4638_), .Y(w_mem_inst__abc_19396_new_n4639_));
OAI21X1 OAI21X1_2416 ( .A(w_mem_inst__abc_19396_new_n4636_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf38), .C(w_mem_inst__abc_19396_new_n4639_), .Y(w_mem_inst__0w_mem_0__31_0__1_));
OAI21X1 OAI21X1_2417 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf36), .B(w_mem_inst__abc_19396_new_n4642_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf68), .Y(w_mem_inst__abc_19396_new_n4643_));
OAI21X1 OAI21X1_2418 ( .A(w_mem_inst_w_mem_1__2_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf67), .C(w_mem_inst__abc_19396_new_n4643_), .Y(w_mem_inst__abc_19396_new_n4644_));
OAI21X1 OAI21X1_2419 ( .A(w_mem_inst__abc_19396_new_n4641_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf37), .C(w_mem_inst__abc_19396_new_n4644_), .Y(w_mem_inst__0w_mem_0__31_0__2_));
OAI21X1 OAI21X1_242 ( .A(_auto_iopadmap_cc_368_execute_22625_107_), .B(_abc_15497_new_n883__bF_buf6), .C(_abc_15497_new_n870__bF_buf2), .Y(_abc_15497_new_n1854_));
OAI21X1 OAI21X1_2420 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf35), .B(w_mem_inst__abc_19396_new_n4647_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf66), .Y(w_mem_inst__abc_19396_new_n4648_));
OAI21X1 OAI21X1_2421 ( .A(w_mem_inst_w_mem_1__3_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf65), .C(w_mem_inst__abc_19396_new_n4648_), .Y(w_mem_inst__abc_19396_new_n4649_));
OAI21X1 OAI21X1_2422 ( .A(w_mem_inst__abc_19396_new_n4646_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf36), .C(w_mem_inst__abc_19396_new_n4649_), .Y(w_mem_inst__0w_mem_0__31_0__3_));
OAI21X1 OAI21X1_2423 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf34), .B(w_mem_inst__abc_19396_new_n4652_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf64), .Y(w_mem_inst__abc_19396_new_n4653_));
OAI21X1 OAI21X1_2424 ( .A(w_mem_inst_w_mem_1__4_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf63), .C(w_mem_inst__abc_19396_new_n4653_), .Y(w_mem_inst__abc_19396_new_n4654_));
OAI21X1 OAI21X1_2425 ( .A(w_mem_inst__abc_19396_new_n4651_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf35), .C(w_mem_inst__abc_19396_new_n4654_), .Y(w_mem_inst__0w_mem_0__31_0__4_));
OAI21X1 OAI21X1_2426 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf33), .B(w_mem_inst__abc_19396_new_n4657_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf62), .Y(w_mem_inst__abc_19396_new_n4658_));
OAI21X1 OAI21X1_2427 ( .A(w_mem_inst_w_mem_1__5_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf61), .C(w_mem_inst__abc_19396_new_n4658_), .Y(w_mem_inst__abc_19396_new_n4659_));
OAI21X1 OAI21X1_2428 ( .A(w_mem_inst__abc_19396_new_n4656_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf34), .C(w_mem_inst__abc_19396_new_n4659_), .Y(w_mem_inst__0w_mem_0__31_0__5_));
OAI21X1 OAI21X1_2429 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf32), .B(w_mem_inst__abc_19396_new_n4662_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf60), .Y(w_mem_inst__abc_19396_new_n4663_));
OAI21X1 OAI21X1_243 ( .A(_abc_15497_new_n870__bF_buf1), .B(_abc_15497_new_n1853_), .C(_abc_15497_new_n1854_), .Y(_0H1_reg_31_0__11_));
OAI21X1 OAI21X1_2430 ( .A(w_mem_inst_w_mem_1__6_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf59), .C(w_mem_inst__abc_19396_new_n4663_), .Y(w_mem_inst__abc_19396_new_n4664_));
OAI21X1 OAI21X1_2431 ( .A(w_mem_inst__abc_19396_new_n4661_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf33), .C(w_mem_inst__abc_19396_new_n4664_), .Y(w_mem_inst__0w_mem_0__31_0__6_));
OAI21X1 OAI21X1_2432 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf31), .B(w_mem_inst__abc_19396_new_n4667_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf58), .Y(w_mem_inst__abc_19396_new_n4668_));
OAI21X1 OAI21X1_2433 ( .A(w_mem_inst_w_mem_1__7_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf57), .C(w_mem_inst__abc_19396_new_n4668_), .Y(w_mem_inst__abc_19396_new_n4669_));
OAI21X1 OAI21X1_2434 ( .A(w_mem_inst__abc_19396_new_n4666_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf32), .C(w_mem_inst__abc_19396_new_n4669_), .Y(w_mem_inst__0w_mem_0__31_0__7_));
OAI21X1 OAI21X1_2435 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf30), .B(w_mem_inst__abc_19396_new_n4672_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf56), .Y(w_mem_inst__abc_19396_new_n4673_));
OAI21X1 OAI21X1_2436 ( .A(w_mem_inst_w_mem_1__8_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf55), .C(w_mem_inst__abc_19396_new_n4673_), .Y(w_mem_inst__abc_19396_new_n4674_));
OAI21X1 OAI21X1_2437 ( .A(w_mem_inst__abc_19396_new_n4671_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf31), .C(w_mem_inst__abc_19396_new_n4674_), .Y(w_mem_inst__0w_mem_0__31_0__8_));
OAI21X1 OAI21X1_2438 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf29), .B(w_mem_inst__abc_19396_new_n4677_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf54), .Y(w_mem_inst__abc_19396_new_n4678_));
OAI21X1 OAI21X1_2439 ( .A(w_mem_inst_w_mem_1__9_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf53), .C(w_mem_inst__abc_19396_new_n4678_), .Y(w_mem_inst__abc_19396_new_n4679_));
OAI21X1 OAI21X1_244 ( .A(_abc_15497_new_n1838_), .B(_abc_15497_new_n1862_), .C(_abc_15497_new_n1861_), .Y(_abc_15497_new_n1863_));
OAI21X1 OAI21X1_2440 ( .A(w_mem_inst__abc_19396_new_n4676_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf30), .C(w_mem_inst__abc_19396_new_n4679_), .Y(w_mem_inst__0w_mem_0__31_0__9_));
OAI21X1 OAI21X1_2441 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf28), .B(w_mem_inst__abc_19396_new_n4682_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf52), .Y(w_mem_inst__abc_19396_new_n4683_));
OAI21X1 OAI21X1_2442 ( .A(w_mem_inst_w_mem_1__10_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf51), .C(w_mem_inst__abc_19396_new_n4683_), .Y(w_mem_inst__abc_19396_new_n4684_));
OAI21X1 OAI21X1_2443 ( .A(w_mem_inst__abc_19396_new_n4681_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf29), .C(w_mem_inst__abc_19396_new_n4684_), .Y(w_mem_inst__0w_mem_0__31_0__10_));
OAI21X1 OAI21X1_2444 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf27), .B(w_mem_inst__abc_19396_new_n4687_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf50), .Y(w_mem_inst__abc_19396_new_n4688_));
OAI21X1 OAI21X1_2445 ( .A(w_mem_inst_w_mem_1__11_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf49), .C(w_mem_inst__abc_19396_new_n4688_), .Y(w_mem_inst__abc_19396_new_n4689_));
OAI21X1 OAI21X1_2446 ( .A(w_mem_inst__abc_19396_new_n4686_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf28), .C(w_mem_inst__abc_19396_new_n4689_), .Y(w_mem_inst__0w_mem_0__31_0__11_));
OAI21X1 OAI21X1_2447 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf26), .B(w_mem_inst__abc_19396_new_n4692_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf48), .Y(w_mem_inst__abc_19396_new_n4693_));
OAI21X1 OAI21X1_2448 ( .A(w_mem_inst_w_mem_1__12_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf47), .C(w_mem_inst__abc_19396_new_n4693_), .Y(w_mem_inst__abc_19396_new_n4694_));
OAI21X1 OAI21X1_2449 ( .A(w_mem_inst__abc_19396_new_n4691_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf27), .C(w_mem_inst__abc_19396_new_n4694_), .Y(w_mem_inst__0w_mem_0__31_0__12_));
OAI21X1 OAI21X1_245 ( .A(_abc_15497_new_n1857_), .B(_abc_15497_new_n1865_), .C(_abc_15497_new_n1868_), .Y(_abc_15497_new_n1869_));
OAI21X1 OAI21X1_2450 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf25), .B(w_mem_inst__abc_19396_new_n4697_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf46), .Y(w_mem_inst__abc_19396_new_n4698_));
OAI21X1 OAI21X1_2451 ( .A(w_mem_inst_w_mem_1__13_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf45), .C(w_mem_inst__abc_19396_new_n4698_), .Y(w_mem_inst__abc_19396_new_n4699_));
OAI21X1 OAI21X1_2452 ( .A(w_mem_inst__abc_19396_new_n4696_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf26), .C(w_mem_inst__abc_19396_new_n4699_), .Y(w_mem_inst__0w_mem_0__31_0__13_));
OAI21X1 OAI21X1_2453 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf24), .B(w_mem_inst__abc_19396_new_n4702_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf44), .Y(w_mem_inst__abc_19396_new_n4703_));
OAI21X1 OAI21X1_2454 ( .A(w_mem_inst_w_mem_1__14_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf43), .C(w_mem_inst__abc_19396_new_n4703_), .Y(w_mem_inst__abc_19396_new_n4704_));
OAI21X1 OAI21X1_2455 ( .A(w_mem_inst__abc_19396_new_n4701_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf25), .C(w_mem_inst__abc_19396_new_n4704_), .Y(w_mem_inst__0w_mem_0__31_0__14_));
OAI21X1 OAI21X1_2456 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf23), .B(w_mem_inst__abc_19396_new_n4707_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf42), .Y(w_mem_inst__abc_19396_new_n4708_));
OAI21X1 OAI21X1_2457 ( .A(w_mem_inst_w_mem_1__15_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf41), .C(w_mem_inst__abc_19396_new_n4708_), .Y(w_mem_inst__abc_19396_new_n4709_));
OAI21X1 OAI21X1_2458 ( .A(w_mem_inst__abc_19396_new_n4706_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf24), .C(w_mem_inst__abc_19396_new_n4709_), .Y(w_mem_inst__0w_mem_0__31_0__15_));
OAI21X1 OAI21X1_2459 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf22), .B(w_mem_inst__abc_19396_new_n4712_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf40), .Y(w_mem_inst__abc_19396_new_n4713_));
OAI21X1 OAI21X1_246 ( .A(_auto_iopadmap_cc_368_execute_22625_109_), .B(_abc_15497_new_n883__bF_buf5), .C(_abc_15497_new_n870__bF_buf11), .Y(_abc_15497_new_n1872_));
OAI21X1 OAI21X1_2460 ( .A(w_mem_inst_w_mem_1__16_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf39), .C(w_mem_inst__abc_19396_new_n4713_), .Y(w_mem_inst__abc_19396_new_n4714_));
OAI21X1 OAI21X1_2461 ( .A(w_mem_inst__abc_19396_new_n4711_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf23), .C(w_mem_inst__abc_19396_new_n4714_), .Y(w_mem_inst__0w_mem_0__31_0__16_));
OAI21X1 OAI21X1_2462 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf21), .B(w_mem_inst__abc_19396_new_n4717_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf38), .Y(w_mem_inst__abc_19396_new_n4718_));
OAI21X1 OAI21X1_2463 ( .A(w_mem_inst_w_mem_1__17_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf37), .C(w_mem_inst__abc_19396_new_n4718_), .Y(w_mem_inst__abc_19396_new_n4719_));
OAI21X1 OAI21X1_2464 ( .A(w_mem_inst__abc_19396_new_n4716_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf22), .C(w_mem_inst__abc_19396_new_n4719_), .Y(w_mem_inst__0w_mem_0__31_0__17_));
OAI21X1 OAI21X1_2465 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf20), .B(w_mem_inst__abc_19396_new_n4722_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf36), .Y(w_mem_inst__abc_19396_new_n4723_));
OAI21X1 OAI21X1_2466 ( .A(w_mem_inst_w_mem_1__18_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf35), .C(w_mem_inst__abc_19396_new_n4723_), .Y(w_mem_inst__abc_19396_new_n4724_));
OAI21X1 OAI21X1_2467 ( .A(w_mem_inst__abc_19396_new_n4721_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf21), .C(w_mem_inst__abc_19396_new_n4724_), .Y(w_mem_inst__0w_mem_0__31_0__18_));
OAI21X1 OAI21X1_2468 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf19), .B(w_mem_inst__abc_19396_new_n4727_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf34), .Y(w_mem_inst__abc_19396_new_n4728_));
OAI21X1 OAI21X1_2469 ( .A(w_mem_inst_w_mem_1__19_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf33), .C(w_mem_inst__abc_19396_new_n4728_), .Y(w_mem_inst__abc_19396_new_n4729_));
OAI21X1 OAI21X1_247 ( .A(_abc_15497_new_n870__bF_buf10), .B(_abc_15497_new_n1871_), .C(_abc_15497_new_n1872_), .Y(_0H1_reg_31_0__13_));
OAI21X1 OAI21X1_2470 ( .A(w_mem_inst__abc_19396_new_n4726_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf20), .C(w_mem_inst__abc_19396_new_n4729_), .Y(w_mem_inst__0w_mem_0__31_0__19_));
OAI21X1 OAI21X1_2471 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf18), .B(w_mem_inst__abc_19396_new_n4732_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf32), .Y(w_mem_inst__abc_19396_new_n4733_));
OAI21X1 OAI21X1_2472 ( .A(w_mem_inst_w_mem_1__20_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf31), .C(w_mem_inst__abc_19396_new_n4733_), .Y(w_mem_inst__abc_19396_new_n4734_));
OAI21X1 OAI21X1_2473 ( .A(w_mem_inst__abc_19396_new_n4731_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf19), .C(w_mem_inst__abc_19396_new_n4734_), .Y(w_mem_inst__0w_mem_0__31_0__20_));
OAI21X1 OAI21X1_2474 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf17), .B(w_mem_inst__abc_19396_new_n4737_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf30), .Y(w_mem_inst__abc_19396_new_n4738_));
OAI21X1 OAI21X1_2475 ( .A(w_mem_inst_w_mem_1__21_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf29), .C(w_mem_inst__abc_19396_new_n4738_), .Y(w_mem_inst__abc_19396_new_n4739_));
OAI21X1 OAI21X1_2476 ( .A(w_mem_inst__abc_19396_new_n4736_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf18), .C(w_mem_inst__abc_19396_new_n4739_), .Y(w_mem_inst__0w_mem_0__31_0__21_));
OAI21X1 OAI21X1_2477 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf16), .B(w_mem_inst__abc_19396_new_n4742_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf28), .Y(w_mem_inst__abc_19396_new_n4743_));
OAI21X1 OAI21X1_2478 ( .A(w_mem_inst_w_mem_1__22_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf27), .C(w_mem_inst__abc_19396_new_n4743_), .Y(w_mem_inst__abc_19396_new_n4744_));
OAI21X1 OAI21X1_2479 ( .A(w_mem_inst__abc_19396_new_n4741_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf17), .C(w_mem_inst__abc_19396_new_n4744_), .Y(w_mem_inst__0w_mem_0__31_0__22_));
OAI21X1 OAI21X1_248 ( .A(_abc_15497_new_n1880_), .B(_abc_15497_new_n1881_), .C(_abc_15497_new_n1868_), .Y(_abc_15497_new_n1882_));
OAI21X1 OAI21X1_2480 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf15), .B(w_mem_inst__abc_19396_new_n4747_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf26), .Y(w_mem_inst__abc_19396_new_n4748_));
OAI21X1 OAI21X1_2481 ( .A(w_mem_inst_w_mem_1__23_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf25), .C(w_mem_inst__abc_19396_new_n4748_), .Y(w_mem_inst__abc_19396_new_n4749_));
OAI21X1 OAI21X1_2482 ( .A(w_mem_inst__abc_19396_new_n4746_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf16), .C(w_mem_inst__abc_19396_new_n4749_), .Y(w_mem_inst__0w_mem_0__31_0__23_));
OAI21X1 OAI21X1_2483 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf14), .B(w_mem_inst__abc_19396_new_n4752_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf24), .Y(w_mem_inst__abc_19396_new_n4753_));
OAI21X1 OAI21X1_2484 ( .A(w_mem_inst_w_mem_1__24_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf23), .C(w_mem_inst__abc_19396_new_n4753_), .Y(w_mem_inst__abc_19396_new_n4754_));
OAI21X1 OAI21X1_2485 ( .A(w_mem_inst__abc_19396_new_n4751_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf15), .C(w_mem_inst__abc_19396_new_n4754_), .Y(w_mem_inst__0w_mem_0__31_0__24_));
OAI21X1 OAI21X1_2486 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf13), .B(w_mem_inst__abc_19396_new_n4757_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf22), .Y(w_mem_inst__abc_19396_new_n4758_));
OAI21X1 OAI21X1_2487 ( .A(w_mem_inst_w_mem_1__25_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf21), .C(w_mem_inst__abc_19396_new_n4758_), .Y(w_mem_inst__abc_19396_new_n4759_));
OAI21X1 OAI21X1_2488 ( .A(w_mem_inst__abc_19396_new_n4756_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf14), .C(w_mem_inst__abc_19396_new_n4759_), .Y(w_mem_inst__0w_mem_0__31_0__25_));
OAI21X1 OAI21X1_2489 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf12), .B(w_mem_inst__abc_19396_new_n4762_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf20), .Y(w_mem_inst__abc_19396_new_n4763_));
OAI21X1 OAI21X1_249 ( .A(_auto_iopadmap_cc_368_execute_22625_109_), .B(b_reg_13_), .C(_abc_15497_new_n1882_), .Y(_abc_15497_new_n1883_));
OAI21X1 OAI21X1_2490 ( .A(w_mem_inst_w_mem_1__26_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf19), .C(w_mem_inst__abc_19396_new_n4763_), .Y(w_mem_inst__abc_19396_new_n4764_));
OAI21X1 OAI21X1_2491 ( .A(w_mem_inst__abc_19396_new_n4761_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf13), .C(w_mem_inst__abc_19396_new_n4764_), .Y(w_mem_inst__0w_mem_0__31_0__26_));
OAI21X1 OAI21X1_2492 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf11), .B(w_mem_inst__abc_19396_new_n4767_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf18), .Y(w_mem_inst__abc_19396_new_n4768_));
OAI21X1 OAI21X1_2493 ( .A(w_mem_inst_w_mem_1__27_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf17), .C(w_mem_inst__abc_19396_new_n4768_), .Y(w_mem_inst__abc_19396_new_n4769_));
OAI21X1 OAI21X1_2494 ( .A(w_mem_inst__abc_19396_new_n4766_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf12), .C(w_mem_inst__abc_19396_new_n4769_), .Y(w_mem_inst__0w_mem_0__31_0__27_));
OAI21X1 OAI21X1_2495 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf10), .B(w_mem_inst__abc_19396_new_n4772_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf16), .Y(w_mem_inst__abc_19396_new_n4773_));
OAI21X1 OAI21X1_2496 ( .A(w_mem_inst_w_mem_1__28_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf15), .C(w_mem_inst__abc_19396_new_n4773_), .Y(w_mem_inst__abc_19396_new_n4774_));
OAI21X1 OAI21X1_2497 ( .A(w_mem_inst__abc_19396_new_n4771_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf11), .C(w_mem_inst__abc_19396_new_n4774_), .Y(w_mem_inst__0w_mem_0__31_0__28_));
OAI21X1 OAI21X1_2498 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf9), .B(w_mem_inst__abc_19396_new_n4777_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf14), .Y(w_mem_inst__abc_19396_new_n4778_));
OAI21X1 OAI21X1_2499 ( .A(w_mem_inst_w_mem_1__29_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf13), .C(w_mem_inst__abc_19396_new_n4778_), .Y(w_mem_inst__abc_19396_new_n4779_));
OAI21X1 OAI21X1_25 ( .A(e_reg_0_), .B(_auto_iopadmap_cc_368_execute_22625_0_), .C(digest_update_bF_buf4), .Y(_abc_15497_new_n939_));
OAI21X1 OAI21X1_250 ( .A(_abc_15497_new_n1879_), .B(_abc_15497_new_n1886_), .C(digest_update_bF_buf4), .Y(_abc_15497_new_n1888_));
OAI21X1 OAI21X1_2500 ( .A(w_mem_inst__abc_19396_new_n4776_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf10), .C(w_mem_inst__abc_19396_new_n4779_), .Y(w_mem_inst__0w_mem_0__31_0__29_));
OAI21X1 OAI21X1_2501 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf8), .B(w_mem_inst__abc_19396_new_n4782_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf12), .Y(w_mem_inst__abc_19396_new_n4783_));
OAI21X1 OAI21X1_2502 ( .A(w_mem_inst_w_mem_1__30_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf11), .C(w_mem_inst__abc_19396_new_n4783_), .Y(w_mem_inst__abc_19396_new_n4784_));
OAI21X1 OAI21X1_2503 ( .A(w_mem_inst__abc_19396_new_n4781_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf9), .C(w_mem_inst__abc_19396_new_n4784_), .Y(w_mem_inst__0w_mem_0__31_0__30_));
OAI21X1 OAI21X1_2504 ( .A(w_mem_inst__abc_19396_new_n2420__bF_buf7), .B(w_mem_inst__abc_19396_new_n4787_), .C(w_mem_inst__abc_19396_new_n2422__bF_buf10), .Y(w_mem_inst__abc_19396_new_n4788_));
OAI21X1 OAI21X1_2505 ( .A(w_mem_inst_w_mem_1__31_), .B(w_mem_inst__abc_19396_new_n2422__bF_buf9), .C(w_mem_inst__abc_19396_new_n4788_), .Y(w_mem_inst__abc_19396_new_n4789_));
OAI21X1 OAI21X1_2506 ( .A(w_mem_inst__abc_19396_new_n4786_), .B(w_mem_inst__abc_19396_new_n2421__bF_buf8), .C(w_mem_inst__abc_19396_new_n4789_), .Y(w_mem_inst__0w_mem_0__31_0__31_));
OAI21X1 OAI21X1_2507 ( .A(w_mem_inst__abc_19396_new_n1626_), .B(w_mem_inst__abc_19396_new_n4791_), .C(w_mem_inst__abc_19396_new_n4792_), .Y(w_mem_inst__0w_ctr_reg_6_0__0_));
OAI21X1 OAI21X1_2508 ( .A(w_mem_inst__abc_19396_new_n1594__bF_buf6), .B(w_mem_inst__abc_19396_new_n1635__bF_buf2), .C(round_ctr_inc_bF_buf13), .Y(w_mem_inst__abc_19396_new_n4794_));
OAI21X1 OAI21X1_2509 ( .A(w_mem_inst__abc_19396_new_n1592_), .B(w_mem_inst__abc_19396_new_n4791_), .C(w_mem_inst__abc_19396_new_n4794_), .Y(w_mem_inst__0w_ctr_reg_6_0__1_));
OAI21X1 OAI21X1_251 ( .A(_abc_15497_new_n1879_), .B(_abc_15497_new_n1886_), .C(_abc_15497_new_n1890_), .Y(_abc_15497_new_n1891_));
OAI21X1 OAI21X1_2510 ( .A(round_ctr_inc_bF_buf12), .B(w_mem_inst__abc_19396_new_n2420__bF_buf5), .C(w_mem_inst_w_ctr_reg_2_), .Y(w_mem_inst__abc_19396_new_n4796_));
OAI21X1 OAI21X1_2511 ( .A(round_ctr_inc_bF_buf10), .B(w_mem_inst__abc_19396_new_n2420__bF_buf4), .C(w_mem_inst_w_ctr_reg_3_), .Y(w_mem_inst__abc_19396_new_n4799_));
OAI21X1 OAI21X1_2512 ( .A(w_mem_inst__abc_19396_new_n1602_), .B(w_mem_inst__abc_19396_new_n4797_), .C(w_mem_inst__abc_19396_new_n4799_), .Y(w_mem_inst__abc_19396_new_n4800_));
OAI21X1 OAI21X1_2513 ( .A(round_ctr_inc_bF_buf8), .B(w_mem_inst__abc_19396_new_n2420__bF_buf3), .C(w_mem_inst_w_ctr_reg_4_), .Y(w_mem_inst__abc_19396_new_n4803_));
OAI21X1 OAI21X1_252 ( .A(_auto_iopadmap_cc_368_execute_22625_111_), .B(_abc_15497_new_n883__bF_buf4), .C(_abc_15497_new_n870__bF_buf9), .Y(_abc_15497_new_n1897_));
OAI21X1 OAI21X1_253 ( .A(_abc_15497_new_n870__bF_buf8), .B(_abc_15497_new_n1896_), .C(_abc_15497_new_n1897_), .Y(_0H1_reg_31_0__15_));
OAI21X1 OAI21X1_254 ( .A(_abc_15497_new_n1900_), .B(_abc_15497_new_n1883_), .C(_abc_15497_new_n1899_), .Y(_abc_15497_new_n1901_));
OAI21X1 OAI21X1_255 ( .A(_abc_15497_new_n1904_), .B(_abc_15497_new_n1824_), .C(_abc_15497_new_n1903_), .Y(_abc_15497_new_n1905_));
OAI21X1 OAI21X1_256 ( .A(_auto_iopadmap_cc_368_execute_22625_112_), .B(_abc_15497_new_n883__bF_buf3), .C(_abc_15497_new_n870__bF_buf7), .Y(_abc_15497_new_n1914_));
OAI21X1 OAI21X1_257 ( .A(_abc_15497_new_n1911_), .B(_abc_15497_new_n1913_), .C(_abc_15497_new_n1914_), .Y(_0H1_reg_31_0__16_));
OAI21X1 OAI21X1_258 ( .A(_abc_15497_new_n1907_), .B(_abc_15497_new_n1908_), .C(_abc_15497_new_n1912_), .Y(_abc_15497_new_n1921_));
OAI21X1 OAI21X1_259 ( .A(_abc_15497_new_n1916_), .B(_abc_15497_new_n1918_), .C(_abc_15497_new_n1926_), .Y(_abc_15497_new_n1927_));
OAI21X1 OAI21X1_26 ( .A(_abc_15497_new_n938_), .B(_abc_15497_new_n942_), .C(_abc_15497_new_n943_), .Y(_abc_15497_new_n944_));
OAI21X1 OAI21X1_260 ( .A(_abc_15497_new_n1927_), .B(_abc_15497_new_n1925_), .C(_abc_15497_new_n1932_), .Y(_abc_15497_new_n1934_));
OAI21X1 OAI21X1_261 ( .A(_auto_iopadmap_cc_368_execute_22625_114_), .B(_abc_15497_new_n883__bF_buf2), .C(_abc_15497_new_n870__bF_buf5), .Y(_abc_15497_new_n1936_));
OAI21X1 OAI21X1_262 ( .A(_abc_15497_new_n1935_), .B(_abc_15497_new_n1933_), .C(_abc_15497_new_n1936_), .Y(_0H1_reg_31_0__18_));
OAI21X1 OAI21X1_263 ( .A(_abc_15497_new_n1945_), .B(_abc_15497_new_n1944_), .C(digest_update_bF_buf1), .Y(_abc_15497_new_n1946_));
OAI21X1 OAI21X1_264 ( .A(_auto_iopadmap_cc_368_execute_22625_115_), .B(_abc_15497_new_n883__bF_buf1), .C(_abc_15497_new_n870__bF_buf4), .Y(_abc_15497_new_n1947_));
OAI21X1 OAI21X1_265 ( .A(_abc_15497_new_n1951_), .B(_abc_15497_new_n1950_), .C(_abc_15497_new_n1952_), .Y(_abc_15497_new_n1953_));
OAI21X1 OAI21X1_266 ( .A(_abc_15497_new_n1961_), .B(_abc_15497_new_n1956_), .C(digest_update_bF_buf0), .Y(_abc_15497_new_n1963_));
OAI21X1 OAI21X1_267 ( .A(_abc_15497_new_n1957_), .B(_abc_15497_new_n1956_), .C(_abc_15497_new_n1970_), .Y(_abc_15497_new_n1971_));
OAI21X1 OAI21X1_268 ( .A(_abc_15497_new_n1976_), .B(_abc_15497_new_n1956_), .C(_abc_15497_new_n1977_), .Y(_abc_15497_new_n1978_));
OAI21X1 OAI21X1_269 ( .A(_auto_iopadmap_cc_368_execute_22625_118_), .B(_abc_15497_new_n883__bF_buf0), .C(_abc_15497_new_n870__bF_buf2), .Y(_abc_15497_new_n1984_));
OAI21X1 OAI21X1_27 ( .A(_abc_15497_new_n941_), .B(_abc_15497_new_n873__bF_buf3), .C(_abc_15497_new_n944_), .Y(_0H4_reg_31_0__1_));
OAI21X1 OAI21X1_270 ( .A(_abc_15497_new_n870__bF_buf1), .B(_abc_15497_new_n1983_), .C(_abc_15497_new_n1984_), .Y(_0H1_reg_31_0__22_));
OAI21X1 OAI21X1_271 ( .A(_auto_iopadmap_cc_368_execute_22625_119_), .B(_abc_15497_new_n883__bF_buf13), .C(_abc_15497_new_n870__bF_buf0), .Y(_abc_15497_new_n1992_));
OAI21X1 OAI21X1_272 ( .A(_abc_15497_new_n870__bF_buf11), .B(_abc_15497_new_n1991_), .C(_abc_15497_new_n1992_), .Y(_0H1_reg_31_0__23_));
OAI21X1 OAI21X1_273 ( .A(_abc_15497_new_n1994_), .B(_abc_15497_new_n1977_), .C(_abc_15497_new_n1998_), .Y(_abc_15497_new_n1999_));
OAI21X1 OAI21X1_274 ( .A(_abc_15497_new_n2009_), .B(_abc_15497_new_n2003_), .C(digest_update_bF_buf8), .Y(_abc_15497_new_n2011_));
OAI21X1 OAI21X1_275 ( .A(_auto_iopadmap_cc_368_execute_22625_120_), .B(_abc_15497_new_n883__bF_buf12), .C(_abc_15497_new_n870__bF_buf10), .Y(_abc_15497_new_n2012_));
OAI21X1 OAI21X1_276 ( .A(_abc_15497_new_n2010_), .B(_abc_15497_new_n2011_), .C(_abc_15497_new_n2012_), .Y(_0H1_reg_31_0__24_));
OAI21X1 OAI21X1_277 ( .A(_abc_15497_new_n2004_), .B(_abc_15497_new_n2003_), .C(_abc_15497_new_n2014_), .Y(_abc_15497_new_n2015_));
OAI21X1 OAI21X1_278 ( .A(_auto_iopadmap_cc_368_execute_22625_121_), .B(_abc_15497_new_n883__bF_buf11), .C(_abc_15497_new_n870__bF_buf9), .Y(_abc_15497_new_n2021_));
OAI21X1 OAI21X1_279 ( .A(_abc_15497_new_n870__bF_buf8), .B(_abc_15497_new_n2020_), .C(_abc_15497_new_n2021_), .Y(_0H1_reg_31_0__25_));
OAI21X1 OAI21X1_28 ( .A(_abc_15497_new_n947_), .B(_abc_15497_new_n941_), .C(_abc_15497_new_n948_), .Y(_abc_15497_new_n949_));
OAI21X1 OAI21X1_280 ( .A(_abc_15497_new_n2016_), .B(_abc_15497_new_n2014_), .C(_abc_15497_new_n2017_), .Y(_abc_15497_new_n2026_));
OAI21X1 OAI21X1_281 ( .A(_abc_15497_new_n2025_), .B(_abc_15497_new_n2003_), .C(_abc_15497_new_n2027_), .Y(_abc_15497_new_n2028_));
OAI21X1 OAI21X1_282 ( .A(_auto_iopadmap_cc_368_execute_22625_122_), .B(_abc_15497_new_n883__bF_buf10), .C(_abc_15497_new_n870__bF_buf7), .Y(_abc_15497_new_n2037_));
OAI21X1 OAI21X1_283 ( .A(_abc_15497_new_n2034_), .B(_abc_15497_new_n2036_), .C(_abc_15497_new_n2037_), .Y(_0H1_reg_31_0__26_));
OAI21X1 OAI21X1_284 ( .A(_abc_15497_new_n2030_), .B(_abc_15497_new_n2031_), .C(_abc_15497_new_n2035_), .Y(_abc_15497_new_n2039_));
OAI21X1 OAI21X1_285 ( .A(_auto_iopadmap_cc_368_execute_22625_123_), .B(_abc_15497_new_n883__bF_buf9), .C(_abc_15497_new_n870__bF_buf6), .Y(_abc_15497_new_n2045_));
OAI21X1 OAI21X1_286 ( .A(_abc_15497_new_n870__bF_buf5), .B(_abc_15497_new_n2044_), .C(_abc_15497_new_n2045_), .Y(_0H1_reg_31_0__27_));
OAI21X1 OAI21X1_287 ( .A(_abc_15497_new_n2040_), .B(_abc_15497_new_n2050_), .C(_abc_15497_new_n2041_), .Y(_abc_15497_new_n2051_));
OAI21X1 OAI21X1_288 ( .A(_abc_15497_new_n2049_), .B(_abc_15497_new_n2003_), .C(_abc_15497_new_n2052_), .Y(_abc_15497_new_n2053_));
OAI21X1 OAI21X1_289 ( .A(_abc_15497_new_n2059_), .B(_abc_15497_new_n2058_), .C(digest_update_bF_buf6), .Y(_abc_15497_new_n2060_));
OAI21X1 OAI21X1_29 ( .A(_abc_15497_new_n950_), .B(_abc_15497_new_n949_), .C(digest_update_bF_buf3), .Y(_abc_15497_new_n953_));
OAI21X1 OAI21X1_290 ( .A(_abc_15497_new_n2059_), .B(_abc_15497_new_n2058_), .C(_abc_15497_new_n2056_), .Y(_abc_15497_new_n2063_));
OAI21X1 OAI21X1_291 ( .A(_abc_15497_new_n2056_), .B(_abc_15497_new_n2064_), .C(_abc_15497_new_n2065_), .Y(_abc_15497_new_n2074_));
OAI21X1 OAI21X1_292 ( .A(_auto_iopadmap_cc_368_execute_22625_126_), .B(_abc_15497_new_n883__bF_buf7), .C(_abc_15497_new_n870__bF_buf2), .Y(_abc_15497_new_n2080_));
OAI21X1 OAI21X1_293 ( .A(_abc_15497_new_n870__bF_buf1), .B(_abc_15497_new_n2079_), .C(_abc_15497_new_n2080_), .Y(_0H1_reg_31_0__30_));
OAI21X1 OAI21X1_294 ( .A(_abc_15497_new_n2073_), .B(_abc_15497_new_n2076_), .C(_abc_15497_new_n2082_), .Y(_abc_15497_new_n2085_));
OAI21X1 OAI21X1_295 ( .A(_auto_iopadmap_cc_368_execute_22625_127_), .B(_abc_15497_new_n883__bF_buf6), .C(_abc_15497_new_n870__bF_buf0), .Y(_abc_15497_new_n2089_));
OAI21X1 OAI21X1_296 ( .A(_abc_15497_new_n2092_), .B(_abc_15497_new_n2093_), .C(digest_update_bF_buf4), .Y(_abc_15497_new_n2094_));
OAI21X1 OAI21X1_297 ( .A(_auto_iopadmap_cc_368_execute_22625_128_), .B(_abc_15497_new_n883__bF_buf5), .C(_abc_15497_new_n870__bF_buf11), .Y(_abc_15497_new_n2095_));
OAI21X1 OAI21X1_298 ( .A(_abc_15497_new_n2091_), .B(_abc_15497_new_n2094_), .C(_abc_15497_new_n2095_), .Y(_0H0_reg_31_0__0_));
OAI21X1 OAI21X1_299 ( .A(_abc_15497_new_n2098_), .B(_abc_15497_new_n2099_), .C(_abc_15497_new_n2100_), .Y(_abc_15497_new_n2101_));
OAI21X1 OAI21X1_3 ( .A(_abc_15497_new_n763_), .B(_abc_15497_new_n781_), .C(_abc_15497_new_n762_), .Y(_abc_15497_new_n782_));
OAI21X1 OAI21X1_30 ( .A(_abc_15497_new_n956_), .B(_abc_15497_new_n946_), .C(_abc_15497_new_n951_), .Y(_abc_15497_new_n957_));
OAI21X1 OAI21X1_300 ( .A(_abc_15497_new_n2097_), .B(_abc_15497_new_n873__bF_buf6), .C(_abc_15497_new_n2101_), .Y(_0H0_reg_31_0__1_));
OAI21X1 OAI21X1_301 ( .A(_abc_15497_new_n2097_), .B(_abc_15497_new_n2104_), .C(_abc_15497_new_n2105_), .Y(_abc_15497_new_n2106_));
OAI21X1 OAI21X1_302 ( .A(_abc_15497_new_n2107_), .B(_abc_15497_new_n2106_), .C(digest_update_bF_buf3), .Y(_abc_15497_new_n2110_));
OAI21X1 OAI21X1_303 ( .A(_abc_15497_new_n2103_), .B(_abc_15497_new_n2113_), .C(_abc_15497_new_n2108_), .Y(_abc_15497_new_n2114_));
OAI21X1 OAI21X1_304 ( .A(_abc_15497_new_n2133_), .B(_abc_15497_new_n2135_), .C(_abc_15497_new_n2132_), .Y(_abc_15497_new_n2136_));
OAI21X1 OAI21X1_305 ( .A(_abc_15497_new_n2131_), .B(_abc_15497_new_n2125_), .C(_abc_15497_new_n2137_), .Y(_abc_15497_new_n2138_));
OAI21X1 OAI21X1_306 ( .A(_abc_15497_new_n2129_), .B(_abc_15497_new_n2134_), .C(_abc_15497_new_n2138_), .Y(_abc_15497_new_n2142_));
OAI21X1 OAI21X1_307 ( .A(_abc_15497_new_n2141_), .B(_abc_15497_new_n2144_), .C(_abc_15497_new_n2148_), .Y(_abc_15497_new_n2155_));
OAI21X1 OAI21X1_308 ( .A(_abc_15497_new_n2152_), .B(_abc_15497_new_n2155_), .C(_abc_15497_new_n2156_), .Y(_abc_15497_new_n2157_));
OAI21X1 OAI21X1_309 ( .A(_abc_15497_new_n2151_), .B(_abc_15497_new_n2159_), .C(_abc_15497_new_n2160_), .Y(_abc_15497_new_n2161_));
OAI21X1 OAI21X1_31 ( .A(_abc_15497_new_n979_), .B(_abc_15497_new_n976_), .C(digest_update_bF_buf2), .Y(_abc_15497_new_n981_));
OAI21X1 OAI21X1_310 ( .A(_abc_15497_new_n2170_), .B(_abc_15497_new_n2162_), .C(digest_update_bF_buf0), .Y(_abc_15497_new_n2171_));
OAI21X1 OAI21X1_311 ( .A(_auto_iopadmap_cc_368_execute_22625_136_), .B(_abc_15497_new_n883__bF_buf4), .C(_abc_15497_new_n870__bF_buf6), .Y(_abc_15497_new_n2172_));
OAI21X1 OAI21X1_312 ( .A(_abc_15497_new_n2171_), .B(_abc_15497_new_n2169_), .C(_abc_15497_new_n2172_), .Y(_0H0_reg_31_0__8_));
OAI21X1 OAI21X1_313 ( .A(_abc_15497_new_n2164_), .B(_abc_15497_new_n2162_), .C(_abc_15497_new_n2174_), .Y(_abc_15497_new_n2175_));
OAI21X1 OAI21X1_314 ( .A(_auto_iopadmap_cc_368_execute_22625_137_), .B(_abc_15497_new_n883__bF_buf3), .C(_abc_15497_new_n870__bF_buf5), .Y(_abc_15497_new_n2178_));
OAI21X1 OAI21X1_315 ( .A(_abc_15497_new_n870__bF_buf4), .B(_abc_15497_new_n2177_), .C(_abc_15497_new_n2178_), .Y(_0H0_reg_31_0__9_));
OAI21X1 OAI21X1_316 ( .A(_abc_15497_new_n2186_), .B(_abc_15497_new_n2187_), .C(_abc_15497_new_n2174_), .Y(_abc_15497_new_n2188_));
OAI21X1 OAI21X1_317 ( .A(_auto_iopadmap_cc_368_execute_22625_137_), .B(a_reg_9_), .C(_abc_15497_new_n2188_), .Y(_abc_15497_new_n2189_));
OAI21X1 OAI21X1_318 ( .A(_abc_15497_new_n2185_), .B(_abc_15497_new_n2193_), .C(digest_update_bF_buf8), .Y(_abc_15497_new_n2195_));
OAI21X1 OAI21X1_319 ( .A(_abc_15497_new_n2181_), .B(_abc_15497_new_n2193_), .C(_abc_15497_new_n2198_), .Y(_abc_15497_new_n2199_));
OAI21X1 OAI21X1_32 ( .A(_auto_iopadmap_cc_368_execute_22625_5_), .B(_abc_15497_new_n883__bF_buf9), .C(_abc_15497_new_n870__bF_buf0), .Y(_abc_15497_new_n982_));
OAI21X1 OAI21X1_320 ( .A(_abc_15497_new_n2197_), .B(_abc_15497_new_n2207_), .C(_abc_15497_new_n2198_), .Y(_abc_15497_new_n2208_));
OAI21X1 OAI21X1_321 ( .A(_auto_iopadmap_cc_368_execute_22625_139_), .B(a_reg_11_), .C(_abc_15497_new_n2208_), .Y(_abc_15497_new_n2209_));
OAI21X1 OAI21X1_322 ( .A(_abc_15497_new_n2204_), .B(_abc_15497_new_n2189_), .C(_abc_15497_new_n2209_), .Y(_abc_15497_new_n2210_));
OAI21X1 OAI21X1_323 ( .A(_abc_15497_new_n2206_), .B(_abc_15497_new_n2162_), .C(_abc_15497_new_n2211_), .Y(_abc_15497_new_n2212_));
OAI21X1 OAI21X1_324 ( .A(_abc_15497_new_n2203_), .B(_abc_15497_new_n2214_), .C(_abc_15497_new_n2218_), .Y(_abc_15497_new_n2221_));
OAI21X1 OAI21X1_325 ( .A(_auto_iopadmap_cc_368_execute_22625_141_), .B(_abc_15497_new_n883__bF_buf2), .C(_abc_15497_new_n870__bF_buf2), .Y(_abc_15497_new_n2226_));
OAI21X1 OAI21X1_326 ( .A(_abc_15497_new_n870__bF_buf1), .B(_abc_15497_new_n2225_), .C(_abc_15497_new_n2226_), .Y(_0H0_reg_31_0__13_));
OAI21X1 OAI21X1_327 ( .A(_abc_15497_new_n2235_), .B(_abc_15497_new_n2233_), .C(_abc_15497_new_n2234_), .Y(_abc_15497_new_n2236_));
OAI21X1 OAI21X1_328 ( .A(_abc_15497_new_n2228_), .B(_abc_15497_new_n2230_), .C(_abc_15497_new_n2238_), .Y(_abc_15497_new_n2242_));
OAI21X1 OAI21X1_329 ( .A(_abc_15497_new_n2250_), .B(_abc_15497_new_n2234_), .C(_abc_15497_new_n2249_), .Y(_abc_15497_new_n2251_));
OAI21X1 OAI21X1_33 ( .A(_abc_15497_new_n980_), .B(_abc_15497_new_n981_), .C(_abc_15497_new_n982_), .Y(_0H4_reg_31_0__5_));
OAI21X1 OAI21X1_330 ( .A(_abc_15497_new_n2254_), .B(_abc_15497_new_n2162_), .C(_abc_15497_new_n2253_), .Y(_abc_15497_new_n2255_));
OAI21X1 OAI21X1_331 ( .A(_abc_15497_new_n2263_), .B(_abc_15497_new_n2262_), .C(digest_update_bF_buf5), .Y(_abc_15497_new_n2264_));
OAI21X1 OAI21X1_332 ( .A(_auto_iopadmap_cc_368_execute_22625_144_), .B(_abc_15497_new_n883__bF_buf1), .C(_abc_15497_new_n870__bF_buf11), .Y(_abc_15497_new_n2265_));
OAI21X1 OAI21X1_333 ( .A(_abc_15497_new_n2261_), .B(_abc_15497_new_n2264_), .C(_abc_15497_new_n2265_), .Y(_0H0_reg_31_0__16_));
OAI21X1 OAI21X1_334 ( .A(_abc_15497_new_n2257_), .B(_abc_15497_new_n2258_), .C(_abc_15497_new_n2273_), .Y(_abc_15497_new_n2274_));
OAI21X1 OAI21X1_335 ( .A(_abc_15497_new_n2259_), .B(_abc_15497_new_n2268_), .C(_abc_15497_new_n2272_), .Y(_abc_15497_new_n2275_));
OAI21X1 OAI21X1_336 ( .A(_abc_15497_new_n2268_), .B(_abc_15497_new_n2274_), .C(_abc_15497_new_n2275_), .Y(_abc_15497_new_n2276_));
OAI21X1 OAI21X1_337 ( .A(_abc_15497_new_n2279_), .B(_abc_15497_new_n2262_), .C(_abc_15497_new_n2280_), .Y(_abc_15497_new_n2281_));
OAI21X1 OAI21X1_338 ( .A(_abc_15497_new_n2281_), .B(_abc_15497_new_n2286_), .C(_abc_15497_new_n2288_), .Y(_abc_15497_new_n2289_));
OAI21X1 OAI21X1_339 ( .A(_abc_15497_new_n871__bF_buf4), .B(_abc_15497_new_n872__bF_buf0), .C(_abc_15497_new_n2283_), .Y(_abc_15497_new_n2290_));
OAI21X1 OAI21X1_34 ( .A(_abc_15497_new_n986_), .B(_abc_15497_new_n985_), .C(digest_update_bF_buf1), .Y(_abc_15497_new_n988_));
OAI21X1 OAI21X1_340 ( .A(digest_update_bF_buf4), .B(_abc_15497_new_n2291_), .C(_abc_15497_new_n2289_), .Y(_0H0_reg_31_0__18_));
OAI21X1 OAI21X1_341 ( .A(_abc_15497_new_n2299_), .B(_abc_15497_new_n2294_), .C(digest_update_bF_buf3), .Y(_abc_15497_new_n2301_));
OAI21X1 OAI21X1_342 ( .A(_abc_15497_new_n2304_), .B(_abc_15497_new_n2280_), .C(_abc_15497_new_n2306_), .Y(_abc_15497_new_n2307_));
OAI21X1 OAI21X1_343 ( .A(_abc_15497_new_n2313_), .B(_abc_15497_new_n2308_), .C(digest_update_bF_buf2), .Y(_abc_15497_new_n2315_));
OAI21X1 OAI21X1_344 ( .A(_abc_15497_new_n2320_), .B(_abc_15497_new_n2322_), .C(_abc_15497_new_n2319_), .Y(_abc_15497_new_n2323_));
OAI21X1 OAI21X1_345 ( .A(_abc_15497_new_n2311_), .B(_abc_15497_new_n2318_), .C(_abc_15497_new_n2324_), .Y(_abc_15497_new_n2325_));
OAI21X1 OAI21X1_346 ( .A(_abc_15497_new_n2318_), .B(_abc_15497_new_n2323_), .C(_abc_15497_new_n2325_), .Y(_abc_15497_new_n2326_));
OAI21X1 OAI21X1_347 ( .A(_auto_iopadmap_cc_368_execute_22625_150_), .B(_abc_15497_new_n883__bF_buf0), .C(_abc_15497_new_n870__bF_buf7), .Y(_abc_15497_new_n2336_));
OAI21X1 OAI21X1_348 ( .A(_abc_15497_new_n870__bF_buf6), .B(_abc_15497_new_n2335_), .C(_abc_15497_new_n2336_), .Y(_0H0_reg_31_0__22_));
OAI21X1 OAI21X1_349 ( .A(_abc_15497_new_n2339_), .B(_abc_15497_new_n2338_), .C(digest_update_bF_buf1), .Y(_abc_15497_new_n2343_));
OAI21X1 OAI21X1_35 ( .A(_auto_iopadmap_cc_368_execute_22625_6_), .B(_abc_15497_new_n883__bF_buf8), .C(_abc_15497_new_n870__bF_buf11), .Y(_abc_15497_new_n989_));
OAI21X1 OAI21X1_350 ( .A(_abc_15497_new_n2340_), .B(_abc_15497_new_n2343_), .C(_abc_15497_new_n2342_), .Y(_0H0_reg_31_0__23_));
OAI21X1 OAI21X1_351 ( .A(_abc_15497_new_n2320_), .B(_abc_15497_new_n2319_), .C(_abc_15497_new_n2328_), .Y(_abc_15497_new_n2346_));
OAI21X1 OAI21X1_352 ( .A(_auto_iopadmap_cc_368_execute_22625_151_), .B(a_reg_23_), .C(_abc_15497_new_n2333_), .Y(_abc_15497_new_n2350_));
OAI21X1 OAI21X1_353 ( .A(_abc_15497_new_n2341_), .B(_abc_15497_new_n2349_), .C(_abc_15497_new_n2350_), .Y(_abc_15497_new_n2351_));
OAI21X1 OAI21X1_354 ( .A(_abc_15497_new_n2353_), .B(_abc_15497_new_n2345_), .C(_abc_15497_new_n2352_), .Y(_abc_15497_new_n2354_));
OAI21X1 OAI21X1_355 ( .A(_abc_15497_new_n2363_), .B(_abc_15497_new_n2357_), .C(digest_update_bF_buf0), .Y(_abc_15497_new_n2365_));
OAI21X1 OAI21X1_356 ( .A(_auto_iopadmap_cc_368_execute_22625_152_), .B(_abc_15497_new_n883__bF_buf13), .C(_abc_15497_new_n870__bF_buf5), .Y(_abc_15497_new_n2366_));
OAI21X1 OAI21X1_357 ( .A(_abc_15497_new_n2364_), .B(_abc_15497_new_n2365_), .C(_abc_15497_new_n2366_), .Y(_0H0_reg_31_0__24_));
OAI21X1 OAI21X1_358 ( .A(_abc_15497_new_n2358_), .B(_abc_15497_new_n2357_), .C(_abc_15497_new_n2368_), .Y(_abc_15497_new_n2369_));
OAI21X1 OAI21X1_359 ( .A(_auto_iopadmap_cc_368_execute_22625_153_), .B(_abc_15497_new_n883__bF_buf12), .C(_abc_15497_new_n870__bF_buf4), .Y(_abc_15497_new_n2376_));
OAI21X1 OAI21X1_36 ( .A(_abc_15497_new_n987_), .B(_abc_15497_new_n988_), .C(_abc_15497_new_n989_), .Y(_0H4_reg_31_0__6_));
OAI21X1 OAI21X1_360 ( .A(_abc_15497_new_n870__bF_buf3), .B(_abc_15497_new_n2375_), .C(_abc_15497_new_n2376_), .Y(_0H0_reg_31_0__25_));
OAI21X1 OAI21X1_361 ( .A(_abc_15497_new_n2380_), .B(_abc_15497_new_n2357_), .C(_abc_15497_new_n2381_), .Y(_abc_15497_new_n2382_));
OAI21X1 OAI21X1_362 ( .A(_auto_iopadmap_cc_368_execute_22625_154_), .B(_abc_15497_new_n883__bF_buf11), .C(_abc_15497_new_n870__bF_buf2), .Y(_abc_15497_new_n2391_));
OAI21X1 OAI21X1_363 ( .A(_abc_15497_new_n2388_), .B(_abc_15497_new_n2390_), .C(_abc_15497_new_n2391_), .Y(_0H0_reg_31_0__26_));
OAI21X1 OAI21X1_364 ( .A(_abc_15497_new_n2384_), .B(_abc_15497_new_n2385_), .C(_abc_15497_new_n2389_), .Y(_abc_15497_new_n2398_));
OAI21X1 OAI21X1_365 ( .A(_abc_15497_new_n2403_), .B(_abc_15497_new_n2357_), .C(_abc_15497_new_n2407_), .Y(_abc_15497_new_n2408_));
OAI21X1 OAI21X1_366 ( .A(_abc_15497_new_n2401_), .B(_abc_15497_new_n2414_), .C(_abc_15497_new_n2411_), .Y(_abc_15497_new_n2415_));
OAI21X1 OAI21X1_367 ( .A(_abc_15497_new_n2420_), .B(_abc_15497_new_n2415_), .C(digest_update_bF_buf6), .Y(_abc_15497_new_n2422_));
OAI21X1 OAI21X1_368 ( .A(_auto_iopadmap_cc_368_execute_22625_157_), .B(_abc_15497_new_n883__bF_buf10), .C(_abc_15497_new_n870__bF_buf0), .Y(_abc_15497_new_n2423_));
OAI21X1 OAI21X1_369 ( .A(_abc_15497_new_n2421_), .B(_abc_15497_new_n2422_), .C(_abc_15497_new_n2423_), .Y(_0H0_reg_31_0__29_));
OAI21X1 OAI21X1_37 ( .A(_abc_15497_new_n1001_), .B(_abc_15497_new_n1000_), .C(digest_update_bF_buf0), .Y(_abc_15497_new_n1002_));
OAI21X1 OAI21X1_370 ( .A(_abc_15497_new_n2417_), .B(_abc_15497_new_n2418_), .C(_abc_15497_new_n2430_), .Y(_abc_15497_new_n2431_));
OAI21X1 OAI21X1_371 ( .A(_abc_15497_new_n2429_), .B(_abc_15497_new_n2433_), .C(digest_update_bF_buf5), .Y(_abc_15497_new_n2435_));
OAI21X1 OAI21X1_372 ( .A(_auto_iopadmap_cc_368_execute_22625_158_), .B(_abc_15497_new_n883__bF_buf9), .C(_abc_15497_new_n870__bF_buf11), .Y(_abc_15497_new_n2436_));
OAI21X1 OAI21X1_373 ( .A(_abc_15497_new_n2434_), .B(_abc_15497_new_n2435_), .C(_abc_15497_new_n2436_), .Y(_0H0_reg_31_0__30_));
OAI21X1 OAI21X1_374 ( .A(_abc_15497_new_n2429_), .B(_abc_15497_new_n2433_), .C(_abc_15497_new_n2428_), .Y(_abc_15497_new_n2439_));
OAI21X1 OAI21X1_375 ( .A(_abc_15497_new_n2440_), .B(_abc_15497_new_n2439_), .C(digest_update_bF_buf4), .Y(_abc_15497_new_n2442_));
OAI21X1 OAI21X1_376 ( .A(_abc_15497_new_n871__bF_buf3), .B(_abc_15497_new_n872__bF_buf4), .C(_abc_15497_new_n1751_), .Y(_abc_15497_new_n2444_));
OAI21X1 OAI21X1_377 ( .A(_abc_15497_new_n1752_), .B(_abc_15497_new_n1648__bF_buf4), .C(_abc_15497_new_n2445_), .Y(_0b_reg_31_0__0_));
OAI21X1 OAI21X1_378 ( .A(_abc_15497_new_n1763_), .B(_abc_15497_new_n1648__bF_buf3), .C(_abc_15497_new_n2448_), .Y(_0b_reg_31_0__1_));
OAI21X1 OAI21X1_379 ( .A(_abc_15497_new_n1771_), .B(_abc_15497_new_n1648__bF_buf2), .C(_abc_15497_new_n2451_), .Y(_0b_reg_31_0__2_));
OAI21X1 OAI21X1_38 ( .A(_auto_iopadmap_cc_368_execute_22625_7_), .B(_abc_15497_new_n883__bF_buf7), .C(_abc_15497_new_n870__bF_buf10), .Y(_abc_15497_new_n1003_));
OAI21X1 OAI21X1_380 ( .A(_auto_iopadmap_cc_368_execute_22625_99_), .B(_abc_15497_new_n883__bF_buf6), .C(round_ctr_rst_bF_buf7), .Y(_abc_15497_new_n2453_));
OAI21X1 OAI21X1_381 ( .A(round_ctr_inc_bF_buf7), .B(_abc_15497_new_n2453_), .C(_abc_15497_new_n2454_), .Y(_0b_reg_31_0__3_));
OAI21X1 OAI21X1_382 ( .A(_abc_15497_new_n1788_), .B(_abc_15497_new_n1648__bF_buf1), .C(_abc_15497_new_n2457_), .Y(_0b_reg_31_0__4_));
OAI21X1 OAI21X1_383 ( .A(_abc_15497_new_n1792_), .B(_abc_15497_new_n1648__bF_buf0), .C(_abc_15497_new_n2460_), .Y(_0b_reg_31_0__5_));
OAI21X1 OAI21X1_384 ( .A(_abc_15497_new_n1802_), .B(_abc_15497_new_n1648__bF_buf8), .C(_abc_15497_new_n2463_), .Y(_0b_reg_31_0__6_));
OAI21X1 OAI21X1_385 ( .A(_auto_iopadmap_cc_368_execute_22625_103_), .B(_abc_15497_new_n883__bF_buf2), .C(round_ctr_rst_bF_buf6), .Y(_abc_15497_new_n2465_));
OAI21X1 OAI21X1_386 ( .A(round_ctr_inc_bF_buf2), .B(_abc_15497_new_n2465_), .C(_abc_15497_new_n2466_), .Y(_0b_reg_31_0__7_));
OAI21X1 OAI21X1_387 ( .A(_abc_15497_new_n871__bF_buf2), .B(_abc_15497_new_n872__bF_buf3), .C(_abc_15497_new_n1819_), .Y(_abc_15497_new_n2468_));
OAI21X1 OAI21X1_388 ( .A(_abc_15497_new_n1820_), .B(_abc_15497_new_n1648__bF_buf7), .C(_abc_15497_new_n2469_), .Y(_0b_reg_31_0__8_));
OAI21X1 OAI21X1_389 ( .A(_auto_iopadmap_cc_368_execute_22625_105_), .B(_abc_15497_new_n883__bF_buf1), .C(round_ctr_rst_bF_buf5), .Y(_abc_15497_new_n2471_));
OAI21X1 OAI21X1_39 ( .A(_abc_15497_new_n978_), .B(_abc_15497_new_n1014_), .C(_abc_15497_new_n1010_), .Y(_abc_15497_new_n1015_));
OAI21X1 OAI21X1_390 ( .A(round_ctr_inc_bF_buf13), .B(_abc_15497_new_n2471_), .C(_abc_15497_new_n2472_), .Y(_0b_reg_31_0__9_));
OAI21X1 OAI21X1_391 ( .A(_abc_15497_new_n1841_), .B(_abc_15497_new_n1648__bF_buf6), .C(_abc_15497_new_n2475_), .Y(_0b_reg_31_0__10_));
OAI21X1 OAI21X1_392 ( .A(_auto_iopadmap_cc_368_execute_22625_107_), .B(_abc_15497_new_n883__bF_buf13), .C(round_ctr_rst_bF_buf4), .Y(_abc_15497_new_n2477_));
OAI21X1 OAI21X1_393 ( .A(round_ctr_inc_bF_buf10), .B(_abc_15497_new_n2477_), .C(_abc_15497_new_n2478_), .Y(_0b_reg_31_0__11_));
OAI21X1 OAI21X1_394 ( .A(_abc_15497_new_n1858_), .B(_abc_15497_new_n1648__bF_buf5), .C(_abc_15497_new_n2481_), .Y(_0b_reg_31_0__12_));
OAI21X1 OAI21X1_395 ( .A(_abc_15497_new_n871__bF_buf1), .B(_abc_15497_new_n872__bF_buf2), .C(_abc_15497_new_n1880_), .Y(_abc_15497_new_n2483_));
OAI21X1 OAI21X1_396 ( .A(_abc_15497_new_n1881_), .B(_abc_15497_new_n1648__bF_buf4), .C(_abc_15497_new_n2484_), .Y(_0b_reg_31_0__13_));
OAI21X1 OAI21X1_397 ( .A(_abc_15497_new_n1876_), .B(_abc_15497_new_n1648__bF_buf3), .C(_abc_15497_new_n2487_), .Y(_0b_reg_31_0__14_));
OAI21X1 OAI21X1_398 ( .A(_auto_iopadmap_cc_368_execute_22625_111_), .B(_abc_15497_new_n883__bF_buf10), .C(round_ctr_rst_bF_buf3), .Y(_abc_15497_new_n2489_));
OAI21X1 OAI21X1_399 ( .A(round_ctr_inc_bF_buf5), .B(_abc_15497_new_n2489_), .C(_abc_15497_new_n2490_), .Y(_0b_reg_31_0__15_));
OAI21X1 OAI21X1_4 ( .A(_abc_15497_new_n789_), .B(_abc_15497_new_n783_), .C(_abc_15497_new_n746_), .Y(_abc_15497_new_n790_));
OAI21X1 OAI21X1_40 ( .A(_abc_15497_new_n1005_), .B(_abc_15497_new_n1008_), .C(_abc_15497_new_n1017_), .Y(_abc_15497_new_n1018_));
OAI21X1 OAI21X1_400 ( .A(_abc_15497_new_n871__bF_buf0), .B(_abc_15497_new_n872__bF_buf1), .C(_abc_15497_new_n1907_), .Y(_abc_15497_new_n2492_));
OAI21X1 OAI21X1_401 ( .A(_abc_15497_new_n1908_), .B(_abc_15497_new_n1648__bF_buf2), .C(_abc_15497_new_n2493_), .Y(_0b_reg_31_0__16_));
OAI21X1 OAI21X1_402 ( .A(_abc_15497_new_n1918_), .B(_abc_15497_new_n1648__bF_buf1), .C(_abc_15497_new_n2496_), .Y(_0b_reg_31_0__17_));
OAI21X1 OAI21X1_403 ( .A(_auto_iopadmap_cc_368_execute_22625_114_), .B(_abc_15497_new_n883__bF_buf8), .C(round_ctr_rst_bF_buf2), .Y(_abc_15497_new_n2498_));
OAI21X1 OAI21X1_404 ( .A(round_ctr_inc_bF_buf1), .B(_abc_15497_new_n2498_), .C(_abc_15497_new_n2499_), .Y(_0b_reg_31_0__18_));
OAI21X1 OAI21X1_405 ( .A(_auto_iopadmap_cc_368_execute_22625_115_), .B(_abc_15497_new_n883__bF_buf7), .C(round_ctr_rst_bF_buf1), .Y(_abc_15497_new_n2501_));
OAI21X1 OAI21X1_406 ( .A(round_ctr_inc_bF_buf13), .B(_abc_15497_new_n2501_), .C(_abc_15497_new_n2502_), .Y(_0b_reg_31_0__19_));
OAI21X1 OAI21X1_407 ( .A(_abc_15497_new_n1958_), .B(_abc_15497_new_n1648__bF_buf0), .C(_abc_15497_new_n2505_), .Y(_0b_reg_31_0__20_));
OAI21X1 OAI21X1_408 ( .A(_abc_15497_new_n1967_), .B(_abc_15497_new_n1648__bF_buf8), .C(_abc_15497_new_n2508_), .Y(_0b_reg_31_0__21_));
OAI21X1 OAI21X1_409 ( .A(_auto_iopadmap_cc_368_execute_22625_118_), .B(_abc_15497_new_n883__bF_buf4), .C(round_ctr_rst_bF_buf0), .Y(_abc_15497_new_n2510_));
OAI21X1 OAI21X1_41 ( .A(_abc_15497_new_n1016_), .B(_abc_15497_new_n1012_), .C(_abc_15497_new_n1019_), .Y(_abc_15497_new_n1020_));
OAI21X1 OAI21X1_410 ( .A(round_ctr_inc_bF_buf9), .B(_abc_15497_new_n2510_), .C(_abc_15497_new_n2511_), .Y(_0b_reg_31_0__22_));
OAI21X1 OAI21X1_411 ( .A(_auto_iopadmap_cc_368_execute_22625_119_), .B(_abc_15497_new_n883__bF_buf3), .C(round_ctr_rst_bF_buf8), .Y(_abc_15497_new_n2513_));
OAI21X1 OAI21X1_412 ( .A(round_ctr_inc_bF_buf7), .B(_abc_15497_new_n2513_), .C(_abc_15497_new_n2514_), .Y(_0b_reg_31_0__23_));
OAI21X1 OAI21X1_413 ( .A(_abc_15497_new_n871__bF_buf4), .B(_abc_15497_new_n872__bF_buf0), .C(_abc_15497_new_n2005_), .Y(_abc_15497_new_n2516_));
OAI21X1 OAI21X1_414 ( .A(_abc_15497_new_n2006_), .B(_abc_15497_new_n1648__bF_buf7), .C(_abc_15497_new_n2517_), .Y(_0b_reg_31_0__24_));
OAI21X1 OAI21X1_415 ( .A(_auto_iopadmap_cc_368_execute_22625_121_), .B(_abc_15497_new_n883__bF_buf2), .C(round_ctr_rst_bF_buf7), .Y(_abc_15497_new_n2519_));
OAI21X1 OAI21X1_416 ( .A(round_ctr_inc_bF_buf4), .B(_abc_15497_new_n2519_), .C(_abc_15497_new_n2520_), .Y(_0b_reg_31_0__25_));
OAI21X1 OAI21X1_417 ( .A(_abc_15497_new_n871__bF_buf3), .B(_abc_15497_new_n872__bF_buf4), .C(_abc_15497_new_n2030_), .Y(_abc_15497_new_n2522_));
OAI21X1 OAI21X1_418 ( .A(_abc_15497_new_n2031_), .B(_abc_15497_new_n1648__bF_buf6), .C(_abc_15497_new_n2523_), .Y(_0b_reg_31_0__26_));
OAI21X1 OAI21X1_419 ( .A(_auto_iopadmap_cc_368_execute_22625_123_), .B(_abc_15497_new_n883__bF_buf1), .C(round_ctr_rst_bF_buf6), .Y(_abc_15497_new_n2525_));
OAI21X1 OAI21X1_42 ( .A(_auto_iopadmap_cc_368_execute_22625_8_), .B(_abc_15497_new_n883__bF_buf6), .C(_abc_15497_new_n870__bF_buf9), .Y(_abc_15497_new_n1022_));
OAI21X1 OAI21X1_420 ( .A(round_ctr_inc_bF_buf1), .B(_abc_15497_new_n2525_), .C(_abc_15497_new_n2526_), .Y(_0b_reg_31_0__27_));
OAI21X1 OAI21X1_421 ( .A(_abc_15497_new_n2054_), .B(_abc_15497_new_n1648__bF_buf5), .C(_abc_15497_new_n2529_), .Y(_0b_reg_31_0__28_));
OAI21X1 OAI21X1_422 ( .A(_auto_iopadmap_cc_368_execute_22625_125_), .B(_abc_15497_new_n883__bF_buf13), .C(round_ctr_rst_bF_buf5), .Y(_abc_15497_new_n2531_));
OAI21X1 OAI21X1_423 ( .A(round_ctr_inc_bF_buf12), .B(_abc_15497_new_n2531_), .C(_abc_15497_new_n2532_), .Y(_0b_reg_31_0__29_));
OAI21X1 OAI21X1_424 ( .A(_auto_iopadmap_cc_368_execute_22625_126_), .B(_abc_15497_new_n883__bF_buf12), .C(round_ctr_rst_bF_buf4), .Y(_abc_15497_new_n2534_));
OAI21X1 OAI21X1_425 ( .A(round_ctr_inc_bF_buf10), .B(_abc_15497_new_n2534_), .C(_abc_15497_new_n2535_), .Y(_0b_reg_31_0__30_));
OAI21X1 OAI21X1_426 ( .A(_auto_iopadmap_cc_368_execute_22625_127_), .B(_abc_15497_new_n883__bF_buf11), .C(round_ctr_rst_bF_buf3), .Y(_abc_15497_new_n2537_));
OAI21X1 OAI21X1_427 ( .A(round_ctr_inc_bF_buf8), .B(_abc_15497_new_n2537_), .C(_abc_15497_new_n2538_), .Y(_0b_reg_31_0__31_));
OAI21X1 OAI21X1_428 ( .A(_abc_15497_new_n1299_), .B(_abc_15497_new_n1648__bF_buf4), .C(_abc_15497_new_n2541_), .Y(_0d_reg_31_0__0_));
OAI21X1 OAI21X1_429 ( .A(_abc_15497_new_n871__bF_buf2), .B(_abc_15497_new_n872__bF_buf3), .C(_abc_15497_new_n1307_), .Y(_abc_15497_new_n2543_));
OAI21X1 OAI21X1_43 ( .A(_abc_15497_new_n870__bF_buf8), .B(_abc_15497_new_n1021_), .C(_abc_15497_new_n1022_), .Y(_0H4_reg_31_0__8_));
OAI21X1 OAI21X1_430 ( .A(_abc_15497_new_n1308_), .B(_abc_15497_new_n1648__bF_buf3), .C(_abc_15497_new_n2544_), .Y(_0d_reg_31_0__1_));
OAI21X1 OAI21X1_431 ( .A(_auto_iopadmap_cc_368_execute_22625_34_), .B(_abc_15497_new_n883__bF_buf9), .C(round_ctr_rst_bF_buf2), .Y(_abc_15497_new_n2546_));
OAI21X1 OAI21X1_432 ( .A(round_ctr_inc_bF_buf4), .B(_abc_15497_new_n2546_), .C(_abc_15497_new_n2547_), .Y(_0d_reg_31_0__2_));
OAI21X1 OAI21X1_433 ( .A(_abc_15497_new_n1320_), .B(_abc_15497_new_n1648__bF_buf2), .C(_abc_15497_new_n2550_), .Y(_0d_reg_31_0__3_));
OAI21X1 OAI21X1_434 ( .A(_abc_15497_new_n871__bF_buf1), .B(_abc_15497_new_n872__bF_buf2), .C(_abc_15497_new_n1332_), .Y(_abc_15497_new_n2552_));
OAI21X1 OAI21X1_435 ( .A(_abc_15497_new_n1333_), .B(_abc_15497_new_n1648__bF_buf1), .C(_abc_15497_new_n2553_), .Y(_0d_reg_31_0__4_));
OAI21X1 OAI21X1_436 ( .A(_abc_15497_new_n871__bF_buf0), .B(_abc_15497_new_n872__bF_buf1), .C(_abc_15497_new_n1342_), .Y(_abc_15497_new_n2555_));
OAI21X1 OAI21X1_437 ( .A(_abc_15497_new_n1343_), .B(_abc_15497_new_n1648__bF_buf0), .C(_abc_15497_new_n2556_), .Y(_0d_reg_31_0__5_));
OAI21X1 OAI21X1_438 ( .A(_abc_15497_new_n871__bF_buf4), .B(_abc_15497_new_n872__bF_buf0), .C(_abc_15497_new_n1356_), .Y(_abc_15497_new_n2558_));
OAI21X1 OAI21X1_439 ( .A(_abc_15497_new_n1357_), .B(_abc_15497_new_n1648__bF_buf8), .C(_abc_15497_new_n2559_), .Y(_0d_reg_31_0__6_));
OAI21X1 OAI21X1_44 ( .A(_abc_15497_new_n1006_), .B(_abc_15497_new_n1007_), .C(_abc_15497_new_n1020_), .Y(_abc_15497_new_n1029_));
OAI21X1 OAI21X1_440 ( .A(_abc_15497_new_n1353_), .B(_abc_15497_new_n1648__bF_buf7), .C(_abc_15497_new_n2562_), .Y(_0d_reg_31_0__7_));
OAI21X1 OAI21X1_441 ( .A(_abc_15497_new_n1364_), .B(_abc_15497_new_n1648__bF_buf6), .C(_abc_15497_new_n2565_), .Y(_0d_reg_31_0__8_));
OAI21X1 OAI21X1_442 ( .A(_abc_15497_new_n1374_), .B(_abc_15497_new_n1648__bF_buf5), .C(_abc_15497_new_n2568_), .Y(_0d_reg_31_0__9_));
OAI21X1 OAI21X1_443 ( .A(_auto_iopadmap_cc_368_execute_22625_42_), .B(_abc_15497_new_n883__bF_buf4), .C(round_ctr_rst_bF_buf1), .Y(_abc_15497_new_n2570_));
OAI21X1 OAI21X1_444 ( .A(round_ctr_inc_bF_buf9), .B(_abc_15497_new_n2570_), .C(_abc_15497_new_n2571_), .Y(_0d_reg_31_0__10_));
OAI21X1 OAI21X1_445 ( .A(_abc_15497_new_n1398_), .B(_abc_15497_new_n1648__bF_buf4), .C(_abc_15497_new_n2574_), .Y(_0d_reg_31_0__11_));
OAI21X1 OAI21X1_446 ( .A(_abc_15497_new_n871__bF_buf3), .B(_abc_15497_new_n872__bF_buf4), .C(_abc_15497_new_n1413_), .Y(_abc_15497_new_n2576_));
OAI21X1 OAI21X1_447 ( .A(_abc_15497_new_n1414_), .B(_abc_15497_new_n1648__bF_buf3), .C(_abc_15497_new_n2577_), .Y(_0d_reg_31_0__12_));
OAI21X1 OAI21X1_448 ( .A(_abc_15497_new_n1425_), .B(_abc_15497_new_n1648__bF_buf2), .C(_abc_15497_new_n2580_), .Y(_0d_reg_31_0__13_));
OAI21X1 OAI21X1_449 ( .A(_auto_iopadmap_cc_368_execute_22625_46_), .B(_abc_15497_new_n883__bF_buf1), .C(round_ctr_rst_bF_buf0), .Y(_abc_15497_new_n2582_));
OAI21X1 OAI21X1_45 ( .A(_abc_15497_new_n1025_), .B(_abc_15497_new_n1029_), .C(_abc_15497_new_n1030_), .Y(_abc_15497_new_n1031_));
OAI21X1 OAI21X1_450 ( .A(round_ctr_inc_bF_buf4), .B(_abc_15497_new_n2582_), .C(_abc_15497_new_n2583_), .Y(_0d_reg_31_0__14_));
OAI21X1 OAI21X1_451 ( .A(_abc_15497_new_n1447_), .B(_abc_15497_new_n1648__bF_buf1), .C(_abc_15497_new_n2586_), .Y(_0d_reg_31_0__15_));
OAI21X1 OAI21X1_452 ( .A(_abc_15497_new_n1462_), .B(_abc_15497_new_n1648__bF_buf0), .C(_abc_15497_new_n2589_), .Y(_0d_reg_31_0__16_));
OAI21X1 OAI21X1_453 ( .A(_auto_iopadmap_cc_368_execute_22625_49_), .B(_abc_15497_new_n883__bF_buf12), .C(round_ctr_rst_bF_buf8), .Y(_abc_15497_new_n2591_));
OAI21X1 OAI21X1_454 ( .A(round_ctr_inc_bF_buf0), .B(_abc_15497_new_n2591_), .C(_abc_15497_new_n2592_), .Y(_0d_reg_31_0__17_));
OAI21X1 OAI21X1_455 ( .A(_abc_15497_new_n1485_), .B(_abc_15497_new_n1648__bF_buf8), .C(_abc_15497_new_n2595_), .Y(_0d_reg_31_0__18_));
OAI21X1 OAI21X1_456 ( .A(_abc_15497_new_n1495_), .B(_abc_15497_new_n1648__bF_buf7), .C(_abc_15497_new_n2598_), .Y(_0d_reg_31_0__19_));
OAI21X1 OAI21X1_457 ( .A(_abc_15497_new_n871__bF_buf2), .B(_abc_15497_new_n872__bF_buf3), .C(_abc_15497_new_n1510_), .Y(_abc_15497_new_n2600_));
OAI21X1 OAI21X1_458 ( .A(_abc_15497_new_n1511_), .B(_abc_15497_new_n1648__bF_buf6), .C(_abc_15497_new_n2601_), .Y(_0d_reg_31_0__20_));
OAI21X1 OAI21X1_459 ( .A(_auto_iopadmap_cc_368_execute_22625_53_), .B(_abc_15497_new_n883__bF_buf9), .C(round_ctr_rst_bF_buf7), .Y(_abc_15497_new_n2603_));
OAI21X1 OAI21X1_46 ( .A(_abc_15497_new_n1034_), .B(_abc_15497_new_n1024_), .C(_abc_15497_new_n1035_), .Y(_abc_15497_new_n1036_));
OAI21X1 OAI21X1_460 ( .A(round_ctr_inc_bF_buf9), .B(_abc_15497_new_n2603_), .C(_abc_15497_new_n2604_), .Y(_0d_reg_31_0__21_));
OAI21X1 OAI21X1_461 ( .A(_abc_15497_new_n1530_), .B(_abc_15497_new_n1648__bF_buf5), .C(_abc_15497_new_n2607_), .Y(_0d_reg_31_0__22_));
OAI21X1 OAI21X1_462 ( .A(_abc_15497_new_n1543_), .B(_abc_15497_new_n1648__bF_buf4), .C(_abc_15497_new_n2610_), .Y(_0d_reg_31_0__23_));
OAI21X1 OAI21X1_463 ( .A(_abc_15497_new_n1562_), .B(_abc_15497_new_n1648__bF_buf3), .C(_abc_15497_new_n2613_), .Y(_0d_reg_31_0__24_));
OAI21X1 OAI21X1_464 ( .A(_abc_15497_new_n1572_), .B(_abc_15497_new_n1648__bF_buf2), .C(_abc_15497_new_n2616_), .Y(_0d_reg_31_0__25_));
OAI21X1 OAI21X1_465 ( .A(_abc_15497_new_n1586_), .B(_abc_15497_new_n1648__bF_buf1), .C(_abc_15497_new_n2619_), .Y(_0d_reg_31_0__26_));
OAI21X1 OAI21X1_466 ( .A(_abc_15497_new_n1596_), .B(_abc_15497_new_n1648__bF_buf0), .C(_abc_15497_new_n2622_), .Y(_0d_reg_31_0__27_));
OAI21X1 OAI21X1_467 ( .A(_auto_iopadmap_cc_368_execute_22625_60_), .B(_abc_15497_new_n883__bF_buf2), .C(round_ctr_rst_bF_buf6), .Y(_abc_15497_new_n2624_));
OAI21X1 OAI21X1_468 ( .A(round_ctr_inc_bF_buf1), .B(_abc_15497_new_n2624_), .C(_abc_15497_new_n2625_), .Y(_0d_reg_31_0__28_));
OAI21X1 OAI21X1_469 ( .A(_abc_15497_new_n1622_), .B(_abc_15497_new_n1648__bF_buf8), .C(_abc_15497_new_n2628_), .Y(_0d_reg_31_0__29_));
OAI21X1 OAI21X1_47 ( .A(_abc_15497_new_n1026_), .B(_abc_15497_new_n1017_), .C(_abc_15497_new_n1037_), .Y(_abc_15497_new_n1038_));
OAI21X1 OAI21X1_470 ( .A(_abc_15497_new_n2630_), .B(_abc_15497_new_n1648__bF_buf7), .C(_abc_15497_new_n2632_), .Y(_0d_reg_31_0__30_));
OAI21X1 OAI21X1_471 ( .A(_abc_15497_new_n769_), .B(_abc_15497_new_n1648__bF_buf6), .C(_abc_15497_new_n2640_), .Y(_0c_reg_31_0__0_));
OAI21X1 OAI21X1_472 ( .A(_auto_iopadmap_cc_368_execute_22625_65_), .B(_abc_15497_new_n883__bF_buf11), .C(round_ctr_rst_bF_buf5), .Y(_abc_15497_new_n2642_));
OAI21X1 OAI21X1_473 ( .A(round_ctr_inc_bF_buf9), .B(_abc_15497_new_n2642_), .C(_abc_15497_new_n2643_), .Y(_0c_reg_31_0__1_));
OAI21X1 OAI21X1_474 ( .A(_auto_iopadmap_cc_368_execute_22625_66_), .B(_abc_15497_new_n883__bF_buf10), .C(round_ctr_rst_bF_buf4), .Y(_abc_15497_new_n2645_));
OAI21X1 OAI21X1_475 ( .A(round_ctr_inc_bF_buf7), .B(_abc_15497_new_n2645_), .C(_abc_15497_new_n2646_), .Y(_0c_reg_31_0__2_));
OAI21X1 OAI21X1_476 ( .A(_auto_iopadmap_cc_368_execute_22625_67_), .B(_abc_15497_new_n883__bF_buf9), .C(round_ctr_rst_bF_buf3), .Y(_abc_15497_new_n2648_));
OAI21X1 OAI21X1_477 ( .A(round_ctr_inc_bF_buf5), .B(_abc_15497_new_n2648_), .C(_abc_15497_new_n2649_), .Y(_0c_reg_31_0__3_));
OAI21X1 OAI21X1_478 ( .A(_auto_iopadmap_cc_368_execute_22625_68_), .B(_abc_15497_new_n883__bF_buf8), .C(round_ctr_rst_bF_buf2), .Y(_abc_15497_new_n2651_));
OAI21X1 OAI21X1_479 ( .A(round_ctr_inc_bF_buf3), .B(_abc_15497_new_n2651_), .C(_abc_15497_new_n2652_), .Y(_0c_reg_31_0__4_));
OAI21X1 OAI21X1_48 ( .A(_abc_15497_new_n1036_), .B(_abc_15497_new_n1028_), .C(_abc_15497_new_n1043_), .Y(_abc_15497_new_n1045_));
OAI21X1 OAI21X1_480 ( .A(_abc_15497_new_n871__bF_buf1), .B(_abc_15497_new_n872__bF_buf2), .C(_abc_15497_new_n760_), .Y(_abc_15497_new_n2654_));
OAI21X1 OAI21X1_481 ( .A(_abc_15497_new_n759_), .B(_abc_15497_new_n1648__bF_buf5), .C(_abc_15497_new_n2655_), .Y(_0c_reg_31_0__5_));
OAI21X1 OAI21X1_482 ( .A(_abc_15497_new_n871__bF_buf0), .B(_abc_15497_new_n872__bF_buf1), .C(_abc_15497_new_n749_), .Y(_abc_15497_new_n2657_));
OAI21X1 OAI21X1_483 ( .A(_abc_15497_new_n748_), .B(_abc_15497_new_n1648__bF_buf4), .C(_abc_15497_new_n2658_), .Y(_0c_reg_31_0__6_));
OAI21X1 OAI21X1_484 ( .A(_auto_iopadmap_cc_368_execute_22625_71_), .B(_abc_15497_new_n883__bF_buf7), .C(round_ctr_rst_bF_buf1), .Y(_abc_15497_new_n2660_));
OAI21X1 OAI21X1_485 ( .A(round_ctr_inc_bF_buf13), .B(_abc_15497_new_n2660_), .C(_abc_15497_new_n2661_), .Y(_0c_reg_31_0__7_));
OAI21X1 OAI21X1_486 ( .A(_abc_15497_new_n741_), .B(_abc_15497_new_n1648__bF_buf3), .C(_abc_15497_new_n2664_), .Y(_0c_reg_31_0__8_));
OAI21X1 OAI21X1_487 ( .A(_abc_15497_new_n738_), .B(_abc_15497_new_n1648__bF_buf2), .C(_abc_15497_new_n2667_), .Y(_0c_reg_31_0__9_));
OAI21X1 OAI21X1_488 ( .A(_abc_15497_new_n871__bF_buf4), .B(_abc_15497_new_n872__bF_buf0), .C(_abc_15497_new_n728_), .Y(_abc_15497_new_n2669_));
OAI21X1 OAI21X1_489 ( .A(_abc_15497_new_n727_), .B(_abc_15497_new_n1648__bF_buf1), .C(_abc_15497_new_n2670_), .Y(_0c_reg_31_0__10_));
OAI21X1 OAI21X1_49 ( .A(_abc_15497_new_n1049_), .B(_abc_15497_new_n1033_), .C(_abc_15497_new_n1045_), .Y(_abc_15497_new_n1050_));
OAI21X1 OAI21X1_490 ( .A(_auto_iopadmap_cc_368_execute_22625_75_), .B(_abc_15497_new_n883__bF_buf4), .C(round_ctr_rst_bF_buf0), .Y(_abc_15497_new_n2672_));
OAI21X1 OAI21X1_491 ( .A(round_ctr_inc_bF_buf8), .B(_abc_15497_new_n2672_), .C(_abc_15497_new_n2673_), .Y(_0c_reg_31_0__11_));
OAI21X1 OAI21X1_492 ( .A(_auto_iopadmap_cc_368_execute_22625_76_), .B(_abc_15497_new_n883__bF_buf3), .C(round_ctr_rst_bF_buf8), .Y(_abc_15497_new_n2675_));
OAI21X1 OAI21X1_493 ( .A(round_ctr_inc_bF_buf6), .B(_abc_15497_new_n2675_), .C(_abc_15497_new_n2676_), .Y(_0c_reg_31_0__12_));
OAI21X1 OAI21X1_494 ( .A(_abc_15497_new_n708_), .B(_abc_15497_new_n1648__bF_buf0), .C(_abc_15497_new_n2679_), .Y(_0c_reg_31_0__13_));
OAI21X1 OAI21X1_495 ( .A(_abc_15497_new_n871__bF_buf3), .B(_abc_15497_new_n872__bF_buf4), .C(_abc_15497_new_n703_), .Y(_abc_15497_new_n2681_));
OAI21X1 OAI21X1_496 ( .A(_abc_15497_new_n702_), .B(_abc_15497_new_n1648__bF_buf8), .C(_abc_15497_new_n2682_), .Y(_0c_reg_31_0__14_));
OAI21X1 OAI21X1_497 ( .A(_auto_iopadmap_cc_368_execute_22625_79_), .B(_abc_15497_new_n883__bF_buf1), .C(round_ctr_rst_bF_buf7), .Y(_abc_15497_new_n2684_));
OAI21X1 OAI21X1_498 ( .A(round_ctr_inc_bF_buf2), .B(_abc_15497_new_n2684_), .C(_abc_15497_new_n2685_), .Y(_0c_reg_31_0__15_));
OAI21X1 OAI21X1_499 ( .A(_abc_15497_new_n832_), .B(_abc_15497_new_n1648__bF_buf7), .C(_abc_15497_new_n2688_), .Y(_0c_reg_31_0__16_));
OAI21X1 OAI21X1_5 ( .A(_abc_15497_new_n725_), .B(_abc_15497_new_n791_), .C(_abc_15497_new_n717_), .Y(_abc_15497_new_n792_));
OAI21X1 OAI21X1_50 ( .A(_abc_15497_new_n1040_), .B(_abc_15497_new_n1051_), .C(_abc_15497_new_n1053_), .Y(_abc_15497_new_n1060_));
OAI21X1 OAI21X1_500 ( .A(_auto_iopadmap_cc_368_execute_22625_81_), .B(_abc_15497_new_n883__bF_buf13), .C(round_ctr_rst_bF_buf6), .Y(_abc_15497_new_n2690_));
OAI21X1 OAI21X1_501 ( .A(round_ctr_inc_bF_buf13), .B(_abc_15497_new_n2690_), .C(_abc_15497_new_n2691_), .Y(_0c_reg_31_0__17_));
OAI21X1 OAI21X1_502 ( .A(_abc_15497_new_n823_), .B(_abc_15497_new_n1648__bF_buf6), .C(_abc_15497_new_n2694_), .Y(_0c_reg_31_0__18_));
OAI21X1 OAI21X1_503 ( .A(_auto_iopadmap_cc_368_execute_22625_83_), .B(_abc_15497_new_n883__bF_buf11), .C(round_ctr_rst_bF_buf5), .Y(_abc_15497_new_n2696_));
OAI21X1 OAI21X1_504 ( .A(round_ctr_inc_bF_buf10), .B(_abc_15497_new_n2696_), .C(_abc_15497_new_n2697_), .Y(_0c_reg_31_0__19_));
OAI21X1 OAI21X1_505 ( .A(_auto_iopadmap_cc_368_execute_22625_84_), .B(_abc_15497_new_n883__bF_buf10), .C(round_ctr_rst_bF_buf4), .Y(_abc_15497_new_n2699_));
OAI21X1 OAI21X1_506 ( .A(round_ctr_inc_bF_buf8), .B(_abc_15497_new_n2699_), .C(_abc_15497_new_n2700_), .Y(_0c_reg_31_0__20_));
OAI21X1 OAI21X1_507 ( .A(_auto_iopadmap_cc_368_execute_22625_85_), .B(_abc_15497_new_n883__bF_buf9), .C(round_ctr_rst_bF_buf3), .Y(_abc_15497_new_n2702_));
OAI21X1 OAI21X1_508 ( .A(round_ctr_inc_bF_buf6), .B(_abc_15497_new_n2702_), .C(_abc_15497_new_n2703_), .Y(_0c_reg_31_0__21_));
OAI21X1 OAI21X1_509 ( .A(_abc_15497_new_n798_), .B(_abc_15497_new_n1648__bF_buf5), .C(_abc_15497_new_n2706_), .Y(_0c_reg_31_0__22_));
OAI21X1 OAI21X1_51 ( .A(_abc_15497_new_n1059_), .B(_abc_15497_new_n1027_), .C(_abc_15497_new_n1061_), .Y(_abc_15497_new_n1062_));
OAI21X1 OAI21X1_510 ( .A(_auto_iopadmap_cc_368_execute_22625_87_), .B(_abc_15497_new_n883__bF_buf7), .C(round_ctr_rst_bF_buf2), .Y(_abc_15497_new_n2708_));
OAI21X1 OAI21X1_511 ( .A(round_ctr_inc_bF_buf3), .B(_abc_15497_new_n2708_), .C(_abc_15497_new_n2709_), .Y(_0c_reg_31_0__23_));
OAI21X1 OAI21X1_512 ( .A(_abc_15497_new_n855_), .B(_abc_15497_new_n1648__bF_buf4), .C(_abc_15497_new_n2712_), .Y(_0c_reg_31_0__24_));
OAI21X1 OAI21X1_513 ( .A(_abc_15497_new_n849_), .B(_abc_15497_new_n1648__bF_buf3), .C(_abc_15497_new_n2715_), .Y(_0c_reg_31_0__25_));
OAI21X1 OAI21X1_514 ( .A(_abc_15497_new_n866_), .B(_abc_15497_new_n1648__bF_buf2), .C(_abc_15497_new_n2718_), .Y(_0c_reg_31_0__26_));
OAI21X1 OAI21X1_515 ( .A(_auto_iopadmap_cc_368_execute_22625_91_), .B(_abc_15497_new_n883__bF_buf3), .C(round_ctr_rst_bF_buf1), .Y(_abc_15497_new_n2720_));
OAI21X1 OAI21X1_516 ( .A(round_ctr_inc_bF_buf12), .B(_abc_15497_new_n2720_), .C(_abc_15497_new_n2721_), .Y(_0c_reg_31_0__27_));
OAI21X1 OAI21X1_517 ( .A(_auto_iopadmap_cc_368_execute_22625_92_), .B(_abc_15497_new_n883__bF_buf2), .C(round_ctr_rst_bF_buf0), .Y(_abc_15497_new_n2723_));
OAI21X1 OAI21X1_518 ( .A(round_ctr_inc_bF_buf10), .B(_abc_15497_new_n2723_), .C(_abc_15497_new_n2724_), .Y(_0c_reg_31_0__28_));
OAI21X1 OAI21X1_519 ( .A(_abc_15497_new_n904_), .B(_abc_15497_new_n1648__bF_buf1), .C(_abc_15497_new_n2727_), .Y(_0c_reg_31_0__29_));
OAI21X1 OAI21X1_52 ( .A(_abc_15497_new_n1064_), .B(_abc_15497_new_n1057_), .C(_abc_15497_new_n1068_), .Y(_abc_15497_new_n1071_));
OAI21X1 OAI21X1_520 ( .A(_abc_15497_new_n912_), .B(_abc_15497_new_n1648__bF_buf0), .C(_abc_15497_new_n2730_), .Y(_0c_reg_31_0__30_));
OAI21X1 OAI21X1_521 ( .A(_auto_iopadmap_cc_368_execute_22625_95_), .B(_abc_15497_new_n883__bF_buf13), .C(round_ctr_rst_bF_buf8), .Y(_abc_15497_new_n2732_));
OAI21X1 OAI21X1_522 ( .A(round_ctr_inc_bF_buf6), .B(_abc_15497_new_n2732_), .C(_abc_15497_new_n2733_), .Y(_0c_reg_31_0__31_));
OAI21X1 OAI21X1_523 ( .A(round_ctr_reg_3_), .B(round_ctr_reg_2_), .C(round_ctr_reg_4_), .Y(_abc_15497_new_n2741_));
OAI21X1 OAI21X1_524 ( .A(_abc_15497_new_n1752_), .B(_abc_15497_new_n769_), .C(_abc_15497_new_n1299_), .Y(_abc_15497_new_n2744_));
OAI21X1 OAI21X1_525 ( .A(_abc_15497_new_n1752_), .B(c_reg_0_), .C(_abc_15497_new_n2744_), .Y(_abc_15497_new_n2745_));
OAI21X1 OAI21X1_526 ( .A(_abc_15497_new_n1299_), .B(_abc_15497_new_n2746_), .C(_abc_15497_new_n2748_), .Y(_abc_15497_new_n2749_));
OAI21X1 OAI21X1_527 ( .A(_abc_15497_new_n1299_), .B(_abc_15497_new_n2748_), .C(_abc_15497_new_n2749_), .Y(_abc_15497_new_n2750_));
OAI21X1 OAI21X1_528 ( .A(_abc_15497_new_n2738_), .B(_abc_15497_new_n2751_), .C(_abc_15497_new_n2755_), .Y(_abc_15497_new_n2756_));
OAI21X1 OAI21X1_529 ( .A(round_ctr_reg_4_), .B(round_ctr_reg_3_), .C(round_ctr_reg_5_), .Y(_abc_15497_new_n2758_));
OAI21X1 OAI21X1_53 ( .A(_auto_iopadmap_cc_368_execute_22625_13_), .B(_abc_15497_new_n883__bF_buf5), .C(_abc_15497_new_n870__bF_buf5), .Y(_abc_15497_new_n1077_));
OAI21X1 OAI21X1_530 ( .A(_abc_15497_new_n2739_), .B(_abc_15497_new_n2773_), .C(_abc_15497_new_n2775_), .Y(_abc_15497_new_n2776_));
OAI21X1 OAI21X1_531 ( .A(_auto_iopadmap_cc_368_execute_22625_128_), .B(_abc_15497_new_n883__bF_buf12), .C(_abc_15497_new_n1650__bF_buf7), .Y(_abc_15497_new_n2777_));
OAI21X1 OAI21X1_532 ( .A(_abc_15497_new_n2093_), .B(_abc_15497_new_n1648__bF_buf8), .C(_abc_15497_new_n2778_), .Y(_0a_reg_31_0__0_));
OAI21X1 OAI21X1_533 ( .A(_abc_15497_new_n2737_), .B(_abc_15497_new_n2753_), .C(_abc_15497_new_n2735_), .Y(_abc_15497_new_n2780_));
OAI21X1 OAI21X1_534 ( .A(_abc_15497_new_n2780__bF_buf3), .B(_abc_15497_new_n2781__bF_buf3), .C(_abc_15497_new_n2786_), .Y(_abc_15497_new_n2787_));
OAI21X1 OAI21X1_535 ( .A(b_reg_1_), .B(_abc_15497_new_n1308_), .C(_abc_15497_new_n2783_), .Y(_abc_15497_new_n2788_));
OAI21X1 OAI21X1_536 ( .A(_abc_15497_new_n2762_), .B(_abc_15497_new_n2763_), .C(_abc_15497_new_n2764_), .Y(_abc_15497_new_n2791_));
OAI21X1 OAI21X1_537 ( .A(_abc_15497_new_n2793_), .B(_abc_15497_new_n2795_), .C(_abc_15497_new_n2792_), .Y(_abc_15497_new_n2796_));
OAI21X1 OAI21X1_538 ( .A(_abc_15497_new_n2802_), .B(_abc_15497_new_n2801_), .C(_abc_15497_new_n2800_), .Y(_abc_15497_new_n2803_));
OAI21X1 OAI21X1_539 ( .A(_abc_15497_new_n2812_), .B(_abc_15497_new_n2809_), .C(_abc_15497_new_n2780__bF_buf2), .Y(_abc_15497_new_n2813_));
OAI21X1 OAI21X1_54 ( .A(_abc_15497_new_n870__bF_buf4), .B(_abc_15497_new_n1076_), .C(_abc_15497_new_n1077_), .Y(_0H4_reg_31_0__13_));
OAI21X1 OAI21X1_540 ( .A(_abc_15497_new_n2815_), .B(_abc_15497_new_n2814_), .C(_abc_15497_new_n2755_), .Y(_abc_15497_new_n2816_));
OAI21X1 OAI21X1_541 ( .A(_abc_15497_new_n2815_), .B(_abc_15497_new_n2814_), .C(_abc_15497_new_n2780__bF_buf1), .Y(_abc_15497_new_n2819_));
OAI21X1 OAI21X1_542 ( .A(_abc_15497_new_n2812_), .B(_abc_15497_new_n2809_), .C(_abc_15497_new_n2755_), .Y(_abc_15497_new_n2820_));
OAI21X1 OAI21X1_543 ( .A(_abc_15497_new_n2818_), .B(_abc_15497_new_n2822_), .C(_abc_15497_new_n2824_), .Y(_0a_reg_31_0__1_));
OAI21X1 OAI21X1_544 ( .A(_abc_15497_new_n2804_), .B(_abc_15497_new_n2806_), .C(_abc_15497_new_n2799_), .Y(_abc_15497_new_n2828_));
OAI21X1 OAI21X1_545 ( .A(_abc_15497_new_n2780__bF_buf3), .B(_abc_15497_new_n2781__bF_buf2), .C(_abc_15497_new_n2834_), .Y(_abc_15497_new_n2835_));
OAI21X1 OAI21X1_546 ( .A(b_reg_2_), .B(_abc_15497_new_n2829_), .C(_abc_15497_new_n2831_), .Y(_abc_15497_new_n2836_));
OAI21X1 OAI21X1_547 ( .A(_abc_15497_new_n2792_), .B(_abc_15497_new_n2793_), .C(_abc_15497_new_n2794_), .Y(_abc_15497_new_n2839_));
OAI21X1 OAI21X1_548 ( .A(_abc_15497_new_n2841_), .B(_abc_15497_new_n2843_), .C(_abc_15497_new_n2840_), .Y(_abc_15497_new_n2844_));
OAI21X1 OAI21X1_549 ( .A(_abc_15497_new_n2755_), .B(_abc_15497_new_n2812_), .C(_abc_15497_new_n2868_), .Y(_abc_15497_new_n2869_));
OAI21X1 OAI21X1_55 ( .A(_abc_15497_new_n1086_), .B(_abc_15497_new_n1084_), .C(_abc_15497_new_n1085_), .Y(_abc_15497_new_n1087_));
OAI21X1 OAI21X1_550 ( .A(_abc_15497_new_n2872_), .B(_abc_15497_new_n2867_), .C(_abc_15497_new_n2821_), .Y(_abc_15497_new_n2873_));
OAI21X1 OAI21X1_551 ( .A(_abc_15497_new_n2866_), .B(_abc_15497_new_n2862_), .C(_abc_15497_new_n2827_), .Y(_abc_15497_new_n2877_));
OAI21X1 OAI21X1_552 ( .A(_abc_15497_new_n1646_), .B(_abc_15497_new_n2879_), .C(_abc_15497_new_n2881_), .Y(_0a_reg_31_0__2_));
OAI21X1 OAI21X1_553 ( .A(_abc_15497_new_n2821_), .B(_abc_15497_new_n2872_), .C(_abc_15497_new_n2876_), .Y(_abc_15497_new_n2883_));
OAI21X1 OAI21X1_554 ( .A(_abc_15497_new_n2889_), .B(_abc_15497_new_n2891_), .C(_abc_15497_new_n1320_), .Y(_abc_15497_new_n2892_));
OAI21X1 OAI21X1_555 ( .A(b_reg_3_), .B(_abc_15497_new_n1320_), .C(_abc_15497_new_n2890_), .Y(_abc_15497_new_n2895_));
OAI21X1 OAI21X1_556 ( .A(_abc_15497_new_n2840_), .B(_abc_15497_new_n2841_), .C(_abc_15497_new_n2842_), .Y(_abc_15497_new_n2898_));
OAI21X1 OAI21X1_557 ( .A(_abc_15497_new_n2901_), .B(_abc_15497_new_n2908_), .C(_abc_15497_new_n2907_), .Y(_abc_15497_new_n2909_));
OAI21X1 OAI21X1_558 ( .A(_abc_15497_new_n2901_), .B(_abc_15497_new_n2908_), .C(_abc_15497_new_n2898_), .Y(_abc_15497_new_n2914_));
OAI21X1 OAI21X1_559 ( .A(_abc_15497_new_n2854_), .B(_abc_15497_new_n2853_), .C(_abc_15497_new_n2847_), .Y(_abc_15497_new_n2918_));
OAI21X1 OAI21X1_56 ( .A(_auto_iopadmap_cc_368_execute_22625_14_), .B(_abc_15497_new_n883__bF_buf4), .C(_abc_15497_new_n870__bF_buf3), .Y(_abc_15497_new_n1091_));
OAI21X1 OAI21X1_560 ( .A(_abc_15497_new_n2917_), .B(_abc_15497_new_n2921_), .C(_abc_15497_new_n2756__bF_buf2), .Y(_abc_15497_new_n2922_));
OAI21X1 OAI21X1_561 ( .A(_abc_15497_new_n2863_), .B(_abc_15497_new_n2923_), .C(_abc_15497_new_n2738_), .Y(_abc_15497_new_n2924_));
OAI21X1 OAI21X1_562 ( .A(_abc_15497_new_n2930_), .B(_abc_15497_new_n2933_), .C(_abc_15497_new_n2885_), .Y(_abc_15497_new_n2934_));
OAI21X1 OAI21X1_563 ( .A(_abc_15497_new_n1646_), .B(_abc_15497_new_n2936_), .C(_abc_15497_new_n2938_), .Y(_0a_reg_31_0__3_));
OAI21X1 OAI21X1_564 ( .A(_abc_15497_new_n2878_), .B(_abc_15497_new_n2935_), .C(_abc_15497_new_n2941_), .Y(_abc_15497_new_n2942_));
OAI21X1 OAI21X1_565 ( .A(_abc_15497_new_n2910_), .B(_abc_15497_new_n2912_), .C(_abc_15497_new_n2906_), .Y(_abc_15497_new_n2945_));
OAI21X1 OAI21X1_566 ( .A(_abc_15497_new_n1333_), .B(_abc_15497_new_n2948_), .C(_abc_15497_new_n2949_), .Y(_abc_15497_new_n2950_));
OAI21X1 OAI21X1_567 ( .A(b_reg_4_), .B(_abc_15497_new_n1333_), .C(_abc_15497_new_n2948_), .Y(_abc_15497_new_n2952_));
OAI21X1 OAI21X1_568 ( .A(_abc_15497_new_n2925__bF_buf0), .B(_abc_15497_new_n2951_), .C(_abc_15497_new_n2953_), .Y(_abc_15497_new_n2954_));
OAI21X1 OAI21X1_569 ( .A(_abc_15497_new_n2903_), .B(_abc_15497_new_n2955_), .C(_abc_15497_new_n2900_), .Y(_abc_15497_new_n2956_));
OAI21X1 OAI21X1_57 ( .A(_abc_15497_new_n1088_), .B(_abc_15497_new_n1090_), .C(_abc_15497_new_n1091_), .Y(_0H4_reg_31_0__14_));
OAI21X1 OAI21X1_570 ( .A(_abc_15497_new_n2958_), .B(_abc_15497_new_n2960_), .C(_abc_15497_new_n2957_), .Y(_abc_15497_new_n2961_));
OAI21X1 OAI21X1_571 ( .A(_abc_15497_new_n2972_), .B(_abc_15497_new_n2970_), .C(_abc_15497_new_n2945_), .Y(_abc_15497_new_n2973_));
OAI21X1 OAI21X1_572 ( .A(_abc_15497_new_n2983_), .B(_abc_15497_new_n2981_), .C(_abc_15497_new_n2975_), .Y(_abc_15497_new_n2984_));
OAI21X1 OAI21X1_573 ( .A(_abc_15497_new_n2983_), .B(_abc_15497_new_n2981_), .C(_abc_15497_new_n2945_), .Y(_abc_15497_new_n2986_));
OAI21X1 OAI21X1_574 ( .A(_abc_15497_new_n2972_), .B(_abc_15497_new_n2970_), .C(_abc_15497_new_n2975_), .Y(_abc_15497_new_n2987_));
OAI21X1 OAI21X1_575 ( .A(_abc_15497_new_n2756__bF_buf4), .B(_abc_15497_new_n2921_), .C(_abc_15497_new_n2926_), .Y(_abc_15497_new_n2990_));
OAI21X1 OAI21X1_576 ( .A(_abc_15497_new_n2997_), .B(_abc_15497_new_n2996_), .C(round_ctr_inc_bF_buf4), .Y(_abc_15497_new_n2998_));
OAI21X1 OAI21X1_577 ( .A(_abc_15497_new_n2995_), .B(_abc_15497_new_n2998_), .C(_abc_15497_new_n3000_), .Y(_0a_reg_31_0__4_));
OAI21X1 OAI21X1_578 ( .A(_abc_15497_new_n2781__bF_buf3), .B(_abc_15497_new_n3005_), .C(_abc_15497_new_n2986_), .Y(_abc_15497_new_n3006_));
OAI21X1 OAI21X1_579 ( .A(_abc_15497_new_n2982_), .B(_abc_15497_new_n2980_), .C(_abc_15497_new_n2964_), .Y(_abc_15497_new_n3007_));
OAI21X1 OAI21X1_58 ( .A(_abc_15497_new_n1080_), .B(_abc_15497_new_n1081_), .C(_abc_15497_new_n1089_), .Y(_abc_15497_new_n1093_));
OAI21X1 OAI21X1_580 ( .A(_abc_15497_new_n2780__bF_buf2), .B(_abc_15497_new_n2781__bF_buf2), .C(_abc_15497_new_n3012_), .Y(_abc_15497_new_n3013_));
OAI21X1 OAI21X1_581 ( .A(b_reg_5_), .B(_abc_15497_new_n1343_), .C(_abc_15497_new_n3009_), .Y(_abc_15497_new_n3014_));
OAI21X1 OAI21X1_582 ( .A(_abc_15497_new_n2957_), .B(_abc_15497_new_n2958_), .C(_abc_15497_new_n2959_), .Y(_abc_15497_new_n3017_));
OAI21X1 OAI21X1_583 ( .A(_abc_15497_new_n3019_), .B(_abc_15497_new_n3021_), .C(_abc_15497_new_n3018_), .Y(_abc_15497_new_n3022_));
OAI21X1 OAI21X1_584 ( .A(_abc_15497_new_n3028_), .B(_abc_15497_new_n3027_), .C(_abc_15497_new_n3026_), .Y(_abc_15497_new_n3029_));
OAI21X1 OAI21X1_585 ( .A(_abc_15497_new_n3040_), .B(_abc_15497_new_n3035_), .C(_abc_15497_new_n2944_), .Y(_abc_15497_new_n3041_));
OAI21X1 OAI21X1_586 ( .A(_abc_15497_new_n3049_), .B(_abc_15497_new_n3050_), .C(_abc_15497_new_n3048_), .Y(_abc_15497_new_n3051_));
OAI21X1 OAI21X1_587 ( .A(_abc_15497_new_n3052_), .B(_abc_15497_new_n3003_), .C(round_ctr_inc_bF_buf3), .Y(_abc_15497_new_n3054_));
OAI21X1 OAI21X1_588 ( .A(_abc_15497_new_n3053_), .B(_abc_15497_new_n3054_), .C(_abc_15497_new_n3056_), .Y(_0a_reg_31_0__5_));
OAI21X1 OAI21X1_589 ( .A(_abc_15497_new_n2993_), .B(_abc_15497_new_n3060_), .C(_abc_15497_new_n3045_), .Y(_abc_15497_new_n3061_));
OAI21X1 OAI21X1_59 ( .A(_auto_iopadmap_cc_368_execute_22625_15_), .B(_abc_15497_new_n883__bF_buf3), .C(_abc_15497_new_n870__bF_buf2), .Y(_abc_15497_new_n1099_));
OAI21X1 OAI21X1_590 ( .A(_abc_15497_new_n3033_), .B(_abc_15497_new_n3032_), .C(_abc_15497_new_n3025_), .Y(_abc_15497_new_n3065_));
OAI21X1 OAI21X1_591 ( .A(_abc_15497_new_n2780__bF_buf1), .B(_abc_15497_new_n2781__bF_buf2), .C(_abc_15497_new_n3070_), .Y(_abc_15497_new_n3071_));
OAI21X1 OAI21X1_592 ( .A(b_reg_6_), .B(_abc_15497_new_n1357_), .C(_abc_15497_new_n3067_), .Y(_abc_15497_new_n3072_));
OAI21X1 OAI21X1_593 ( .A(_abc_15497_new_n3018_), .B(_abc_15497_new_n3019_), .C(_abc_15497_new_n3020_), .Y(_abc_15497_new_n3075_));
OAI21X1 OAI21X1_594 ( .A(_abc_15497_new_n3077_), .B(_abc_15497_new_n3079_), .C(_abc_15497_new_n3076_), .Y(_abc_15497_new_n3080_));
OAI21X1 OAI21X1_595 ( .A(_abc_15497_new_n3086_), .B(_abc_15497_new_n3085_), .C(_abc_15497_new_n3084_), .Y(_abc_15497_new_n3087_));
OAI21X1 OAI21X1_596 ( .A(_abc_15497_new_n3098_), .B(_abc_15497_new_n3093_), .C(_abc_15497_new_n2739_), .Y(_abc_15497_new_n3099_));
OAI21X1 OAI21X1_597 ( .A(_abc_15497_new_n3105_), .B(_abc_15497_new_n3106_), .C(_abc_15497_new_n3104_), .Y(_abc_15497_new_n3107_));
OAI21X1 OAI21X1_598 ( .A(_abc_15497_new_n3111_), .B(_abc_15497_new_n3110_), .C(round_ctr_inc_bF_buf2), .Y(_abc_15497_new_n3112_));
OAI21X1 OAI21X1_599 ( .A(_abc_15497_new_n3109_), .B(_abc_15497_new_n3112_), .C(_abc_15497_new_n3114_), .Y(_0a_reg_31_0__6_));
OAI21X1 OAI21X1_6 ( .A(_abc_15497_new_n810_), .B(_abc_15497_new_n805_), .C(_abc_15497_new_n811_), .Y(_abc_15497_new_n812_));
OAI21X1 OAI21X1_60 ( .A(_abc_15497_new_n870__bF_buf1), .B(_abc_15497_new_n1098_), .C(_abc_15497_new_n1099_), .Y(_0H4_reg_31_0__15_));
OAI21X1 OAI21X1_600 ( .A(_abc_15497_new_n3111_), .B(_abc_15497_new_n3110_), .C(_abc_15497_new_n3116_), .Y(_abc_15497_new_n3117_));
OAI21X1 OAI21X1_601 ( .A(_abc_15497_new_n2739_), .B(_abc_15497_new_n3093_), .C(_abc_15497_new_n3101_), .Y(_abc_15497_new_n3118_));
OAI21X1 OAI21X1_602 ( .A(_abc_15497_new_n3091_), .B(_abc_15497_new_n3090_), .C(_abc_15497_new_n3083_), .Y(_abc_15497_new_n3119_));
OAI21X1 OAI21X1_603 ( .A(b_reg_7_), .B(_abc_15497_new_n1353_), .C(_abc_15497_new_n3121_), .Y(_abc_15497_new_n3126_));
OAI21X1 OAI21X1_604 ( .A(_abc_15497_new_n3076_), .B(_abc_15497_new_n3077_), .C(_abc_15497_new_n3078_), .Y(_abc_15497_new_n3130_));
OAI21X1 OAI21X1_605 ( .A(_abc_15497_new_n3132_), .B(_abc_15497_new_n3134_), .C(_abc_15497_new_n3131_), .Y(_abc_15497_new_n3135_));
OAI21X1 OAI21X1_606 ( .A(_abc_15497_new_n3141_), .B(_abc_15497_new_n3140_), .C(_abc_15497_new_n3139_), .Y(_abc_15497_new_n3142_));
OAI21X1 OAI21X1_607 ( .A(_abc_15497_new_n2780__bF_buf0), .B(_abc_15497_new_n2781__bF_buf1), .C(_abc_15497_new_n3124_), .Y(_abc_15497_new_n3145_));
OAI21X1 OAI21X1_608 ( .A(_abc_15497_new_n3141_), .B(_abc_15497_new_n3140_), .C(_abc_15497_new_n3130_), .Y(_abc_15497_new_n3149_));
OAI21X1 OAI21X1_609 ( .A(_abc_15497_new_n3151_), .B(_abc_15497_new_n3144_), .C(_abc_15497_new_n3119_), .Y(_abc_15497_new_n3152_));
OAI21X1 OAI21X1_61 ( .A(_abc_15497_new_n1103_), .B(_abc_15497_new_n1085_), .C(_abc_15497_new_n1105_), .Y(_abc_15497_new_n1106_));
OAI21X1 OAI21X1_610 ( .A(_abc_15497_new_n3156_), .B(_abc_15497_new_n3155_), .C(_abc_15497_new_n3154_), .Y(_abc_15497_new_n3157_));
OAI21X1 OAI21X1_611 ( .A(_abc_15497_new_n2159_), .B(_abc_15497_new_n1648__bF_buf7), .C(_abc_15497_new_n3165_), .Y(_0a_reg_31_0__7_));
OAI21X1 OAI21X1_612 ( .A(_abc_15497_new_n3151_), .B(_abc_15497_new_n3144_), .C(_abc_15497_new_n3154_), .Y(_abc_15497_new_n3167_));
OAI21X1 OAI21X1_613 ( .A(_abc_15497_new_n3143_), .B(_abc_15497_new_n3129_), .C(_abc_15497_new_n3138_), .Y(_abc_15497_new_n3169_));
OAI21X1 OAI21X1_614 ( .A(_abc_15497_new_n2780__bF_buf3), .B(_abc_15497_new_n2781__bF_buf0), .C(_abc_15497_new_n3174_), .Y(_abc_15497_new_n3175_));
OAI21X1 OAI21X1_615 ( .A(b_reg_8_), .B(_abc_15497_new_n1364_), .C(_abc_15497_new_n3171_), .Y(_abc_15497_new_n3176_));
OAI21X1 OAI21X1_616 ( .A(_abc_15497_new_n3131_), .B(_abc_15497_new_n3132_), .C(_abc_15497_new_n3133_), .Y(_abc_15497_new_n3178_));
OAI21X1 OAI21X1_617 ( .A(_abc_15497_new_n3180_), .B(_abc_15497_new_n3182_), .C(_abc_15497_new_n3179_), .Y(_abc_15497_new_n3183_));
OAI21X1 OAI21X1_618 ( .A(_abc_15497_new_n3134_), .B(_abc_15497_new_n3141_), .C(_abc_15497_new_n3186_), .Y(_abc_15497_new_n3188_));
OAI21X1 OAI21X1_619 ( .A(_abc_15497_new_n3194_), .B(_abc_15497_new_n3189_), .C(_abc_15497_new_n3169_), .Y(_abc_15497_new_n3195_));
OAI21X1 OAI21X1_62 ( .A(_abc_15497_new_n1109_), .B(_abc_15497_new_n1017_), .C(_abc_15497_new_n1107_), .Y(_abc_15497_new_n1110_));
OAI21X1 OAI21X1_620 ( .A(_abc_15497_new_n3194_), .B(_abc_15497_new_n3189_), .C(_abc_15497_new_n3197_), .Y(_abc_15497_new_n3205_));
OAI21X1 OAI21X1_621 ( .A(_abc_15497_new_n3209_), .B(_abc_15497_new_n3208_), .C(_abc_15497_new_n3167_), .Y(_abc_15497_new_n3210_));
OAI21X1 OAI21X1_622 ( .A(_abc_15497_new_n3116_), .B(_abc_15497_new_n3162_), .C(_abc_15497_new_n3159_), .Y(_abc_15497_new_n3215_));
OAI21X1 OAI21X1_623 ( .A(_abc_15497_new_n2996_), .B(_abc_15497_new_n3214_), .C(_abc_15497_new_n3216_), .Y(_abc_15497_new_n3217_));
OAI21X1 OAI21X1_624 ( .A(_abc_15497_new_n3211_), .B(_abc_15497_new_n3217_), .C(_abc_15497_new_n3219_), .Y(_abc_15497_new_n3220_));
OAI21X1 OAI21X1_625 ( .A(_auto_iopadmap_cc_368_execute_22625_136_), .B(_abc_15497_new_n883__bF_buf4), .C(_abc_15497_new_n1650__bF_buf9), .Y(_abc_15497_new_n3221_));
OAI21X1 OAI21X1_626 ( .A(_abc_15497_new_n2166_), .B(_abc_15497_new_n1648__bF_buf6), .C(_abc_15497_new_n3222_), .Y(_0a_reg_31_0__8_));
OAI21X1 OAI21X1_627 ( .A(_abc_15497_new_n871__bF_buf2), .B(_abc_15497_new_n872__bF_buf3), .C(_abc_15497_new_n2186_), .Y(_abc_15497_new_n3224_));
OAI21X1 OAI21X1_628 ( .A(_abc_15497_new_n2759__bF_buf0), .B(_abc_15497_new_n3228_), .C(_abc_15497_new_n3204_), .Y(_abc_15497_new_n3229_));
OAI21X1 OAI21X1_629 ( .A(_abc_15497_new_n3200_), .B(_abc_15497_new_n3199_), .C(_abc_15497_new_n3191_), .Y(_abc_15497_new_n3230_));
OAI21X1 OAI21X1_63 ( .A(_abc_15497_new_n1112_), .B(_abc_15497_new_n1101_), .C(_abc_15497_new_n1116_), .Y(_abc_15497_new_n1119_));
OAI21X1 OAI21X1_630 ( .A(d_reg_9_), .B(_abc_15497_new_n3231_), .C(_abc_15497_new_n3233_), .Y(_abc_15497_new_n3234_));
OAI21X1 OAI21X1_631 ( .A(_abc_15497_new_n3235_), .B(_abc_15497_new_n3231_), .C(_abc_15497_new_n1374_), .Y(_abc_15497_new_n3236_));
OAI21X1 OAI21X1_632 ( .A(_abc_15497_new_n3231_), .B(_abc_15497_new_n3234_), .C(_abc_15497_new_n3236_), .Y(_abc_15497_new_n3237_));
OAI21X1 OAI21X1_633 ( .A(_abc_15497_new_n3179_), .B(_abc_15497_new_n3180_), .C(_abc_15497_new_n3181_), .Y(_abc_15497_new_n3241_));
OAI21X1 OAI21X1_634 ( .A(_abc_15497_new_n3243_), .B(_abc_15497_new_n3245_), .C(_abc_15497_new_n3242_), .Y(_abc_15497_new_n3246_));
OAI21X1 OAI21X1_635 ( .A(_abc_15497_new_n3260_), .B(_abc_15497_new_n3261_), .C(_abc_15497_new_n3251_), .Y(_abc_15497_new_n3262_));
OAI21X1 OAI21X1_636 ( .A(_abc_15497_new_n3240_), .B(_abc_15497_new_n3238_), .C(_abc_15497_new_n3263_), .Y(_abc_15497_new_n3266_));
OAI21X1 OAI21X1_637 ( .A(_abc_15497_new_n3250_), .B(_abc_15497_new_n3252_), .C(_abc_15497_new_n3258_), .Y(_abc_15497_new_n3267_));
OAI21X1 OAI21X1_638 ( .A(_abc_15497_new_n3268_), .B(_abc_15497_new_n3265_), .C(_abc_15497_new_n2944_), .Y(_abc_15497_new_n3269_));
OAI21X1 OAI21X1_639 ( .A(_abc_15497_new_n3276_), .B(_abc_15497_new_n3277_), .C(_abc_15497_new_n3275_), .Y(_abc_15497_new_n3278_));
OAI21X1 OAI21X1_64 ( .A(_auto_iopadmap_cc_368_execute_22625_17_), .B(_abc_15497_new_n883__bF_buf2), .C(_abc_15497_new_n870__bF_buf0), .Y(_abc_15497_new_n1126_));
OAI21X1 OAI21X1_640 ( .A(_abc_15497_new_n2187_), .B(_abc_15497_new_n1648__bF_buf5), .C(_abc_15497_new_n3281_), .Y(_0a_reg_31_0__9_));
OAI21X1 OAI21X1_641 ( .A(_abc_15497_new_n3225_), .B(_abc_15497_new_n3283_), .C(_abc_15497_new_n3274_), .Y(_abc_15497_new_n3284_));
OAI21X1 OAI21X1_642 ( .A(_abc_15497_new_n3263_), .B(_abc_15497_new_n3258_), .C(_abc_15497_new_n3259_), .Y(_abc_15497_new_n3289_));
OAI21X1 OAI21X1_643 ( .A(_abc_15497_new_n2780__bF_buf2), .B(_abc_15497_new_n2781__bF_buf0), .C(_abc_15497_new_n3295_), .Y(_abc_15497_new_n3296_));
OAI21X1 OAI21X1_644 ( .A(b_reg_10_), .B(_abc_15497_new_n3290_), .C(_abc_15497_new_n3292_), .Y(_abc_15497_new_n3297_));
OAI21X1 OAI21X1_645 ( .A(_abc_15497_new_n3242_), .B(_abc_15497_new_n3243_), .C(_abc_15497_new_n3244_), .Y(_abc_15497_new_n3300_));
OAI21X1 OAI21X1_646 ( .A(_abc_15497_new_n3303_), .B(_abc_15497_new_n3305_), .C(_abc_15497_new_n3302_), .Y(_abc_15497_new_n3306_));
OAI21X1 OAI21X1_647 ( .A(_abc_15497_new_n3311_), .B(_abc_15497_new_n3310_), .C(_abc_15497_new_n3300_), .Y(_abc_15497_new_n3312_));
OAI21X1 OAI21X1_648 ( .A(_abc_15497_new_n3311_), .B(_abc_15497_new_n3310_), .C(_abc_15497_new_n3301_), .Y(_abc_15497_new_n3320_));
OAI21X1 OAI21X1_649 ( .A(_abc_15497_new_n3326_), .B(_abc_15497_new_n3323_), .C(_abc_15497_new_n2924__bF_buf2), .Y(_abc_15497_new_n3327_));
OAI21X1 OAI21X1_65 ( .A(_abc_15497_new_n870__bF_buf11), .B(_abc_15497_new_n1125_), .C(_abc_15497_new_n1126_), .Y(_0H4_reg_31_0__17_));
OAI21X1 OAI21X1_650 ( .A(_abc_15497_new_n3237_), .B(_abc_15497_new_n2925__bF_buf3), .C(_abc_15497_new_n3329_), .Y(_abc_15497_new_n3330_));
OAI21X1 OAI21X1_651 ( .A(_abc_15497_new_n2944_), .B(_abc_15497_new_n3265_), .C(_abc_15497_new_n3272_), .Y(_abc_15497_new_n3337_));
OAI21X1 OAI21X1_652 ( .A(_abc_15497_new_n3338_), .B(_abc_15497_new_n3339_), .C(_abc_15497_new_n3337_), .Y(_abc_15497_new_n3340_));
OAI21X1 OAI21X1_653 ( .A(_abc_15497_new_n3342_), .B(_abc_15497_new_n3287_), .C(round_ctr_inc_bF_buf13), .Y(_abc_15497_new_n3344_));
OAI21X1 OAI21X1_654 ( .A(_abc_15497_new_n3343_), .B(_abc_15497_new_n3344_), .C(_abc_15497_new_n3346_), .Y(_0a_reg_31_0__10_));
OAI21X1 OAI21X1_655 ( .A(_abc_15497_new_n3342_), .B(_abc_15497_new_n3287_), .C(_abc_15497_new_n3348_), .Y(_abc_15497_new_n3349_));
OAI21X1 OAI21X1_656 ( .A(_abc_15497_new_n2924__bF_buf0), .B(_abc_15497_new_n3323_), .C(_abc_15497_new_n3334_), .Y(_abc_15497_new_n3350_));
OAI21X1 OAI21X1_657 ( .A(_abc_15497_new_n3321_), .B(_abc_15497_new_n3318_), .C(_abc_15497_new_n3319_), .Y(_abc_15497_new_n3351_));
OAI21X1 OAI21X1_658 ( .A(_abc_15497_new_n2780__bF_buf1), .B(_abc_15497_new_n2781__bF_buf3), .C(_abc_15497_new_n3356_), .Y(_abc_15497_new_n3357_));
OAI21X1 OAI21X1_659 ( .A(b_reg_11_), .B(_abc_15497_new_n1398_), .C(_abc_15497_new_n3353_), .Y(_abc_15497_new_n3358_));
OAI21X1 OAI21X1_66 ( .A(_abc_15497_new_n1121_), .B(_abc_15497_new_n1122_), .C(_abc_15497_new_n1136_), .Y(_abc_15497_new_n1137_));
OAI21X1 OAI21X1_660 ( .A(_abc_15497_new_n3302_), .B(_abc_15497_new_n3303_), .C(_abc_15497_new_n3304_), .Y(_abc_15497_new_n3360_));
OAI21X1 OAI21X1_661 ( .A(_abc_15497_new_n3362_), .B(_abc_15497_new_n3363_), .C(_abc_15497_new_n3361_), .Y(_abc_15497_new_n3364_));
OAI21X1 OAI21X1_662 ( .A(_abc_15497_new_n3371_), .B(_abc_15497_new_n3370_), .C(_abc_15497_new_n3369_), .Y(_abc_15497_new_n3372_));
OAI21X1 OAI21X1_663 ( .A(_abc_15497_new_n3371_), .B(_abc_15497_new_n3370_), .C(_abc_15497_new_n3360_), .Y(_abc_15497_new_n3377_));
OAI21X1 OAI21X1_664 ( .A(_abc_15497_new_n3374_), .B(_abc_15497_new_n3379_), .C(_abc_15497_new_n3351_), .Y(_abc_15497_new_n3380_));
OAI21X1 OAI21X1_665 ( .A(_abc_15497_new_n3383_), .B(_abc_15497_new_n3384_), .C(_abc_15497_new_n3382_), .Y(_abc_15497_new_n3385_));
OAI21X1 OAI21X1_666 ( .A(_abc_15497_new_n3383_), .B(_abc_15497_new_n3384_), .C(_abc_15497_new_n3351_), .Y(_abc_15497_new_n3387_));
OAI21X1 OAI21X1_667 ( .A(_abc_15497_new_n3374_), .B(_abc_15497_new_n3379_), .C(_abc_15497_new_n3382_), .Y(_abc_15497_new_n3388_));
OAI21X1 OAI21X1_668 ( .A(_abc_15497_new_n3394_), .B(_abc_15497_new_n3395_), .C(_abc_15497_new_n3391_), .Y(_abc_15497_new_n3396_));
OAI21X1 OAI21X1_669 ( .A(_abc_15497_new_n3397_), .B(_abc_15497_new_n3349_), .C(round_ctr_inc_bF_buf12), .Y(_abc_15497_new_n3399_));
OAI21X1 OAI21X1_67 ( .A(_abc_15497_new_n1137_), .B(_abc_15497_new_n1134_), .C(_abc_15497_new_n1135_), .Y(_abc_15497_new_n1138_));
OAI21X1 OAI21X1_670 ( .A(_abc_15497_new_n3398_), .B(_abc_15497_new_n3399_), .C(_abc_15497_new_n3401_), .Y(_0a_reg_31_0__11_));
OAI21X1 OAI21X1_671 ( .A(_abc_15497_new_n3348_), .B(_abc_15497_new_n3404_), .C(_abc_15497_new_n3390_), .Y(_abc_15497_new_n3406_));
OAI21X1 OAI21X1_672 ( .A(_abc_15497_new_n3408_), .B(_abc_15497_new_n3403_), .C(_abc_15497_new_n3407_), .Y(_abc_15497_new_n3409_));
OAI21X1 OAI21X1_673 ( .A(_abc_15497_new_n3373_), .B(_abc_15497_new_n3414_), .C(_abc_15497_new_n3368_), .Y(_abc_15497_new_n3418_));
OAI21X1 OAI21X1_674 ( .A(_abc_15497_new_n2780__bF_buf3), .B(_abc_15497_new_n2781__bF_buf2), .C(_abc_15497_new_n3424_), .Y(_abc_15497_new_n3425_));
OAI21X1 OAI21X1_675 ( .A(b_reg_12_), .B(_abc_15497_new_n1414_), .C(_abc_15497_new_n3420_), .Y(_abc_15497_new_n3426_));
OAI21X1 OAI21X1_676 ( .A(_abc_15497_new_n3361_), .B(_abc_15497_new_n3362_), .C(_abc_15497_new_n3366_), .Y(_abc_15497_new_n3429_));
OAI21X1 OAI21X1_677 ( .A(_abc_15497_new_n3432_), .B(_abc_15497_new_n3434_), .C(_abc_15497_new_n3431_), .Y(_abc_15497_new_n3435_));
OAI21X1 OAI21X1_678 ( .A(_abc_15497_new_n3439_), .B(_abc_15497_new_n3440_), .C(_abc_15497_new_n3429_), .Y(_abc_15497_new_n3441_));
OAI21X1 OAI21X1_679 ( .A(b_reg_12_), .B(c_reg_12_), .C(_abc_15497_new_n3444_), .Y(_abc_15497_new_n3445_));
OAI21X1 OAI21X1_68 ( .A(_abc_15497_new_n1133_), .B(_abc_15497_new_n1138_), .C(digest_update_bF_buf4), .Y(_abc_15497_new_n1140_));
OAI21X1 OAI21X1_680 ( .A(_abc_15497_new_n3439_), .B(_abc_15497_new_n3440_), .C(_abc_15497_new_n3430_), .Y(_abc_15497_new_n3450_));
OAI21X1 OAI21X1_681 ( .A(_abc_15497_new_n3458_), .B(_abc_15497_new_n3453_), .C(_abc_15497_new_n2925__bF_buf2), .Y(_abc_15497_new_n3459_));
OAI21X1 OAI21X1_682 ( .A(_abc_15497_new_n2780__bF_buf2), .B(_abc_15497_new_n3466_), .C(_abc_15497_new_n3387_), .Y(_abc_15497_new_n3467_));
OAI21X1 OAI21X1_683 ( .A(_abc_15497_new_n3458_), .B(_abc_15497_new_n3453_), .C(_abc_15497_new_n2756__bF_buf2), .Y(_abc_15497_new_n3469_));
OAI21X1 OAI21X1_684 ( .A(_abc_15497_new_n3472_), .B(_abc_15497_new_n3474_), .C(_abc_15497_new_n3476_), .Y(_0a_reg_31_0__12_));
OAI21X1 OAI21X1_685 ( .A(_abc_15497_new_n2756__bF_buf1), .B(_abc_15497_new_n3453_), .C(_abc_15497_new_n3461_), .Y(_abc_15497_new_n3479_));
OAI21X1 OAI21X1_686 ( .A(_abc_15497_new_n3451_), .B(_abc_15497_new_n3448_), .C(_abc_15497_new_n3449_), .Y(_abc_15497_new_n3480_));
OAI21X1 OAI21X1_687 ( .A(_abc_15497_new_n3481_), .B(_abc_15497_new_n3482_), .C(_abc_15497_new_n1425_), .Y(_abc_15497_new_n3483_));
OAI21X1 OAI21X1_688 ( .A(d_reg_13_), .B(_abc_15497_new_n3482_), .C(_abc_15497_new_n3484_), .Y(_abc_15497_new_n3489_));
OAI21X1 OAI21X1_689 ( .A(b_reg_13_), .B(_abc_15497_new_n1425_), .C(_abc_15497_new_n3485_), .Y(_abc_15497_new_n3490_));
OAI21X1 OAI21X1_69 ( .A(_abc_15497_new_n1129_), .B(_abc_15497_new_n1138_), .C(_abc_15497_new_n1143_), .Y(_abc_15497_new_n1144_));
OAI21X1 OAI21X1_690 ( .A(_abc_15497_new_n3431_), .B(_abc_15497_new_n3432_), .C(_abc_15497_new_n3433_), .Y(_abc_15497_new_n3493_));
OAI21X1 OAI21X1_691 ( .A(_abc_15497_new_n3495_), .B(_abc_15497_new_n3496_), .C(_abc_15497_new_n3494_), .Y(_abc_15497_new_n3497_));
OAI21X1 OAI21X1_692 ( .A(_abc_15497_new_n3488_), .B(_abc_15497_new_n3492_), .C(_abc_15497_new_n3510_), .Y(_abc_15497_new_n3513_));
OAI21X1 OAI21X1_693 ( .A(_abc_15497_new_n3502_), .B(_abc_15497_new_n3504_), .C(_abc_15497_new_n3507_), .Y(_abc_15497_new_n3514_));
OAI21X1 OAI21X1_694 ( .A(_abc_15497_new_n3515_), .B(_abc_15497_new_n3512_), .C(_abc_15497_new_n2780__bF_buf1), .Y(_abc_15497_new_n3516_));
OAI21X1 OAI21X1_695 ( .A(_abc_15497_new_n3524_), .B(_abc_15497_new_n3525_), .C(_abc_15497_new_n3523_), .Y(_abc_15497_new_n3526_));
OAI21X1 OAI21X1_696 ( .A(_abc_15497_new_n3528_), .B(_abc_15497_new_n3478_), .C(round_ctr_inc_bF_buf10), .Y(_abc_15497_new_n3529_));
OAI21X1 OAI21X1_697 ( .A(_auto_iopadmap_cc_368_execute_22625_141_), .B(_abc_15497_new_n883__bF_buf0), .C(_abc_15497_new_n1650__bF_buf4), .Y(_abc_15497_new_n3532_));
OAI21X1 OAI21X1_698 ( .A(_abc_15497_new_n3531_), .B(_abc_15497_new_n1648__bF_buf4), .C(_abc_15497_new_n3532_), .Y(_abc_15497_new_n3533_));
OAI21X1 OAI21X1_699 ( .A(_abc_15497_new_n3510_), .B(_abc_15497_new_n3507_), .C(_abc_15497_new_n3508_), .Y(_abc_15497_new_n3542_));
OAI21X1 OAI21X1_7 ( .A(_abc_15497_new_n835_), .B(_abc_15497_new_n828_), .C(_abc_15497_new_n836_), .Y(_abc_15497_new_n837_));
OAI21X1 OAI21X1_70 ( .A(e_reg_17_), .B(_auto_iopadmap_cc_368_execute_22625_17_), .C(_abc_15497_new_n1137_), .Y(_abc_15497_new_n1151_));
OAI21X1 OAI21X1_700 ( .A(_abc_15497_new_n3544_), .B(_abc_15497_new_n3545_), .C(_abc_15497_new_n3543_), .Y(_abc_15497_new_n3546_));
OAI21X1 OAI21X1_701 ( .A(b_reg_14_), .B(_abc_15497_new_n3543_), .C(_abc_15497_new_n3548_), .Y(_abc_15497_new_n3554_));
OAI21X1 OAI21X1_702 ( .A(_abc_15497_new_n3494_), .B(_abc_15497_new_n3495_), .C(_abc_15497_new_n3499_), .Y(_abc_15497_new_n3557_));
OAI21X1 OAI21X1_703 ( .A(_abc_15497_new_n3560_), .B(_abc_15497_new_n3561_), .C(_abc_15497_new_n3559_), .Y(_abc_15497_new_n3562_));
OAI21X1 OAI21X1_704 ( .A(_abc_15497_new_n3568_), .B(_abc_15497_new_n3567_), .C(_abc_15497_new_n3557_), .Y(_abc_15497_new_n3569_));
OAI21X1 OAI21X1_705 ( .A(_abc_15497_new_n3551_), .B(_abc_15497_new_n3556_), .C(_abc_15497_new_n3570_), .Y(_abc_15497_new_n3571_));
OAI21X1 OAI21X1_706 ( .A(_abc_15497_new_n3568_), .B(_abc_15497_new_n3567_), .C(_abc_15497_new_n3558_), .Y(_abc_15497_new_n3575_));
OAI21X1 OAI21X1_707 ( .A(_abc_15497_new_n3551_), .B(_abc_15497_new_n3556_), .C(_abc_15497_new_n3576_), .Y(_abc_15497_new_n3579_));
OAI21X1 OAI21X1_708 ( .A(_abc_15497_new_n3581_), .B(_abc_15497_new_n3578_), .C(_abc_15497_new_n2759__bF_buf4), .Y(_abc_15497_new_n3582_));
OAI21X1 OAI21X1_709 ( .A(_abc_15497_new_n3487_), .B(_abc_15497_new_n2925__bF_buf3), .C(_abc_15497_new_n3584_), .Y(_abc_15497_new_n3585_));
OAI21X1 OAI21X1_71 ( .A(_abc_15497_new_n1153_), .B(_abc_15497_new_n1151_), .C(_abc_15497_new_n1152_), .Y(_abc_15497_new_n1154_));
OAI21X1 OAI21X1_710 ( .A(_abc_15497_new_n2780__bF_buf3), .B(_abc_15497_new_n3512_), .C(_abc_15497_new_n3520_), .Y(_abc_15497_new_n3592_));
OAI21X1 OAI21X1_711 ( .A(_abc_15497_new_n3593_), .B(_abc_15497_new_n3594_), .C(_abc_15497_new_n3592_), .Y(_abc_15497_new_n3595_));
OAI21X1 OAI21X1_712 ( .A(_abc_15497_new_n3597_), .B(_abc_15497_new_n3599_), .C(_abc_15497_new_n3601_), .Y(_0a_reg_31_0__14_));
OAI21X1 OAI21X1_713 ( .A(_abc_15497_new_n2759__bF_buf1), .B(_abc_15497_new_n3578_), .C(_abc_15497_new_n3589_), .Y(_abc_15497_new_n3605_));
OAI21X1 OAI21X1_714 ( .A(_abc_15497_new_n3576_), .B(_abc_15497_new_n3573_), .C(_abc_15497_new_n3574_), .Y(_abc_15497_new_n3606_));
OAI21X1 OAI21X1_715 ( .A(d_reg_15_), .B(_abc_15497_new_n3607_), .C(_abc_15497_new_n3610_), .Y(_abc_15497_new_n3611_));
OAI21X1 OAI21X1_716 ( .A(_abc_15497_new_n3612_), .B(_abc_15497_new_n3607_), .C(_abc_15497_new_n1447_), .Y(_abc_15497_new_n3613_));
OAI21X1 OAI21X1_717 ( .A(_abc_15497_new_n3607_), .B(_abc_15497_new_n3611_), .C(_abc_15497_new_n3613_), .Y(_abc_15497_new_n3614_));
OAI21X1 OAI21X1_718 ( .A(b_reg_15_), .B(_abc_15497_new_n1447_), .C(_abc_15497_new_n3616_), .Y(_abc_15497_new_n3617_));
OAI21X1 OAI21X1_719 ( .A(_abc_15497_new_n2924__bF_buf3), .B(_abc_15497_new_n3611_), .C(_abc_15497_new_n3618_), .Y(_abc_15497_new_n3619_));
OAI21X1 OAI21X1_72 ( .A(_abc_15497_new_n1154_), .B(_abc_15497_new_n1158_), .C(_abc_15497_new_n1165_), .Y(_abc_15497_new_n1167_));
OAI21X1 OAI21X1_720 ( .A(_abc_15497_new_n3559_), .B(_abc_15497_new_n3560_), .C(_abc_15497_new_n3564_), .Y(_abc_15497_new_n3620_));
OAI21X1 OAI21X1_721 ( .A(_abc_15497_new_n3623_), .B(_abc_15497_new_n3625_), .C(_abc_15497_new_n3622_), .Y(_abc_15497_new_n3626_));
OAI21X1 OAI21X1_722 ( .A(_abc_15497_new_n3630_), .B(_abc_15497_new_n3631_), .C(_abc_15497_new_n3620_), .Y(_abc_15497_new_n3632_));
OAI21X1 OAI21X1_723 ( .A(_abc_15497_new_n3619_), .B(_abc_15497_new_n3615_), .C(_abc_15497_new_n3633_), .Y(_abc_15497_new_n3634_));
OAI21X1 OAI21X1_724 ( .A(_abc_15497_new_n3608_), .B(_abc_15497_new_n3609_), .C(_abc_15497_new_n3635_), .Y(_abc_15497_new_n3636_));
OAI21X1 OAI21X1_725 ( .A(_abc_15497_new_n3630_), .B(_abc_15497_new_n3631_), .C(_abc_15497_new_n3621_), .Y(_abc_15497_new_n3640_));
OAI21X1 OAI21X1_726 ( .A(_abc_15497_new_n3619_), .B(_abc_15497_new_n3615_), .C(_abc_15497_new_n3641_), .Y(_abc_15497_new_n3644_));
OAI21X1 OAI21X1_727 ( .A(_abc_15497_new_n3646_), .B(_abc_15497_new_n3643_), .C(_abc_15497_new_n2743__bF_buf0), .Y(_abc_15497_new_n3647_));
OAI21X1 OAI21X1_728 ( .A(_abc_15497_new_n3550_), .B(_abc_15497_new_n2925__bF_buf1), .C(_abc_15497_new_n3648_), .Y(_abc_15497_new_n3649_));
OAI21X1 OAI21X1_729 ( .A(_abc_15497_new_n3657_), .B(_abc_15497_new_n3658_), .C(_abc_15497_new_n3656_), .Y(_abc_15497_new_n3659_));
OAI21X1 OAI21X1_73 ( .A(_auto_iopadmap_cc_368_execute_22625_20_), .B(_abc_15497_new_n883__bF_buf1), .C(_abc_15497_new_n870__bF_buf9), .Y(_abc_15497_new_n1169_));
OAI21X1 OAI21X1_730 ( .A(_abc_15497_new_n3541_), .B(_abc_15497_new_n3603_), .C(_abc_15497_new_n3598_), .Y(_abc_15497_new_n3662_));
OAI21X1 OAI21X1_731 ( .A(_abc_15497_new_n3663_), .B(_abc_15497_new_n3662_), .C(round_ctr_inc_bF_buf8), .Y(_abc_15497_new_n3664_));
OAI21X1 OAI21X1_732 ( .A(_abc_15497_new_n3661_), .B(_abc_15497_new_n3664_), .C(_abc_15497_new_n3666_), .Y(_0a_reg_31_0__15_));
OAI21X1 OAI21X1_733 ( .A(_abc_15497_new_n3604_), .B(_abc_15497_new_n3660_), .C(_abc_15497_new_n3655_), .Y(_abc_15497_new_n3671_));
OAI21X1 OAI21X1_734 ( .A(_abc_15497_new_n3669_), .B(_abc_15497_new_n3407_), .C(_abc_15497_new_n3672_), .Y(_abc_15497_new_n3673_));
OAI21X1 OAI21X1_735 ( .A(_abc_15497_new_n2738_), .B(_abc_15497_new_n2751_), .C(_abc_15497_new_n2924__bF_buf1), .Y(_abc_15497_new_n3678_));
OAI21X1 OAI21X1_736 ( .A(_abc_15497_new_n3683_), .B(_abc_15497_new_n3684_), .C(_abc_15497_new_n2756__bF_buf2), .Y(_abc_15497_new_n3685_));
OAI21X1 OAI21X1_737 ( .A(d_reg_16_), .B(b_reg_16_), .C(c_reg_16_), .Y(_abc_15497_new_n3686_));
OAI21X1 OAI21X1_738 ( .A(_abc_15497_new_n1462_), .B(b_reg_16_), .C(_abc_15497_new_n3686_), .Y(_abc_15497_new_n3687_));
OAI21X1 OAI21X1_739 ( .A(_abc_15497_new_n1462_), .B(_abc_15497_new_n1908_), .C(_abc_15497_new_n3686_), .Y(_abc_15497_new_n3688_));
OAI21X1 OAI21X1_74 ( .A(_abc_15497_new_n1168_), .B(_abc_15497_new_n1166_), .C(_abc_15497_new_n1169_), .Y(_0H4_reg_31_0__20_));
OAI21X1 OAI21X1_740 ( .A(_abc_15497_new_n3622_), .B(_abc_15497_new_n3623_), .C(_abc_15497_new_n3624_), .Y(_abc_15497_new_n3691_));
OAI21X1 OAI21X1_741 ( .A(_abc_15497_new_n3707_), .B(_abc_15497_new_n3708_), .C(_abc_15497_new_n3678_), .Y(_abc_15497_new_n3709_));
OAI21X1 OAI21X1_742 ( .A(_abc_15497_new_n3676_), .B(_abc_15497_new_n3713_), .C(_abc_15497_new_n3716_), .Y(_abc_15497_new_n3717_));
OAI21X1 OAI21X1_743 ( .A(_auto_iopadmap_cc_368_execute_22625_144_), .B(_abc_15497_new_n883__bF_buf11), .C(_abc_15497_new_n1650__bF_buf1), .Y(_abc_15497_new_n3718_));
OAI21X1 OAI21X1_744 ( .A(_abc_15497_new_n2258_), .B(_abc_15497_new_n1648__bF_buf3), .C(_abc_15497_new_n3719_), .Y(_0a_reg_31_0__16_));
OAI21X1 OAI21X1_745 ( .A(_abc_15497_new_n3679_), .B(_abc_15497_new_n3707_), .C(_abc_15497_new_n3705_), .Y(_abc_15497_new_n3722_));
OAI21X1 OAI21X1_746 ( .A(_abc_15497_new_n3625_), .B(_abc_15497_new_n3631_), .C(_abc_15497_new_n3723_), .Y(_abc_15497_new_n3724_));
OAI21X1 OAI21X1_747 ( .A(_abc_15497_new_n3699_), .B(_abc_15497_new_n3697_), .C(_abc_15497_new_n3724_), .Y(_abc_15497_new_n3725_));
OAI21X1 OAI21X1_748 ( .A(_abc_15497_new_n3726_), .B(_abc_15497_new_n3729_), .C(_abc_15497_new_n3730_), .Y(_abc_15497_new_n3731_));
OAI21X1 OAI21X1_749 ( .A(b_reg_17_), .B(_abc_15497_new_n3726_), .C(_abc_15497_new_n3729_), .Y(_abc_15497_new_n3733_));
OAI21X1 OAI21X1_75 ( .A(_abc_15497_new_n1162_), .B(_abc_15497_new_n1163_), .C(_abc_15497_new_n1167_), .Y(_abc_15497_new_n1176_));
OAI21X1 OAI21X1_750 ( .A(_abc_15497_new_n2925__bF_buf0), .B(_abc_15497_new_n3732_), .C(_abc_15497_new_n3734_), .Y(_abc_15497_new_n3735_));
OAI21X1 OAI21X1_751 ( .A(_abc_15497_new_n3739_), .B(_abc_15497_new_n3740_), .C(_abc_15497_new_n3738_), .Y(_abc_15497_new_n3741_));
OAI21X1 OAI21X1_752 ( .A(_abc_15497_new_n3736_), .B(_abc_15497_new_n3737_), .C(_abc_15497_new_n3744_), .Y(_abc_15497_new_n3745_));
OAI21X1 OAI21X1_753 ( .A(_abc_15497_new_n3754_), .B(_abc_15497_new_n3759_), .C(_abc_15497_new_n2944_), .Y(_abc_15497_new_n3760_));
OAI21X1 OAI21X1_754 ( .A(_abc_15497_new_n3757_), .B(_abc_15497_new_n3758_), .C(_abc_15497_new_n3756_), .Y(_abc_15497_new_n3761_));
OAI21X1 OAI21X1_755 ( .A(_abc_15497_new_n3754_), .B(_abc_15497_new_n3759_), .C(_abc_15497_new_n2781__bF_buf0), .Y(_abc_15497_new_n3767_));
OAI21X1 OAI21X1_756 ( .A(_abc_15497_new_n3770_), .B(_abc_15497_new_n3721_), .C(round_ctr_inc_bF_buf7), .Y(_abc_15497_new_n3771_));
OAI21X1 OAI21X1_757 ( .A(_abc_15497_new_n2270_), .B(_abc_15497_new_n1648__bF_buf2), .C(_abc_15497_new_n3774_), .Y(_0a_reg_31_0__17_));
OAI21X1 OAI21X1_758 ( .A(_abc_15497_new_n2781__bF_buf3), .B(_abc_15497_new_n3754_), .C(_abc_15497_new_n3762_), .Y(_abc_15497_new_n3782_));
OAI21X1 OAI21X1_759 ( .A(_abc_15497_new_n3751_), .B(_abc_15497_new_n3752_), .C(_abc_15497_new_n3745_), .Y(_abc_15497_new_n3783_));
OAI21X1 OAI21X1_76 ( .A(_abc_15497_new_n1173_), .B(_abc_15497_new_n1171_), .C(_abc_15497_new_n1181_), .Y(_abc_15497_new_n1182_));
OAI21X1 OAI21X1_760 ( .A(d_reg_18_), .B(b_reg_18_), .C(_abc_15497_new_n3784_), .Y(_abc_15497_new_n3790_));
OAI21X1 OAI21X1_761 ( .A(d_reg_18_), .B(b_reg_18_), .C(c_reg_18_), .Y(_abc_15497_new_n3791_));
OAI21X1 OAI21X1_762 ( .A(_abc_15497_new_n1485_), .B(_abc_15497_new_n3785_), .C(_abc_15497_new_n3791_), .Y(_abc_15497_new_n3792_));
OAI21X1 OAI21X1_763 ( .A(_abc_15497_new_n2742__bF_buf1), .B(_abc_15497_new_n3790_), .C(_abc_15497_new_n3793_), .Y(_abc_15497_new_n3794_));
OAI21X1 OAI21X1_764 ( .A(_abc_15497_new_n1121_), .B(_abc_15497_new_n2214_), .C(_abc_15497_new_n3743_), .Y(_abc_15497_new_n3796_));
OAI21X1 OAI21X1_765 ( .A(_abc_15497_new_n3819_), .B(_abc_15497_new_n3781_), .C(round_ctr_inc_bF_buf6), .Y(_abc_15497_new_n3821_));
OAI21X1 OAI21X1_766 ( .A(_abc_15497_new_n3820_), .B(_abc_15497_new_n3821_), .C(_abc_15497_new_n3822_), .Y(_0a_reg_31_0__18_));
OAI21X1 OAI21X1_767 ( .A(_abc_15497_new_n3819_), .B(_abc_15497_new_n3781_), .C(_abc_15497_new_n3825_), .Y(_abc_15497_new_n3826_));
OAI21X1 OAI21X1_768 ( .A(_abc_15497_new_n3833_), .B(c_reg_19_), .C(_abc_15497_new_n3834_), .Y(_abc_15497_new_n3835_));
OAI21X1 OAI21X1_769 ( .A(d_reg_19_), .B(b_reg_19_), .C(c_reg_19_), .Y(_abc_15497_new_n3836_));
OAI21X1 OAI21X1_77 ( .A(_abc_15497_new_n1188_), .B(_abc_15497_new_n1183_), .C(digest_update_bF_buf2), .Y(_abc_15497_new_n1190_));
OAI21X1 OAI21X1_770 ( .A(_abc_15497_new_n1495_), .B(_abc_15497_new_n3833_), .C(_abc_15497_new_n3836_), .Y(_abc_15497_new_n3837_));
OAI21X1 OAI21X1_771 ( .A(_abc_15497_new_n2742__bF_buf0), .B(_abc_15497_new_n3835_), .C(_abc_15497_new_n3838_), .Y(_abc_15497_new_n3839_));
OAI21X1 OAI21X1_772 ( .A(_abc_15497_new_n1130_), .B(_abc_15497_new_n3531_), .C(_abc_15497_new_n3800_), .Y(_abc_15497_new_n3840_));
OAI21X1 OAI21X1_773 ( .A(_abc_15497_new_n3832_), .B(_abc_15497_new_n3839_), .C(_abc_15497_new_n3846_), .Y(_abc_15497_new_n3847_));
OAI21X1 OAI21X1_774 ( .A(_abc_15497_new_n3795_), .B(_abc_15497_new_n3802_), .C(_abc_15497_new_n3806_), .Y(_abc_15497_new_n3852_));
OAI21X1 OAI21X1_775 ( .A(_abc_15497_new_n3832_), .B(_abc_15497_new_n3839_), .C(_abc_15497_new_n3849_), .Y(_abc_15497_new_n3853_));
OAI21X1 OAI21X1_776 ( .A(_abc_15497_new_n3858_), .B(_abc_15497_new_n3857_), .C(_abc_15497_new_n3678_), .Y(_abc_15497_new_n3859_));
OAI21X1 OAI21X1_777 ( .A(_abc_15497_new_n3858_), .B(_abc_15497_new_n3857_), .C(_abc_15497_new_n3679_), .Y(_abc_15497_new_n3862_));
OAI21X1 OAI21X1_778 ( .A(_abc_15497_new_n3864_), .B(_abc_15497_new_n3826_), .C(round_ctr_inc_bF_buf5), .Y(_abc_15497_new_n3866_));
OAI21X1 OAI21X1_779 ( .A(_abc_15497_new_n3865_), .B(_abc_15497_new_n3866_), .C(_abc_15497_new_n3868_), .Y(_0a_reg_31_0__19_));
OAI21X1 OAI21X1_78 ( .A(_auto_iopadmap_cc_368_execute_22625_22_), .B(_abc_15497_new_n883__bF_buf0), .C(_abc_15497_new_n870__bF_buf7), .Y(_abc_15497_new_n1191_));
OAI21X1 OAI21X1_780 ( .A(_abc_15497_new_n3811_), .B(_abc_15497_new_n3812_), .C(_abc_15497_new_n3878_), .Y(_abc_15497_new_n3879_));
OAI21X1 OAI21X1_781 ( .A(_abc_15497_new_n3877_), .B(_abc_15497_new_n3824_), .C(_abc_15497_new_n3879_), .Y(_abc_15497_new_n3880_));
OAI21X1 OAI21X1_782 ( .A(_abc_15497_new_n3876_), .B(_abc_15497_new_n3779_), .C(_abc_15497_new_n3880_), .Y(_abc_15497_new_n3881_));
OAI21X1 OAI21X1_783 ( .A(_abc_15497_new_n3884_), .B(_abc_15497_new_n3675_), .C(_abc_15497_new_n3882_), .Y(_abc_15497_new_n3885_));
OAI21X1 OAI21X1_784 ( .A(_abc_15497_new_n3679_), .B(_abc_15497_new_n3857_), .C(_abc_15497_new_n3855_), .Y(_abc_15497_new_n3886_));
OAI21X1 OAI21X1_785 ( .A(_abc_15497_new_n3888_), .B(_abc_15497_new_n3889_), .C(_abc_15497_new_n3890_), .Y(_abc_15497_new_n3891_));
OAI21X1 OAI21X1_786 ( .A(_abc_15497_new_n3895_), .B(_abc_15497_new_n3896_), .C(_abc_15497_new_n2756__bF_buf1), .Y(_abc_15497_new_n3897_));
OAI21X1 OAI21X1_787 ( .A(d_reg_20_), .B(b_reg_20_), .C(c_reg_20_), .Y(_abc_15497_new_n3898_));
OAI21X1 OAI21X1_788 ( .A(_abc_15497_new_n1511_), .B(b_reg_20_), .C(_abc_15497_new_n3898_), .Y(_abc_15497_new_n3899_));
OAI21X1 OAI21X1_789 ( .A(_abc_15497_new_n1511_), .B(_abc_15497_new_n1958_), .C(_abc_15497_new_n3898_), .Y(_abc_15497_new_n3900_));
OAI21X1 OAI21X1_79 ( .A(_abc_15497_new_n1189_), .B(_abc_15497_new_n1190_), .C(_abc_15497_new_n1191_), .Y(_0H4_reg_31_0__22_));
OAI21X1 OAI21X1_790 ( .A(_abc_15497_new_n1146_), .B(_abc_15497_new_n2230_), .C(_abc_15497_new_n3844_), .Y(_abc_15497_new_n3903_));
OAI21X1 OAI21X1_791 ( .A(_abc_15497_new_n3848_), .B(_abc_15497_new_n3846_), .C(_abc_15497_new_n3891_), .Y(_abc_15497_new_n3915_));
OAI21X1 OAI21X1_792 ( .A(_abc_15497_new_n3920_), .B(_abc_15497_new_n3921_), .C(_abc_15497_new_n3678_), .Y(_abc_15497_new_n3922_));
OAI21X1 OAI21X1_793 ( .A(_abc_15497_new_n3920_), .B(_abc_15497_new_n3921_), .C(_abc_15497_new_n3679_), .Y(_abc_15497_new_n3926_));
OAI21X1 OAI21X1_794 ( .A(_abc_15497_new_n3929_), .B(_abc_15497_new_n3931_), .C(_abc_15497_new_n3933_), .Y(_0a_reg_31_0__20_));
OAI21X1 OAI21X1_795 ( .A(_abc_15497_new_n3679_), .B(_abc_15497_new_n3920_), .C(_abc_15497_new_n3918_), .Y(_abc_15497_new_n3937_));
OAI21X1 OAI21X1_796 ( .A(_abc_15497_new_n3938_), .B(_abc_15497_new_n3939_), .C(_abc_15497_new_n3940_), .Y(_abc_15497_new_n3941_));
OAI21X1 OAI21X1_797 ( .A(_abc_15497_new_n3945_), .B(_abc_15497_new_n3946_), .C(_abc_15497_new_n2756__bF_buf0), .Y(_abc_15497_new_n3947_));
OAI21X1 OAI21X1_798 ( .A(d_reg_21_), .B(b_reg_21_), .C(c_reg_21_), .Y(_abc_15497_new_n3949_));
OAI21X1 OAI21X1_799 ( .A(_abc_15497_new_n3948_), .B(b_reg_21_), .C(_abc_15497_new_n3949_), .Y(_abc_15497_new_n3950_));
OAI21X1 OAI21X1_8 ( .A(_abc_15497_new_n862_), .B(_abc_15497_new_n848_), .C(_abc_15497_new_n863_), .Y(_abc_15497_new_n864_));
OAI21X1 OAI21X1_80 ( .A(_abc_15497_new_n1184_), .B(_abc_15497_new_n1183_), .C(_abc_15497_new_n1185_), .Y(_abc_15497_new_n1193_));
OAI21X1 OAI21X1_800 ( .A(_abc_15497_new_n3948_), .B(_abc_15497_new_n1967_), .C(_abc_15497_new_n3949_), .Y(_abc_15497_new_n3951_));
OAI21X1 OAI21X1_801 ( .A(_abc_15497_new_n1162_), .B(_abc_15497_new_n2244_), .C(_abc_15497_new_n3907_), .Y(_abc_15497_new_n3954_));
OAI21X1 OAI21X1_802 ( .A(_abc_15497_new_n3911_), .B(_abc_15497_new_n3909_), .C(_abc_15497_new_n3941_), .Y(_abc_15497_new_n3966_));
OAI21X1 OAI21X1_803 ( .A(_abc_15497_new_n3971_), .B(_abc_15497_new_n3972_), .C(_abc_15497_new_n2780__bF_buf2), .Y(_abc_15497_new_n3973_));
OAI21X1 OAI21X1_804 ( .A(_abc_15497_new_n3971_), .B(_abc_15497_new_n3972_), .C(_abc_15497_new_n2755_), .Y(_abc_15497_new_n3977_));
OAI21X1 OAI21X1_805 ( .A(_abc_15497_new_n3980_), .B(_abc_15497_new_n3936_), .C(round_ctr_inc_bF_buf3), .Y(_abc_15497_new_n3982_));
OAI21X1 OAI21X1_806 ( .A(_abc_15497_new_n3981_), .B(_abc_15497_new_n3982_), .C(_abc_15497_new_n3984_), .Y(_0a_reg_31_0__21_));
OAI21X1 OAI21X1_807 ( .A(_abc_15497_new_n2755_), .B(_abc_15497_new_n3971_), .C(_abc_15497_new_n3969_), .Y(_abc_15497_new_n3992_));
OAI21X1 OAI21X1_808 ( .A(_abc_15497_new_n3993_), .B(_abc_15497_new_n3994_), .C(_abc_15497_new_n3995_), .Y(_abc_15497_new_n3996_));
OAI21X1 OAI21X1_809 ( .A(_abc_15497_new_n4000_), .B(_abc_15497_new_n4001_), .C(_abc_15497_new_n2756__bF_buf4), .Y(_abc_15497_new_n4002_));
OAI21X1 OAI21X1_81 ( .A(_auto_iopadmap_cc_368_execute_22625_23_), .B(_abc_15497_new_n883__bF_buf13), .C(_abc_15497_new_n870__bF_buf6), .Y(_abc_15497_new_n1199_));
OAI21X1 OAI21X1_810 ( .A(d_reg_22_), .B(b_reg_22_), .C(c_reg_22_), .Y(_abc_15497_new_n4003_));
OAI21X1 OAI21X1_811 ( .A(_abc_15497_new_n1530_), .B(b_reg_22_), .C(_abc_15497_new_n4003_), .Y(_abc_15497_new_n4004_));
OAI21X1 OAI21X1_812 ( .A(_abc_15497_new_n1530_), .B(_abc_15497_new_n4005_), .C(_abc_15497_new_n4003_), .Y(_abc_15497_new_n4006_));
OAI21X1 OAI21X1_813 ( .A(_abc_15497_new_n1173_), .B(_abc_15497_new_n2258_), .C(_abc_15497_new_n3958_), .Y(_abc_15497_new_n4009_));
OAI21X1 OAI21X1_814 ( .A(_abc_15497_new_n3962_), .B(_abc_15497_new_n3960_), .C(_abc_15497_new_n3996_), .Y(_abc_15497_new_n4021_));
OAI21X1 OAI21X1_815 ( .A(_abc_15497_new_n4026_), .B(_abc_15497_new_n4027_), .C(_abc_15497_new_n2756__bF_buf3), .Y(_abc_15497_new_n4028_));
OAI21X1 OAI21X1_816 ( .A(_abc_15497_new_n4026_), .B(_abc_15497_new_n4027_), .C(_abc_15497_new_n2925__bF_buf0), .Y(_abc_15497_new_n4032_));
OAI21X1 OAI21X1_817 ( .A(_abc_15497_new_n4035_), .B(_abc_15497_new_n3991_), .C(round_ctr_inc_bF_buf2), .Y(_abc_15497_new_n4037_));
OAI21X1 OAI21X1_818 ( .A(_abc_15497_new_n871__bF_buf1), .B(_abc_15497_new_n872__bF_buf2), .C(_abc_15497_new_n2331_), .Y(_abc_15497_new_n4038_));
OAI21X1 OAI21X1_819 ( .A(_abc_15497_new_n4036_), .B(_abc_15497_new_n4037_), .C(_abc_15497_new_n4039_), .Y(_0a_reg_31_0__22_));
OAI21X1 OAI21X1_82 ( .A(_abc_15497_new_n870__bF_buf5), .B(_abc_15497_new_n1198_), .C(_abc_15497_new_n1199_), .Y(_0H4_reg_31_0__23_));
OAI21X1 OAI21X1_820 ( .A(_abc_15497_new_n2925__bF_buf3), .B(_abc_15497_new_n4026_), .C(_abc_15497_new_n4024_), .Y(_abc_15497_new_n4044_));
OAI21X1 OAI21X1_821 ( .A(_abc_15497_new_n4045_), .B(_abc_15497_new_n4046_), .C(_abc_15497_new_n4047_), .Y(_abc_15497_new_n4048_));
OAI21X1 OAI21X1_822 ( .A(_abc_15497_new_n4017_), .B(_abc_15497_new_n4015_), .C(_abc_15497_new_n4048_), .Y(_abc_15497_new_n4049_));
OAI21X1 OAI21X1_823 ( .A(_abc_15497_new_n1543_), .B(_abc_15497_new_n4052_), .C(_abc_15497_new_n4053_), .Y(_abc_15497_new_n4054_));
OAI21X1 OAI21X1_824 ( .A(b_reg_23_), .B(_abc_15497_new_n1543_), .C(_abc_15497_new_n4052_), .Y(_abc_15497_new_n4056_));
OAI21X1 OAI21X1_825 ( .A(_abc_15497_new_n2925__bF_buf2), .B(_abc_15497_new_n4055_), .C(_abc_15497_new_n4057_), .Y(_abc_15497_new_n4058_));
OAI21X1 OAI21X1_826 ( .A(_abc_15497_new_n4010_), .B(_abc_15497_new_n4011_), .C(_abc_15497_new_n4062_), .Y(_abc_15497_new_n4063_));
OAI21X1 OAI21X1_827 ( .A(_abc_15497_new_n4074_), .B(_abc_15497_new_n4079_), .C(_abc_15497_new_n2739_), .Y(_abc_15497_new_n4080_));
OAI21X1 OAI21X1_828 ( .A(_abc_15497_new_n4074_), .B(_abc_15497_new_n4079_), .C(_abc_15497_new_n2738_), .Y(_abc_15497_new_n4087_));
OAI21X1 OAI21X1_829 ( .A(_abc_15497_new_n4041_), .B(_abc_15497_new_n4042_), .C(_abc_15497_new_n4089_), .Y(_abc_15497_new_n4092_));
OAI21X1 OAI21X1_83 ( .A(_abc_15497_new_n1201_), .B(_abc_15497_new_n1205_), .C(_abc_15497_new_n1206_), .Y(_abc_15497_new_n1207_));
OAI21X1 OAI21X1_830 ( .A(_abc_15497_new_n4093_), .B(_abc_15497_new_n4091_), .C(_abc_15497_new_n4095_), .Y(_0a_reg_31_0__23_));
OAI21X1 OAI21X1_831 ( .A(_abc_15497_new_n3990_), .B(_abc_15497_new_n4099_), .C(_abc_15497_new_n4102_), .Y(_abc_15497_new_n4103_));
OAI21X1 OAI21X1_832 ( .A(_abc_15497_new_n4105_), .B(_abc_15497_new_n3675_), .C(_abc_15497_new_n4104_), .Y(_abc_15497_new_n4106_));
OAI21X1 OAI21X1_833 ( .A(_abc_15497_new_n2738_), .B(_abc_15497_new_n4074_), .C(_abc_15497_new_n4082_), .Y(_abc_15497_new_n4107_));
OAI21X1 OAI21X1_834 ( .A(_abc_15497_new_n4059_), .B(_abc_15497_new_n4071_), .C(_abc_15497_new_n4068_), .Y(_abc_15497_new_n4108_));
OAI21X1 OAI21X1_835 ( .A(_abc_15497_new_n4109_), .B(_abc_15497_new_n4111_), .C(_abc_15497_new_n1562_), .Y(_abc_15497_new_n4112_));
OAI21X1 OAI21X1_836 ( .A(_abc_15497_new_n2006_), .B(_abc_15497_new_n855_), .C(_abc_15497_new_n4111_), .Y(_abc_15497_new_n4113_));
OAI21X1 OAI21X1_837 ( .A(b_reg_24_), .B(_abc_15497_new_n1562_), .C(_abc_15497_new_n4110_), .Y(_abc_15497_new_n4115_));
OAI21X1 OAI21X1_838 ( .A(_abc_15497_new_n4064_), .B(_abc_15497_new_n4065_), .C(_abc_15497_new_n4120_), .Y(_abc_15497_new_n4121_));
OAI21X1 OAI21X1_839 ( .A(_abc_15497_new_n4123_), .B(_abc_15497_new_n4124_), .C(_abc_15497_new_n4122_), .Y(_abc_15497_new_n4125_));
OAI21X1 OAI21X1_84 ( .A(_abc_15497_new_n1218_), .B(_abc_15497_new_n1210_), .C(digest_update_bF_buf1), .Y(_abc_15497_new_n1219_));
OAI21X1 OAI21X1_840 ( .A(_abc_15497_new_n4133_), .B(_abc_15497_new_n4135_), .C(_abc_15497_new_n2924__bF_buf0), .Y(_abc_15497_new_n4138_));
OAI21X1 OAI21X1_841 ( .A(_abc_15497_new_n4106_), .B(_abc_15497_new_n4143_), .C(_abc_15497_new_n4144_), .Y(_abc_15497_new_n4145_));
OAI21X1 OAI21X1_842 ( .A(_auto_iopadmap_cc_368_execute_22625_152_), .B(_abc_15497_new_n883__bF_buf5), .C(_abc_15497_new_n1650__bF_buf3), .Y(_abc_15497_new_n4146_));
OAI21X1 OAI21X1_843 ( .A(_abc_15497_new_n2360_), .B(_abc_15497_new_n1648__bF_buf1), .C(_abc_15497_new_n4147_), .Y(_0a_reg_31_0__24_));
OAI21X1 OAI21X1_844 ( .A(_abc_15497_new_n2924__bF_buf4), .B(_abc_15497_new_n4133_), .C(_abc_15497_new_n4134_), .Y(_abc_15497_new_n4151_));
OAI21X1 OAI21X1_845 ( .A(_abc_15497_new_n4152_), .B(_abc_15497_new_n4131_), .C(_abc_15497_new_n4128_), .Y(_abc_15497_new_n4153_));
OAI21X1 OAI21X1_846 ( .A(_abc_15497_new_n1572_), .B(_abc_15497_new_n4156_), .C(_abc_15497_new_n4157_), .Y(_abc_15497_new_n4158_));
OAI21X1 OAI21X1_847 ( .A(d_reg_25_), .B(_abc_15497_new_n4155_), .C(_abc_15497_new_n4158_), .Y(_abc_15497_new_n4159_));
OAI21X1 OAI21X1_848 ( .A(b_reg_25_), .B(_abc_15497_new_n1572_), .C(_abc_15497_new_n4156_), .Y(_abc_15497_new_n4160_));
OAI21X1 OAI21X1_849 ( .A(_abc_15497_new_n2925__bF_buf1), .B(_abc_15497_new_n4159_), .C(_abc_15497_new_n4161_), .Y(_abc_15497_new_n4162_));
OAI21X1 OAI21X1_85 ( .A(_auto_iopadmap_cc_368_execute_22625_24_), .B(_abc_15497_new_n883__bF_buf12), .C(_abc_15497_new_n870__bF_buf4), .Y(_abc_15497_new_n1220_));
OAI21X1 OAI21X1_850 ( .A(_abc_15497_new_n4141_), .B(_abc_15497_new_n4139_), .C(_abc_15497_new_n4150_), .Y(_abc_15497_new_n4181_));
OAI21X1 OAI21X1_851 ( .A(_abc_15497_new_n4182_), .B(_abc_15497_new_n4181_), .C(round_ctr_inc_bF_buf0), .Y(_abc_15497_new_n4183_));
OAI21X1 OAI21X1_852 ( .A(_abc_15497_new_n871__bF_buf0), .B(_abc_15497_new_n872__bF_buf1), .C(_abc_15497_new_n2371_), .Y(_abc_15497_new_n4184_));
OAI21X1 OAI21X1_853 ( .A(_abc_15497_new_n4180_), .B(_abc_15497_new_n4183_), .C(_abc_15497_new_n4185_), .Y(_0a_reg_31_0__25_));
OAI21X1 OAI21X1_854 ( .A(_abc_15497_new_n4141_), .B(_abc_15497_new_n4139_), .C(_abc_15497_new_n4178_), .Y(_abc_15497_new_n4187_));
OAI21X1 OAI21X1_855 ( .A(_abc_15497_new_n4151_), .B(_abc_15497_new_n4176_), .C(_abc_15497_new_n4187_), .Y(_abc_15497_new_n4188_));
OAI21X1 OAI21X1_856 ( .A(_abc_15497_new_n4163_), .B(_abc_15497_new_n4168_), .C(_abc_15497_new_n4192_), .Y(_abc_15497_new_n4193_));
OAI21X1 OAI21X1_857 ( .A(_abc_15497_new_n4196_), .B(_abc_15497_new_n4198_), .C(_abc_15497_new_n2756__bF_buf4), .Y(_abc_15497_new_n4199_));
OAI21X1 OAI21X1_858 ( .A(b_reg_26_), .B(_abc_15497_new_n1586_), .C(_abc_15497_new_n4194_), .Y(_abc_15497_new_n4200_));
OAI21X1 OAI21X1_859 ( .A(_abc_15497_new_n866_), .B(_abc_15497_new_n2031_), .C(_abc_15497_new_n1586_), .Y(_abc_15497_new_n4201_));
OAI21X1 OAI21X1_86 ( .A(_abc_15497_new_n1219_), .B(_abc_15497_new_n1217_), .C(_abc_15497_new_n1220_), .Y(_0H4_reg_31_0__24_));
OAI21X1 OAI21X1_860 ( .A(_abc_15497_new_n4165_), .B(_abc_15497_new_n2310_), .C(_abc_15497_new_n4205_), .Y(_abc_15497_new_n4206_));
OAI21X1 OAI21X1_861 ( .A(_abc_15497_new_n4208_), .B(_abc_15497_new_n4209_), .C(_abc_15497_new_n4207_), .Y(_abc_15497_new_n4210_));
OAI21X1 OAI21X1_862 ( .A(_abc_15497_new_n4216_), .B(_abc_15497_new_n4217_), .C(_abc_15497_new_n3679_), .Y(_abc_15497_new_n4220_));
OAI21X1 OAI21X1_863 ( .A(_abc_15497_new_n4221_), .B(_abc_15497_new_n4219_), .C(_abc_15497_new_n4174_), .Y(_abc_15497_new_n4222_));
OAI21X1 OAI21X1_864 ( .A(_abc_15497_new_n2781__bF_buf2), .B(_abc_15497_new_n2759__bF_buf4), .C(_abc_15497_new_n4218_), .Y(_abc_15497_new_n4223_));
OAI21X1 OAI21X1_865 ( .A(_abc_15497_new_n4191_), .B(_abc_15497_new_n4225_), .C(_abc_15497_new_n4226_), .Y(_abc_15497_new_n4227_));
OAI21X1 OAI21X1_866 ( .A(_auto_iopadmap_cc_368_execute_22625_154_), .B(_abc_15497_new_n883__bF_buf4), .C(_abc_15497_new_n1650__bF_buf1), .Y(_abc_15497_new_n4228_));
OAI21X1 OAI21X1_867 ( .A(_abc_15497_new_n2385_), .B(_abc_15497_new_n1648__bF_buf0), .C(_abc_15497_new_n4229_), .Y(_0a_reg_31_0__26_));
OAI21X1 OAI21X1_868 ( .A(_abc_15497_new_n4173_), .B(_abc_15497_new_n4231_), .C(_abc_15497_new_n4232_), .Y(_abc_15497_new_n4233_));
OAI21X1 OAI21X1_869 ( .A(_abc_15497_new_n3679_), .B(_abc_15497_new_n4216_), .C(_abc_15497_new_n4234_), .Y(_abc_15497_new_n4235_));
OAI21X1 OAI21X1_87 ( .A(_abc_15497_new_n1212_), .B(_abc_15497_new_n1210_), .C(_abc_15497_new_n1222_), .Y(_abc_15497_new_n1223_));
OAI21X1 OAI21X1_870 ( .A(_abc_15497_new_n4236_), .B(_abc_15497_new_n4214_), .C(_abc_15497_new_n4237_), .Y(_abc_15497_new_n4238_));
OAI21X1 OAI21X1_871 ( .A(_abc_15497_new_n4239_), .B(_abc_15497_new_n4240_), .C(_abc_15497_new_n1596_), .Y(_abc_15497_new_n4241_));
OAI21X1 OAI21X1_872 ( .A(c_reg_27_), .B(b_reg_27_), .C(_abc_15497_new_n4241_), .Y(_abc_15497_new_n4242_));
OAI21X1 OAI21X1_873 ( .A(b_reg_27_), .B(_abc_15497_new_n1596_), .C(_abc_15497_new_n4243_), .Y(_abc_15497_new_n4247_));
OAI21X1 OAI21X1_874 ( .A(_abc_15497_new_n2924__bF_buf3), .B(_abc_15497_new_n4242_), .C(_abc_15497_new_n4248_), .Y(_abc_15497_new_n4249_));
OAI21X1 OAI21X1_875 ( .A(_abc_15497_new_n4263_), .B(_abc_15497_new_n4233_), .C(round_ctr_inc_bF_buf13), .Y(_abc_15497_new_n4265_));
OAI21X1 OAI21X1_876 ( .A(_abc_15497_new_n4264_), .B(_abc_15497_new_n4265_), .C(_abc_15497_new_n4267_), .Y(_0a_reg_31_0__27_));
OAI21X1 OAI21X1_877 ( .A(_abc_15497_new_n4188_), .B(_abc_15497_new_n4270_), .C(_abc_15497_new_n4273_), .Y(_abc_15497_new_n4274_));
OAI21X1 OAI21X1_878 ( .A(_abc_15497_new_n4250_), .B(_abc_15497_new_n4255_), .C(_abc_15497_new_n4278_), .Y(_abc_15497_new_n4279_));
OAI21X1 OAI21X1_879 ( .A(_abc_15497_new_n2925__bF_buf0), .B(_abc_15497_new_n4284_), .C(_abc_15497_new_n4288_), .Y(_abc_15497_new_n4289_));
OAI21X1 OAI21X1_88 ( .A(_auto_iopadmap_cc_368_execute_22625_25_), .B(_abc_15497_new_n883__bF_buf11), .C(_abc_15497_new_n870__bF_buf3), .Y(_abc_15497_new_n1229_));
OAI21X1 OAI21X1_880 ( .A(_abc_15497_new_n4302_), .B(_abc_15497_new_n4303_), .C(_abc_15497_new_n4275_), .Y(_abc_15497_new_n4304_));
OAI21X1 OAI21X1_881 ( .A(_abc_15497_new_n3673_), .B(_abc_15497_new_n4312_), .C(_abc_15497_new_n4314_), .Y(_abc_15497_new_n4315_));
OAI21X1 OAI21X1_882 ( .A(_abc_15497_new_n4274_), .B(_abc_15497_new_n4317_), .C(_abc_15497_new_n4318_), .Y(_abc_15497_new_n4319_));
OAI21X1 OAI21X1_883 ( .A(_abc_15497_new_n1646_), .B(_abc_15497_new_n4320_), .C(_abc_15497_new_n4322_), .Y(_0a_reg_31_0__28_));
OAI21X1 OAI21X1_884 ( .A(_abc_15497_new_n4302_), .B(_abc_15497_new_n4275_), .C(_abc_15497_new_n4324_), .Y(_abc_15497_new_n4325_));
OAI21X1 OAI21X1_885 ( .A(_abc_15497_new_n4291_), .B(_abc_15497_new_n4295_), .C(_abc_15497_new_n4328_), .Y(_abc_15497_new_n4329_));
OAI21X1 OAI21X1_886 ( .A(_abc_15497_new_n4334_), .B(_abc_15497_new_n4331_), .C(d_reg_29_), .Y(_abc_15497_new_n4337_));
OAI21X1 OAI21X1_887 ( .A(d_reg_29_), .B(_abc_15497_new_n4331_), .C(_abc_15497_new_n4339_), .Y(_abc_15497_new_n4340_));
OAI21X1 OAI21X1_888 ( .A(_abc_15497_new_n2924__bF_buf2), .B(_abc_15497_new_n4340_), .C(_abc_15497_new_n2742__bF_buf2), .Y(_abc_15497_new_n4341_));
OAI21X1 OAI21X1_889 ( .A(_abc_15497_new_n4341_), .B(_abc_15497_new_n4338_), .C(_abc_15497_new_n4333_), .Y(_abc_15497_new_n4342_));
OAI21X1 OAI21X1_89 ( .A(_abc_15497_new_n870__bF_buf2), .B(_abc_15497_new_n1228_), .C(_abc_15497_new_n1229_), .Y(_0H4_reg_31_0__25_));
OAI21X1 OAI21X1_890 ( .A(_abc_15497_new_n2738_), .B(_abc_15497_new_n2743__bF_buf2), .C(_abc_15497_new_n4353_), .Y(_abc_15497_new_n4354_));
OAI21X1 OAI21X1_891 ( .A(_abc_15497_new_n4359_), .B(_abc_15497_new_n4325_), .C(round_ctr_inc_bF_buf12), .Y(_abc_15497_new_n4361_));
OAI21X1 OAI21X1_892 ( .A(_abc_15497_new_n871__bF_buf4), .B(_abc_15497_new_n872__bF_buf0), .C(_abc_15497_new_n2417_), .Y(_abc_15497_new_n4362_));
OAI21X1 OAI21X1_893 ( .A(_abc_15497_new_n4360_), .B(_abc_15497_new_n4361_), .C(_abc_15497_new_n4363_), .Y(_0a_reg_31_0__29_));
OAI21X1 OAI21X1_894 ( .A(_abc_15497_new_n4365_), .B(_abc_15497_new_n4275_), .C(_abc_15497_new_n4367_), .Y(_abc_15497_new_n4368_));
OAI21X1 OAI21X1_895 ( .A(_abc_15497_new_n2944_), .B(_abc_15497_new_n4353_), .C(_abc_15497_new_n4369_), .Y(_abc_15497_new_n4370_));
OAI21X1 OAI21X1_896 ( .A(_abc_15497_new_n4343_), .B(_abc_15497_new_n4347_), .C(_abc_15497_new_n4350_), .Y(_abc_15497_new_n4371_));
OAI21X1 OAI21X1_897 ( .A(_abc_15497_new_n4376_), .B(_abc_15497_new_n4373_), .C(d_reg_30_), .Y(_abc_15497_new_n4379_));
OAI21X1 OAI21X1_898 ( .A(d_reg_30_), .B(_abc_15497_new_n4373_), .C(_abc_15497_new_n4381_), .Y(_abc_15497_new_n4382_));
OAI21X1 OAI21X1_899 ( .A(_abc_15497_new_n2924__bF_buf1), .B(_abc_15497_new_n4382_), .C(_abc_15497_new_n2742__bF_buf1), .Y(_abc_15497_new_n4383_));
OAI21X1 OAI21X1_9 ( .A(_abc_15497_new_n871__bF_buf4), .B(_abc_15497_new_n872__bF_buf4), .C(_abc_15497_new_n870__bF_buf11), .Y(_abc_15497_new_n873_));
OAI21X1 OAI21X1_90 ( .A(_abc_15497_new_n1224_), .B(_abc_15497_new_n1222_), .C(_abc_15497_new_n1225_), .Y(_abc_15497_new_n1235_));
OAI21X1 OAI21X1_900 ( .A(_abc_15497_new_n4383_), .B(_abc_15497_new_n4380_), .C(_abc_15497_new_n4375_), .Y(_abc_15497_new_n4384_));
OAI21X1 OAI21X1_901 ( .A(_abc_15497_new_n1273_), .B(_abc_15497_new_n2360_), .C(_abc_15497_new_n4385_), .Y(_abc_15497_new_n4386_));
OAI21X1 OAI21X1_902 ( .A(_abc_15497_new_n871__bF_buf3), .B(_abc_15497_new_n872__bF_buf4), .C(_abc_15497_new_n2425_), .Y(_abc_15497_new_n4403_));
OAI21X1 OAI21X1_903 ( .A(_abc_15497_new_n1646_), .B(_abc_15497_new_n4402_), .C(_abc_15497_new_n4404_), .Y(_0a_reg_31_0__30_));
OAI21X1 OAI21X1_904 ( .A(_abc_15497_new_n4274_), .B(_abc_15497_new_n4317_), .C(_abc_15497_new_n4407_), .Y(_abc_15497_new_n4408_));
OAI21X1 OAI21X1_905 ( .A(_abc_15497_new_n2759__bF_buf2), .B(_abc_15497_new_n4412_), .C(_abc_15497_new_n4411_), .Y(_abc_15497_new_n4413_));
OAI21X1 OAI21X1_906 ( .A(_abc_15497_new_n4384_), .B(_abc_15497_new_n4395_), .C(_abc_15497_new_n4414_), .Y(_abc_15497_new_n4415_));
OAI21X1 OAI21X1_907 ( .A(d_reg_31_), .B(_abc_15497_new_n4418_), .C(_abc_15497_new_n4422_), .Y(_abc_15497_new_n4423_));
OAI21X1 OAI21X1_908 ( .A(_abc_15497_new_n2743__bF_buf5), .B(_abc_15497_new_n4424_), .C(_abc_15497_new_n4417_), .Y(_abc_15497_new_n4425_));
OAI21X1 OAI21X1_909 ( .A(_abc_15497_new_n4388_), .B(_abc_15497_new_n2372_), .C(_abc_15497_new_n4392_), .Y(_abc_15497_new_n4426_));
OAI21X1 OAI21X1_91 ( .A(_abc_15497_new_n1234_), .B(_abc_15497_new_n1210_), .C(_abc_15497_new_n1236_), .Y(_abc_15497_new_n1237_));
OAI21X1 OAI21X1_910 ( .A(_abc_15497_new_n4436_), .B(_abc_15497_new_n4435_), .C(round_ctr_inc_bF_buf11), .Y(_abc_15497_new_n4437_));
OAI21X1 OAI21X1_911 ( .A(_abc_15497_new_n4434_), .B(_abc_15497_new_n4437_), .C(_abc_15497_new_n4439_), .Y(_0a_reg_31_0__31_));
OAI21X1 OAI21X1_912 ( .A(_abc_15497_new_n871__bF_buf2), .B(_abc_15497_new_n4449_), .C(_abc_15497_new_n870__bF_buf10), .Y(_abc_15497_abc_9717_auto_fsm_map_cc_170_map_fsm_844_0_));
OAI21X1 OAI21X1_913 ( .A(_abc_15497_new_n1646_), .B(_abc_15497_new_n4447_), .C(_abc_15497_new_n870__bF_buf9), .Y(_abc_15497_new_n4451_));
OAI21X1 OAI21X1_914 ( .A(_abc_15497_new_n1646_), .B(_abc_15497_new_n4451_), .C(_abc_15497_new_n1644_), .Y(_abc_15497_abc_9717_auto_fsm_map_cc_170_map_fsm_844_2_));
OAI21X1 OAI21X1_915 ( .A(_abc_15497_new_n4443_), .B(_abc_15497_new_n1648__bF_buf8), .C(_abc_15497_new_n4453_), .Y(_0round_ctr_reg_6_0__0_));
OAI21X1 OAI21X1_916 ( .A(_abc_15497_new_n4442_), .B(_abc_15497_new_n4443_), .C(round_ctr_inc_bF_buf8), .Y(_abc_15497_new_n4456_));
OAI21X1 OAI21X1_917 ( .A(round_ctr_inc_bF_buf6), .B(_abc_15497_new_n1644_), .C(round_ctr_reg_3_), .Y(_abc_15497_new_n4462_));
OAI21X1 OAI21X1_918 ( .A(round_ctr_inc_bF_buf5), .B(_abc_15497_new_n1644_), .C(round_ctr_reg_4_), .Y(_abc_15497_new_n4466_));
OAI21X1 OAI21X1_919 ( .A(round_ctr_inc_bF_buf4), .B(_abc_15497_new_n1644_), .C(round_ctr_reg_5_), .Y(_abc_15497_new_n4469_));
OAI21X1 OAI21X1_92 ( .A(_abc_15497_new_n1244_), .B(_abc_15497_new_n1243_), .C(digest_update_bF_buf0), .Y(_abc_15497_new_n1245_));
OAI21X1 OAI21X1_920 ( .A(round_ctr_inc_bF_buf3), .B(_abc_15497_new_n1644_), .C(round_ctr_reg_6_), .Y(_abc_15497_new_n4472_));
OAI21X1 OAI21X1_921 ( .A(_abc_15497_new_n4474_), .B(round_ctr_rst_bF_buf7), .C(_abc_15497_new_n870__bF_buf8), .Y(_0digest_valid_reg_0_0_));
OAI21X1 OAI21X1_922 ( .A(_abc_15497_new_n769_), .B(_abc_15497_new_n770_), .C(digest_update_bF_buf3), .Y(_abc_15497_new_n4477_));
OAI21X1 OAI21X1_923 ( .A(_auto_iopadmap_cc_368_execute_22625_67_), .B(_abc_15497_new_n883__bF_buf12), .C(_abc_15497_new_n870__bF_buf7), .Y(_abc_15497_new_n4488_));
OAI21X1 OAI21X1_924 ( .A(_abc_15497_new_n870__bF_buf6), .B(_abc_15497_new_n4487_), .C(_abc_15497_new_n4488_), .Y(_0H2_reg_31_0__3_));
OAI21X1 OAI21X1_925 ( .A(_abc_15497_new_n4495_), .B(_abc_15497_new_n4494_), .C(digest_update_bF_buf8), .Y(_abc_15497_new_n4496_));
OAI21X1 OAI21X1_926 ( .A(_auto_iopadmap_cc_368_execute_22625_69_), .B(_abc_15497_new_n883__bF_buf10), .C(_abc_15497_new_n870__bF_buf5), .Y(_abc_15497_new_n4497_));
OAI21X1 OAI21X1_927 ( .A(_abc_15497_new_n750_), .B(_abc_15497_new_n755_), .C(_abc_15497_new_n4501_), .Y(_abc_15497_new_n4502_));
OAI21X1 OAI21X1_928 ( .A(_auto_iopadmap_cc_368_execute_22625_70_), .B(_abc_15497_new_n883__bF_buf9), .C(_abc_15497_new_n870__bF_buf4), .Y(_abc_15497_new_n4505_));
OAI21X1 OAI21X1_929 ( .A(_abc_15497_new_n870__bF_buf3), .B(_abc_15497_new_n4504_), .C(_abc_15497_new_n4505_), .Y(_0H2_reg_31_0__6_));
OAI21X1 OAI21X1_93 ( .A(_abc_15497_new_n1239_), .B(_abc_15497_new_n1231_), .C(_abc_15497_new_n1253_), .Y(_abc_15497_new_n1254_));
OAI21X1 OAI21X1_930 ( .A(_abc_15497_new_n748_), .B(_abc_15497_new_n749_), .C(_abc_15497_new_n4503_), .Y(_abc_15497_new_n4507_));
OAI21X1 OAI21X1_931 ( .A(_auto_iopadmap_cc_368_execute_22625_71_), .B(_abc_15497_new_n883__bF_buf8), .C(_abc_15497_new_n870__bF_buf2), .Y(_abc_15497_new_n4509_));
OAI21X1 OAI21X1_932 ( .A(_abc_15497_new_n870__bF_buf1), .B(_abc_15497_new_n4508_), .C(_abc_15497_new_n4509_), .Y(_0H2_reg_31_0__7_));
OAI21X1 OAI21X1_933 ( .A(_abc_15497_new_n757_), .B(_abc_15497_new_n4501_), .C(_abc_15497_new_n753_), .Y(_abc_15497_new_n4511_));
OAI21X1 OAI21X1_934 ( .A(_abc_15497_new_n787_), .B(_abc_15497_new_n783_), .C(digest_update_bF_buf7), .Y(_abc_15497_new_n4513_));
OAI21X1 OAI21X1_935 ( .A(_abc_15497_new_n784_), .B(_abc_15497_new_n4515_), .C(digest_update_bF_buf6), .Y(_abc_15497_new_n4517_));
OAI21X1 OAI21X1_936 ( .A(_abc_15497_new_n729_), .B(_abc_15497_new_n734_), .C(_abc_15497_new_n4520_), .Y(_abc_15497_new_n4521_));
OAI21X1 OAI21X1_937 ( .A(_auto_iopadmap_cc_368_execute_22625_74_), .B(_abc_15497_new_n883__bF_buf7), .C(_abc_15497_new_n870__bF_buf0), .Y(_abc_15497_new_n4524_));
OAI21X1 OAI21X1_938 ( .A(_abc_15497_new_n870__bF_buf11), .B(_abc_15497_new_n4523_), .C(_abc_15497_new_n4524_), .Y(_0H2_reg_31_0__10_));
OAI21X1 OAI21X1_939 ( .A(_abc_15497_new_n727_), .B(_abc_15497_new_n728_), .C(_abc_15497_new_n4522_), .Y(_abc_15497_new_n4526_));
OAI21X1 OAI21X1_94 ( .A(_abc_15497_new_n1240_), .B(_abc_15497_new_n1248_), .C(_abc_15497_new_n1252_), .Y(_abc_15497_new_n1255_));
OAI21X1 OAI21X1_940 ( .A(_auto_iopadmap_cc_368_execute_22625_75_), .B(_abc_15497_new_n883__bF_buf6), .C(_abc_15497_new_n870__bF_buf10), .Y(_abc_15497_new_n4528_));
OAI21X1 OAI21X1_941 ( .A(_abc_15497_new_n870__bF_buf9), .B(_abc_15497_new_n4527_), .C(_abc_15497_new_n4528_), .Y(_0H2_reg_31_0__11_));
OAI21X1 OAI21X1_942 ( .A(_abc_15497_new_n736_), .B(_abc_15497_new_n4520_), .C(_abc_15497_new_n732_), .Y(_abc_15497_new_n4530_));
OAI21X1 OAI21X1_943 ( .A(_abc_15497_new_n721_), .B(_abc_15497_new_n791_), .C(digest_update_bF_buf5), .Y(_abc_15497_new_n4532_));
OAI21X1 OAI21X1_944 ( .A(_auto_iopadmap_cc_368_execute_22625_76_), .B(_abc_15497_new_n883__bF_buf5), .C(_abc_15497_new_n870__bF_buf8), .Y(_abc_15497_new_n4533_));
OAI21X1 OAI21X1_945 ( .A(_abc_15497_new_n4531_), .B(_abc_15497_new_n4532_), .C(_abc_15497_new_n4533_), .Y(_0H2_reg_31_0__12_));
OAI21X1 OAI21X1_946 ( .A(_abc_15497_new_n718_), .B(_abc_15497_new_n4535_), .C(digest_update_bF_buf4), .Y(_abc_15497_new_n4537_));
OAI21X1 OAI21X1_947 ( .A(_abc_15497_new_n723_), .B(_abc_15497_new_n791_), .C(_abc_15497_new_n714_), .Y(_abc_15497_new_n4539_));
OAI21X1 OAI21X1_948 ( .A(_auto_iopadmap_cc_368_execute_22625_78_), .B(_abc_15497_new_n883__bF_buf4), .C(_abc_15497_new_n870__bF_buf7), .Y(_abc_15497_new_n4543_));
OAI21X1 OAI21X1_949 ( .A(_abc_15497_new_n4540_), .B(_abc_15497_new_n4542_), .C(_abc_15497_new_n4543_), .Y(_0H2_reg_31_0__14_));
OAI21X1 OAI21X1_95 ( .A(_abc_15497_new_n1248_), .B(_abc_15497_new_n1254_), .C(_abc_15497_new_n1255_), .Y(_abc_15497_new_n1256_));
OAI21X1 OAI21X1_950 ( .A(_abc_15497_new_n702_), .B(_abc_15497_new_n703_), .C(_abc_15497_new_n4541_), .Y(_abc_15497_new_n4545_));
OAI21X1 OAI21X1_951 ( .A(_auto_iopadmap_cc_368_execute_22625_79_), .B(_abc_15497_new_n883__bF_buf3), .C(_abc_15497_new_n870__bF_buf6), .Y(_abc_15497_new_n4547_));
OAI21X1 OAI21X1_952 ( .A(_abc_15497_new_n870__bF_buf5), .B(_abc_15497_new_n4546_), .C(_abc_15497_new_n4547_), .Y(_0H2_reg_31_0__15_));
OAI21X1 OAI21X1_953 ( .A(_abc_15497_new_n843_), .B(_abc_15497_new_n4550_), .C(digest_update_bF_buf2), .Y(_abc_15497_new_n4551_));
OAI21X1 OAI21X1_954 ( .A(_auto_iopadmap_cc_368_execute_22625_81_), .B(_abc_15497_new_n883__bF_buf2), .C(_abc_15497_new_n870__bF_buf4), .Y(_abc_15497_new_n4555_));
OAI21X1 OAI21X1_955 ( .A(_abc_15497_new_n870__bF_buf3), .B(_abc_15497_new_n4554_), .C(_abc_15497_new_n4555_), .Y(_0H2_reg_31_0__17_));
OAI21X1 OAI21X1_956 ( .A(_abc_15497_new_n845_), .B(_abc_15497_new_n4550_), .C(_abc_15497_new_n835_), .Y(_abc_15497_new_n4557_));
OAI21X1 OAI21X1_957 ( .A(_auto_iopadmap_cc_368_execute_22625_83_), .B(_abc_15497_new_n883__bF_buf1), .C(_abc_15497_new_n870__bF_buf1), .Y(_abc_15497_new_n4562_));
OAI21X1 OAI21X1_958 ( .A(_abc_15497_new_n870__bF_buf0), .B(_abc_15497_new_n4561_), .C(_abc_15497_new_n4562_), .Y(_0H2_reg_31_0__19_));
OAI21X1 OAI21X1_959 ( .A(_abc_15497_new_n816_), .B(_abc_15497_new_n4567_), .C(digest_update_bF_buf1), .Y(_abc_15497_new_n4568_));
OAI21X1 OAI21X1_96 ( .A(_abc_15497_new_n1250_), .B(_abc_15497_new_n1247_), .C(_abc_15497_new_n1261_), .Y(_abc_15497_new_n1262_));
OAI21X1 OAI21X1_960 ( .A(_auto_iopadmap_cc_368_execute_22625_84_), .B(_abc_15497_new_n883__bF_buf0), .C(_abc_15497_new_n870__bF_buf11), .Y(_abc_15497_new_n4569_));
OAI21X1 OAI21X1_961 ( .A(_abc_15497_new_n4568_), .B(_abc_15497_new_n4566_), .C(_abc_15497_new_n4569_), .Y(_0H2_reg_31_0__20_));
OAI21X1 OAI21X1_962 ( .A(_abc_15497_new_n4573_), .B(_abc_15497_new_n4572_), .C(digest_update_bF_buf0), .Y(_abc_15497_new_n4574_));
OAI21X1 OAI21X1_963 ( .A(_auto_iopadmap_cc_368_execute_22625_85_), .B(_abc_15497_new_n883__bF_buf13), .C(_abc_15497_new_n870__bF_buf10), .Y(_abc_15497_new_n4575_));
OAI21X1 OAI21X1_964 ( .A(_abc_15497_new_n818_), .B(_abc_15497_new_n4567_), .C(_abc_15497_new_n810_), .Y(_abc_15497_new_n4577_));
OAI21X1 OAI21X1_965 ( .A(_abc_15497_new_n803_), .B(_abc_15497_new_n4579_), .C(digest_update_bF_buf8), .Y(_abc_15497_new_n4580_));
OAI21X1 OAI21X1_966 ( .A(_abc_15497_new_n801_), .B(_abc_15497_new_n4579_), .C(_abc_15497_new_n4583_), .Y(_abc_15497_new_n4584_));
OAI21X1 OAI21X1_967 ( .A(_abc_15497_new_n860_), .B(_abc_15497_new_n848_), .C(digest_update_bF_buf7), .Y(_abc_15497_new_n4589_));
OAI21X1 OAI21X1_968 ( .A(_abc_15497_new_n854_), .B(_abc_15497_new_n4592_), .C(digest_update_bF_buf6), .Y(_abc_15497_new_n4594_));
OAI21X1 OAI21X1_969 ( .A(w_mem_inst__abc_19396_new_n1591_), .B(w_mem_inst__abc_19396_new_n1598__bF_buf4), .C(w_mem_inst__abc_19396_new_n1586__bF_buf3), .Y(w_mem_inst__abc_19396_new_n1599_));
OAI21X1 OAI21X1_97 ( .A(_abc_15497_new_n1262_), .B(_abc_15497_new_n1260_), .C(_abc_15497_new_n1264_), .Y(_abc_15497_new_n1266_));
OAI21X1 OAI21X1_970 ( .A(w_mem_inst__abc_19396_new_n1600_), .B(w_mem_inst__abc_19396_new_n1604__bF_buf4), .C(w_mem_inst__abc_19396_new_n1607_), .Y(w_mem_inst__abc_19396_new_n1608_));
OAI21X1 OAI21X1_971 ( .A(w_mem_inst__abc_19396_new_n1609_), .B(w_mem_inst__abc_19396_new_n1611__bF_buf4), .C(w_mem_inst__abc_19396_new_n1614_), .Y(w_mem_inst__abc_19396_new_n1615_));
OAI21X1 OAI21X1_972 ( .A(w_mem_inst__abc_19396_new_n1646_), .B(w_mem_inst__abc_19396_new_n1598__bF_buf3), .C(w_mem_inst__abc_19396_new_n1586__bF_buf2), .Y(w_mem_inst__abc_19396_new_n1647_));
OAI21X1 OAI21X1_973 ( .A(w_mem_inst__abc_19396_new_n1648_), .B(w_mem_inst__abc_19396_new_n1604__bF_buf3), .C(w_mem_inst__abc_19396_new_n1649_), .Y(w_mem_inst__abc_19396_new_n1650_));
OAI21X1 OAI21X1_974 ( .A(w_mem_inst__abc_19396_new_n1651_), .B(w_mem_inst__abc_19396_new_n1611__bF_buf3), .C(w_mem_inst__abc_19396_new_n1652_), .Y(w_mem_inst__abc_19396_new_n1653_));
OAI21X1 OAI21X1_975 ( .A(w_mem_inst__abc_19396_new_n1671_), .B(w_mem_inst__abc_19396_new_n1598__bF_buf2), .C(w_mem_inst__abc_19396_new_n1586__bF_buf1), .Y(w_mem_inst__abc_19396_new_n1672_));
OAI21X1 OAI21X1_976 ( .A(w_mem_inst__abc_19396_new_n1673_), .B(w_mem_inst__abc_19396_new_n1604__bF_buf2), .C(w_mem_inst__abc_19396_new_n1674_), .Y(w_mem_inst__abc_19396_new_n1675_));
OAI21X1 OAI21X1_977 ( .A(w_mem_inst__abc_19396_new_n1676_), .B(w_mem_inst__abc_19396_new_n1611__bF_buf2), .C(w_mem_inst__abc_19396_new_n1677_), .Y(w_mem_inst__abc_19396_new_n1678_));
OAI21X1 OAI21X1_978 ( .A(w_mem_inst__abc_19396_new_n1696_), .B(w_mem_inst__abc_19396_new_n1598__bF_buf1), .C(w_mem_inst__abc_19396_new_n1586__bF_buf0), .Y(w_mem_inst__abc_19396_new_n1697_));
OAI21X1 OAI21X1_979 ( .A(w_mem_inst__abc_19396_new_n1698_), .B(w_mem_inst__abc_19396_new_n1604__bF_buf1), .C(w_mem_inst__abc_19396_new_n1699_), .Y(w_mem_inst__abc_19396_new_n1700_));
OAI21X1 OAI21X1_98 ( .A(_abc_15497_new_n871__bF_buf2), .B(_abc_15497_new_n872__bF_buf2), .C(_auto_iopadmap_cc_368_execute_22625_29_), .Y(_abc_15497_new_n1269_));
OAI21X1 OAI21X1_980 ( .A(w_mem_inst__abc_19396_new_n1701_), .B(w_mem_inst__abc_19396_new_n1611__bF_buf1), .C(w_mem_inst__abc_19396_new_n1702_), .Y(w_mem_inst__abc_19396_new_n1703_));
OAI21X1 OAI21X1_981 ( .A(w_mem_inst__abc_19396_new_n1721_), .B(w_mem_inst__abc_19396_new_n1598__bF_buf0), .C(w_mem_inst__abc_19396_new_n1586__bF_buf4), .Y(w_mem_inst__abc_19396_new_n1722_));
OAI21X1 OAI21X1_982 ( .A(w_mem_inst__abc_19396_new_n1723_), .B(w_mem_inst__abc_19396_new_n1604__bF_buf0), .C(w_mem_inst__abc_19396_new_n1724_), .Y(w_mem_inst__abc_19396_new_n1725_));
OAI21X1 OAI21X1_983 ( .A(w_mem_inst__abc_19396_new_n1726_), .B(w_mem_inst__abc_19396_new_n1611__bF_buf0), .C(w_mem_inst__abc_19396_new_n1727_), .Y(w_mem_inst__abc_19396_new_n1728_));
OAI21X1 OAI21X1_984 ( .A(w_mem_inst__abc_19396_new_n1746_), .B(w_mem_inst__abc_19396_new_n1598__bF_buf4), .C(w_mem_inst__abc_19396_new_n1586__bF_buf3), .Y(w_mem_inst__abc_19396_new_n1747_));
OAI21X1 OAI21X1_985 ( .A(w_mem_inst__abc_19396_new_n1748_), .B(w_mem_inst__abc_19396_new_n1604__bF_buf4), .C(w_mem_inst__abc_19396_new_n1749_), .Y(w_mem_inst__abc_19396_new_n1750_));
OAI21X1 OAI21X1_986 ( .A(w_mem_inst__abc_19396_new_n1751_), .B(w_mem_inst__abc_19396_new_n1611__bF_buf4), .C(w_mem_inst__abc_19396_new_n1752_), .Y(w_mem_inst__abc_19396_new_n1753_));
OAI21X1 OAI21X1_987 ( .A(w_mem_inst__abc_19396_new_n1771_), .B(w_mem_inst__abc_19396_new_n1598__bF_buf3), .C(w_mem_inst__abc_19396_new_n1586__bF_buf2), .Y(w_mem_inst__abc_19396_new_n1772_));
OAI21X1 OAI21X1_988 ( .A(w_mem_inst__abc_19396_new_n1773_), .B(w_mem_inst__abc_19396_new_n1604__bF_buf3), .C(w_mem_inst__abc_19396_new_n1774_), .Y(w_mem_inst__abc_19396_new_n1775_));
OAI21X1 OAI21X1_989 ( .A(w_mem_inst__abc_19396_new_n1776_), .B(w_mem_inst__abc_19396_new_n1611__bF_buf3), .C(w_mem_inst__abc_19396_new_n1777_), .Y(w_mem_inst__abc_19396_new_n1778_));
OAI21X1 OAI21X1_99 ( .A(_abc_15497_new_n1276_), .B(_abc_15497_new_n1271_), .C(digest_update_bF_buf7), .Y(_abc_15497_new_n1277_));
OAI21X1 OAI21X1_990 ( .A(w_mem_inst__abc_19396_new_n1796_), .B(w_mem_inst__abc_19396_new_n1598__bF_buf2), .C(w_mem_inst__abc_19396_new_n1586__bF_buf1), .Y(w_mem_inst__abc_19396_new_n1797_));
OAI21X1 OAI21X1_991 ( .A(w_mem_inst__abc_19396_new_n1798_), .B(w_mem_inst__abc_19396_new_n1604__bF_buf2), .C(w_mem_inst__abc_19396_new_n1799_), .Y(w_mem_inst__abc_19396_new_n1800_));
OAI21X1 OAI21X1_992 ( .A(w_mem_inst__abc_19396_new_n1801_), .B(w_mem_inst__abc_19396_new_n1611__bF_buf2), .C(w_mem_inst__abc_19396_new_n1802_), .Y(w_mem_inst__abc_19396_new_n1803_));
OAI21X1 OAI21X1_993 ( .A(w_mem_inst__abc_19396_new_n1821_), .B(w_mem_inst__abc_19396_new_n1598__bF_buf1), .C(w_mem_inst__abc_19396_new_n1586__bF_buf0), .Y(w_mem_inst__abc_19396_new_n1822_));
OAI21X1 OAI21X1_994 ( .A(w_mem_inst__abc_19396_new_n1823_), .B(w_mem_inst__abc_19396_new_n1604__bF_buf1), .C(w_mem_inst__abc_19396_new_n1824_), .Y(w_mem_inst__abc_19396_new_n1825_));
OAI21X1 OAI21X1_995 ( .A(w_mem_inst__abc_19396_new_n1826_), .B(w_mem_inst__abc_19396_new_n1611__bF_buf1), .C(w_mem_inst__abc_19396_new_n1827_), .Y(w_mem_inst__abc_19396_new_n1828_));
OAI21X1 OAI21X1_996 ( .A(w_mem_inst__abc_19396_new_n1846_), .B(w_mem_inst__abc_19396_new_n1598__bF_buf0), .C(w_mem_inst__abc_19396_new_n1586__bF_buf4), .Y(w_mem_inst__abc_19396_new_n1847_));
OAI21X1 OAI21X1_997 ( .A(w_mem_inst__abc_19396_new_n1848_), .B(w_mem_inst__abc_19396_new_n1604__bF_buf0), .C(w_mem_inst__abc_19396_new_n1849_), .Y(w_mem_inst__abc_19396_new_n1850_));
OAI21X1 OAI21X1_998 ( .A(w_mem_inst__abc_19396_new_n1851_), .B(w_mem_inst__abc_19396_new_n1611__bF_buf0), .C(w_mem_inst__abc_19396_new_n1852_), .Y(w_mem_inst__abc_19396_new_n1853_));
OAI21X1 OAI21X1_999 ( .A(w_mem_inst__abc_19396_new_n1871_), .B(w_mem_inst__abc_19396_new_n1598__bF_buf4), .C(w_mem_inst__abc_19396_new_n1586__bF_buf3), .Y(w_mem_inst__abc_19396_new_n1872_));
OAI22X1 OAI22X1_1 ( .A(_abc_15497_new_n698_), .B(_abc_15497_new_n873__bF_buf7), .C(_abc_15497_new_n869_), .D(_abc_15497_new_n875_), .Y(_0H2_reg_31_0__26_));
OAI22X1 OAI22X1_10 ( .A(_abc_15497_new_n1057_), .B(_abc_15497_new_n873__bF_buf5), .C(_abc_15497_new_n1067_), .D(_abc_15497_new_n1069_), .Y(_0H4_reg_31_0__12_));
OAI22X1 OAI22X1_11 ( .A(_abc_15497_new_n1101_), .B(_abc_15497_new_n873__bF_buf4), .C(_abc_15497_new_n1115_), .D(_abc_15497_new_n1117_), .Y(_0H4_reg_31_0__16_));
OAI22X1 OAI22X1_12 ( .A(_abc_15497_new_n1128_), .B(_abc_15497_new_n873__bF_buf3), .C(_abc_15497_new_n1139_), .D(_abc_15497_new_n1140_), .Y(_0H4_reg_31_0__18_));
OAI22X1 OAI22X1_13 ( .A(_abc_15497_new_n1142_), .B(_abc_15497_new_n873__bF_buf2), .C(_abc_15497_new_n870__bF_buf10), .D(_abc_15497_new_n1149_), .Y(_0H4_reg_31_0__19_));
OAI22X1 OAI22X1_14 ( .A(_abc_15497_new_n1171_), .B(_abc_15497_new_n873__bF_buf1), .C(_abc_15497_new_n870__bF_buf8), .D(_abc_15497_new_n1177_), .Y(_0H4_reg_31_0__21_));
OAI22X1 OAI22X1_15 ( .A(_abc_15497_new_n1231_), .B(_abc_15497_new_n873__bF_buf0), .C(_abc_15497_new_n1242_), .D(_abc_15497_new_n1245_), .Y(_0H4_reg_31_0__26_));
OAI22X1 OAI22X1_16 ( .A(_abc_15497_new_n1247_), .B(_abc_15497_new_n873__bF_buf7), .C(_abc_15497_new_n870__bF_buf1), .D(_abc_15497_new_n1256_), .Y(_0H4_reg_31_0__27_));
OAI22X1 OAI22X1_17 ( .A(_abc_15497_new_n1258_), .B(_abc_15497_new_n873__bF_buf6), .C(_abc_15497_new_n1267_), .D(_abc_15497_new_n1265_), .Y(_0H4_reg_31_0__28_));
OAI22X1 OAI22X1_18 ( .A(_abc_15497_new_n1300_), .B(_abc_15497_new_n1301_), .C(_abc_15497_new_n1298_), .D(_abc_15497_new_n873__bF_buf5), .Y(_0H3_reg_31_0__0_));
OAI22X1 OAI22X1_19 ( .A(_abc_15497_new_n1317_), .B(_abc_15497_new_n873__bF_buf4), .C(_abc_15497_new_n1323_), .D(_abc_15497_new_n1324_), .Y(_0H3_reg_31_0__3_));
OAI22X1 OAI22X1_2 ( .A(_abc_15497_new_n901_), .B(_abc_15497_new_n873__bF_buf6), .C(_abc_15497_new_n908_), .D(_abc_15497_new_n909_), .Y(_0H2_reg_31_0__29_));
OAI22X1 OAI22X1_20 ( .A(_abc_15497_new_n1351_), .B(_abc_15497_new_n873__bF_buf3), .C(_abc_15497_new_n870__bF_buf7), .D(_abc_15497_new_n1359_), .Y(_0H3_reg_31_0__7_));
OAI22X1 OAI22X1_21 ( .A(_abc_15497_new_n1361_), .B(_abc_15497_new_n873__bF_buf2), .C(_abc_15497_new_n1368_), .D(_abc_15497_new_n1369_), .Y(_0H3_reg_31_0__8_));
OAI22X1 OAI22X1_22 ( .A(_abc_15497_new_n1371_), .B(_abc_15497_new_n873__bF_buf1), .C(_abc_15497_new_n870__bF_buf6), .D(_abc_15497_new_n1380_), .Y(_0H3_reg_31_0__9_));
OAI22X1 OAI22X1_23 ( .A(_abc_15497_new_n1395_), .B(_abc_15497_new_n873__bF_buf0), .C(_abc_15497_new_n1402_), .D(_abc_15497_new_n1403_), .Y(_0H3_reg_31_0__11_));
OAI22X1 OAI22X1_24 ( .A(_abc_15497_new_n1422_), .B(_abc_15497_new_n873__bF_buf7), .C(_abc_15497_new_n870__bF_buf2), .D(_abc_15497_new_n1430_), .Y(_0H3_reg_31_0__13_));
OAI22X1 OAI22X1_25 ( .A(_abc_15497_new_n1444_), .B(_abc_15497_new_n873__bF_buf6), .C(_abc_15497_new_n870__bF_buf0), .D(_abc_15497_new_n1450_), .Y(_0H3_reg_31_0__15_));
OAI22X1 OAI22X1_26 ( .A(_abc_15497_new_n1452_), .B(_abc_15497_new_n873__bF_buf5), .C(_abc_15497_new_n870__bF_buf11), .D(_abc_15497_new_n1465_), .Y(_0H3_reg_31_0__16_));
OAI22X1 OAI22X1_27 ( .A(_abc_15497_new_n1477_), .B(_abc_15497_new_n873__bF_buf4), .C(_abc_15497_new_n1490_), .D(_abc_15497_new_n1488_), .Y(_0H3_reg_31_0__18_));
OAI22X1 OAI22X1_28 ( .A(_abc_15497_new_n1492_), .B(_abc_15497_new_n873__bF_buf3), .C(_abc_15497_new_n1499_), .D(_abc_15497_new_n1500_), .Y(_0H3_reg_31_0__19_));
OAI22X1 OAI22X1_29 ( .A(_abc_15497_new_n1528_), .B(_abc_15497_new_n873__bF_buf2), .C(_abc_15497_new_n1537_), .D(_abc_15497_new_n1538_), .Y(_0H3_reg_31_0__22_));
OAI22X1 OAI22X1_3 ( .A(_abc_15497_new_n911_), .B(_abc_15497_new_n873__bF_buf5), .C(_abc_15497_new_n920_), .D(_abc_15497_new_n923_), .Y(_0H2_reg_31_0__30_));
OAI22X1 OAI22X1_30 ( .A(_abc_15497_new_n1540_), .B(_abc_15497_new_n873__bF_buf1), .C(_abc_15497_new_n1547_), .D(_abc_15497_new_n1548_), .Y(_0H3_reg_31_0__23_));
OAI22X1 OAI22X1_31 ( .A(_abc_15497_new_n1550_), .B(_abc_15497_new_n873__bF_buf0), .C(_abc_15497_new_n1567_), .D(_abc_15497_new_n1565_), .Y(_0H3_reg_31_0__24_));
OAI22X1 OAI22X1_32 ( .A(_abc_15497_new_n1569_), .B(_abc_15497_new_n873__bF_buf7), .C(_abc_15497_new_n870__bF_buf6), .D(_abc_15497_new_n1578_), .Y(_0H3_reg_31_0__25_));
OAI22X1 OAI22X1_33 ( .A(_abc_15497_new_n1580_), .B(_abc_15497_new_n873__bF_buf6), .C(_abc_15497_new_n1590_), .D(_abc_15497_new_n1591_), .Y(_0H3_reg_31_0__26_));
OAI22X1 OAI22X1_34 ( .A(_abc_15497_new_n1593_), .B(_abc_15497_new_n873__bF_buf5), .C(_abc_15497_new_n870__bF_buf5), .D(_abc_15497_new_n1602_), .Y(_0H3_reg_31_0__27_));
OAI22X1 OAI22X1_35 ( .A(_abc_15497_new_n1628_), .B(_abc_15497_new_n873__bF_buf4), .C(_abc_15497_new_n870__bF_buf2), .D(_abc_15497_new_n1635_), .Y(_0H3_reg_31_0__30_));
OAI22X1 OAI22X1_36 ( .A(_abc_15497_new_n1637_), .B(_abc_15497_new_n873__bF_buf3), .C(_abc_15497_new_n1641_), .D(_abc_15497_new_n1642_), .Y(_0H3_reg_31_0__31_));
OAI22X1 OAI22X1_37 ( .A(_abc_15497_new_n1762_), .B(_abc_15497_new_n873__bF_buf1), .C(_abc_15497_new_n1769_), .D(_abc_15497_new_n1768_), .Y(_0H1_reg_31_0__2_));
OAI22X1 OAI22X1_38 ( .A(_abc_15497_new_n1779_), .B(_abc_15497_new_n873__bF_buf0), .C(_abc_15497_new_n1783_), .D(_abc_15497_new_n1785_), .Y(_0H1_reg_31_0__4_));
OAI22X1 OAI22X1_39 ( .A(_abc_15497_new_n1787_), .B(_abc_15497_new_n873__bF_buf7), .C(_abc_15497_new_n870__bF_buf9), .D(_abc_15497_new_n1797_), .Y(_0H1_reg_31_0__5_));
OAI22X1 OAI22X1_4 ( .A(_abc_15497_new_n938_), .B(_abc_15497_new_n939_), .C(_abc_15497_new_n936_), .D(_abc_15497_new_n873__bF_buf4), .Y(_0H4_reg_31_0__0_));
OAI22X1 OAI22X1_40 ( .A(_abc_15497_new_n1799_), .B(_abc_15497_new_n873__bF_buf6), .C(_abc_15497_new_n870__bF_buf8), .D(_abc_15497_new_n1805_), .Y(_0H1_reg_31_0__6_));
OAI22X1 OAI22X1_41 ( .A(_abc_15497_new_n1836_), .B(_abc_15497_new_n873__bF_buf5), .C(_abc_15497_new_n1844_), .D(_abc_15497_new_n1846_), .Y(_0H1_reg_31_0__10_));
OAI22X1 OAI22X1_42 ( .A(_abc_15497_new_n1856_), .B(_abc_15497_new_n873__bF_buf4), .C(_abc_15497_new_n870__bF_buf0), .D(_abc_15497_new_n1866_), .Y(_0H1_reg_31_0__12_));
OAI22X1 OAI22X1_43 ( .A(_abc_15497_new_n1874_), .B(_abc_15497_new_n873__bF_buf3), .C(_abc_15497_new_n1887_), .D(_abc_15497_new_n1888_), .Y(_0H1_reg_31_0__14_));
OAI22X1 OAI22X1_44 ( .A(_abc_15497_new_n1916_), .B(_abc_15497_new_n873__bF_buf2), .C(_abc_15497_new_n870__bF_buf6), .D(_abc_15497_new_n1922_), .Y(_0H1_reg_31_0__17_));
OAI22X1 OAI22X1_45 ( .A(_abc_15497_new_n1949_), .B(_abc_15497_new_n873__bF_buf1), .C(_abc_15497_new_n1962_), .D(_abc_15497_new_n1963_), .Y(_0H1_reg_31_0__20_));
OAI22X1 OAI22X1_46 ( .A(_abc_15497_new_n1965_), .B(_abc_15497_new_n873__bF_buf0), .C(_abc_15497_new_n870__bF_buf3), .D(_abc_15497_new_n1972_), .Y(_0H1_reg_31_0__21_));
OAI22X1 OAI22X1_47 ( .A(_abc_15497_new_n2047_), .B(_abc_15497_new_n873__bF_buf7), .C(_abc_15497_new_n2057_), .D(_abc_15497_new_n2060_), .Y(_0H1_reg_31_0__28_));
OAI22X1 OAI22X1_48 ( .A(_abc_15497_new_n2103_), .B(_abc_15497_new_n873__bF_buf5), .C(_abc_15497_new_n2110_), .D(_abc_15497_new_n2109_), .Y(_0H0_reg_31_0__2_));
OAI22X1 OAI22X1_49 ( .A(_abc_15497_new_n2112_), .B(_abc_15497_new_n873__bF_buf4), .C(_abc_15497_new_n870__bF_buf9), .D(_abc_15497_new_n2120_), .Y(_0H0_reg_31_0__3_));
OAI22X1 OAI22X1_5 ( .A(_abc_15497_new_n946_), .B(_abc_15497_new_n873__bF_buf2), .C(_abc_15497_new_n953_), .D(_abc_15497_new_n952_), .Y(_0H4_reg_31_0__2_));
OAI22X1 OAI22X1_50 ( .A(_abc_15497_new_n2122_), .B(_abc_15497_new_n873__bF_buf3), .C(_abc_15497_new_n2125_), .D(_abc_15497_new_n2127_), .Y(_0H0_reg_31_0__4_));
OAI22X1 OAI22X1_51 ( .A(_abc_15497_new_n2129_), .B(_abc_15497_new_n873__bF_buf2), .C(_abc_15497_new_n870__bF_buf8), .D(_abc_15497_new_n2139_), .Y(_0H0_reg_31_0__5_));
OAI22X1 OAI22X1_52 ( .A(_abc_15497_new_n2141_), .B(_abc_15497_new_n873__bF_buf1), .C(_abc_15497_new_n2147_), .D(_abc_15497_new_n2149_), .Y(_0H0_reg_31_0__6_));
OAI22X1 OAI22X1_53 ( .A(_abc_15497_new_n2151_), .B(_abc_15497_new_n873__bF_buf0), .C(_abc_15497_new_n2154_), .D(_abc_15497_new_n2157_), .Y(_0H0_reg_31_0__7_));
OAI22X1 OAI22X1_54 ( .A(_abc_15497_new_n2180_), .B(_abc_15497_new_n873__bF_buf7), .C(_abc_15497_new_n2194_), .D(_abc_15497_new_n2195_), .Y(_0H0_reg_31_0__10_));
OAI22X1 OAI22X1_55 ( .A(_abc_15497_new_n2197_), .B(_abc_15497_new_n873__bF_buf6), .C(_abc_15497_new_n870__bF_buf3), .D(_abc_15497_new_n2201_), .Y(_0H0_reg_31_0__11_));
OAI22X1 OAI22X1_56 ( .A(_abc_15497_new_n2203_), .B(_abc_15497_new_n873__bF_buf5), .C(_abc_15497_new_n2217_), .D(_abc_15497_new_n2219_), .Y(_0H0_reg_31_0__12_));
OAI22X1 OAI22X1_57 ( .A(_abc_15497_new_n2228_), .B(_abc_15497_new_n873__bF_buf4), .C(_abc_15497_new_n2237_), .D(_abc_15497_new_n2239_), .Y(_0H0_reg_31_0__14_));
OAI22X1 OAI22X1_58 ( .A(_abc_15497_new_n2241_), .B(_abc_15497_new_n873__bF_buf3), .C(_abc_15497_new_n870__bF_buf0), .D(_abc_15497_new_n2247_), .Y(_0H0_reg_31_0__15_));
OAI22X1 OAI22X1_59 ( .A(_abc_15497_new_n2267_), .B(_abc_15497_new_n873__bF_buf2), .C(_abc_15497_new_n870__bF_buf10), .D(_abc_15497_new_n2276_), .Y(_0H0_reg_31_0__17_));
OAI22X1 OAI22X1_6 ( .A(_abc_15497_new_n955_), .B(_abc_15497_new_n873__bF_buf1), .C(_abc_15497_new_n870__bF_buf3), .D(_abc_15497_new_n964_), .Y(_0H4_reg_31_0__3_));
OAI22X1 OAI22X1_60 ( .A(_abc_15497_new_n2293_), .B(_abc_15497_new_n873__bF_buf1), .C(_abc_15497_new_n2300_), .D(_abc_15497_new_n2301_), .Y(_0H0_reg_31_0__19_));
OAI22X1 OAI22X1_61 ( .A(_abc_15497_new_n2303_), .B(_abc_15497_new_n873__bF_buf0), .C(_abc_15497_new_n2314_), .D(_abc_15497_new_n2315_), .Y(_0H0_reg_31_0__20_));
OAI22X1 OAI22X1_62 ( .A(_abc_15497_new_n2317_), .B(_abc_15497_new_n873__bF_buf7), .C(_abc_15497_new_n870__bF_buf8), .D(_abc_15497_new_n2326_), .Y(_0H0_reg_31_0__21_));
OAI22X1 OAI22X1_63 ( .A(_abc_15497_new_n2393_), .B(_abc_15497_new_n873__bF_buf5), .C(_abc_15497_new_n870__bF_buf1), .D(_abc_15497_new_n2399_), .Y(_0H0_reg_31_0__27_));
OAI22X1 OAI22X1_64 ( .A(_abc_15497_new_n2401_), .B(_abc_15497_new_n873__bF_buf4), .C(_abc_15497_new_n2410_), .D(_abc_15497_new_n2412_), .Y(_0H0_reg_31_0__28_));
OAI22X1 OAI22X1_65 ( .A(_abc_15497_new_n2438_), .B(_abc_15497_new_n873__bF_buf3), .C(_abc_15497_new_n2441_), .D(_abc_15497_new_n2442_), .Y(_0H0_reg_31_0__31_));
OAI22X1 OAI22X1_66 ( .A(_abc_15497_new_n2742__bF_buf0), .B(_abc_15497_new_n2978_), .C(_abc_15497_new_n2924__bF_buf3), .D(_abc_15497_new_n2977_), .Y(_abc_15497_new_n2979_));
OAI22X1 OAI22X1_67 ( .A(_abc_15497_new_n2742__bF_buf3), .B(_abc_15497_new_n3127_), .C(_abc_15497_new_n2924__bF_buf2), .D(_abc_15497_new_n3125_), .Y(_abc_15497_new_n3128_));
OAI22X1 OAI22X1_68 ( .A(_abc_15497_new_n2742__bF_buf2), .B(_abc_15497_new_n3239_), .C(_abc_15497_new_n3234_), .D(_abc_15497_new_n2924__bF_buf4), .Y(_abc_15497_new_n3240_));
OAI22X1 OAI22X1_69 ( .A(_abc_15497_new_n3252_), .B(_abc_15497_new_n3250_), .C(_abc_15497_new_n3240_), .D(_abc_15497_new_n3238_), .Y(_abc_15497_new_n3253_));
OAI22X1 OAI22X1_7 ( .A(_abc_15497_new_n1024_), .B(_abc_15497_new_n873__bF_buf0), .C(_abc_15497_new_n1028_), .D(_abc_15497_new_n1031_), .Y(_0H4_reg_31_0__9_));
OAI22X1 OAI22X1_70 ( .A(_abc_15497_new_n2742__bF_buf1), .B(_abc_15497_new_n3316_), .C(_abc_15497_new_n2924__bF_buf3), .D(_abc_15497_new_n3315_), .Y(_abc_15497_new_n3317_));
OAI22X1 OAI22X1_71 ( .A(_abc_15497_new_n2742__bF_buf3), .B(_abc_15497_new_n3412_), .C(_abc_15497_new_n2924__bF_buf4), .D(_abc_15497_new_n3411_), .Y(_abc_15497_new_n3413_));
OAI22X1 OAI22X1_72 ( .A(_abc_15497_new_n2742__bF_buf2), .B(_abc_15497_new_n3446_), .C(_abc_15497_new_n3445_), .D(_abc_15497_new_n2924__bF_buf3), .Y(_abc_15497_new_n3447_));
OAI22X1 OAI22X1_73 ( .A(_abc_15497_new_n2742__bF_buf1), .B(_abc_15497_new_n3491_), .C(_abc_15497_new_n3489_), .D(_abc_15497_new_n2924__bF_buf2), .Y(_abc_15497_new_n3492_));
OAI22X1 OAI22X1_74 ( .A(_abc_15497_new_n3502_), .B(_abc_15497_new_n3504_), .C(_abc_15497_new_n3492_), .D(_abc_15497_new_n3488_), .Y(_abc_15497_new_n3505_));
OAI22X1 OAI22X1_75 ( .A(_abc_15497_new_n2742__bF_buf0), .B(_abc_15497_new_n3555_), .C(_abc_15497_new_n2924__bF_buf1), .D(_abc_15497_new_n3553_), .Y(_abc_15497_new_n3556_));
OAI22X1 OAI22X1_76 ( .A(_abc_15497_new_n3873_), .B(_abc_15497_new_n3870_), .C(_abc_15497_new_n3874_), .D(_abc_15497_new_n3875_), .Y(_abc_15497_new_n3876_));
OAI22X1 OAI22X1_77 ( .A(_abc_15497_new_n2924__bF_buf4), .B(_abc_15497_new_n4423_), .C(_abc_15497_new_n2925__bF_buf1), .D(_abc_15497_new_n4421_), .Y(_abc_15497_new_n4424_));
OAI22X1 OAI22X1_78 ( .A(_abc_15497_new_n770_), .B(_abc_15497_new_n873__bF_buf2), .C(_abc_15497_new_n4476_), .D(_abc_15497_new_n4477_), .Y(_0H2_reg_31_0__0_));
OAI22X1 OAI22X1_79 ( .A(_abc_15497_new_n742_), .B(_abc_15497_new_n873__bF_buf1), .C(_abc_15497_new_n4512_), .D(_abc_15497_new_n4513_), .Y(_0H2_reg_31_0__8_));
OAI22X1 OAI22X1_8 ( .A(_abc_15497_new_n1033_), .B(_abc_15497_new_n873__bF_buf7), .C(_abc_15497_new_n1044_), .D(_abc_15497_new_n1046_), .Y(_0H4_reg_31_0__10_));
OAI22X1 OAI22X1_80 ( .A(_abc_15497_new_n739_), .B(_abc_15497_new_n873__bF_buf0), .C(_abc_15497_new_n4516_), .D(_abc_15497_new_n4517_), .Y(_0H2_reg_31_0__9_));
OAI22X1 OAI22X1_81 ( .A(_abc_15497_new_n709_), .B(_abc_15497_new_n873__bF_buf7), .C(_abc_15497_new_n4536_), .D(_abc_15497_new_n4537_), .Y(_0H2_reg_31_0__13_));
OAI22X1 OAI22X1_82 ( .A(_abc_15497_new_n833_), .B(_abc_15497_new_n873__bF_buf6), .C(_abc_15497_new_n4551_), .D(_abc_15497_new_n4549_), .Y(_0H2_reg_31_0__16_));
OAI22X1 OAI22X1_83 ( .A(_abc_15497_new_n824_), .B(_abc_15497_new_n873__bF_buf5), .C(_abc_15497_new_n870__bF_buf2), .D(_abc_15497_new_n4558_), .Y(_0H2_reg_31_0__18_));
OAI22X1 OAI22X1_84 ( .A(_abc_15497_new_n799_), .B(_abc_15497_new_n873__bF_buf4), .C(_abc_15497_new_n4578_), .D(_abc_15497_new_n4580_), .Y(_0H2_reg_31_0__22_));
OAI22X1 OAI22X1_85 ( .A(_abc_15497_new_n856_), .B(_abc_15497_new_n873__bF_buf3), .C(_abc_15497_new_n4588_), .D(_abc_15497_new_n4589_), .Y(_0H2_reg_31_0__24_));
OAI22X1 OAI22X1_86 ( .A(_abc_15497_new_n850_), .B(_abc_15497_new_n873__bF_buf2), .C(_abc_15497_new_n4593_), .D(_abc_15497_new_n4594_), .Y(_0H2_reg_31_0__25_));
OAI22X1 OAI22X1_9 ( .A(_abc_15497_new_n1048_), .B(_abc_15497_new_n873__bF_buf6), .C(_abc_15497_new_n870__bF_buf6), .D(_abc_15497_new_n1055_), .Y(_0H4_reg_31_0__11_));
OR2X2 OR2X2_1 ( .A(e_reg_4_), .B(_auto_iopadmap_cc_368_execute_22625_4_), .Y(_abc_15497_new_n966_));
OR2X2 OR2X2_10 ( .A(_abc_15497_new_n2063_), .B(_abc_15497_new_n2068_), .Y(_abc_15497_new_n2069_));
OR2X2 OR2X2_11 ( .A(_abc_15497_new_n2076_), .B(_abc_15497_new_n2073_), .Y(_abc_15497_new_n2078_));
OR2X2 OR2X2_12 ( .A(_abc_15497_new_n873__bF_buf6), .B(_abc_15497_new_n2341_), .Y(_abc_15497_new_n2342_));
OR2X2 OR2X2_13 ( .A(_abc_15497_new_n2783_), .B(_abc_15497_new_n1308_), .Y(_abc_15497_new_n2785_));
OR2X2 OR2X2_14 ( .A(_abc_15497_new_n2831_), .B(_abc_15497_new_n2829_), .Y(_abc_15497_new_n2833_));
OR2X2 OR2X2_15 ( .A(_abc_15497_new_n2904_), .B(_abc_15497_new_n2903_), .Y(_abc_15497_new_n2905_));
OR2X2 OR2X2_16 ( .A(_abc_15497_new_n3009_), .B(_abc_15497_new_n1343_), .Y(_abc_15497_new_n3011_));
OR2X2 OR2X2_17 ( .A(_abc_15497_new_n3067_), .B(_abc_15497_new_n1357_), .Y(_abc_15497_new_n3069_));
OR2X2 OR2X2_18 ( .A(_abc_15497_new_n3171_), .B(_abc_15497_new_n1364_), .Y(_abc_15497_new_n3173_));
OR2X2 OR2X2_19 ( .A(_abc_15497_new_n3186_), .B(_abc_15497_new_n3178_), .Y(_abc_15497_new_n3187_));
OR2X2 OR2X2_2 ( .A(_abc_15497_new_n978_), .B(_abc_15497_new_n977_), .Y(_abc_15497_new_n979_));
OR2X2 OR2X2_20 ( .A(_abc_15497_new_n3292_), .B(_abc_15497_new_n3290_), .Y(_abc_15497_new_n3294_));
OR2X2 OR2X2_21 ( .A(e_reg_13_), .B(a_reg_8_), .Y(_abc_15497_new_n3498_));
OR2X2 OR2X2_22 ( .A(_abc_15497_new_n3530_), .B(_abc_15497_new_n3533_), .Y(_0a_reg_31_0__13_));
OR2X2 OR2X2_23 ( .A(_abc_15497_new_n3603_), .B(_abc_15497_new_n3541_), .Y(_abc_15497_new_n3604_));
OR2X2 OR2X2_24 ( .A(e_reg_15_), .B(a_reg_10_), .Y(_abc_15497_new_n3627_));
OR2X2 OR2X2_25 ( .A(_abc_15497_new_n3693_), .B(_abc_15497_new_n3692_), .Y(_abc_15497_new_n3695_));
OR2X2 OR2X2_26 ( .A(_abc_15497_new_n3798_), .B(_abc_15497_new_n3797_), .Y(_abc_15497_new_n3800_));
OR2X2 OR2X2_27 ( .A(_abc_15497_new_n3789_), .B(_abc_15497_new_n3794_), .Y(_abc_15497_new_n3804_));
OR2X2 OR2X2_28 ( .A(_abc_15497_new_n3805_), .B(_abc_15497_new_n3796_), .Y(_abc_15497_new_n3807_));
OR2X2 OR2X2_29 ( .A(_abc_15497_new_n3842_), .B(_abc_15497_new_n3841_), .Y(_abc_15497_new_n3844_));
OR2X2 OR2X2_3 ( .A(_abc_15497_new_n1017_), .B(_abc_15497_new_n1026_), .Y(_abc_15497_new_n1027_));
OR2X2 OR2X2_30 ( .A(_abc_15497_new_n3832_), .B(_abc_15497_new_n3839_), .Y(_abc_15497_new_n3887_));
OR2X2 OR2X2_31 ( .A(_abc_15497_new_n3905_), .B(_abc_15497_new_n3904_), .Y(_abc_15497_new_n3907_));
OR2X2 OR2X2_32 ( .A(_abc_15497_new_n3956_), .B(_abc_15497_new_n3955_), .Y(_abc_15497_new_n3958_));
OR2X2 OR2X2_33 ( .A(_abc_15497_new_n4011_), .B(_abc_15497_new_n4010_), .Y(_abc_15497_new_n4013_));
OR2X2 OR2X2_34 ( .A(_abc_15497_new_n4065_), .B(_abc_15497_new_n4064_), .Y(_abc_15497_new_n4067_));
OR2X2 OR2X2_35 ( .A(_abc_15497_new_n4071_), .B(_abc_15497_new_n4059_), .Y(_abc_15497_new_n4072_));
OR2X2 OR2X2_36 ( .A(_abc_15497_new_n4071_), .B(_abc_15497_new_n4058_), .Y(_abc_15497_new_n4078_));
OR2X2 OR2X2_37 ( .A(_abc_15497_new_n4168_), .B(_abc_15497_new_n4163_), .Y(_abc_15497_new_n4169_));
OR2X2 OR2X2_38 ( .A(_abc_15497_new_n4176_), .B(_abc_15497_new_n4151_), .Y(_abc_15497_new_n4177_));
OR2X2 OR2X2_39 ( .A(_abc_15497_new_n4253_), .B(_abc_15497_new_n4252_), .Y(_abc_15497_new_n4254_));
OR2X2 OR2X2_4 ( .A(_abc_15497_new_n1041_), .B(_abc_15497_new_n1039_), .Y(_abc_15497_new_n1042_));
OR2X2 OR2X2_40 ( .A(_abc_15497_new_n4255_), .B(_abc_15497_new_n4250_), .Y(_abc_15497_new_n4256_));
OR2X2 OR2X2_41 ( .A(_abc_15497_new_n4291_), .B(_abc_15497_new_n4295_), .Y(_abc_15497_new_n4296_));
OR2X2 OR2X2_42 ( .A(_abc_15497_new_n4349_), .B(_abc_15497_new_n4342_), .Y(_abc_15497_new_n4350_));
OR2X2 OR2X2_43 ( .A(_abc_15497_new_n4353_), .B(_abc_15497_new_n2944_), .Y(_abc_15497_new_n4355_));
OR2X2 OR2X2_44 ( .A(_abc_15497_new_n4356_), .B(_abc_15497_new_n4327_), .Y(_abc_15497_new_n4358_));
OR2X2 OR2X2_45 ( .A(_abc_15497_new_n4390_), .B(w_30_), .Y(_abc_15497_new_n4391_));
OR2X2 OR2X2_46 ( .A(_abc_15497_new_n4395_), .B(_abc_15497_new_n4384_), .Y(_abc_15497_new_n4396_));
OR2X2 OR2X2_47 ( .A(_abc_15497_new_n4459_), .B(_abc_15497_new_n1646_), .Y(_abc_15497_new_n4463_));
OR2X2 OR2X2_48 ( .A(_abc_15497_new_n4564_), .B(_abc_15497_new_n837_), .Y(_abc_15497_new_n4565_));
OR2X2 OR2X2_49 ( .A(_abc_15497_new_n4584_), .B(_abc_15497_new_n797_), .Y(_abc_15497_new_n4585_));
OR2X2 OR2X2_5 ( .A(_abc_15497_new_n1260_), .B(_abc_15497_new_n1262_), .Y(_abc_15497_new_n1263_));
OR2X2 OR2X2_50 ( .A(w_mem_inst_w_ctr_reg_4_), .B(w_mem_inst_w_ctr_reg_6_), .Y(w_mem_inst__abc_19396_new_n1585_));
OR2X2 OR2X2_51 ( .A(w_mem_inst_w_ctr_reg_1_), .B(w_mem_inst_w_ctr_reg_0_), .Y(w_mem_inst__abc_19396_new_n1601_));
OR2X2 OR2X2_52 ( .A(w_mem_inst__abc_19396_new_n1603_), .B(w_mem_inst__abc_19396_new_n1601_), .Y(w_mem_inst__abc_19396_new_n1604_));
OR2X2 OR2X2_6 ( .A(_abc_15497_new_n1321_), .B(_abc_15497_new_n1319_), .Y(_abc_15497_new_n1322_));
OR2X2 OR2X2_7 ( .A(_abc_15497_new_n1427_), .B(_abc_15497_new_n1415_), .Y(_abc_15497_new_n1428_));
OR2X2 OR2X2_8 ( .A(_abc_15497_new_n1865_), .B(_abc_15497_new_n1884_), .Y(_abc_15497_new_n1885_));
OR2X2 OR2X2_9 ( .A(_abc_15497_new_n1925_), .B(_abc_15497_new_n1927_), .Y(_abc_15497_new_n1928_));
XNOR2X1 XNOR2X1_1 ( .A(_abc_15497_new_n877_), .B(_abc_15497_new_n881_), .Y(_abc_15497_new_n882_));
XNOR2X1 XNOR2X1_10 ( .A(_abc_15497_new_n1223_), .B(_abc_15497_new_n1227_), .Y(_abc_15497_new_n1228_));
XNOR2X1 XNOR2X1_100 ( .A(w_mem_inst_w_mem_13__2_), .B(w_mem_inst_w_mem_8__2_), .Y(w_mem_inst__abc_19396_new_n1693_));
XNOR2X1 XNOR2X1_101 ( .A(w_mem_inst_w_mem_2__2_), .B(w_mem_inst_w_mem_0__2_), .Y(w_mem_inst__abc_19396_new_n1694_));
XNOR2X1 XNOR2X1_102 ( .A(w_mem_inst__abc_19396_new_n1693_), .B(w_mem_inst__abc_19396_new_n1694_), .Y(w_mem_inst__abc_19396_new_n1695_));
XNOR2X1 XNOR2X1_103 ( .A(w_mem_inst_w_mem_13__3_), .B(w_mem_inst_w_mem_8__3_), .Y(w_mem_inst__abc_19396_new_n1718_));
XNOR2X1 XNOR2X1_104 ( .A(w_mem_inst_w_mem_2__3_), .B(w_mem_inst_w_mem_0__3_), .Y(w_mem_inst__abc_19396_new_n1719_));
XNOR2X1 XNOR2X1_105 ( .A(w_mem_inst__abc_19396_new_n1718_), .B(w_mem_inst__abc_19396_new_n1719_), .Y(w_mem_inst__abc_19396_new_n1720_));
XNOR2X1 XNOR2X1_106 ( .A(w_mem_inst_w_mem_13__4_), .B(w_mem_inst_w_mem_8__4_), .Y(w_mem_inst__abc_19396_new_n1743_));
XNOR2X1 XNOR2X1_107 ( .A(w_mem_inst_w_mem_2__4_), .B(w_mem_inst_w_mem_0__4_), .Y(w_mem_inst__abc_19396_new_n1744_));
XNOR2X1 XNOR2X1_108 ( .A(w_mem_inst__abc_19396_new_n1743_), .B(w_mem_inst__abc_19396_new_n1744_), .Y(w_mem_inst__abc_19396_new_n1745_));
XNOR2X1 XNOR2X1_109 ( .A(w_mem_inst_w_mem_13__5_), .B(w_mem_inst_w_mem_8__5_), .Y(w_mem_inst__abc_19396_new_n1768_));
XNOR2X1 XNOR2X1_11 ( .A(e_reg_31_), .B(_auto_iopadmap_cc_368_execute_22625_31_), .Y(_abc_15497_new_n1292_));
XNOR2X1 XNOR2X1_110 ( .A(w_mem_inst_w_mem_2__5_), .B(w_mem_inst_w_mem_0__5_), .Y(w_mem_inst__abc_19396_new_n1769_));
XNOR2X1 XNOR2X1_111 ( .A(w_mem_inst__abc_19396_new_n1768_), .B(w_mem_inst__abc_19396_new_n1769_), .Y(w_mem_inst__abc_19396_new_n1770_));
XNOR2X1 XNOR2X1_112 ( .A(w_mem_inst_w_mem_13__6_), .B(w_mem_inst_w_mem_8__6_), .Y(w_mem_inst__abc_19396_new_n1793_));
XNOR2X1 XNOR2X1_113 ( .A(w_mem_inst_w_mem_2__6_), .B(w_mem_inst_w_mem_0__6_), .Y(w_mem_inst__abc_19396_new_n1794_));
XNOR2X1 XNOR2X1_114 ( .A(w_mem_inst__abc_19396_new_n1793_), .B(w_mem_inst__abc_19396_new_n1794_), .Y(w_mem_inst__abc_19396_new_n1795_));
XNOR2X1 XNOR2X1_115 ( .A(w_mem_inst_w_mem_13__7_), .B(w_mem_inst_w_mem_8__7_), .Y(w_mem_inst__abc_19396_new_n1818_));
XNOR2X1 XNOR2X1_116 ( .A(w_mem_inst_w_mem_2__7_), .B(w_mem_inst_w_mem_0__7_), .Y(w_mem_inst__abc_19396_new_n1819_));
XNOR2X1 XNOR2X1_117 ( .A(w_mem_inst__abc_19396_new_n1818_), .B(w_mem_inst__abc_19396_new_n1819_), .Y(w_mem_inst__abc_19396_new_n1820_));
XNOR2X1 XNOR2X1_118 ( .A(w_mem_inst_w_mem_13__8_), .B(w_mem_inst_w_mem_8__8_), .Y(w_mem_inst__abc_19396_new_n1843_));
XNOR2X1 XNOR2X1_119 ( .A(w_mem_inst_w_mem_2__8_), .B(w_mem_inst_w_mem_0__8_), .Y(w_mem_inst__abc_19396_new_n1844_));
XNOR2X1 XNOR2X1_12 ( .A(_abc_15497_new_n1303_), .B(_abc_15497_new_n1300_), .Y(_abc_15497_new_n1304_));
XNOR2X1 XNOR2X1_120 ( .A(w_mem_inst__abc_19396_new_n1843_), .B(w_mem_inst__abc_19396_new_n1844_), .Y(w_mem_inst__abc_19396_new_n1845_));
XNOR2X1 XNOR2X1_121 ( .A(w_mem_inst_w_mem_13__9_), .B(w_mem_inst_w_mem_8__9_), .Y(w_mem_inst__abc_19396_new_n1868_));
XNOR2X1 XNOR2X1_122 ( .A(w_mem_inst_w_mem_2__9_), .B(w_mem_inst_w_mem_0__9_), .Y(w_mem_inst__abc_19396_new_n1869_));
XNOR2X1 XNOR2X1_123 ( .A(w_mem_inst__abc_19396_new_n1868_), .B(w_mem_inst__abc_19396_new_n1869_), .Y(w_mem_inst__abc_19396_new_n1870_));
XNOR2X1 XNOR2X1_124 ( .A(w_mem_inst_w_mem_13__10_), .B(w_mem_inst_w_mem_8__10_), .Y(w_mem_inst__abc_19396_new_n1893_));
XNOR2X1 XNOR2X1_125 ( .A(w_mem_inst_w_mem_2__10_), .B(w_mem_inst_w_mem_0__10_), .Y(w_mem_inst__abc_19396_new_n1894_));
XNOR2X1 XNOR2X1_126 ( .A(w_mem_inst__abc_19396_new_n1893_), .B(w_mem_inst__abc_19396_new_n1894_), .Y(w_mem_inst__abc_19396_new_n1895_));
XNOR2X1 XNOR2X1_127 ( .A(w_mem_inst_w_mem_13__11_), .B(w_mem_inst_w_mem_8__11_), .Y(w_mem_inst__abc_19396_new_n1918_));
XNOR2X1 XNOR2X1_128 ( .A(w_mem_inst_w_mem_2__11_), .B(w_mem_inst_w_mem_0__11_), .Y(w_mem_inst__abc_19396_new_n1919_));
XNOR2X1 XNOR2X1_129 ( .A(w_mem_inst__abc_19396_new_n1918_), .B(w_mem_inst__abc_19396_new_n1919_), .Y(w_mem_inst__abc_19396_new_n1920_));
XNOR2X1 XNOR2X1_13 ( .A(_abc_15497_new_n1310_), .B(_abc_15497_new_n1313_), .Y(_abc_15497_new_n1314_));
XNOR2X1 XNOR2X1_130 ( .A(w_mem_inst_w_mem_13__12_), .B(w_mem_inst_w_mem_8__12_), .Y(w_mem_inst__abc_19396_new_n1943_));
XNOR2X1 XNOR2X1_131 ( .A(w_mem_inst_w_mem_2__12_), .B(w_mem_inst_w_mem_0__12_), .Y(w_mem_inst__abc_19396_new_n1944_));
XNOR2X1 XNOR2X1_132 ( .A(w_mem_inst__abc_19396_new_n1943_), .B(w_mem_inst__abc_19396_new_n1944_), .Y(w_mem_inst__abc_19396_new_n1945_));
XNOR2X1 XNOR2X1_133 ( .A(w_mem_inst_w_mem_13__13_), .B(w_mem_inst_w_mem_8__13_), .Y(w_mem_inst__abc_19396_new_n1968_));
XNOR2X1 XNOR2X1_134 ( .A(w_mem_inst_w_mem_2__13_), .B(w_mem_inst_w_mem_0__13_), .Y(w_mem_inst__abc_19396_new_n1969_));
XNOR2X1 XNOR2X1_135 ( .A(w_mem_inst__abc_19396_new_n1968_), .B(w_mem_inst__abc_19396_new_n1969_), .Y(w_mem_inst__abc_19396_new_n1970_));
XNOR2X1 XNOR2X1_136 ( .A(w_mem_inst_w_mem_13__14_), .B(w_mem_inst_w_mem_8__14_), .Y(w_mem_inst__abc_19396_new_n1993_));
XNOR2X1 XNOR2X1_137 ( .A(w_mem_inst_w_mem_2__14_), .B(w_mem_inst_w_mem_0__14_), .Y(w_mem_inst__abc_19396_new_n1994_));
XNOR2X1 XNOR2X1_138 ( .A(w_mem_inst__abc_19396_new_n1993_), .B(w_mem_inst__abc_19396_new_n1994_), .Y(w_mem_inst__abc_19396_new_n1995_));
XNOR2X1 XNOR2X1_139 ( .A(w_mem_inst_w_mem_13__15_), .B(w_mem_inst_w_mem_8__15_), .Y(w_mem_inst__abc_19396_new_n2018_));
XNOR2X1 XNOR2X1_14 ( .A(_abc_15497_new_n1328_), .B(_abc_15497_new_n1326_), .Y(_abc_15497_new_n1329_));
XNOR2X1 XNOR2X1_140 ( .A(w_mem_inst_w_mem_2__15_), .B(w_mem_inst_w_mem_0__15_), .Y(w_mem_inst__abc_19396_new_n2019_));
XNOR2X1 XNOR2X1_141 ( .A(w_mem_inst__abc_19396_new_n2018_), .B(w_mem_inst__abc_19396_new_n2019_), .Y(w_mem_inst__abc_19396_new_n2020_));
XNOR2X1 XNOR2X1_142 ( .A(w_mem_inst_w_mem_13__16_), .B(w_mem_inst_w_mem_8__16_), .Y(w_mem_inst__abc_19396_new_n2043_));
XNOR2X1 XNOR2X1_143 ( .A(w_mem_inst_w_mem_2__16_), .B(w_mem_inst_w_mem_0__16_), .Y(w_mem_inst__abc_19396_new_n2044_));
XNOR2X1 XNOR2X1_144 ( .A(w_mem_inst__abc_19396_new_n2043_), .B(w_mem_inst__abc_19396_new_n2044_), .Y(w_mem_inst__abc_19396_new_n2045_));
XNOR2X1 XNOR2X1_145 ( .A(w_mem_inst_w_mem_13__17_), .B(w_mem_inst_w_mem_8__17_), .Y(w_mem_inst__abc_19396_new_n2068_));
XNOR2X1 XNOR2X1_146 ( .A(w_mem_inst_w_mem_2__17_), .B(w_mem_inst_w_mem_0__17_), .Y(w_mem_inst__abc_19396_new_n2069_));
XNOR2X1 XNOR2X1_147 ( .A(w_mem_inst__abc_19396_new_n2068_), .B(w_mem_inst__abc_19396_new_n2069_), .Y(w_mem_inst__abc_19396_new_n2070_));
XNOR2X1 XNOR2X1_148 ( .A(w_mem_inst_w_mem_13__18_), .B(w_mem_inst_w_mem_8__18_), .Y(w_mem_inst__abc_19396_new_n2093_));
XNOR2X1 XNOR2X1_149 ( .A(w_mem_inst_w_mem_2__18_), .B(w_mem_inst_w_mem_0__18_), .Y(w_mem_inst__abc_19396_new_n2094_));
XNOR2X1 XNOR2X1_15 ( .A(_abc_15497_new_n1358_), .B(_abc_15497_new_n1355_), .Y(_abc_15497_new_n1359_));
XNOR2X1 XNOR2X1_150 ( .A(w_mem_inst__abc_19396_new_n2093_), .B(w_mem_inst__abc_19396_new_n2094_), .Y(w_mem_inst__abc_19396_new_n2095_));
XNOR2X1 XNOR2X1_151 ( .A(w_mem_inst_w_mem_13__19_), .B(w_mem_inst_w_mem_8__19_), .Y(w_mem_inst__abc_19396_new_n2118_));
XNOR2X1 XNOR2X1_152 ( .A(w_mem_inst_w_mem_2__19_), .B(w_mem_inst_w_mem_0__19_), .Y(w_mem_inst__abc_19396_new_n2119_));
XNOR2X1 XNOR2X1_153 ( .A(w_mem_inst__abc_19396_new_n2118_), .B(w_mem_inst__abc_19396_new_n2119_), .Y(w_mem_inst__abc_19396_new_n2120_));
XNOR2X1 XNOR2X1_154 ( .A(w_mem_inst_w_mem_13__20_), .B(w_mem_inst_w_mem_8__20_), .Y(w_mem_inst__abc_19396_new_n2143_));
XNOR2X1 XNOR2X1_155 ( .A(w_mem_inst_w_mem_2__20_), .B(w_mem_inst_w_mem_0__20_), .Y(w_mem_inst__abc_19396_new_n2144_));
XNOR2X1 XNOR2X1_156 ( .A(w_mem_inst__abc_19396_new_n2143_), .B(w_mem_inst__abc_19396_new_n2144_), .Y(w_mem_inst__abc_19396_new_n2145_));
XNOR2X1 XNOR2X1_157 ( .A(w_mem_inst_w_mem_13__21_), .B(w_mem_inst_w_mem_8__21_), .Y(w_mem_inst__abc_19396_new_n2168_));
XNOR2X1 XNOR2X1_158 ( .A(w_mem_inst_w_mem_2__21_), .B(w_mem_inst_w_mem_0__21_), .Y(w_mem_inst__abc_19396_new_n2169_));
XNOR2X1 XNOR2X1_159 ( .A(w_mem_inst__abc_19396_new_n2168_), .B(w_mem_inst__abc_19396_new_n2169_), .Y(w_mem_inst__abc_19396_new_n2170_));
XNOR2X1 XNOR2X1_16 ( .A(_abc_15497_new_n1445_), .B(_abc_15497_new_n1449_), .Y(_abc_15497_new_n1450_));
XNOR2X1 XNOR2X1_160 ( .A(w_mem_inst_w_mem_13__22_), .B(w_mem_inst_w_mem_8__22_), .Y(w_mem_inst__abc_19396_new_n2193_));
XNOR2X1 XNOR2X1_161 ( .A(w_mem_inst_w_mem_2__22_), .B(w_mem_inst_w_mem_0__22_), .Y(w_mem_inst__abc_19396_new_n2194_));
XNOR2X1 XNOR2X1_162 ( .A(w_mem_inst__abc_19396_new_n2193_), .B(w_mem_inst__abc_19396_new_n2194_), .Y(w_mem_inst__abc_19396_new_n2195_));
XNOR2X1 XNOR2X1_163 ( .A(w_mem_inst_w_mem_13__23_), .B(w_mem_inst_w_mem_8__23_), .Y(w_mem_inst__abc_19396_new_n2218_));
XNOR2X1 XNOR2X1_164 ( .A(w_mem_inst_w_mem_2__23_), .B(w_mem_inst_w_mem_0__23_), .Y(w_mem_inst__abc_19396_new_n2219_));
XNOR2X1 XNOR2X1_165 ( .A(w_mem_inst__abc_19396_new_n2218_), .B(w_mem_inst__abc_19396_new_n2219_), .Y(w_mem_inst__abc_19396_new_n2220_));
XNOR2X1 XNOR2X1_166 ( .A(w_mem_inst_w_mem_13__24_), .B(w_mem_inst_w_mem_8__24_), .Y(w_mem_inst__abc_19396_new_n2243_));
XNOR2X1 XNOR2X1_167 ( .A(w_mem_inst_w_mem_2__24_), .B(w_mem_inst_w_mem_0__24_), .Y(w_mem_inst__abc_19396_new_n2244_));
XNOR2X1 XNOR2X1_168 ( .A(w_mem_inst__abc_19396_new_n2243_), .B(w_mem_inst__abc_19396_new_n2244_), .Y(w_mem_inst__abc_19396_new_n2245_));
XNOR2X1 XNOR2X1_169 ( .A(w_mem_inst_w_mem_13__25_), .B(w_mem_inst_w_mem_8__25_), .Y(w_mem_inst__abc_19396_new_n2268_));
XNOR2X1 XNOR2X1_17 ( .A(_abc_15497_new_n1460_), .B(_abc_15497_new_n1464_), .Y(_abc_15497_new_n1465_));
XNOR2X1 XNOR2X1_170 ( .A(w_mem_inst_w_mem_2__25_), .B(w_mem_inst_w_mem_0__25_), .Y(w_mem_inst__abc_19396_new_n2269_));
XNOR2X1 XNOR2X1_171 ( .A(w_mem_inst__abc_19396_new_n2268_), .B(w_mem_inst__abc_19396_new_n2269_), .Y(w_mem_inst__abc_19396_new_n2270_));
XNOR2X1 XNOR2X1_172 ( .A(w_mem_inst_w_mem_13__26_), .B(w_mem_inst_w_mem_8__26_), .Y(w_mem_inst__abc_19396_new_n2293_));
XNOR2X1 XNOR2X1_173 ( .A(w_mem_inst_w_mem_2__26_), .B(w_mem_inst_w_mem_0__26_), .Y(w_mem_inst__abc_19396_new_n2294_));
XNOR2X1 XNOR2X1_174 ( .A(w_mem_inst__abc_19396_new_n2293_), .B(w_mem_inst__abc_19396_new_n2294_), .Y(w_mem_inst__abc_19396_new_n2295_));
XNOR2X1 XNOR2X1_175 ( .A(w_mem_inst_w_mem_13__27_), .B(w_mem_inst_w_mem_8__27_), .Y(w_mem_inst__abc_19396_new_n2318_));
XNOR2X1 XNOR2X1_176 ( .A(w_mem_inst_w_mem_2__27_), .B(w_mem_inst_w_mem_0__27_), .Y(w_mem_inst__abc_19396_new_n2319_));
XNOR2X1 XNOR2X1_177 ( .A(w_mem_inst__abc_19396_new_n2318_), .B(w_mem_inst__abc_19396_new_n2319_), .Y(w_mem_inst__abc_19396_new_n2320_));
XNOR2X1 XNOR2X1_178 ( .A(w_mem_inst_w_mem_13__28_), .B(w_mem_inst_w_mem_8__28_), .Y(w_mem_inst__abc_19396_new_n2343_));
XNOR2X1 XNOR2X1_179 ( .A(w_mem_inst_w_mem_2__28_), .B(w_mem_inst_w_mem_0__28_), .Y(w_mem_inst__abc_19396_new_n2344_));
XNOR2X1 XNOR2X1_18 ( .A(_abc_15497_new_n1634_), .B(_abc_15497_new_n1630_), .Y(_abc_15497_new_n1635_));
XNOR2X1 XNOR2X1_180 ( .A(w_mem_inst__abc_19396_new_n2343_), .B(w_mem_inst__abc_19396_new_n2344_), .Y(w_mem_inst__abc_19396_new_n2345_));
XNOR2X1 XNOR2X1_181 ( .A(w_mem_inst_w_mem_13__29_), .B(w_mem_inst_w_mem_8__29_), .Y(w_mem_inst__abc_19396_new_n2368_));
XNOR2X1 XNOR2X1_182 ( .A(w_mem_inst_w_mem_2__29_), .B(w_mem_inst_w_mem_0__29_), .Y(w_mem_inst__abc_19396_new_n2369_));
XNOR2X1 XNOR2X1_183 ( .A(w_mem_inst__abc_19396_new_n2368_), .B(w_mem_inst__abc_19396_new_n2369_), .Y(w_mem_inst__abc_19396_new_n2370_));
XNOR2X1 XNOR2X1_184 ( .A(w_mem_inst_w_mem_13__30_), .B(w_mem_inst_w_mem_8__30_), .Y(w_mem_inst__abc_19396_new_n2393_));
XNOR2X1 XNOR2X1_185 ( .A(w_mem_inst_w_mem_2__30_), .B(w_mem_inst_w_mem_0__30_), .Y(w_mem_inst__abc_19396_new_n2394_));
XNOR2X1 XNOR2X1_186 ( .A(w_mem_inst__abc_19396_new_n2393_), .B(w_mem_inst__abc_19396_new_n2394_), .Y(w_mem_inst__abc_19396_new_n2395_));
XNOR2X1 XNOR2X1_19 ( .A(_abc_15497_new_n1772_), .B(_abc_15497_new_n1775_), .Y(_abc_15497_new_n1776_));
XNOR2X1 XNOR2X1_2 ( .A(_auto_iopadmap_cc_368_execute_22625_95_), .B(c_reg_31_), .Y(_abc_15497_new_n929_));
XNOR2X1 XNOR2X1_20 ( .A(_auto_iopadmap_cc_368_execute_22625_100_), .B(b_reg_4_), .Y(_abc_15497_new_n1780_));
XNOR2X1 XNOR2X1_21 ( .A(_abc_15497_new_n1800_), .B(_abc_15497_new_n1804_), .Y(_abc_15497_new_n1805_));
XNOR2X1 XNOR2X1_22 ( .A(_abc_15497_new_n1825_), .B(_abc_15497_new_n1822_), .Y(_abc_15497_new_n1826_));
XNOR2X1 XNOR2X1_23 ( .A(_abc_15497_new_n1848_), .B(_abc_15497_new_n1852_), .Y(_abc_15497_new_n1853_));
XNOR2X1 XNOR2X1_24 ( .A(_abc_15497_new_n1869_), .B(_abc_15497_new_n1870_), .Y(_abc_15497_new_n1871_));
XNOR2X1 XNOR2X1_25 ( .A(_abc_15497_new_n1891_), .B(_abc_15497_new_n1895_), .Y(_abc_15497_new_n1896_));
XNOR2X1 XNOR2X1_26 ( .A(_abc_15497_new_n1921_), .B(_abc_15497_new_n1920_), .Y(_abc_15497_new_n1922_));
XNOR2X1 XNOR2X1_27 ( .A(_abc_15497_new_n1971_), .B(_abc_15497_new_n1969_), .Y(_abc_15497_new_n1972_));
XNOR2X1 XNOR2X1_28 ( .A(_abc_15497_new_n1978_), .B(_abc_15497_new_n1982_), .Y(_abc_15497_new_n1983_));
XNOR2X1 XNOR2X1_29 ( .A(_abc_15497_new_n2015_), .B(_abc_15497_new_n2019_), .Y(_abc_15497_new_n2020_));
XNOR2X1 XNOR2X1_3 ( .A(e_reg_6_), .B(_auto_iopadmap_cc_368_execute_22625_6_), .Y(_abc_15497_new_n986_));
XNOR2X1 XNOR2X1_30 ( .A(_abc_15497_new_n2039_), .B(_abc_15497_new_n2043_), .Y(_abc_15497_new_n2044_));
XNOR2X1 XNOR2X1_31 ( .A(_auto_iopadmap_cc_368_execute_22625_127_), .B(b_reg_31_), .Y(_abc_15497_new_n2083_));
XNOR2X1 XNOR2X1_32 ( .A(_auto_iopadmap_cc_368_execute_22625_132_), .B(a_reg_4_), .Y(_abc_15497_new_n2123_));
XNOR2X1 XNOR2X1_33 ( .A(_abc_15497_new_n2175_), .B(_abc_15497_new_n2176_), .Y(_abc_15497_new_n2177_));
XNOR2X1 XNOR2X1_34 ( .A(_abc_15497_new_n2199_), .B(_abc_15497_new_n2200_), .Y(_abc_15497_new_n2201_));
XNOR2X1 XNOR2X1_35 ( .A(_abc_15497_new_n2221_), .B(_abc_15497_new_n2224_), .Y(_abc_15497_new_n2225_));
XNOR2X1 XNOR2X1_36 ( .A(_abc_15497_new_n2242_), .B(_abc_15497_new_n2246_), .Y(_abc_15497_new_n2247_));
XNOR2X1 XNOR2X1_37 ( .A(_abc_15497_new_n2329_), .B(_abc_15497_new_n2334_), .Y(_abc_15497_new_n2335_));
XNOR2X1 XNOR2X1_38 ( .A(_auto_iopadmap_cc_368_execute_22625_151_), .B(a_reg_23_), .Y(_abc_15497_new_n2339_));
XNOR2X1 XNOR2X1_39 ( .A(_abc_15497_new_n2369_), .B(_abc_15497_new_n2374_), .Y(_abc_15497_new_n2375_));
XNOR2X1 XNOR2X1_4 ( .A(_abc_15497_new_n1071_), .B(_abc_15497_new_n1075_), .Y(_abc_15497_new_n1076_));
XNOR2X1 XNOR2X1_40 ( .A(_abc_15497_new_n2398_), .B(_abc_15497_new_n2397_), .Y(_abc_15497_new_n2399_));
XNOR2X1 XNOR2X1_41 ( .A(_abc_15497_new_n2766_), .B(_abc_15497_new_n2762_), .Y(_abc_15497_new_n2767_));
XNOR2X1 XNOR2X1_42 ( .A(_abc_15497_new_n3117_), .B(_abc_15497_new_n3162_), .Y(_abc_15497_new_n3163_));
XNOR2X1 XNOR2X1_43 ( .A(_abc_15497_new_n3227_), .B(_abc_15497_new_n3279_), .Y(_abc_15497_new_n3280_));
XNOR2X1 XNOR2X1_44 ( .A(d_reg_16_), .B(b_reg_16_), .Y(_abc_15497_new_n3682_));
XNOR2X1 XNOR2X1_45 ( .A(e_reg_16_), .B(a_reg_11_), .Y(_abc_15497_new_n3693_));
XNOR2X1 XNOR2X1_46 ( .A(_abc_15497_new_n3696_), .B(_abc_15497_new_n3691_), .Y(_abc_15497_new_n3700_));
XNOR2X1 XNOR2X1_47 ( .A(_abc_15497_new_n3787_), .B(d_reg_18_), .Y(_abc_15497_new_n3788_));
XNOR2X1 XNOR2X1_48 ( .A(e_reg_18_), .B(a_reg_13_), .Y(_abc_15497_new_n3798_));
XNOR2X1 XNOR2X1_49 ( .A(b_reg_19_), .B(c_reg_19_), .Y(_abc_15497_new_n3830_));
XNOR2X1 XNOR2X1_5 ( .A(_abc_15497_new_n1093_), .B(_abc_15497_new_n1097_), .Y(_abc_15497_new_n1098_));
XNOR2X1 XNOR2X1_50 ( .A(_abc_15497_new_n3830_), .B(_abc_15497_new_n1495_), .Y(_abc_15497_new_n3831_));
XNOR2X1 XNOR2X1_51 ( .A(e_reg_19_), .B(a_reg_14_), .Y(_abc_15497_new_n3842_));
XNOR2X1 XNOR2X1_52 ( .A(_abc_15497_new_n3840_), .B(_abc_15497_new_n3845_), .Y(_abc_15497_new_n3849_));
XNOR2X1 XNOR2X1_53 ( .A(d_reg_20_), .B(b_reg_20_), .Y(_abc_15497_new_n3894_));
XNOR2X1 XNOR2X1_54 ( .A(e_reg_20_), .B(a_reg_15_), .Y(_abc_15497_new_n3905_));
XNOR2X1 XNOR2X1_55 ( .A(_abc_15497_new_n3903_), .B(_abc_15497_new_n3908_), .Y(_abc_15497_new_n3912_));
XNOR2X1 XNOR2X1_56 ( .A(d_reg_21_), .B(b_reg_21_), .Y(_abc_15497_new_n3944_));
XNOR2X1 XNOR2X1_57 ( .A(e_reg_21_), .B(a_reg_16_), .Y(_abc_15497_new_n3956_));
XNOR2X1 XNOR2X1_58 ( .A(_abc_15497_new_n3954_), .B(_abc_15497_new_n3959_), .Y(_abc_15497_new_n3963_));
XNOR2X1 XNOR2X1_59 ( .A(d_reg_22_), .B(b_reg_22_), .Y(_abc_15497_new_n3999_));
XNOR2X1 XNOR2X1_6 ( .A(_abc_15497_new_n1119_), .B(_abc_15497_new_n1124_), .Y(_abc_15497_new_n1125_));
XNOR2X1 XNOR2X1_60 ( .A(e_reg_22_), .B(a_reg_17_), .Y(_abc_15497_new_n4011_));
XNOR2X1 XNOR2X1_61 ( .A(_abc_15497_new_n4009_), .B(_abc_15497_new_n4014_), .Y(_abc_15497_new_n4018_));
XNOR2X1 XNOR2X1_62 ( .A(e_reg_23_), .B(a_reg_18_), .Y(_abc_15497_new_n4065_));
XNOR2X1 XNOR2X1_63 ( .A(_abc_15497_new_n4131_), .B(_abc_15497_new_n4117_), .Y(_abc_15497_new_n4132_));
XNOR2X1 XNOR2X1_64 ( .A(_abc_15497_new_n4167_), .B(w_25_), .Y(_abc_15497_new_n4168_));
XNOR2X1 XNOR2X1_65 ( .A(_abc_15497_new_n4171_), .B(_abc_15497_new_n4162_), .Y(_abc_15497_new_n4172_));
XNOR2X1 XNOR2X1_66 ( .A(_abc_15497_new_n4214_), .B(_abc_15497_new_n4204_), .Y(_abc_15497_new_n4215_));
XNOR2X1 XNOR2X1_67 ( .A(_abc_15497_new_n4245_), .B(d_reg_27_), .Y(_abc_15497_new_n4246_));
XNOR2X1 XNOR2X1_68 ( .A(_abc_15497_new_n4254_), .B(_abc_15497_new_n4251_), .Y(_abc_15497_new_n4255_));
XNOR2X1 XNOR2X1_69 ( .A(_abc_15497_new_n4283_), .B(d_reg_28_), .Y(_abc_15497_new_n4284_));
XNOR2X1 XNOR2X1_7 ( .A(_abc_15497_new_n1144_), .B(_abc_15497_new_n1148_), .Y(_abc_15497_new_n1149_));
XNOR2X1 XNOR2X1_70 ( .A(_abc_15497_new_n4294_), .B(w_28_), .Y(_abc_15497_new_n4295_));
XNOR2X1 XNOR2X1_71 ( .A(_abc_15497_new_n4299_), .B(_abc_15497_new_n4279_), .Y(_abc_15497_new_n4300_));
XNOR2X1 XNOR2X1_72 ( .A(_abc_15497_new_n4300_), .B(_abc_15497_new_n2742__bF_buf3), .Y(_abc_15497_new_n4301_));
XNOR2X1 XNOR2X1_73 ( .A(_abc_15497_new_n4346_), .B(w_29_), .Y(_abc_15497_new_n4347_));
XNOR2X1 XNOR2X1_74 ( .A(_abc_15497_new_n4398_), .B(_abc_15497_new_n4371_), .Y(_abc_15497_new_n4399_));
XNOR2X1 XNOR2X1_75 ( .A(_abc_15497_new_n4399_), .B(_abc_15497_new_n2924__bF_buf0), .Y(_abc_15497_new_n4400_));
XNOR2X1 XNOR2X1_76 ( .A(_abc_15497_new_n4400_), .B(_abc_15497_new_n4370_), .Y(_abc_15497_new_n4401_));
XNOR2X1 XNOR2X1_77 ( .A(_abc_15497_new_n4368_), .B(_abc_15497_new_n4401_), .Y(_abc_15497_new_n4402_));
XNOR2X1 XNOR2X1_78 ( .A(_abc_15497_new_n4420_), .B(d_reg_31_), .Y(_abc_15497_new_n4421_));
XNOR2X1 XNOR2X1_79 ( .A(e_reg_31_), .B(w_31_), .Y(_abc_15497_new_n4427_));
XNOR2X1 XNOR2X1_8 ( .A(_abc_15497_new_n1176_), .B(_abc_15497_new_n1175_), .Y(_abc_15497_new_n1177_));
XNOR2X1 XNOR2X1_80 ( .A(_abc_15497_new_n4427_), .B(a_reg_26_), .Y(_abc_15497_new_n4428_));
XNOR2X1 XNOR2X1_81 ( .A(_abc_15497_new_n4431_), .B(_abc_15497_new_n2739_), .Y(_abc_15497_new_n4432_));
XNOR2X1 XNOR2X1_82 ( .A(_abc_15497_new_n4413_), .B(_abc_15497_new_n4432_), .Y(_abc_15497_new_n4433_));
XNOR2X1 XNOR2X1_83 ( .A(_abc_15497_new_n772_), .B(_abc_15497_new_n771_), .Y(_abc_15497_new_n4480_));
XNOR2X1 XNOR2X1_84 ( .A(_abc_15497_new_n774_), .B(_abc_15497_new_n776_), .Y(_abc_15497_new_n4483_));
XNOR2X1 XNOR2X1_85 ( .A(_abc_15497_new_n778_), .B(_abc_15497_new_n779_), .Y(_abc_15497_new_n4491_));
XNOR2X1 XNOR2X1_86 ( .A(_abc_15497_new_n4507_), .B(_abc_15497_new_n752_), .Y(_abc_15497_new_n4508_));
XNOR2X1 XNOR2X1_87 ( .A(_abc_15497_new_n4526_), .B(_abc_15497_new_n731_), .Y(_abc_15497_new_n4527_));
XNOR2X1 XNOR2X1_88 ( .A(_abc_15497_new_n4545_), .B(_abc_15497_new_n701_), .Y(_abc_15497_new_n4546_));
XNOR2X1 XNOR2X1_89 ( .A(_abc_15497_new_n4553_), .B(_abc_15497_new_n840_), .Y(_abc_15497_new_n4554_));
XNOR2X1 XNOR2X1_9 ( .A(_abc_15497_new_n1193_), .B(_abc_15497_new_n1197_), .Y(_abc_15497_new_n1198_));
XNOR2X1 XNOR2X1_90 ( .A(_abc_15497_new_n4557_), .B(_abc_15497_new_n827_), .Y(_abc_15497_new_n4558_));
XNOR2X1 XNOR2X1_91 ( .A(w_mem_inst_w_mem_8__31_), .B(w_mem_inst_w_mem_13__31_), .Y(w_mem_inst__abc_19396_new_n1588_));
XNOR2X1 XNOR2X1_92 ( .A(w_mem_inst_w_mem_2__31_), .B(w_mem_inst_w_mem_0__31_), .Y(w_mem_inst__abc_19396_new_n1589_));
XNOR2X1 XNOR2X1_93 ( .A(w_mem_inst__abc_19396_new_n1588_), .B(w_mem_inst__abc_19396_new_n1589_), .Y(w_mem_inst__abc_19396_new_n1590_));
XNOR2X1 XNOR2X1_94 ( .A(w_mem_inst_w_mem_13__0_), .B(w_mem_inst_w_mem_8__0_), .Y(w_mem_inst__abc_19396_new_n1643_));
XNOR2X1 XNOR2X1_95 ( .A(w_mem_inst_w_mem_2__0_), .B(w_mem_inst_w_mem_0__0_), .Y(w_mem_inst__abc_19396_new_n1644_));
XNOR2X1 XNOR2X1_96 ( .A(w_mem_inst__abc_19396_new_n1643_), .B(w_mem_inst__abc_19396_new_n1644_), .Y(w_mem_inst__abc_19396_new_n1645_));
XNOR2X1 XNOR2X1_97 ( .A(w_mem_inst_w_mem_13__1_), .B(w_mem_inst_w_mem_8__1_), .Y(w_mem_inst__abc_19396_new_n1668_));
XNOR2X1 XNOR2X1_98 ( .A(w_mem_inst_w_mem_2__1_), .B(w_mem_inst_w_mem_0__1_), .Y(w_mem_inst__abc_19396_new_n1669_));
XNOR2X1 XNOR2X1_99 ( .A(w_mem_inst__abc_19396_new_n1668_), .B(w_mem_inst__abc_19396_new_n1669_), .Y(w_mem_inst__abc_19396_new_n1670_));
XOR2X1 XOR2X1_1 ( .A(c_reg_1_), .B(_auto_iopadmap_cc_368_execute_22625_65_), .Y(_abc_15497_new_n772_));
XOR2X1 XOR2X1_10 ( .A(_auto_iopadmap_cc_368_execute_22625_33_), .B(d_reg_1_), .Y(_abc_15497_new_n1303_));
XOR2X1 XOR2X1_11 ( .A(_auto_iopadmap_cc_368_execute_22625_36_), .B(d_reg_4_), .Y(_abc_15497_new_n1326_));
XOR2X1 XOR2X1_12 ( .A(_auto_iopadmap_cc_368_execute_22625_37_), .B(d_reg_5_), .Y(_abc_15497_new_n1336_));
XOR2X1 XOR2X1_13 ( .A(_auto_iopadmap_cc_368_execute_22625_38_), .B(d_reg_6_), .Y(_abc_15497_new_n1345_));
XOR2X1 XOR2X1_14 ( .A(_abc_15497_new_n1520_), .B(_abc_15497_new_n1524_), .Y(_abc_15497_new_n1525_));
XOR2X1 XOR2X1_15 ( .A(_auto_iopadmap_cc_368_execute_22625_60_), .B(d_reg_28_), .Y(_abc_15497_new_n1611_));
XOR2X1 XOR2X1_16 ( .A(_auto_iopadmap_cc_368_execute_22625_62_), .B(d_reg_30_), .Y(_abc_15497_new_n1629_));
XOR2X1 XOR2X1_17 ( .A(_auto_iopadmap_cc_368_execute_22625_63_), .B(d_reg_31_), .Y(_abc_15497_new_n1640_));
XOR2X1 XOR2X1_18 ( .A(_auto_iopadmap_cc_368_execute_22625_97_), .B(b_reg_1_), .Y(_abc_15497_new_n1758_));
XOR2X1 XOR2X1_19 ( .A(_auto_iopadmap_cc_368_execute_22625_98_), .B(b_reg_2_), .Y(_abc_15497_new_n1766_));
XOR2X1 XOR2X1_2 ( .A(c_reg_4_), .B(_auto_iopadmap_cc_368_execute_22625_68_), .Y(_abc_15497_new_n779_));
XOR2X1 XOR2X1_20 ( .A(_abc_15497_new_n1829_), .B(_abc_15497_new_n1832_), .Y(_abc_15497_new_n1833_));
XOR2X1 XOR2X1_21 ( .A(_abc_15497_new_n1865_), .B(_abc_15497_new_n1860_), .Y(_abc_15497_new_n1866_));
XOR2X1 XOR2X1_22 ( .A(_auto_iopadmap_cc_368_execute_22625_109_), .B(b_reg_13_), .Y(_abc_15497_new_n1870_));
XOR2X1 XOR2X1_23 ( .A(_abc_15497_new_n1986_), .B(_abc_15497_new_n1990_), .Y(_abc_15497_new_n1991_));
XOR2X1 XOR2X1_24 ( .A(_auto_iopadmap_cc_368_execute_22625_126_), .B(b_reg_30_), .Y(_abc_15497_new_n2072_));
XOR2X1 XOR2X1_25 ( .A(_auto_iopadmap_cc_368_execute_22625_129_), .B(a_reg_1_), .Y(_abc_15497_new_n2099_));
XOR2X1 XOR2X1_26 ( .A(_auto_iopadmap_cc_368_execute_22625_130_), .B(a_reg_2_), .Y(_abc_15497_new_n2107_));
XOR2X1 XOR2X1_27 ( .A(_abc_15497_new_n2114_), .B(_abc_15497_new_n2119_), .Y(_abc_15497_new_n2120_));
XOR2X1 XOR2X1_28 ( .A(_auto_iopadmap_cc_368_execute_22625_135_), .B(a_reg_7_), .Y(_abc_15497_new_n2152_));
XOR2X1 XOR2X1_29 ( .A(_auto_iopadmap_cc_368_execute_22625_137_), .B(a_reg_9_), .Y(_abc_15497_new_n2176_));
XOR2X1 XOR2X1_3 ( .A(e_reg_1_), .B(_auto_iopadmap_cc_368_execute_22625_1_), .Y(_abc_15497_new_n942_));
XOR2X1 XOR2X1_30 ( .A(_auto_iopadmap_cc_368_execute_22625_139_), .B(a_reg_11_), .Y(_abc_15497_new_n2200_));
XOR2X1 XOR2X1_31 ( .A(_auto_iopadmap_cc_368_execute_22625_156_), .B(a_reg_28_), .Y(_abc_15497_new_n2409_));
XOR2X1 XOR2X1_32 ( .A(_auto_iopadmap_cc_368_execute_22625_159_), .B(a_reg_31_), .Y(_abc_15497_new_n2440_));
XOR2X1 XOR2X1_33 ( .A(_abc_15497_new_n2935_), .B(_abc_15497_new_n2883_), .Y(_abc_15497_new_n2936_));
XOR2X1 XOR2X1_34 ( .A(_abc_15497_new_n3696_), .B(_abc_15497_new_n3691_), .Y(_abc_15497_new_n3697_));
XOR2X1 XOR2X1_35 ( .A(_abc_15497_new_n3796_), .B(_abc_15497_new_n3801_), .Y(_abc_15497_new_n3802_));
XOR2X1 XOR2X1_36 ( .A(_abc_15497_new_n3840_), .B(_abc_15497_new_n3845_), .Y(_abc_15497_new_n3846_));
XOR2X1 XOR2X1_37 ( .A(_abc_15497_new_n3903_), .B(_abc_15497_new_n3908_), .Y(_abc_15497_new_n3909_));
XOR2X1 XOR2X1_38 ( .A(_abc_15497_new_n3954_), .B(_abc_15497_new_n3959_), .Y(_abc_15497_new_n3960_));
XOR2X1 XOR2X1_39 ( .A(_abc_15497_new_n4009_), .B(_abc_15497_new_n4014_), .Y(_abc_15497_new_n4015_));
XOR2X1 XOR2X1_4 ( .A(e_reg_2_), .B(_auto_iopadmap_cc_368_execute_22625_2_), .Y(_abc_15497_new_n950_));
XOR2X1 XOR2X1_40 ( .A(_abc_15497_new_n4206_), .B(_abc_15497_new_n4213_), .Y(_abc_15497_new_n4214_));
XOR2X1 XOR2X1_41 ( .A(_abc_15497_new_n4258_), .B(_abc_15497_new_n4249_), .Y(_abc_15497_new_n4259_));
XOR2X1 XOR2X1_42 ( .A(_abc_15497_new_n4259_), .B(_abc_15497_new_n4238_), .Y(_abc_15497_new_n4260_));
XOR2X1 XOR2X1_43 ( .A(_abc_15497_new_n4298_), .B(_abc_15497_new_n4289_), .Y(_abc_15497_new_n4299_));
XOR2X1 XOR2X1_44 ( .A(_abc_15497_new_n4347_), .B(_abc_15497_new_n4343_), .Y(_abc_15497_new_n4348_));
XOR2X1 XOR2X1_45 ( .A(_abc_15497_new_n4352_), .B(_abc_15497_new_n4329_), .Y(_abc_15497_new_n4353_));
XOR2X1 XOR2X1_46 ( .A(_abc_15497_new_n4393_), .B(_abc_15497_new_n4386_), .Y(_abc_15497_new_n4394_));
XOR2X1 XOR2X1_47 ( .A(_abc_15497_new_n4426_), .B(_abc_15497_new_n4428_), .Y(_abc_15497_new_n4429_));
XOR2X1 XOR2X1_48 ( .A(_abc_15497_new_n4425_), .B(_abc_15497_new_n4429_), .Y(_abc_15497_new_n4430_));
XOR2X1 XOR2X1_49 ( .A(_abc_15497_new_n4415_), .B(_abc_15497_new_n4430_), .Y(_abc_15497_new_n4431_));
XOR2X1 XOR2X1_5 ( .A(_abc_15497_new_n957_), .B(_abc_15497_new_n963_), .Y(_abc_15497_new_n964_));
XOR2X1 XOR2X1_50 ( .A(_abc_15497_new_n777_), .B(_abc_15497_new_n4486_), .Y(_abc_15497_new_n4487_));
XOR2X1 XOR2X1_51 ( .A(_abc_15497_new_n4560_), .B(_abc_15497_new_n822_), .Y(_abc_15497_new_n4561_));
XOR2X1 XOR2X1_6 ( .A(e_reg_9_), .B(_auto_iopadmap_cc_368_execute_22625_9_), .Y(_abc_15497_new_n1025_));
XOR2X1 XOR2X1_7 ( .A(_abc_15497_new_n1050_), .B(_abc_15497_new_n1054_), .Y(_abc_15497_new_n1055_));
XOR2X1 XOR2X1_8 ( .A(e_reg_28_), .B(_auto_iopadmap_cc_368_execute_22625_28_), .Y(_abc_15497_new_n1264_));
XOR2X1 XOR2X1_9 ( .A(e_reg_30_), .B(_auto_iopadmap_cc_368_execute_22625_30_), .Y(_abc_15497_new_n1280_));


endmodule