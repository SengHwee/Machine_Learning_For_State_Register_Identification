module b01_reset(clock, RESET_G, nRESET_G, LINE1, LINE2, OUTP_REG, OVERFLW_REG);

input LINE1;
input LINE2;
output OUTP_REG;
output OVERFLW_REG;
input RESET_G;
wire STATO_REG_0_; 
wire STATO_REG_1_; 
wire STATO_REG_2_; 
wire _abc_289_new_n12_; 
wire _abc_289_new_n13_; 
wire _abc_289_new_n15_; 
wire _abc_289_new_n16_; 
wire _abc_289_new_n17_; 
wire _abc_289_new_n18_; 
wire _abc_289_new_n19_; 
wire _abc_289_new_n20_; 
wire _abc_289_new_n21_; 
wire _abc_289_new_n22_; 
wire _abc_289_new_n23_; 
wire _abc_289_new_n24_; 
wire _abc_289_new_n25_; 
wire _abc_289_new_n26_; 
wire _abc_289_new_n27_; 
wire _abc_289_new_n28_; 
wire _abc_289_new_n29_; 
wire _abc_289_new_n30_; 
wire _abc_289_new_n32_; 
wire _abc_289_new_n33_; 
wire _abc_289_new_n34_; 
wire _abc_289_new_n35_; 
wire _abc_289_new_n36_; 
wire _abc_289_new_n37_; 
wire _abc_289_new_n38_; 
wire _abc_289_new_n40_; 
wire _abc_289_new_n41_; 
wire _abc_289_new_n42_; 
wire _abc_289_new_n43_; 
wire _abc_289_new_n45_; 
wire _abc_289_new_n46_; 
wire _abc_289_new_n47_; 
input clock;
wire n14; 
wire n18; 
wire n23; 
wire n28; 
wire n33; 
input nRESET_G;
AOI21X1 AOI21X1_1 ( .A(_abc_289_new_n15_), .B(STATO_REG_1_), .C(_abc_289_new_n24_), .Y(_abc_289_new_n25_));
AOI21X1 AOI21X1_2 ( .A(_abc_289_new_n25_), .B(_abc_289_new_n23_), .C(_abc_289_new_n12_), .Y(_abc_289_new_n26_));
AOI21X1 AOI21X1_3 ( .A(n14), .B(_abc_289_new_n27_), .C(_abc_289_new_n29_), .Y(_abc_289_new_n30_));
AOI21X1 AOI21X1_4 ( .A(LINE2), .B(LINE1), .C(_abc_289_new_n15_), .Y(_abc_289_new_n35_));
AOI22X1 AOI22X1_1 ( .A(_abc_289_new_n28_), .B(_abc_289_new_n35_), .C(_abc_289_new_n36_), .D(_abc_289_new_n37_), .Y(_abc_289_new_n38_));
DFFPOSX1 DFFPOSX1_1 ( .CLK(clock), .D(n18), .Q(STATO_REG_2_));
DFFPOSX1 DFFPOSX1_2 ( .CLK(clock), .D(n14), .Q(OVERFLW_REG));
DFFPOSX1 DFFPOSX1_3 ( .CLK(clock), .D(n28), .Q(STATO_REG_0_));
DFFPOSX1 DFFPOSX1_4 ( .CLK(clock), .D(n33), .Q(OUTP_REG));
DFFPOSX1 DFFPOSX1_5 ( .CLK(clock), .D(n23), .Q(STATO_REG_1_));
INVX1 INVX1_1 ( .A(nRESET_G), .Y(_abc_289_new_n12_));
INVX1 INVX1_2 ( .A(STATO_REG_0_), .Y(_abc_289_new_n15_));
INVX1 INVX1_3 ( .A(LINE2), .Y(_abc_289_new_n17_));
INVX1 INVX1_4 ( .A(LINE1), .Y(_abc_289_new_n18_));
INVX1 INVX1_5 ( .A(_abc_289_new_n22_), .Y(_abc_289_new_n23_));
INVX1 INVX1_6 ( .A(STATO_REG_2_), .Y(_abc_289_new_n24_));
INVX1 INVX1_7 ( .A(STATO_REG_1_), .Y(_abc_289_new_n28_));
INVX1 INVX1_8 ( .A(_abc_289_new_n27_), .Y(_abc_289_new_n42_));
NAND2X1 NAND2X1_1 ( .A(STATO_REG_0_), .B(STATO_REG_1_), .Y(_abc_289_new_n13_));
NAND2X1 NAND2X1_2 ( .A(LINE2), .B(LINE1), .Y(_abc_289_new_n27_));
NAND2X1 NAND2X1_3 ( .A(STATO_REG_1_), .B(_abc_289_new_n22_), .Y(_abc_289_new_n33_));
NAND3X1 NAND3X1_1 ( .A(LINE2), .B(LINE1), .C(_abc_289_new_n15_), .Y(_abc_289_new_n16_));
NAND3X1 NAND3X1_2 ( .A(_abc_289_new_n20_), .B(_abc_289_new_n16_), .C(_abc_289_new_n19_), .Y(_abc_289_new_n21_));
NAND3X1 NAND3X1_3 ( .A(_abc_289_new_n21_), .B(_abc_289_new_n26_), .C(_abc_289_new_n30_), .Y(n28));
NAND3X1 NAND3X1_4 ( .A(STATO_REG_2_), .B(_abc_289_new_n32_), .C(_abc_289_new_n33_), .Y(_abc_289_new_n34_));
NAND3X1 NAND3X1_5 ( .A(nRESET_G), .B(_abc_289_new_n34_), .C(_abc_289_new_n38_), .Y(n23));
NAND3X1 NAND3X1_6 ( .A(_abc_289_new_n27_), .B(_abc_289_new_n23_), .C(_abc_289_new_n40_), .Y(_abc_289_new_n41_));
NAND3X1 NAND3X1_7 ( .A(nRESET_G), .B(_abc_289_new_n43_), .C(_abc_289_new_n41_), .Y(n33));
NAND3X1 NAND3X1_8 ( .A(nRESET_G), .B(_abc_289_new_n45_), .C(_abc_289_new_n47_), .Y(n18));
NOR2X1 NOR2X1_1 ( .A(STATO_REG_2_), .B(STATO_REG_1_), .Y(_abc_289_new_n20_));
NOR2X1 NOR2X1_2 ( .A(LINE2), .B(LINE1), .Y(_abc_289_new_n22_));
NOR2X1 NOR2X1_3 ( .A(STATO_REG_0_), .B(_abc_289_new_n28_), .Y(_abc_289_new_n36_));
NOR2X1 NOR2X1_4 ( .A(STATO_REG_1_), .B(_abc_289_new_n24_), .Y(_abc_289_new_n46_));
NOR3X1 NOR3X1_1 ( .A(STATO_REG_2_), .B(_abc_289_new_n12_), .C(_abc_289_new_n13_), .Y(n14));
NOR3X1 NOR3X1_2 ( .A(STATO_REG_0_), .B(_abc_289_new_n28_), .C(_abc_289_new_n27_), .Y(_abc_289_new_n29_));
OAI21X1 OAI21X1_1 ( .A(_abc_289_new_n17_), .B(_abc_289_new_n18_), .C(STATO_REG_0_), .Y(_abc_289_new_n19_));
OAI21X1 OAI21X1_2 ( .A(LINE2), .B(LINE1), .C(_abc_289_new_n15_), .Y(_abc_289_new_n32_));
OAI21X1 OAI21X1_3 ( .A(_abc_289_new_n17_), .B(_abc_289_new_n18_), .C(STATO_REG_2_), .Y(_abc_289_new_n37_));
OAI21X1 OAI21X1_4 ( .A(STATO_REG_0_), .B(_abc_289_new_n28_), .C(STATO_REG_2_), .Y(_abc_289_new_n40_));
OAI21X1 OAI21X1_5 ( .A(_abc_289_new_n22_), .B(_abc_289_new_n42_), .C(_abc_289_new_n25_), .Y(_abc_289_new_n43_));
OAI21X1 OAI21X1_6 ( .A(_abc_289_new_n42_), .B(_abc_289_new_n36_), .C(_abc_289_new_n24_), .Y(_abc_289_new_n45_));
OAI21X1 OAI21X1_7 ( .A(STATO_REG_0_), .B(_abc_289_new_n23_), .C(_abc_289_new_n46_), .Y(_abc_289_new_n47_));


endmodule