module b01_reset(clock, RESET_G, nRESET_G, LINE1, LINE2, OUTP_REG, OVERFLW_REG);
  input LINE1;
  input LINE2;
  output OUTP_REG;
  output OVERFLW_REG;
  input RESET_G;
  wire STATO_REG_0_;
  wire STATO_REG_1_;
  wire STATO_REG_2_;
  wire _abc_291_n12;
  wire _abc_291_n13;
  wire _abc_291_n14;
  wire _abc_291_n16;
  wire _abc_291_n17;
  wire _abc_291_n18;
  wire _abc_291_n19;
  wire _abc_291_n20;
  wire _abc_291_n21;
  wire _abc_291_n22;
  wire _abc_291_n23_1;
  wire _abc_291_n24;
  wire _abc_291_n25;
  wire _abc_291_n26;
  wire _abc_291_n27;
  wire _abc_291_n28;
  wire _abc_291_n29;
  wire _abc_291_n30_1;
  wire _abc_291_n31;
  wire _abc_291_n32;
  wire _abc_291_n33;
  wire _abc_291_n34;
  wire _abc_291_n35_1;
  wire _abc_291_n36;
  wire _abc_291_n37;
  wire _abc_291_n39;
  wire _abc_291_n40_1;
  wire _abc_291_n41;
  wire _abc_291_n42;
  wire _abc_291_n43;
  wire _abc_291_n44;
  wire _abc_291_n45;
  wire _abc_291_n46;
  wire _abc_291_n47;
  wire _abc_291_n49;
  wire _abc_291_n50;
  wire _abc_291_n51;
  wire _abc_291_n52;
  wire _abc_291_n53;
  wire _abc_291_n55;
  wire _abc_291_n56;
  wire _abc_291_n57;
  wire _abc_291_n58;
  wire _abc_291_n59;
  wire _abc_291_n60;
  input clock;
  wire n14;
  wire n18;
  wire n23;
  wire n28;
  wire n33;
  input nRESET_G;
  AND2X2 AND2X2_1 ( .A(_abc_291_n12), .B(nRESET_G), .Y(_abc_291_n13) );
  AND2X2 AND2X2_10 ( .A(_abc_291_n12), .B(_abc_291_n30_1), .Y(_abc_291_n31) );
  AND2X2 AND2X2_11 ( .A(_abc_291_n29), .B(_abc_291_n31), .Y(_abc_291_n32) );
  AND2X2 AND2X2_12 ( .A(_abc_291_n32), .B(_abc_291_n27), .Y(_abc_291_n33) );
  AND2X2 AND2X2_13 ( .A(_abc_291_n21), .B(_abc_291_n16), .Y(_abc_291_n35_1) );
  AND2X2 AND2X2_14 ( .A(_abc_291_n26), .B(_abc_291_n30_1), .Y(_abc_291_n39) );
  AND2X2 AND2X2_15 ( .A(_abc_291_n43), .B(STATO_REG_2_), .Y(_abc_291_n44) );
  AND2X2 AND2X2_16 ( .A(_abc_291_n44), .B(_abc_291_n42), .Y(_abc_291_n45) );
  AND2X2 AND2X2_17 ( .A(_abc_291_n21), .B(_abc_291_n12), .Y(_abc_291_n46) );
  AND2X2 AND2X2_18 ( .A(_abc_291_n17), .B(_abc_291_n19), .Y(_abc_291_n49) );
  AND2X2 AND2X2_19 ( .A(_abc_291_n22), .B(_abc_291_n49), .Y(_abc_291_n50) );
  AND2X2 AND2X2_2 ( .A(STATO_REG_0_), .B(STATO_REG_1_), .Y(_abc_291_n14) );
  AND2X2 AND2X2_20 ( .A(_abc_291_n23_1), .B(_abc_291_n51), .Y(_abc_291_n52) );
  AND2X2 AND2X2_21 ( .A(_abc_291_n30_1), .B(STATO_REG_2_), .Y(_abc_291_n56) );
  AND2X2 AND2X2_22 ( .A(_abc_291_n55), .B(_abc_291_n56), .Y(_abc_291_n57) );
  AND2X2 AND2X2_23 ( .A(_abc_291_n58), .B(_abc_291_n12), .Y(_abc_291_n59) );
  AND2X2 AND2X2_3 ( .A(_abc_291_n13), .B(_abc_291_n14), .Y(n14) );
  AND2X2 AND2X2_4 ( .A(LINE2), .B(LINE1), .Y(_abc_291_n16) );
  AND2X2 AND2X2_5 ( .A(n14), .B(_abc_291_n17), .Y(_abc_291_n18) );
  AND2X2 AND2X2_6 ( .A(_abc_291_n20), .B(STATO_REG_1_), .Y(_abc_291_n21) );
  AND2X2 AND2X2_7 ( .A(_abc_291_n23_1), .B(_abc_291_n19), .Y(_abc_291_n24) );
  AND2X2 AND2X2_8 ( .A(_abc_291_n17), .B(STATO_REG_0_), .Y(_abc_291_n26) );
  AND2X2 AND2X2_9 ( .A(_abc_291_n16), .B(_abc_291_n20), .Y(_abc_291_n28) );
  DFFPOSX1 DFFPOSX1_1 ( .CLK(clock), .D(n33), .Q(OUTP_REG) );
  DFFPOSX1 DFFPOSX1_2 ( .CLK(clock), .D(n14), .Q(OVERFLW_REG) );
  DFFPOSX1 DFFPOSX1_3 ( .CLK(clock), .D(n18), .Q(STATO_REG_2_) );
  DFFPOSX1 DFFPOSX1_4 ( .CLK(clock), .D(n23), .Q(STATO_REG_1_) );
  DFFPOSX1 DFFPOSX1_5 ( .CLK(clock), .D(n28), .Q(STATO_REG_0_) );
  INVX1 INVX1_1 ( .A(_abc_291_n16), .Y(_abc_291_n17) );
  INVX1 INVX1_2 ( .A(STATO_REG_0_), .Y(_abc_291_n20) );
  INVX1 INVX1_3 ( .A(_abc_291_n22), .Y(_abc_291_n23_1) );
  INVX1 INVX1_4 ( .A(_abc_291_n26), .Y(_abc_291_n27) );
  INVX1 INVX1_5 ( .A(_abc_291_n28), .Y(_abc_291_n29) );
  INVX1 INVX1_6 ( .A(STATO_REG_1_), .Y(_abc_291_n30_1) );
  INVX1 INVX1_7 ( .A(nRESET_G), .Y(_abc_291_n34) );
  INVX1 INVX1_8 ( .A(_abc_291_n19), .Y(_abc_291_n41) );
  INVX1 INVX1_9 ( .A(_abc_291_n49), .Y(_abc_291_n51) );
  INVX2 INVX2_1 ( .A(STATO_REG_2_), .Y(_abc_291_n12) );
  OR2X2 OR2X2_1 ( .A(LINE2), .B(LINE1), .Y(_abc_291_n19) );
  OR2X2 OR2X2_10 ( .A(_abc_291_n45), .B(_abc_291_n46), .Y(_abc_291_n47) );
  OR2X2 OR2X2_11 ( .A(_abc_291_n47), .B(_abc_291_n40_1), .Y(n23) );
  OR2X2 OR2X2_12 ( .A(_abc_291_n52), .B(_abc_291_n34), .Y(_abc_291_n53) );
  OR2X2 OR2X2_13 ( .A(_abc_291_n53), .B(_abc_291_n50), .Y(n33) );
  OR2X2 OR2X2_14 ( .A(_abc_291_n19), .B(STATO_REG_0_), .Y(_abc_291_n55) );
  OR2X2 OR2X2_15 ( .A(_abc_291_n21), .B(_abc_291_n16), .Y(_abc_291_n58) );
  OR2X2 OR2X2_16 ( .A(_abc_291_n59), .B(_abc_291_n34), .Y(_abc_291_n60) );
  OR2X2 OR2X2_17 ( .A(_abc_291_n60), .B(_abc_291_n57), .Y(n18) );
  OR2X2 OR2X2_2 ( .A(_abc_291_n21), .B(_abc_291_n12), .Y(_abc_291_n22) );
  OR2X2 OR2X2_3 ( .A(_abc_291_n24), .B(_abc_291_n18), .Y(_abc_291_n25) );
  OR2X2 OR2X2_4 ( .A(_abc_291_n35_1), .B(_abc_291_n34), .Y(_abc_291_n36) );
  OR2X2 OR2X2_5 ( .A(_abc_291_n33), .B(_abc_291_n36), .Y(_abc_291_n37) );
  OR2X2 OR2X2_6 ( .A(_abc_291_n37), .B(_abc_291_n25), .Y(n28) );
  OR2X2 OR2X2_7 ( .A(_abc_291_n36), .B(_abc_291_n39), .Y(_abc_291_n40_1) );
  OR2X2 OR2X2_8 ( .A(_abc_291_n41), .B(STATO_REG_0_), .Y(_abc_291_n42) );
  OR2X2 OR2X2_9 ( .A(_abc_291_n19), .B(_abc_291_n30_1), .Y(_abc_291_n43) );
endmodule