module uart(clk, rst, rx, transmit, \tx_byte[0] , \tx_byte[1] , \tx_byte[2] , \tx_byte[3] , \tx_byte[4] , \tx_byte[5] , \tx_byte[6] , \tx_byte[7] , tx, received, \rx_byte[0] , \rx_byte[1] , \rx_byte[2] , \rx_byte[3] , \rx_byte[4] , \rx_byte[5] , \rx_byte[6] , \rx_byte[7] , is_receiving, is_transmitting, recv_error);

wire _0recv_state_2_0__0_; 
wire _0recv_state_2_0__1_; 
wire _0recv_state_2_0__2_; 
wire _0rx_bits_remaining_3_0__0_; 
wire _0rx_bits_remaining_3_0__1_; 
wire _0rx_bits_remaining_3_0__2_; 
wire _0rx_bits_remaining_3_0__3_; 
wire _0rx_clk_divider_10_0__0_; 
wire _0rx_clk_divider_10_0__10_; 
wire _0rx_clk_divider_10_0__1_; 
wire _0rx_clk_divider_10_0__2_; 
wire _0rx_clk_divider_10_0__3_; 
wire _0rx_clk_divider_10_0__4_; 
wire _0rx_clk_divider_10_0__5_; 
wire _0rx_clk_divider_10_0__6_; 
wire _0rx_clk_divider_10_0__7_; 
wire _0rx_clk_divider_10_0__8_; 
wire _0rx_clk_divider_10_0__9_; 
wire _0rx_countdown_5_0__0_; 
wire _0rx_countdown_5_0__1_; 
wire _0rx_countdown_5_0__2_; 
wire _0rx_countdown_5_0__3_; 
wire _0rx_countdown_5_0__4_; 
wire _0rx_countdown_5_0__5_; 
wire _0rx_data_7_0__0_; 
wire _0rx_data_7_0__1_; 
wire _0rx_data_7_0__2_; 
wire _0rx_data_7_0__3_; 
wire _0rx_data_7_0__4_; 
wire _0rx_data_7_0__5_; 
wire _0rx_data_7_0__6_; 
wire _0rx_data_7_0__7_; 
wire _0tx_bits_remaining_3_0__0_; 
wire _0tx_bits_remaining_3_0__1_; 
wire _0tx_bits_remaining_3_0__2_; 
wire _0tx_bits_remaining_3_0__3_; 
wire _0tx_clk_divider_10_0__0_; 
wire _0tx_clk_divider_10_0__10_; 
wire _0tx_clk_divider_10_0__1_; 
wire _0tx_clk_divider_10_0__2_; 
wire _0tx_clk_divider_10_0__3_; 
wire _0tx_clk_divider_10_0__4_; 
wire _0tx_clk_divider_10_0__5_; 
wire _0tx_clk_divider_10_0__6_; 
wire _0tx_clk_divider_10_0__7_; 
wire _0tx_clk_divider_10_0__8_; 
wire _0tx_clk_divider_10_0__9_; 
wire _0tx_countdown_5_0__0_; 
wire _0tx_countdown_5_0__1_; 
wire _0tx_countdown_5_0__2_; 
wire _0tx_countdown_5_0__3_; 
wire _0tx_countdown_5_0__4_; 
wire _0tx_countdown_5_0__5_; 
wire _0tx_data_7_0__0_; 
wire _0tx_data_7_0__1_; 
wire _0tx_data_7_0__2_; 
wire _0tx_data_7_0__3_; 
wire _0tx_data_7_0__4_; 
wire _0tx_data_7_0__5_; 
wire _0tx_data_7_0__6_; 
wire _0tx_data_7_0__7_; 
wire _0tx_out_0_0_; 
wire _0tx_state_1_0__0_; 
wire _0tx_state_1_0__1_; 
wire _abc_2284_new_n144_; 
wire _abc_2284_new_n145_; 
wire _abc_2284_new_n146_; 
wire _abc_2284_new_n147_; 
wire _abc_2284_new_n150_; 
wire _abc_2284_new_n152_; 
wire _abc_2284_new_n153_; 
wire _abc_2284_new_n155_; 
wire _abc_2284_new_n156_; 
wire _abc_2284_new_n157_; 
wire _abc_2284_new_n158_; 
wire _abc_2284_new_n159_; 
wire _abc_2284_new_n160_; 
wire _abc_2284_new_n161_; 
wire _abc_2284_new_n162_; 
wire _abc_2284_new_n163_; 
wire _abc_2284_new_n164_; 
wire _abc_2284_new_n165_; 
wire _abc_2284_new_n166_; 
wire _abc_2284_new_n167_; 
wire _abc_2284_new_n168_; 
wire _abc_2284_new_n169_; 
wire _abc_2284_new_n170_; 
wire _abc_2284_new_n171_; 
wire _abc_2284_new_n172_; 
wire _abc_2284_new_n173_; 
wire _abc_2284_new_n174_; 
wire _abc_2284_new_n175_; 
wire _abc_2284_new_n176_; 
wire _abc_2284_new_n177_; 
wire _abc_2284_new_n178_; 
wire _abc_2284_new_n179_; 
wire _abc_2284_new_n180_; 
wire _abc_2284_new_n181_; 
wire _abc_2284_new_n182_; 
wire _abc_2284_new_n183_; 
wire _abc_2284_new_n184_; 
wire _abc_2284_new_n185_; 
wire _abc_2284_new_n186_; 
wire _abc_2284_new_n187_; 
wire _abc_2284_new_n188_; 
wire _abc_2284_new_n189_; 
wire _abc_2284_new_n190_; 
wire _abc_2284_new_n191_; 
wire _abc_2284_new_n192_; 
wire _abc_2284_new_n193_; 
wire _abc_2284_new_n194_; 
wire _abc_2284_new_n195_; 
wire _abc_2284_new_n196_; 
wire _abc_2284_new_n197_; 
wire _abc_2284_new_n198_; 
wire _abc_2284_new_n199_; 
wire _abc_2284_new_n200_; 
wire _abc_2284_new_n201_; 
wire _abc_2284_new_n202_; 
wire _abc_2284_new_n203_; 
wire _abc_2284_new_n204_; 
wire _abc_2284_new_n205_; 
wire _abc_2284_new_n206_; 
wire _abc_2284_new_n207_; 
wire _abc_2284_new_n208_; 
wire _abc_2284_new_n209_; 
wire _abc_2284_new_n210_; 
wire _abc_2284_new_n211_; 
wire _abc_2284_new_n212_; 
wire _abc_2284_new_n213_; 
wire _abc_2284_new_n214_; 
wire _abc_2284_new_n215_; 
wire _abc_2284_new_n216_; 
wire _abc_2284_new_n217_; 
wire _abc_2284_new_n218_; 
wire _abc_2284_new_n219_; 
wire _abc_2284_new_n220_; 
wire _abc_2284_new_n221_; 
wire _abc_2284_new_n222_; 
wire _abc_2284_new_n223_; 
wire _abc_2284_new_n224_; 
wire _abc_2284_new_n225_; 
wire _abc_2284_new_n226_; 
wire _abc_2284_new_n227_; 
wire _abc_2284_new_n228_; 
wire _abc_2284_new_n229_; 
wire _abc_2284_new_n230_; 
wire _abc_2284_new_n231_; 
wire _abc_2284_new_n232_; 
wire _abc_2284_new_n233_; 
wire _abc_2284_new_n234_; 
wire _abc_2284_new_n235_; 
wire _abc_2284_new_n236_; 
wire _abc_2284_new_n237_; 
wire _abc_2284_new_n238_; 
wire _abc_2284_new_n239_; 
wire _abc_2284_new_n240_; 
wire _abc_2284_new_n241_; 
wire _abc_2284_new_n242_; 
wire _abc_2284_new_n243_; 
wire _abc_2284_new_n244_; 
wire _abc_2284_new_n245_; 
wire _abc_2284_new_n246_; 
wire _abc_2284_new_n247_; 
wire _abc_2284_new_n248_; 
wire _abc_2284_new_n249_; 
wire _abc_2284_new_n250_; 
wire _abc_2284_new_n251_; 
wire _abc_2284_new_n252_; 
wire _abc_2284_new_n253_; 
wire _abc_2284_new_n254_; 
wire _abc_2284_new_n255_; 
wire _abc_2284_new_n256_; 
wire _abc_2284_new_n257_; 
wire _abc_2284_new_n258_; 
wire _abc_2284_new_n259_; 
wire _abc_2284_new_n260_; 
wire _abc_2284_new_n261_; 
wire _abc_2284_new_n262_; 
wire _abc_2284_new_n263_; 
wire _abc_2284_new_n264_; 
wire _abc_2284_new_n265_; 
wire _abc_2284_new_n266_; 
wire _abc_2284_new_n267_; 
wire _abc_2284_new_n268_; 
wire _abc_2284_new_n269_; 
wire _abc_2284_new_n270_; 
wire _abc_2284_new_n271_; 
wire _abc_2284_new_n272_; 
wire _abc_2284_new_n273_; 
wire _abc_2284_new_n274_; 
wire _abc_2284_new_n275_; 
wire _abc_2284_new_n276_; 
wire _abc_2284_new_n277_; 
wire _abc_2284_new_n278_; 
wire _abc_2284_new_n279_; 
wire _abc_2284_new_n280_; 
wire _abc_2284_new_n281_; 
wire _abc_2284_new_n282_; 
wire _abc_2284_new_n283_; 
wire _abc_2284_new_n284_; 
wire _abc_2284_new_n285_; 
wire _abc_2284_new_n286_; 
wire _abc_2284_new_n287_; 
wire _abc_2284_new_n288_; 
wire _abc_2284_new_n289_; 
wire _abc_2284_new_n290_; 
wire _abc_2284_new_n291_; 
wire _abc_2284_new_n292_; 
wire _abc_2284_new_n293_; 
wire _abc_2284_new_n294_; 
wire _abc_2284_new_n295_; 
wire _abc_2284_new_n296_; 
wire _abc_2284_new_n297_; 
wire _abc_2284_new_n298_; 
wire _abc_2284_new_n299_; 
wire _abc_2284_new_n301_; 
wire _abc_2284_new_n302_; 
wire _abc_2284_new_n303_; 
wire _abc_2284_new_n304_; 
wire _abc_2284_new_n305_; 
wire _abc_2284_new_n306_; 
wire _abc_2284_new_n307_; 
wire _abc_2284_new_n309_; 
wire _abc_2284_new_n310_; 
wire _abc_2284_new_n311_; 
wire _abc_2284_new_n312_; 
wire _abc_2284_new_n313_; 
wire _abc_2284_new_n314_; 
wire _abc_2284_new_n315_; 
wire _abc_2284_new_n317_; 
wire _abc_2284_new_n318_; 
wire _abc_2284_new_n319_; 
wire _abc_2284_new_n320_; 
wire _abc_2284_new_n321_; 
wire _abc_2284_new_n322_; 
wire _abc_2284_new_n323_; 
wire _abc_2284_new_n325_; 
wire _abc_2284_new_n326_; 
wire _abc_2284_new_n327_; 
wire _abc_2284_new_n328_; 
wire _abc_2284_new_n329_; 
wire _abc_2284_new_n330_; 
wire _abc_2284_new_n331_; 
wire _abc_2284_new_n333_; 
wire _abc_2284_new_n334_; 
wire _abc_2284_new_n335_; 
wire _abc_2284_new_n336_; 
wire _abc_2284_new_n337_; 
wire _abc_2284_new_n338_; 
wire _abc_2284_new_n339_; 
wire _abc_2284_new_n341_; 
wire _abc_2284_new_n342_; 
wire _abc_2284_new_n343_; 
wire _abc_2284_new_n344_; 
wire _abc_2284_new_n345_; 
wire _abc_2284_new_n346_; 
wire _abc_2284_new_n347_; 
wire _abc_2284_new_n348_; 
wire _abc_2284_new_n350_; 
wire _abc_2284_new_n351_; 
wire _abc_2284_new_n352_; 
wire _abc_2284_new_n354_; 
wire _abc_2284_new_n355_; 
wire _abc_2284_new_n356_; 
wire _abc_2284_new_n357_; 
wire _abc_2284_new_n358_; 
wire _abc_2284_new_n359_; 
wire _abc_2284_new_n360_; 
wire _abc_2284_new_n361_; 
wire _abc_2284_new_n363_; 
wire _abc_2284_new_n364_; 
wire _abc_2284_new_n365_; 
wire _abc_2284_new_n366_; 
wire _abc_2284_new_n367_; 
wire _abc_2284_new_n368_; 
wire _abc_2284_new_n369_; 
wire _abc_2284_new_n370_; 
wire _abc_2284_new_n372_; 
wire _abc_2284_new_n373_; 
wire _abc_2284_new_n374_; 
wire _abc_2284_new_n375_; 
wire _abc_2284_new_n376_; 
wire _abc_2284_new_n377_; 
wire _abc_2284_new_n378_; 
wire _abc_2284_new_n379_; 
wire _abc_2284_new_n381_; 
wire _abc_2284_new_n382_; 
wire _abc_2284_new_n383_; 
wire _abc_2284_new_n385_; 
wire _abc_2284_new_n386_; 
wire _abc_2284_new_n388_; 
wire _abc_2284_new_n390_; 
wire _abc_2284_new_n391_; 
wire _abc_2284_new_n392_; 
wire _abc_2284_new_n394_; 
wire _abc_2284_new_n395_; 
wire _abc_2284_new_n396_; 
wire _abc_2284_new_n397_; 
wire _abc_2284_new_n398_; 
wire _abc_2284_new_n400_; 
wire _abc_2284_new_n402_; 
wire _abc_2284_new_n404_; 
wire _abc_2284_new_n405_; 
wire _abc_2284_new_n406_; 
wire _abc_2284_new_n408_; 
wire _abc_2284_new_n409_; 
wire _abc_2284_new_n410_; 
wire _abc_2284_new_n412_; 
wire _abc_2284_new_n413_; 
wire _abc_2284_new_n414_; 
wire _abc_2284_new_n415_; 
wire _abc_2284_new_n416_; 
wire _abc_2284_new_n417_; 
wire _abc_2284_new_n418_; 
wire _abc_2284_new_n420_; 
wire _abc_2284_new_n421_; 
wire _abc_2284_new_n422_; 
wire _abc_2284_new_n423_; 
wire _abc_2284_new_n424_; 
wire _abc_2284_new_n425_; 
wire _abc_2284_new_n426_; 
wire _abc_2284_new_n427_; 
wire _abc_2284_new_n428_; 
wire _abc_2284_new_n429_; 
wire _abc_2284_new_n430_; 
wire _abc_2284_new_n431_; 
wire _abc_2284_new_n432_; 
wire _abc_2284_new_n433_; 
wire _abc_2284_new_n434_; 
wire _abc_2284_new_n435_; 
wire _abc_2284_new_n436_; 
wire _abc_2284_new_n437_; 
wire _abc_2284_new_n438_; 
wire _abc_2284_new_n439_; 
wire _abc_2284_new_n440_; 
wire _abc_2284_new_n441_; 
wire _abc_2284_new_n442_; 
wire _abc_2284_new_n443_; 
wire _abc_2284_new_n444_; 
wire _abc_2284_new_n445_; 
wire _abc_2284_new_n446_; 
wire _abc_2284_new_n447_; 
wire _abc_2284_new_n448_; 
wire _abc_2284_new_n449_; 
wire _abc_2284_new_n450_; 
wire _abc_2284_new_n451_; 
wire _abc_2284_new_n452_; 
wire _abc_2284_new_n453_; 
wire _abc_2284_new_n454_; 
wire _abc_2284_new_n455_; 
wire _abc_2284_new_n456_; 
wire _abc_2284_new_n457_; 
wire _abc_2284_new_n458_; 
wire _abc_2284_new_n459_; 
wire _abc_2284_new_n460_; 
wire _abc_2284_new_n461_; 
wire _abc_2284_new_n462_; 
wire _abc_2284_new_n463_; 
wire _abc_2284_new_n464_; 
wire _abc_2284_new_n465_; 
wire _abc_2284_new_n466_; 
wire _abc_2284_new_n467_; 
wire _abc_2284_new_n468_; 
wire _abc_2284_new_n469_; 
wire _abc_2284_new_n470_; 
wire _abc_2284_new_n471_; 
wire _abc_2284_new_n472_; 
wire _abc_2284_new_n473_; 
wire _abc_2284_new_n474_; 
wire _abc_2284_new_n475_; 
wire _abc_2284_new_n476_; 
wire _abc_2284_new_n477_; 
wire _abc_2284_new_n479_; 
wire _abc_2284_new_n480_; 
wire _abc_2284_new_n481_; 
wire _abc_2284_new_n482_; 
wire _abc_2284_new_n483_; 
wire _abc_2284_new_n484_; 
wire _abc_2284_new_n485_; 
wire _abc_2284_new_n486_; 
wire _abc_2284_new_n487_; 
wire _abc_2284_new_n488_; 
wire _abc_2284_new_n489_; 
wire _abc_2284_new_n491_; 
wire _abc_2284_new_n492_; 
wire _abc_2284_new_n493_; 
wire _abc_2284_new_n494_; 
wire _abc_2284_new_n495_; 
wire _abc_2284_new_n496_; 
wire _abc_2284_new_n497_; 
wire _abc_2284_new_n498_; 
wire _abc_2284_new_n499_; 
wire _abc_2284_new_n500_; 
wire _abc_2284_new_n501_; 
wire _abc_2284_new_n502_; 
wire _abc_2284_new_n503_; 
wire _abc_2284_new_n504_; 
wire _abc_2284_new_n505_; 
wire _abc_2284_new_n506_; 
wire _abc_2284_new_n507_; 
wire _abc_2284_new_n508_; 
wire _abc_2284_new_n509_; 
wire _abc_2284_new_n510_; 
wire _abc_2284_new_n511_; 
wire _abc_2284_new_n512_; 
wire _abc_2284_new_n513_; 
wire _abc_2284_new_n514_; 
wire _abc_2284_new_n515_; 
wire _abc_2284_new_n516_; 
wire _abc_2284_new_n517_; 
wire _abc_2284_new_n518_; 
wire _abc_2284_new_n519_; 
wire _abc_2284_new_n520_; 
wire _abc_2284_new_n521_; 
wire _abc_2284_new_n522_; 
wire _abc_2284_new_n523_; 
wire _abc_2284_new_n524_; 
wire _abc_2284_new_n525_; 
wire _abc_2284_new_n526_; 
wire _abc_2284_new_n527_; 
wire _abc_2284_new_n528_; 
wire _abc_2284_new_n529_; 
wire _abc_2284_new_n530_; 
wire _abc_2284_new_n531_; 
wire _abc_2284_new_n532_; 
wire _abc_2284_new_n533_; 
wire _abc_2284_new_n534_; 
wire _abc_2284_new_n535_; 
wire _abc_2284_new_n536_; 
wire _abc_2284_new_n537_; 
wire _abc_2284_new_n538_; 
wire _abc_2284_new_n539_; 
wire _abc_2284_new_n540_; 
wire _abc_2284_new_n541_; 
wire _abc_2284_new_n542_; 
wire _abc_2284_new_n543_; 
wire _abc_2284_new_n544_; 
wire _abc_2284_new_n545_; 
wire _abc_2284_new_n546_; 
wire _abc_2284_new_n547_; 
wire _abc_2284_new_n548_; 
wire _abc_2284_new_n549_; 
wire _abc_2284_new_n550_; 
wire _abc_2284_new_n551_; 
wire _abc_2284_new_n552_; 
wire _abc_2284_new_n553_; 
wire _abc_2284_new_n554_; 
wire _abc_2284_new_n556_; 
wire _abc_2284_new_n557_; 
wire _abc_2284_new_n558_; 
wire _abc_2284_new_n560_; 
wire _abc_2284_new_n561_; 
wire _abc_2284_new_n562_; 
wire _abc_2284_new_n563_; 
wire _abc_2284_new_n564_; 
wire _abc_2284_new_n565_; 
wire _abc_2284_new_n566_; 
wire _abc_2284_new_n567_; 
wire _abc_2284_new_n568_; 
wire _abc_2284_new_n569_; 
wire _abc_2284_new_n570_; 
wire _abc_2284_new_n571_; 
wire _abc_2284_new_n572_; 
wire _abc_2284_new_n573_; 
wire _abc_2284_new_n575_; 
wire _abc_2284_new_n577_; 
wire _abc_2284_new_n578_; 
wire _abc_2284_new_n579_; 
wire _abc_2284_new_n580_; 
wire _abc_2284_new_n581_; 
wire _abc_2284_new_n582_; 
wire _abc_2284_new_n583_; 
wire _abc_2284_new_n584_; 
wire _abc_2284_new_n585_; 
wire _abc_2284_new_n586_; 
wire _abc_2284_new_n587_; 
wire _abc_2284_new_n588_; 
wire _abc_2284_new_n589_; 
wire _abc_2284_new_n590_; 
wire _abc_2284_new_n591_; 
wire _abc_2284_new_n592_; 
wire _abc_2284_new_n593_; 
wire _abc_2284_new_n594_; 
wire _abc_2284_new_n595_; 
wire _abc_2284_new_n596_; 
wire _abc_2284_new_n598_; 
wire _abc_2284_new_n599_; 
wire _abc_2284_new_n600_; 
wire _abc_2284_new_n602_; 
wire _abc_2284_new_n603_; 
wire _abc_2284_new_n604_; 
wire _abc_2284_new_n605_; 
wire _abc_2284_new_n606_; 
wire _abc_2284_new_n607_; 
wire _abc_2284_new_n608_; 
wire _abc_2284_new_n609_; 
wire _abc_2284_new_n611_; 
wire _abc_2284_new_n612_; 
wire _abc_2284_new_n613_; 
wire _abc_2284_new_n614_; 
wire _abc_2284_new_n615_; 
wire _abc_2284_new_n616_; 
wire _abc_2284_new_n617_; 
wire _abc_2284_new_n619_; 
wire _abc_2284_new_n620_; 
wire _abc_2284_new_n621_; 
wire _abc_2284_new_n622_; 
wire _abc_2284_new_n623_; 
wire _abc_2284_new_n624_; 
wire _abc_2284_new_n625_; 
wire _abc_2284_new_n627_; 
wire _abc_2284_new_n628_; 
wire _abc_2284_new_n629_; 
wire _abc_2284_new_n630_; 
wire _abc_2284_new_n631_; 
wire _abc_2284_new_n632_; 
wire _abc_2284_new_n634_; 
wire _abc_2284_new_n635_; 
wire _abc_2284_new_n636_; 
wire _abc_2284_new_n637_; 
wire _abc_2284_new_n638_; 
wire _abc_2284_new_n639_; 
wire _abc_2284_new_n640_; 
wire _abc_2284_new_n641_; 
wire _abc_2284_new_n644_; 
wire _abc_2284_new_n645_; 
wire _abc_2284_new_n646_; 
wire _abc_2284_new_n648_; 
wire _abc_2284_new_n649_; 
wire _abc_2284_new_n650_; 
wire _abc_2284_new_n651_; 
wire _abc_2284_new_n653_; 
wire _abc_2284_new_n654_; 
wire _abc_2284_new_n655_; 
wire _abc_2284_new_n657_; 
wire _abc_2284_new_n658_; 
wire _abc_2284_new_n660_; 
wire _abc_2284_new_n662_; 
wire _abc_2284_new_n664_; 
wire _abc_2284_new_n666_; 
wire _abc_2284_new_n667_; 
wire _abc_2284_new_n669_; 
wire _abc_2284_new_n671_; 
wire _abc_2284_new_n672_; 
wire _abc_2284_new_n674_; 
wire _abc_2284_new_n675_; 
wire _abc_2284_new_n677_; 
wire _abc_2284_new_n678_; 
wire _abc_2284_new_n679_; 
wire _abc_2284_new_n680_; 
wire _abc_2284_new_n682_; 
wire _abc_2284_new_n683_; 
wire _abc_2284_new_n684_; 
wire _abc_2284_new_n685_; 
wire _abc_2284_new_n686_; 
wire _abc_2284_new_n688_; 
wire _abc_2284_new_n689_; 
wire _abc_2284_new_n690_; 
wire _abc_2284_new_n692_; 
wire _abc_2284_new_n694_; 
wire _abc_2284_new_n696_; 
wire _abc_2284_new_n698_; 
wire _abc_2284_new_n700_; 
wire _abc_2284_new_n701_; 
wire _abc_2284_new_n703_; 
wire _abc_2284_new_n704_; 
wire _abc_2284_new_n706_; 
wire _abc_2284_new_n707_; 
wire _abc_2284_new_n709_; 
wire _abc_2284_new_n710_; 
wire _abc_2284_new_n711_; 
wire _abc_2284_new_n712_; 
wire _abc_2284_new_n714_; 
wire _abc_2284_new_n715_; 
wire _abc_2284_new_n716_; 
wire _abc_2284_new_n717_; 
wire _abc_2284_new_n719_; 
wire _abc_2284_new_n720_; 
wire _abc_2284_new_n721_; 
wire _abc_2284_new_n722_; 
wire _abc_2284_new_n724_; 
wire _abc_2284_new_n725_; 
wire _abc_2284_new_n726_; 
wire _abc_2284_new_n727_; 
wire _abc_2284_new_n729_; 
wire _abc_2284_new_n730_; 
wire _abc_2284_new_n731_; 
wire _abc_2284_new_n732_; 
wire _abc_2284_new_n734_; 
wire _abc_2284_new_n735_; 
wire _abc_2284_new_n736_; 
wire _abc_2284_new_n737_; 
wire _abc_2284_new_n739_; 
wire _abc_2284_new_n740_; 
wire _abc_2284_new_n741_; 
wire _abc_2284_new_n742_; 
wire _abc_2284_new_n744_; 
wire _abc_2284_new_n745_; 
wire _abc_2284_new_n746_; 
input clk;
output is_receiving;
output is_transmitting;
output received;
output recv_error;
wire recv_state_0_; 
wire recv_state_1_; 
wire recv_state_2_; 
input rst;
input rx;
wire rx_bits_remaining_0_; 
wire rx_bits_remaining_1_; 
wire rx_bits_remaining_2_; 
wire rx_bits_remaining_3_; 
output \rx_byte[0] ;
output \rx_byte[1] ;
output \rx_byte[2] ;
output \rx_byte[3] ;
output \rx_byte[4] ;
output \rx_byte[5] ;
output \rx_byte[6] ;
output \rx_byte[7] ;
wire rx_clk_divider_0_; 
wire rx_clk_divider_10_; 
wire rx_clk_divider_1_; 
wire rx_clk_divider_2_; 
wire rx_clk_divider_3_; 
wire rx_clk_divider_4_; 
wire rx_clk_divider_5_; 
wire rx_clk_divider_6_; 
wire rx_clk_divider_7_; 
wire rx_clk_divider_8_; 
wire rx_clk_divider_9_; 
wire rx_countdown_0_; 
wire rx_countdown_1_; 
wire rx_countdown_2_; 
wire rx_countdown_3_; 
wire rx_countdown_4_; 
wire rx_countdown_5_; 
input transmit;
output tx;
wire tx_bits_remaining_0_; 
wire tx_bits_remaining_1_; 
wire tx_bits_remaining_2_; 
wire tx_bits_remaining_3_; 
input \tx_byte[0] ;
input \tx_byte[1] ;
input \tx_byte[2] ;
input \tx_byte[3] ;
input \tx_byte[4] ;
input \tx_byte[5] ;
input \tx_byte[6] ;
input \tx_byte[7] ;
wire tx_clk_divider_0_; 
wire tx_clk_divider_10_; 
wire tx_clk_divider_1_; 
wire tx_clk_divider_2_; 
wire tx_clk_divider_3_; 
wire tx_clk_divider_4_; 
wire tx_clk_divider_5_; 
wire tx_clk_divider_6_; 
wire tx_clk_divider_7_; 
wire tx_clk_divider_8_; 
wire tx_clk_divider_9_; 
wire tx_countdown_0_; 
wire tx_countdown_1_; 
wire tx_countdown_2_; 
wire tx_countdown_3_; 
wire tx_countdown_4_; 
wire tx_countdown_5_; 
wire tx_data_0_; 
wire tx_data_1_; 
wire tx_data_2_; 
wire tx_data_3_; 
wire tx_data_4_; 
wire tx_data_5_; 
wire tx_data_6_; 
wire tx_data_7_; 
wire tx_state_0_; 
wire tx_state_1_; 
AND2X2 AND2X2_1 ( .A(_abc_2284_new_n144_), .B(_abc_2284_new_n145_), .Y(_abc_2284_new_n146_));
AND2X2 AND2X2_10 ( .A(_abc_2284_new_n164_), .B(_abc_2284_new_n167_), .Y(_abc_2284_new_n168_));
AND2X2 AND2X2_100 ( .A(_abc_2284_new_n293_), .B(\tx_byte[4] ), .Y(_abc_2284_new_n329_));
AND2X2 AND2X2_101 ( .A(_abc_2284_new_n297_), .B(tx_data_4_), .Y(_abc_2284_new_n330_));
AND2X2 AND2X2_102 ( .A(_abc_2284_new_n284_), .B(tx_data_5_), .Y(_abc_2284_new_n333_));
AND2X2 AND2X2_103 ( .A(_abc_2284_new_n283_), .B(tx_data_6_), .Y(_abc_2284_new_n334_));
AND2X2 AND2X2_104 ( .A(_abc_2284_new_n335_), .B(_abc_2284_new_n158_), .Y(_abc_2284_new_n336_));
AND2X2 AND2X2_105 ( .A(_abc_2284_new_n293_), .B(\tx_byte[5] ), .Y(_abc_2284_new_n337_));
AND2X2 AND2X2_106 ( .A(_abc_2284_new_n297_), .B(tx_data_5_), .Y(_abc_2284_new_n338_));
AND2X2 AND2X2_107 ( .A(_abc_2284_new_n158_), .B(tx_data_7_), .Y(_abc_2284_new_n342_));
AND2X2 AND2X2_108 ( .A(_abc_2284_new_n284_), .B(_abc_2284_new_n158_), .Y(_abc_2284_new_n343_));
AND2X2 AND2X2_109 ( .A(_abc_2284_new_n344_), .B(_abc_2284_new_n341_), .Y(_abc_2284_new_n345_));
AND2X2 AND2X2_11 ( .A(_abc_2284_new_n169_), .B(_abc_2284_new_n170_), .Y(_abc_2284_new_n171_));
AND2X2 AND2X2_110 ( .A(_abc_2284_new_n293_), .B(\tx_byte[6] ), .Y(_abc_2284_new_n346_));
AND2X2 AND2X2_111 ( .A(_abc_2284_new_n297_), .B(tx_data_6_), .Y(_abc_2284_new_n347_));
AND2X2 AND2X2_112 ( .A(_abc_2284_new_n293_), .B(\tx_byte[7] ), .Y(_abc_2284_new_n350_));
AND2X2 AND2X2_113 ( .A(_abc_2284_new_n351_), .B(tx_data_7_), .Y(_abc_2284_new_n352_));
AND2X2 AND2X2_114 ( .A(_abc_2284_new_n158_), .B(_abc_2284_new_n282_), .Y(_abc_2284_new_n354_));
AND2X2 AND2X2_115 ( .A(_abc_2284_new_n279_), .B(_abc_2284_new_n355_), .Y(_abc_2284_new_n356_));
AND2X2 AND2X2_116 ( .A(_abc_2284_new_n357_), .B(tx_bits_remaining_0_), .Y(_abc_2284_new_n358_));
AND2X2 AND2X2_117 ( .A(_abc_2284_new_n359_), .B(_abc_2284_new_n354_), .Y(_abc_2284_new_n360_));
AND2X2 AND2X2_118 ( .A(_abc_2284_new_n297_), .B(tx_bits_remaining_0_), .Y(_abc_2284_new_n361_));
AND2X2 AND2X2_119 ( .A(_abc_2284_new_n279_), .B(_abc_2284_new_n363_), .Y(_abc_2284_new_n364_));
AND2X2 AND2X2_12 ( .A(_abc_2284_new_n172_), .B(_abc_2284_new_n173_), .Y(_abc_2284_new_n174_));
AND2X2 AND2X2_120 ( .A(_abc_2284_new_n364_), .B(_abc_2284_new_n281_), .Y(_abc_2284_new_n365_));
AND2X2 AND2X2_121 ( .A(_abc_2284_new_n366_), .B(tx_bits_remaining_1_), .Y(_abc_2284_new_n367_));
AND2X2 AND2X2_122 ( .A(_abc_2284_new_n368_), .B(_abc_2284_new_n158_), .Y(_abc_2284_new_n369_));
AND2X2 AND2X2_123 ( .A(_abc_2284_new_n297_), .B(tx_bits_remaining_1_), .Y(_abc_2284_new_n370_));
AND2X2 AND2X2_124 ( .A(_abc_2284_new_n364_), .B(_abc_2284_new_n372_), .Y(_abc_2284_new_n373_));
AND2X2 AND2X2_125 ( .A(_abc_2284_new_n158_), .B(tx_bits_remaining_3_), .Y(_abc_2284_new_n374_));
AND2X2 AND2X2_126 ( .A(_abc_2284_new_n373_), .B(_abc_2284_new_n374_), .Y(_abc_2284_new_n375_));
AND2X2 AND2X2_127 ( .A(_abc_2284_new_n376_), .B(_abc_2284_new_n158_), .Y(_abc_2284_new_n377_));
AND2X2 AND2X2_128 ( .A(_abc_2284_new_n378_), .B(tx_bits_remaining_2_), .Y(_abc_2284_new_n379_));
AND2X2 AND2X2_129 ( .A(_abc_2284_new_n373_), .B(_abc_2284_new_n158_), .Y(_abc_2284_new_n381_));
AND2X2 AND2X2_13 ( .A(_abc_2284_new_n171_), .B(_abc_2284_new_n174_), .Y(_abc_2284_new_n175_));
AND2X2 AND2X2_130 ( .A(_abc_2284_new_n382_), .B(tx_bits_remaining_3_), .Y(_abc_2284_new_n383_));
AND2X2 AND2X2_131 ( .A(_abc_2284_new_n385_), .B(_abc_2284_new_n386_), .Y(_0tx_countdown_5_0__0_));
AND2X2 AND2X2_132 ( .A(_abc_2284_new_n388_), .B(_abc_2284_new_n386_), .Y(_0tx_countdown_5_0__1_));
AND2X2 AND2X2_133 ( .A(_abc_2284_new_n279_), .B(_abc_2284_new_n354_), .Y(_abc_2284_new_n390_));
AND2X2 AND2X2_134 ( .A(_abc_2284_new_n279_), .B(_abc_2284_new_n395_), .Y(_abc_2284_new_n396_));
AND2X2 AND2X2_135 ( .A(_abc_2284_new_n396_), .B(_abc_2284_new_n158_), .Y(_abc_2284_new_n397_));
AND2X2 AND2X2_136 ( .A(_abc_2284_new_n351_), .B(_abc_2284_new_n398_), .Y(_0tx_countdown_5_0__3_));
AND2X2 AND2X2_137 ( .A(_abc_2284_new_n400_), .B(_abc_2284_new_n386_), .Y(_0tx_countdown_5_0__4_));
AND2X2 AND2X2_138 ( .A(_abc_2284_new_n402_), .B(_abc_2284_new_n386_), .Y(_0tx_countdown_5_0__5_));
AND2X2 AND2X2_139 ( .A(_abc_2284_new_n396_), .B(_abc_2284_new_n155_), .Y(_abc_2284_new_n404_));
AND2X2 AND2X2_14 ( .A(_abc_2284_new_n168_), .B(_abc_2284_new_n175_), .Y(_abc_2284_new_n176_));
AND2X2 AND2X2_140 ( .A(_abc_2284_new_n405_), .B(_abc_2284_new_n157_), .Y(_abc_2284_new_n406_));
AND2X2 AND2X2_141 ( .A(_abc_2284_new_n279_), .B(_abc_2284_new_n289_), .Y(_abc_2284_new_n409_));
AND2X2 AND2X2_142 ( .A(_abc_2284_new_n408_), .B(_abc_2284_new_n410_), .Y(_0tx_state_1_0__1_));
AND2X2 AND2X2_143 ( .A(_abc_2284_new_n283_), .B(_abc_2284_new_n412_), .Y(_abc_2284_new_n413_));
AND2X2 AND2X2_144 ( .A(_abc_2284_new_n415_), .B(_abc_2284_new_n158_), .Y(_abc_2284_new_n416_));
AND2X2 AND2X2_145 ( .A(_abc_2284_new_n414_), .B(_abc_2284_new_n416_), .Y(_abc_2284_new_n417_));
AND2X2 AND2X2_146 ( .A(_abc_2284_new_n297_), .B(tx), .Y(_abc_2284_new_n418_));
AND2X2 AND2X2_147 ( .A(_abc_2284_new_n424_), .B(_abc_2284_new_n425_), .Y(_abc_2284_new_n426_));
AND2X2 AND2X2_148 ( .A(_abc_2284_new_n435_), .B(_abc_2284_new_n436_), .Y(_abc_2284_new_n437_));
AND2X2 AND2X2_149 ( .A(_abc_2284_new_n437_), .B(_abc_2284_new_n434_), .Y(_abc_2284_new_n438_));
AND2X2 AND2X2_15 ( .A(_abc_2284_new_n176_), .B(_abc_2284_new_n161_), .Y(_abc_2284_new_n177_));
AND2X2 AND2X2_150 ( .A(_abc_2284_new_n439_), .B(_abc_2284_new_n432_), .Y(_abc_2284_new_n440_));
AND2X2 AND2X2_151 ( .A(_abc_2284_new_n441_), .B(rx_clk_divider_7_), .Y(_abc_2284_new_n442_));
AND2X2 AND2X2_152 ( .A(_abc_2284_new_n443_), .B(_abc_2284_new_n430_), .Y(_abc_2284_new_n444_));
AND2X2 AND2X2_153 ( .A(_abc_2284_new_n445_), .B(_abc_2284_new_n424_), .Y(_abc_2284_new_n446_));
AND2X2 AND2X2_154 ( .A(_abc_2284_new_n423_), .B(rx_clk_divider_4_), .Y(_abc_2284_new_n447_));
AND2X2 AND2X2_155 ( .A(_abc_2284_new_n451_), .B(rx_clk_divider_0_), .Y(_abc_2284_new_n452_));
AND2X2 AND2X2_156 ( .A(_abc_2284_new_n450_), .B(_abc_2284_new_n452_), .Y(_abc_2284_new_n453_));
AND2X2 AND2X2_157 ( .A(_abc_2284_new_n425_), .B(_abc_2284_new_n454_), .Y(_abc_2284_new_n455_));
AND2X2 AND2X2_158 ( .A(_abc_2284_new_n455_), .B(_abc_2284_new_n434_), .Y(_abc_2284_new_n456_));
AND2X2 AND2X2_159 ( .A(_abc_2284_new_n453_), .B(_abc_2284_new_n456_), .Y(_abc_2284_new_n457_));
AND2X2 AND2X2_16 ( .A(_abc_2284_new_n177_), .B(_abc_2284_new_n160_), .Y(_abc_2284_new_n178_));
AND2X2 AND2X2_160 ( .A(_abc_2284_new_n449_), .B(_abc_2284_new_n457_), .Y(_abc_2284_new_n458_));
AND2X2 AND2X2_161 ( .A(_abc_2284_new_n444_), .B(_abc_2284_new_n458_), .Y(_abc_2284_new_n459_));
AND2X2 AND2X2_162 ( .A(_abc_2284_new_n440_), .B(_abc_2284_new_n459_), .Y(_abc_2284_new_n460_));
AND2X2 AND2X2_163 ( .A(_abc_2284_new_n460_), .B(_abc_2284_new_n420_), .Y(_abc_2284_new_n461_));
AND2X2 AND2X2_164 ( .A(_abc_2284_new_n462_), .B(rx_countdown_0_), .Y(_abc_2284_new_n463_));
AND2X2 AND2X2_165 ( .A(_abc_2284_new_n461_), .B(_abc_2284_new_n464_), .Y(_abc_2284_new_n465_));
AND2X2 AND2X2_166 ( .A(is_receiving), .B(_abc_2284_new_n156_), .Y(_abc_2284_new_n467_));
AND2X2 AND2X2_167 ( .A(_abc_2284_new_n468_), .B(rx), .Y(_abc_2284_new_n469_));
AND2X2 AND2X2_168 ( .A(_abc_2284_new_n156_), .B(recv_state_2_), .Y(_abc_2284_new_n470_));
AND2X2 AND2X2_169 ( .A(_abc_2284_new_n470_), .B(_abc_2284_new_n144_), .Y(_abc_2284_new_n471_));
AND2X2 AND2X2_17 ( .A(_abc_2284_new_n179_), .B(_abc_2284_new_n159_), .Y(_abc_2284_new_n180_));
AND2X2 AND2X2_170 ( .A(_abc_2284_new_n156_), .B(recv_state_1_), .Y(_abc_2284_new_n472_));
AND2X2 AND2X2_171 ( .A(_abc_2284_new_n156_), .B(recv_state_0_), .Y(_abc_2284_new_n473_));
AND2X2 AND2X2_172 ( .A(_abc_2284_new_n473_), .B(_abc_2284_new_n145_), .Y(_abc_2284_new_n474_));
AND2X2 AND2X2_173 ( .A(_abc_2284_new_n466_), .B(_abc_2284_new_n477_), .Y(_0rx_countdown_5_0__0_));
AND2X2 AND2X2_174 ( .A(_abc_2284_new_n468_), .B(_abc_2284_new_n479_), .Y(_abc_2284_new_n480_));
AND2X2 AND2X2_175 ( .A(_abc_2284_new_n481_), .B(rx_countdown_1_), .Y(_abc_2284_new_n482_));
AND2X2 AND2X2_176 ( .A(_abc_2284_new_n465_), .B(_abc_2284_new_n483_), .Y(_abc_2284_new_n484_));
AND2X2 AND2X2_177 ( .A(_abc_2284_new_n153_), .B(_abc_2284_new_n156_), .Y(_abc_2284_new_n486_));
AND2X2 AND2X2_178 ( .A(_abc_2284_new_n486_), .B(_abc_2284_new_n152_), .Y(_abc_2284_new_n487_));
AND2X2 AND2X2_179 ( .A(_abc_2284_new_n485_), .B(_abc_2284_new_n488_), .Y(_abc_2284_new_n489_));
AND2X2 AND2X2_18 ( .A(_abc_2284_new_n178_), .B(tx_clk_divider_10_), .Y(_abc_2284_new_n181_));
AND2X2 AND2X2_180 ( .A(_abc_2284_new_n146_), .B(_abc_2284_new_n472_), .Y(_abc_2284_new_n491_));
AND2X2 AND2X2_181 ( .A(_abc_2284_new_n432_), .B(_abc_2284_new_n420_), .Y(_abc_2284_new_n492_));
AND2X2 AND2X2_182 ( .A(_abc_2284_new_n438_), .B(_abc_2284_new_n433_), .Y(_abc_2284_new_n493_));
AND2X2 AND2X2_183 ( .A(_abc_2284_new_n493_), .B(rx_clk_divider_10_), .Y(_abc_2284_new_n494_));
AND2X2 AND2X2_184 ( .A(_abc_2284_new_n496_), .B(_abc_2284_new_n431_), .Y(_abc_2284_new_n497_));
AND2X2 AND2X2_185 ( .A(_abc_2284_new_n440_), .B(_abc_2284_new_n497_), .Y(_abc_2284_new_n498_));
AND2X2 AND2X2_186 ( .A(_abc_2284_new_n495_), .B(_abc_2284_new_n498_), .Y(_abc_2284_new_n499_));
AND2X2 AND2X2_187 ( .A(_abc_2284_new_n500_), .B(_abc_2284_new_n441_), .Y(_abc_2284_new_n501_));
AND2X2 AND2X2_188 ( .A(_abc_2284_new_n444_), .B(_abc_2284_new_n501_), .Y(_abc_2284_new_n502_));
AND2X2 AND2X2_189 ( .A(_abc_2284_new_n503_), .B(_abc_2284_new_n428_), .Y(_abc_2284_new_n504_));
AND2X2 AND2X2_19 ( .A(_abc_2284_new_n179_), .B(_abc_2284_new_n183_), .Y(_abc_2284_new_n184_));
AND2X2 AND2X2_190 ( .A(_abc_2284_new_n504_), .B(_abc_2284_new_n449_), .Y(_abc_2284_new_n505_));
AND2X2 AND2X2_191 ( .A(_abc_2284_new_n502_), .B(_abc_2284_new_n505_), .Y(_abc_2284_new_n506_));
AND2X2 AND2X2_192 ( .A(_abc_2284_new_n506_), .B(_abc_2284_new_n453_), .Y(_abc_2284_new_n507_));
AND2X2 AND2X2_193 ( .A(_abc_2284_new_n499_), .B(_abc_2284_new_n507_), .Y(_abc_2284_new_n508_));
AND2X2 AND2X2_194 ( .A(_abc_2284_new_n464_), .B(_abc_2284_new_n483_), .Y(_abc_2284_new_n509_));
AND2X2 AND2X2_195 ( .A(_abc_2284_new_n513_), .B(_abc_2284_new_n510_), .Y(_abc_2284_new_n514_));
AND2X2 AND2X2_196 ( .A(_abc_2284_new_n508_), .B(_abc_2284_new_n514_), .Y(_abc_2284_new_n515_));
AND2X2 AND2X2_197 ( .A(_abc_2284_new_n516_), .B(_abc_2284_new_n517_), .Y(_abc_2284_new_n518_));
AND2X2 AND2X2_198 ( .A(_abc_2284_new_n481_), .B(_abc_2284_new_n519_), .Y(_abc_2284_new_n520_));
AND2X2 AND2X2_199 ( .A(_abc_2284_new_n483_), .B(_abc_2284_new_n521_), .Y(_abc_2284_new_n522_));
AND2X2 AND2X2_2 ( .A(recv_state_1_), .B(recv_state_2_), .Y(_abc_2284_new_n150_));
AND2X2 AND2X2_20 ( .A(_abc_2284_new_n185_), .B(_abc_2284_new_n186_), .Y(_abc_2284_new_n187_));
AND2X2 AND2X2_200 ( .A(_abc_2284_new_n520_), .B(_abc_2284_new_n522_), .Y(_abc_2284_new_n523_));
AND2X2 AND2X2_201 ( .A(_abc_2284_new_n518_), .B(_abc_2284_new_n523_), .Y(_abc_2284_new_n524_));
AND2X2 AND2X2_202 ( .A(_abc_2284_new_n528_), .B(_abc_2284_new_n521_), .Y(_abc_2284_new_n529_));
AND2X2 AND2X2_203 ( .A(_abc_2284_new_n531_), .B(_abc_2284_new_n532_), .Y(_abc_2284_new_n533_));
AND2X2 AND2X2_204 ( .A(_abc_2284_new_n508_), .B(_abc_2284_new_n533_), .Y(_abc_2284_new_n534_));
AND2X2 AND2X2_205 ( .A(_abc_2284_new_n535_), .B(_abc_2284_new_n536_), .Y(_abc_2284_new_n537_));
AND2X2 AND2X2_206 ( .A(_abc_2284_new_n526_), .B(rx_countdown_3_), .Y(_abc_2284_new_n538_));
AND2X2 AND2X2_207 ( .A(_abc_2284_new_n508_), .B(_abc_2284_new_n539_), .Y(_abc_2284_new_n540_));
AND2X2 AND2X2_208 ( .A(_abc_2284_new_n541_), .B(_abc_2284_new_n543_), .Y(_abc_2284_new_n544_));
AND2X2 AND2X2_209 ( .A(_abc_2284_new_n537_), .B(_abc_2284_new_n544_), .Y(_abc_2284_new_n545_));
AND2X2 AND2X2_21 ( .A(_abc_2284_new_n184_), .B(_abc_2284_new_n187_), .Y(_abc_2284_new_n188_));
AND2X2 AND2X2_210 ( .A(_abc_2284_new_n545_), .B(_abc_2284_new_n524_), .Y(_abc_2284_new_n546_));
AND2X2 AND2X2_211 ( .A(_abc_2284_new_n546_), .B(_abc_2284_new_n491_), .Y(_abc_2284_new_n547_));
AND2X2 AND2X2_212 ( .A(_abc_2284_new_n474_), .B(_abc_2284_new_n152_), .Y(_abc_2284_new_n550_));
AND2X2 AND2X2_213 ( .A(_abc_2284_new_n546_), .B(_abc_2284_new_n479_), .Y(_abc_2284_new_n551_));
AND2X2 AND2X2_214 ( .A(_abc_2284_new_n551_), .B(_abc_2284_new_n550_), .Y(_abc_2284_new_n552_));
AND2X2 AND2X2_215 ( .A(_abc_2284_new_n553_), .B(_abc_2284_new_n477_), .Y(_abc_2284_new_n554_));
AND2X2 AND2X2_216 ( .A(_abc_2284_new_n557_), .B(_abc_2284_new_n477_), .Y(_abc_2284_new_n558_));
AND2X2 AND2X2_217 ( .A(_abc_2284_new_n450_), .B(rx_clk_divider_0_), .Y(_abc_2284_new_n560_));
AND2X2 AND2X2_218 ( .A(_abc_2284_new_n449_), .B(_abc_2284_new_n451_), .Y(_abc_2284_new_n561_));
AND2X2 AND2X2_219 ( .A(_abc_2284_new_n561_), .B(_abc_2284_new_n560_), .Y(_abc_2284_new_n562_));
AND2X2 AND2X2_22 ( .A(_abc_2284_new_n182_), .B(_abc_2284_new_n188_), .Y(_abc_2284_new_n189_));
AND2X2 AND2X2_220 ( .A(_abc_2284_new_n504_), .B(_abc_2284_new_n454_), .Y(_abc_2284_new_n563_));
AND2X2 AND2X2_221 ( .A(_abc_2284_new_n562_), .B(_abc_2284_new_n563_), .Y(_abc_2284_new_n564_));
AND2X2 AND2X2_222 ( .A(_abc_2284_new_n564_), .B(_abc_2284_new_n444_), .Y(_abc_2284_new_n565_));
AND2X2 AND2X2_223 ( .A(_abc_2284_new_n440_), .B(_abc_2284_new_n434_), .Y(_abc_2284_new_n566_));
AND2X2 AND2X2_224 ( .A(_abc_2284_new_n565_), .B(_abc_2284_new_n566_), .Y(_abc_2284_new_n567_));
AND2X2 AND2X2_225 ( .A(_abc_2284_new_n567_), .B(_abc_2284_new_n495_), .Y(_abc_2284_new_n568_));
AND2X2 AND2X2_226 ( .A(_abc_2284_new_n568_), .B(_abc_2284_new_n528_), .Y(_abc_2284_new_n569_));
AND2X2 AND2X2_227 ( .A(_abc_2284_new_n569_), .B(_abc_2284_new_n521_), .Y(_abc_2284_new_n570_));
AND2X2 AND2X2_228 ( .A(_abc_2284_new_n571_), .B(rx_countdown_4_), .Y(_abc_2284_new_n572_));
AND2X2 AND2X2_229 ( .A(_abc_2284_new_n573_), .B(_abc_2284_new_n477_), .Y(_0rx_countdown_5_0__4_));
AND2X2 AND2X2_23 ( .A(_abc_2284_new_n164_), .B(tx_clk_divider_0_), .Y(_abc_2284_new_n190_));
AND2X2 AND2X2_230 ( .A(_abc_2284_new_n575_), .B(_abc_2284_new_n477_), .Y(_0rx_countdown_5_0__5_));
AND2X2 AND2X2_231 ( .A(_abc_2284_new_n474_), .B(recv_state_1_), .Y(_abc_2284_new_n577_));
AND2X2 AND2X2_232 ( .A(_abc_2284_new_n578_), .B(_abc_2284_new_n473_), .Y(_abc_2284_new_n579_));
AND2X2 AND2X2_233 ( .A(_abc_2284_new_n580_), .B(_abc_2284_new_n577_), .Y(_abc_2284_new_n581_));
AND2X2 AND2X2_234 ( .A(_abc_2284_new_n582_), .B(rx_bits_remaining_0_), .Y(_abc_2284_new_n583_));
AND2X2 AND2X2_235 ( .A(_abc_2284_new_n584_), .B(_abc_2284_new_n585_), .Y(_abc_2284_new_n586_));
AND2X2 AND2X2_236 ( .A(_abc_2284_new_n586_), .B(_abc_2284_new_n583_), .Y(_abc_2284_new_n587_));
AND2X2 AND2X2_237 ( .A(_abc_2284_new_n546_), .B(_abc_2284_new_n587_), .Y(_abc_2284_new_n588_));
AND2X2 AND2X2_238 ( .A(_abc_2284_new_n589_), .B(_abc_2284_new_n491_), .Y(_abc_2284_new_n590_));
AND2X2 AND2X2_239 ( .A(_abc_2284_new_n591_), .B(_abc_2284_new_n550_), .Y(_abc_2284_new_n592_));
AND2X2 AND2X2_24 ( .A(_abc_2284_new_n190_), .B(_abc_2284_new_n165_), .Y(_abc_2284_new_n191_));
AND2X2 AND2X2_240 ( .A(_abc_2284_new_n472_), .B(_abc_2284_new_n153_), .Y(_abc_2284_new_n593_));
AND2X2 AND2X2_241 ( .A(_abc_2284_new_n591_), .B(_abc_2284_new_n577_), .Y(_abc_2284_new_n598_));
AND2X2 AND2X2_242 ( .A(_abc_2284_new_n546_), .B(rx), .Y(_abc_2284_new_n602_));
AND2X2 AND2X2_243 ( .A(_abc_2284_new_n602_), .B(_abc_2284_new_n550_), .Y(_abc_2284_new_n603_));
AND2X2 AND2X2_244 ( .A(_abc_2284_new_n546_), .B(_abc_2284_new_n577_), .Y(_abc_2284_new_n604_));
AND2X2 AND2X2_245 ( .A(_abc_2284_new_n578_), .B(_abc_2284_new_n606_), .Y(_abc_2284_new_n607_));
AND2X2 AND2X2_246 ( .A(_abc_2284_new_n607_), .B(_abc_2284_new_n471_), .Y(_abc_2284_new_n608_));
AND2X2 AND2X2_247 ( .A(_abc_2284_new_n546_), .B(_abc_2284_new_n611_), .Y(_abc_2284_new_n612_));
AND2X2 AND2X2_248 ( .A(_abc_2284_new_n578_), .B(rx_bits_remaining_0_), .Y(_abc_2284_new_n613_));
AND2X2 AND2X2_249 ( .A(_abc_2284_new_n614_), .B(_abc_2284_new_n491_), .Y(_abc_2284_new_n615_));
AND2X2 AND2X2_25 ( .A(_abc_2284_new_n168_), .B(_abc_2284_new_n171_), .Y(_abc_2284_new_n193_));
AND2X2 AND2X2_250 ( .A(_abc_2284_new_n616_), .B(rx_bits_remaining_0_), .Y(_abc_2284_new_n617_));
AND2X2 AND2X2_251 ( .A(_abc_2284_new_n619_), .B(rx_bits_remaining_1_), .Y(_abc_2284_new_n620_));
AND2X2 AND2X2_252 ( .A(_abc_2284_new_n611_), .B(_abc_2284_new_n582_), .Y(_abc_2284_new_n621_));
AND2X2 AND2X2_253 ( .A(_abc_2284_new_n546_), .B(_abc_2284_new_n621_), .Y(_abc_2284_new_n622_));
AND2X2 AND2X2_254 ( .A(_abc_2284_new_n623_), .B(_abc_2284_new_n491_), .Y(_abc_2284_new_n624_));
AND2X2 AND2X2_255 ( .A(_abc_2284_new_n616_), .B(rx_bits_remaining_1_), .Y(_abc_2284_new_n625_));
AND2X2 AND2X2_256 ( .A(_abc_2284_new_n622_), .B(_abc_2284_new_n584_), .Y(_abc_2284_new_n627_));
AND2X2 AND2X2_257 ( .A(_abc_2284_new_n628_), .B(rx_bits_remaining_2_), .Y(_abc_2284_new_n629_));
AND2X2 AND2X2_258 ( .A(_abc_2284_new_n630_), .B(_abc_2284_new_n491_), .Y(_abc_2284_new_n631_));
AND2X2 AND2X2_259 ( .A(_abc_2284_new_n616_), .B(rx_bits_remaining_2_), .Y(_abc_2284_new_n632_));
AND2X2 AND2X2_26 ( .A(_abc_2284_new_n193_), .B(_abc_2284_new_n172_), .Y(_abc_2284_new_n194_));
AND2X2 AND2X2_260 ( .A(_abc_2284_new_n627_), .B(rx_bits_remaining_3_), .Y(_abc_2284_new_n634_));
AND2X2 AND2X2_261 ( .A(_abc_2284_new_n636_), .B(_abc_2284_new_n491_), .Y(_abc_2284_new_n637_));
AND2X2 AND2X2_262 ( .A(_abc_2284_new_n637_), .B(_abc_2284_new_n635_), .Y(_abc_2284_new_n638_));
AND2X2 AND2X2_263 ( .A(_abc_2284_new_n639_), .B(rx_bits_remaining_3_), .Y(_abc_2284_new_n640_));
AND2X2 AND2X2_264 ( .A(_abc_2284_new_n386_), .B(_abc_2284_new_n166_), .Y(_0tx_clk_divider_10_0__0_));
AND2X2 AND2X2_265 ( .A(tx_clk_divider_1_), .B(tx_clk_divider_0_), .Y(_abc_2284_new_n644_));
AND2X2 AND2X2_266 ( .A(_abc_2284_new_n167_), .B(_abc_2284_new_n162_), .Y(_abc_2284_new_n648_));
AND2X2 AND2X2_267 ( .A(_abc_2284_new_n198_), .B(tx_clk_divider_2_), .Y(_abc_2284_new_n649_));
AND2X2 AND2X2_268 ( .A(_abc_2284_new_n653_), .B(tx_clk_divider_3_), .Y(_abc_2284_new_n654_));
AND2X2 AND2X2_269 ( .A(_abc_2284_new_n655_), .B(_abc_2284_new_n386_), .Y(_0tx_clk_divider_10_0__3_));
AND2X2 AND2X2_27 ( .A(_abc_2284_new_n195_), .B(_abc_2284_new_n192_), .Y(_abc_2284_new_n196_));
AND2X2 AND2X2_270 ( .A(_abc_2284_new_n660_), .B(_abc_2284_new_n386_), .Y(_0tx_clk_divider_10_0__5_));
AND2X2 AND2X2_271 ( .A(_abc_2284_new_n662_), .B(_abc_2284_new_n386_), .Y(_0tx_clk_divider_10_0__6_));
AND2X2 AND2X2_272 ( .A(_abc_2284_new_n664_), .B(_abc_2284_new_n386_), .Y(_0tx_clk_divider_10_0__7_));
AND2X2 AND2X2_273 ( .A(_abc_2284_new_n669_), .B(_abc_2284_new_n386_), .Y(_0tx_clk_divider_10_0__9_));
AND2X2 AND2X2_274 ( .A(_abc_2284_new_n675_), .B(_abc_2284_new_n674_), .Y(_0rx_clk_divider_10_0__0_));
AND2X2 AND2X2_275 ( .A(rx_clk_divider_1_), .B(rx_clk_divider_0_), .Y(_abc_2284_new_n678_));
AND2X2 AND2X2_276 ( .A(_abc_2284_new_n677_), .B(_abc_2284_new_n682_), .Y(_abc_2284_new_n683_));
AND2X2 AND2X2_277 ( .A(_abc_2284_new_n422_), .B(rx_clk_divider_2_), .Y(_abc_2284_new_n684_));
AND2X2 AND2X2_278 ( .A(_abc_2284_new_n688_), .B(rx_clk_divider_3_), .Y(_abc_2284_new_n689_));
AND2X2 AND2X2_279 ( .A(_abc_2284_new_n675_), .B(_abc_2284_new_n690_), .Y(_0rx_clk_divider_10_0__3_));
AND2X2 AND2X2_28 ( .A(_abc_2284_new_n203_), .B(_abc_2284_new_n202_), .Y(_abc_2284_new_n204_));
AND2X2 AND2X2_280 ( .A(_abc_2284_new_n694_), .B(_abc_2284_new_n675_), .Y(_0rx_clk_divider_10_0__5_));
AND2X2 AND2X2_281 ( .A(_abc_2284_new_n696_), .B(_abc_2284_new_n675_), .Y(_0rx_clk_divider_10_0__6_));
AND2X2 AND2X2_282 ( .A(_abc_2284_new_n698_), .B(_abc_2284_new_n675_), .Y(_0rx_clk_divider_10_0__7_));
AND2X2 AND2X2_283 ( .A(_abc_2284_new_n431_), .B(rx_clk_divider_9_), .Y(_abc_2284_new_n703_));
AND2X2 AND2X2_284 ( .A(_abc_2284_new_n704_), .B(_abc_2284_new_n675_), .Y(_0rx_clk_divider_10_0__9_));
AND2X2 AND2X2_285 ( .A(_abc_2284_new_n547_), .B(_abc_2284_new_n710_), .Y(_abc_2284_new_n711_));
AND2X2 AND2X2_286 ( .A(_abc_2284_new_n712_), .B(_abc_2284_new_n709_), .Y(_0rx_data_7_0__0_));
AND2X2 AND2X2_287 ( .A(_abc_2284_new_n547_), .B(_abc_2284_new_n715_), .Y(_abc_2284_new_n716_));
AND2X2 AND2X2_288 ( .A(_abc_2284_new_n717_), .B(_abc_2284_new_n714_), .Y(_0rx_data_7_0__1_));
AND2X2 AND2X2_289 ( .A(_abc_2284_new_n547_), .B(_abc_2284_new_n720_), .Y(_abc_2284_new_n721_));
AND2X2 AND2X2_29 ( .A(_abc_2284_new_n196_), .B(_abc_2284_new_n204_), .Y(_abc_2284_new_n205_));
AND2X2 AND2X2_290 ( .A(_abc_2284_new_n722_), .B(_abc_2284_new_n719_), .Y(_0rx_data_7_0__2_));
AND2X2 AND2X2_291 ( .A(_abc_2284_new_n547_), .B(_abc_2284_new_n725_), .Y(_abc_2284_new_n726_));
AND2X2 AND2X2_292 ( .A(_abc_2284_new_n727_), .B(_abc_2284_new_n724_), .Y(_0rx_data_7_0__3_));
AND2X2 AND2X2_293 ( .A(_abc_2284_new_n547_), .B(_abc_2284_new_n730_), .Y(_abc_2284_new_n731_));
AND2X2 AND2X2_294 ( .A(_abc_2284_new_n732_), .B(_abc_2284_new_n729_), .Y(_0rx_data_7_0__4_));
AND2X2 AND2X2_295 ( .A(_abc_2284_new_n547_), .B(_abc_2284_new_n735_), .Y(_abc_2284_new_n736_));
AND2X2 AND2X2_296 ( .A(_abc_2284_new_n737_), .B(_abc_2284_new_n734_), .Y(_0rx_data_7_0__5_));
AND2X2 AND2X2_297 ( .A(_abc_2284_new_n547_), .B(_abc_2284_new_n740_), .Y(_abc_2284_new_n741_));
AND2X2 AND2X2_298 ( .A(_abc_2284_new_n742_), .B(_abc_2284_new_n739_), .Y(_0rx_data_7_0__6_));
AND2X2 AND2X2_299 ( .A(_abc_2284_new_n547_), .B(_abc_2284_new_n479_), .Y(_abc_2284_new_n744_));
AND2X2 AND2X2_3 ( .A(_abc_2284_new_n150_), .B(_abc_2284_new_n144_), .Y(received));
AND2X2 AND2X2_30 ( .A(_abc_2284_new_n168_), .B(_abc_2284_new_n169_), .Y(_abc_2284_new_n206_));
AND2X2 AND2X2_300 ( .A(_abc_2284_new_n745_), .B(_abc_2284_new_n746_), .Y(_0rx_data_7_0__7_));
AND2X2 AND2X2_31 ( .A(_abc_2284_new_n207_), .B(_abc_2284_new_n201_), .Y(_abc_2284_new_n208_));
AND2X2 AND2X2_32 ( .A(_abc_2284_new_n210_), .B(_abc_2284_new_n209_), .Y(_abc_2284_new_n211_));
AND2X2 AND2X2_33 ( .A(_abc_2284_new_n208_), .B(_abc_2284_new_n211_), .Y(_abc_2284_new_n212_));
AND2X2 AND2X2_34 ( .A(_abc_2284_new_n205_), .B(_abc_2284_new_n212_), .Y(_abc_2284_new_n213_));
AND2X2 AND2X2_35 ( .A(_abc_2284_new_n213_), .B(_abc_2284_new_n191_), .Y(_abc_2284_new_n214_));
AND2X2 AND2X2_36 ( .A(_abc_2284_new_n214_), .B(_abc_2284_new_n189_), .Y(_abc_2284_new_n215_));
AND2X2 AND2X2_37 ( .A(_abc_2284_new_n216_), .B(_abc_2284_new_n217_), .Y(_abc_2284_new_n218_));
AND2X2 AND2X2_38 ( .A(tx_countdown_0_), .B(tx_countdown_1_), .Y(_abc_2284_new_n219_));
AND2X2 AND2X2_39 ( .A(_abc_2284_new_n215_), .B(_abc_2284_new_n220_), .Y(_abc_2284_new_n221_));
AND2X2 AND2X2_4 ( .A(recv_state_0_), .B(recv_state_2_), .Y(_abc_2284_new_n153_));
AND2X2 AND2X2_40 ( .A(_abc_2284_new_n222_), .B(_abc_2284_new_n223_), .Y(_abc_2284_new_n224_));
AND2X2 AND2X2_41 ( .A(_abc_2284_new_n211_), .B(_abc_2284_new_n191_), .Y(_abc_2284_new_n225_));
AND2X2 AND2X2_42 ( .A(_abc_2284_new_n208_), .B(_abc_2284_new_n225_), .Y(_abc_2284_new_n226_));
AND2X2 AND2X2_43 ( .A(_abc_2284_new_n204_), .B(_abc_2284_new_n161_), .Y(_abc_2284_new_n227_));
AND2X2 AND2X2_44 ( .A(_abc_2284_new_n226_), .B(_abc_2284_new_n227_), .Y(_abc_2284_new_n228_));
AND2X2 AND2X2_45 ( .A(_abc_2284_new_n228_), .B(_abc_2284_new_n196_), .Y(_abc_2284_new_n229_));
AND2X2 AND2X2_46 ( .A(_abc_2284_new_n229_), .B(_abc_2284_new_n184_), .Y(_abc_2284_new_n230_));
AND2X2 AND2X2_47 ( .A(_abc_2284_new_n230_), .B(_abc_2284_new_n182_), .Y(_abc_2284_new_n231_));
AND2X2 AND2X2_48 ( .A(_abc_2284_new_n231_), .B(_abc_2284_new_n216_), .Y(_abc_2284_new_n232_));
AND2X2 AND2X2_49 ( .A(_abc_2284_new_n233_), .B(_abc_2284_new_n234_), .Y(_abc_2284_new_n235_));
AND2X2 AND2X2_5 ( .A(_abc_2284_new_n153_), .B(_abc_2284_new_n152_), .Y(recv_error));
AND2X2 AND2X2_50 ( .A(_abc_2284_new_n235_), .B(_abc_2284_new_n224_), .Y(_abc_2284_new_n236_));
AND2X2 AND2X2_51 ( .A(_abc_2284_new_n218_), .B(_abc_2284_new_n237_), .Y(_abc_2284_new_n238_));
AND2X2 AND2X2_52 ( .A(_abc_2284_new_n242_), .B(_abc_2284_new_n239_), .Y(_abc_2284_new_n243_));
AND2X2 AND2X2_53 ( .A(_abc_2284_new_n215_), .B(_abc_2284_new_n243_), .Y(_abc_2284_new_n244_));
AND2X2 AND2X2_54 ( .A(_abc_2284_new_n245_), .B(_abc_2284_new_n246_), .Y(_abc_2284_new_n247_));
AND2X2 AND2X2_55 ( .A(_abc_2284_new_n250_), .B(_abc_2284_new_n248_), .Y(_abc_2284_new_n251_));
AND2X2 AND2X2_56 ( .A(_abc_2284_new_n215_), .B(_abc_2284_new_n251_), .Y(_abc_2284_new_n252_));
AND2X2 AND2X2_57 ( .A(_abc_2284_new_n253_), .B(_abc_2284_new_n254_), .Y(_abc_2284_new_n255_));
AND2X2 AND2X2_58 ( .A(_abc_2284_new_n247_), .B(_abc_2284_new_n255_), .Y(_abc_2284_new_n256_));
AND2X2 AND2X2_59 ( .A(_abc_2284_new_n236_), .B(_abc_2284_new_n256_), .Y(_abc_2284_new_n257_));
AND2X2 AND2X2_6 ( .A(_abc_2284_new_n156_), .B(tx_state_0_), .Y(_abc_2284_new_n157_));
AND2X2 AND2X2_60 ( .A(_abc_2284_new_n237_), .B(_abc_2284_new_n240_), .Y(_abc_2284_new_n259_));
AND2X2 AND2X2_61 ( .A(_abc_2284_new_n218_), .B(_abc_2284_new_n259_), .Y(_abc_2284_new_n260_));
AND2X2 AND2X2_62 ( .A(_abc_2284_new_n260_), .B(_abc_2284_new_n258_), .Y(_abc_2284_new_n261_));
AND2X2 AND2X2_63 ( .A(_abc_2284_new_n262_), .B(tx_countdown_5_), .Y(_abc_2284_new_n263_));
AND2X2 AND2X2_64 ( .A(_abc_2284_new_n261_), .B(_abc_2284_new_n264_), .Y(_abc_2284_new_n265_));
AND2X2 AND2X2_65 ( .A(_abc_2284_new_n215_), .B(_abc_2284_new_n266_), .Y(_abc_2284_new_n267_));
AND2X2 AND2X2_66 ( .A(_abc_2284_new_n268_), .B(_abc_2284_new_n269_), .Y(_abc_2284_new_n270_));
AND2X2 AND2X2_67 ( .A(_abc_2284_new_n271_), .B(tx_countdown_4_), .Y(_abc_2284_new_n272_));
AND2X2 AND2X2_68 ( .A(_abc_2284_new_n215_), .B(_abc_2284_new_n273_), .Y(_abc_2284_new_n274_));
AND2X2 AND2X2_69 ( .A(_abc_2284_new_n275_), .B(_abc_2284_new_n276_), .Y(_abc_2284_new_n277_));
AND2X2 AND2X2_7 ( .A(_abc_2284_new_n157_), .B(_abc_2284_new_n155_), .Y(_abc_2284_new_n158_));
AND2X2 AND2X2_70 ( .A(_abc_2284_new_n270_), .B(_abc_2284_new_n277_), .Y(_abc_2284_new_n278_));
AND2X2 AND2X2_71 ( .A(_abc_2284_new_n257_), .B(_abc_2284_new_n278_), .Y(_abc_2284_new_n279_));
AND2X2 AND2X2_72 ( .A(_abc_2284_new_n279_), .B(_abc_2284_new_n282_), .Y(_abc_2284_new_n283_));
AND2X2 AND2X2_73 ( .A(_abc_2284_new_n284_), .B(tx_data_0_), .Y(_abc_2284_new_n285_));
AND2X2 AND2X2_74 ( .A(_abc_2284_new_n283_), .B(tx_data_1_), .Y(_abc_2284_new_n286_));
AND2X2 AND2X2_75 ( .A(_abc_2284_new_n287_), .B(_abc_2284_new_n158_), .Y(_abc_2284_new_n288_));
AND2X2 AND2X2_76 ( .A(_abc_2284_new_n156_), .B(tx_state_1_), .Y(_abc_2284_new_n290_));
AND2X2 AND2X2_77 ( .A(_abc_2284_new_n289_), .B(_abc_2284_new_n291_), .Y(_abc_2284_new_n292_));
AND2X2 AND2X2_78 ( .A(_abc_2284_new_n292_), .B(transmit), .Y(_abc_2284_new_n293_));
AND2X2 AND2X2_79 ( .A(_abc_2284_new_n293_), .B(\tx_byte[0] ), .Y(_abc_2284_new_n294_));
AND2X2 AND2X2_8 ( .A(_abc_2284_new_n162_), .B(_abc_2284_new_n163_), .Y(_abc_2284_new_n164_));
AND2X2 AND2X2_80 ( .A(_abc_2284_new_n292_), .B(_abc_2284_new_n295_), .Y(_abc_2284_new_n296_));
AND2X2 AND2X2_81 ( .A(_abc_2284_new_n297_), .B(tx_data_0_), .Y(_abc_2284_new_n298_));
AND2X2 AND2X2_82 ( .A(_abc_2284_new_n284_), .B(tx_data_1_), .Y(_abc_2284_new_n301_));
AND2X2 AND2X2_83 ( .A(_abc_2284_new_n283_), .B(tx_data_2_), .Y(_abc_2284_new_n302_));
AND2X2 AND2X2_84 ( .A(_abc_2284_new_n303_), .B(_abc_2284_new_n158_), .Y(_abc_2284_new_n304_));
AND2X2 AND2X2_85 ( .A(_abc_2284_new_n293_), .B(\tx_byte[1] ), .Y(_abc_2284_new_n305_));
AND2X2 AND2X2_86 ( .A(_abc_2284_new_n297_), .B(tx_data_1_), .Y(_abc_2284_new_n306_));
AND2X2 AND2X2_87 ( .A(_abc_2284_new_n284_), .B(tx_data_2_), .Y(_abc_2284_new_n309_));
AND2X2 AND2X2_88 ( .A(_abc_2284_new_n283_), .B(tx_data_3_), .Y(_abc_2284_new_n310_));
AND2X2 AND2X2_89 ( .A(_abc_2284_new_n311_), .B(_abc_2284_new_n158_), .Y(_abc_2284_new_n312_));
AND2X2 AND2X2_9 ( .A(_abc_2284_new_n165_), .B(_abc_2284_new_n166_), .Y(_abc_2284_new_n167_));
AND2X2 AND2X2_90 ( .A(_abc_2284_new_n293_), .B(\tx_byte[2] ), .Y(_abc_2284_new_n313_));
AND2X2 AND2X2_91 ( .A(_abc_2284_new_n297_), .B(tx_data_2_), .Y(_abc_2284_new_n314_));
AND2X2 AND2X2_92 ( .A(_abc_2284_new_n284_), .B(tx_data_3_), .Y(_abc_2284_new_n317_));
AND2X2 AND2X2_93 ( .A(_abc_2284_new_n283_), .B(tx_data_4_), .Y(_abc_2284_new_n318_));
AND2X2 AND2X2_94 ( .A(_abc_2284_new_n319_), .B(_abc_2284_new_n158_), .Y(_abc_2284_new_n320_));
AND2X2 AND2X2_95 ( .A(_abc_2284_new_n293_), .B(\tx_byte[3] ), .Y(_abc_2284_new_n321_));
AND2X2 AND2X2_96 ( .A(_abc_2284_new_n297_), .B(tx_data_3_), .Y(_abc_2284_new_n322_));
AND2X2 AND2X2_97 ( .A(_abc_2284_new_n284_), .B(tx_data_4_), .Y(_abc_2284_new_n325_));
AND2X2 AND2X2_98 ( .A(_abc_2284_new_n283_), .B(tx_data_5_), .Y(_abc_2284_new_n326_));
AND2X2 AND2X2_99 ( .A(_abc_2284_new_n327_), .B(_abc_2284_new_n158_), .Y(_abc_2284_new_n328_));
DFFPOSX1 DFFPOSX1_1 ( .CLK(clk), .D(_0rx_clk_divider_10_0__6_), .Q(rx_clk_divider_6_));
DFFPOSX1 DFFPOSX1_10 ( .CLK(clk), .D(_0tx_clk_divider_10_0__4_), .Q(tx_clk_divider_4_));
DFFPOSX1 DFFPOSX1_11 ( .CLK(clk), .D(_0tx_clk_divider_10_0__5_), .Q(tx_clk_divider_5_));
DFFPOSX1 DFFPOSX1_12 ( .CLK(clk), .D(_0tx_clk_divider_10_0__6_), .Q(tx_clk_divider_6_));
DFFPOSX1 DFFPOSX1_13 ( .CLK(clk), .D(_0tx_clk_divider_10_0__7_), .Q(tx_clk_divider_7_));
DFFPOSX1 DFFPOSX1_14 ( .CLK(clk), .D(_0tx_clk_divider_10_0__8_), .Q(tx_clk_divider_8_));
DFFPOSX1 DFFPOSX1_15 ( .CLK(clk), .D(_0tx_clk_divider_10_0__9_), .Q(tx_clk_divider_9_));
DFFPOSX1 DFFPOSX1_16 ( .CLK(clk), .D(_0tx_clk_divider_10_0__10_), .Q(tx_clk_divider_10_));
DFFPOSX1 DFFPOSX1_17 ( .CLK(clk), .D(_0recv_state_2_0__0_), .Q(recv_state_0_));
DFFPOSX1 DFFPOSX1_18 ( .CLK(clk), .D(_0recv_state_2_0__1_), .Q(recv_state_1_));
DFFPOSX1 DFFPOSX1_19 ( .CLK(clk), .D(_0recv_state_2_0__2_), .Q(recv_state_2_));
DFFPOSX1 DFFPOSX1_2 ( .CLK(clk), .D(_0rx_clk_divider_10_0__7_), .Q(rx_clk_divider_7_));
DFFPOSX1 DFFPOSX1_20 ( .CLK(clk), .D(_0rx_countdown_5_0__0_), .Q(rx_countdown_0_));
DFFPOSX1 DFFPOSX1_21 ( .CLK(clk), .D(_0rx_countdown_5_0__1_), .Q(rx_countdown_1_));
DFFPOSX1 DFFPOSX1_22 ( .CLK(clk), .D(_0rx_countdown_5_0__2_), .Q(rx_countdown_2_));
DFFPOSX1 DFFPOSX1_23 ( .CLK(clk), .D(_0rx_countdown_5_0__3_), .Q(rx_countdown_3_));
DFFPOSX1 DFFPOSX1_24 ( .CLK(clk), .D(_0rx_countdown_5_0__4_), .Q(rx_countdown_4_));
DFFPOSX1 DFFPOSX1_25 ( .CLK(clk), .D(_0rx_countdown_5_0__5_), .Q(rx_countdown_5_));
DFFPOSX1 DFFPOSX1_26 ( .CLK(clk), .D(_0rx_bits_remaining_3_0__0_), .Q(rx_bits_remaining_0_));
DFFPOSX1 DFFPOSX1_27 ( .CLK(clk), .D(_0rx_bits_remaining_3_0__1_), .Q(rx_bits_remaining_1_));
DFFPOSX1 DFFPOSX1_28 ( .CLK(clk), .D(_0rx_bits_remaining_3_0__2_), .Q(rx_bits_remaining_2_));
DFFPOSX1 DFFPOSX1_29 ( .CLK(clk), .D(_0rx_bits_remaining_3_0__3_), .Q(rx_bits_remaining_3_));
DFFPOSX1 DFFPOSX1_3 ( .CLK(clk), .D(_0rx_clk_divider_10_0__8_), .Q(rx_clk_divider_8_));
DFFPOSX1 DFFPOSX1_30 ( .CLK(clk), .D(_0rx_data_7_0__0_), .Q(\rx_byte[0] ));
DFFPOSX1 DFFPOSX1_31 ( .CLK(clk), .D(_0rx_data_7_0__1_), .Q(\rx_byte[1] ));
DFFPOSX1 DFFPOSX1_32 ( .CLK(clk), .D(_0rx_data_7_0__2_), .Q(\rx_byte[2] ));
DFFPOSX1 DFFPOSX1_33 ( .CLK(clk), .D(_0rx_data_7_0__3_), .Q(\rx_byte[3] ));
DFFPOSX1 DFFPOSX1_34 ( .CLK(clk), .D(_0rx_data_7_0__4_), .Q(\rx_byte[4] ));
DFFPOSX1 DFFPOSX1_35 ( .CLK(clk), .D(_0rx_data_7_0__5_), .Q(\rx_byte[5] ));
DFFPOSX1 DFFPOSX1_36 ( .CLK(clk), .D(_0rx_data_7_0__6_), .Q(\rx_byte[6] ));
DFFPOSX1 DFFPOSX1_37 ( .CLK(clk), .D(_0rx_data_7_0__7_), .Q(\rx_byte[7] ));
DFFPOSX1 DFFPOSX1_38 ( .CLK(clk), .D(_0tx_out_0_0_), .Q(tx));
DFFPOSX1 DFFPOSX1_39 ( .CLK(clk), .D(_0tx_state_1_0__0_), .Q(tx_state_0_));
DFFPOSX1 DFFPOSX1_4 ( .CLK(clk), .D(_0rx_clk_divider_10_0__9_), .Q(rx_clk_divider_9_));
DFFPOSX1 DFFPOSX1_40 ( .CLK(clk), .D(_0tx_state_1_0__1_), .Q(tx_state_1_));
DFFPOSX1 DFFPOSX1_41 ( .CLK(clk), .D(_0tx_countdown_5_0__0_), .Q(tx_countdown_0_));
DFFPOSX1 DFFPOSX1_42 ( .CLK(clk), .D(_0tx_countdown_5_0__1_), .Q(tx_countdown_1_));
DFFPOSX1 DFFPOSX1_43 ( .CLK(clk), .D(_0tx_countdown_5_0__2_), .Q(tx_countdown_2_));
DFFPOSX1 DFFPOSX1_44 ( .CLK(clk), .D(_0tx_countdown_5_0__3_), .Q(tx_countdown_3_));
DFFPOSX1 DFFPOSX1_45 ( .CLK(clk), .D(_0tx_countdown_5_0__4_), .Q(tx_countdown_4_));
DFFPOSX1 DFFPOSX1_46 ( .CLK(clk), .D(_0tx_countdown_5_0__5_), .Q(tx_countdown_5_));
DFFPOSX1 DFFPOSX1_47 ( .CLK(clk), .D(_0tx_bits_remaining_3_0__0_), .Q(tx_bits_remaining_0_));
DFFPOSX1 DFFPOSX1_48 ( .CLK(clk), .D(_0tx_bits_remaining_3_0__1_), .Q(tx_bits_remaining_1_));
DFFPOSX1 DFFPOSX1_49 ( .CLK(clk), .D(_0tx_bits_remaining_3_0__2_), .Q(tx_bits_remaining_2_));
DFFPOSX1 DFFPOSX1_5 ( .CLK(clk), .D(_0rx_clk_divider_10_0__10_), .Q(rx_clk_divider_10_));
DFFPOSX1 DFFPOSX1_50 ( .CLK(clk), .D(_0tx_bits_remaining_3_0__3_), .Q(tx_bits_remaining_3_));
DFFPOSX1 DFFPOSX1_51 ( .CLK(clk), .D(_0tx_data_7_0__0_), .Q(tx_data_0_));
DFFPOSX1 DFFPOSX1_52 ( .CLK(clk), .D(_0tx_data_7_0__1_), .Q(tx_data_1_));
DFFPOSX1 DFFPOSX1_53 ( .CLK(clk), .D(_0tx_data_7_0__2_), .Q(tx_data_2_));
DFFPOSX1 DFFPOSX1_54 ( .CLK(clk), .D(_0tx_data_7_0__3_), .Q(tx_data_3_));
DFFPOSX1 DFFPOSX1_55 ( .CLK(clk), .D(_0tx_data_7_0__4_), .Q(tx_data_4_));
DFFPOSX1 DFFPOSX1_56 ( .CLK(clk), .D(_0tx_data_7_0__5_), .Q(tx_data_5_));
DFFPOSX1 DFFPOSX1_57 ( .CLK(clk), .D(_0tx_data_7_0__6_), .Q(tx_data_6_));
DFFPOSX1 DFFPOSX1_58 ( .CLK(clk), .D(_0tx_data_7_0__7_), .Q(tx_data_7_));
DFFPOSX1 DFFPOSX1_59 ( .CLK(clk), .D(_0rx_clk_divider_10_0__0_), .Q(rx_clk_divider_0_));
DFFPOSX1 DFFPOSX1_6 ( .CLK(clk), .D(_0tx_clk_divider_10_0__0_), .Q(tx_clk_divider_0_));
DFFPOSX1 DFFPOSX1_60 ( .CLK(clk), .D(_0rx_clk_divider_10_0__1_), .Q(rx_clk_divider_1_));
DFFPOSX1 DFFPOSX1_61 ( .CLK(clk), .D(_0rx_clk_divider_10_0__2_), .Q(rx_clk_divider_2_));
DFFPOSX1 DFFPOSX1_62 ( .CLK(clk), .D(_0rx_clk_divider_10_0__3_), .Q(rx_clk_divider_3_));
DFFPOSX1 DFFPOSX1_63 ( .CLK(clk), .D(_0rx_clk_divider_10_0__4_), .Q(rx_clk_divider_4_));
DFFPOSX1 DFFPOSX1_64 ( .CLK(clk), .D(_0rx_clk_divider_10_0__5_), .Q(rx_clk_divider_5_));
DFFPOSX1 DFFPOSX1_7 ( .CLK(clk), .D(_0tx_clk_divider_10_0__1_), .Q(tx_clk_divider_1_));
DFFPOSX1 DFFPOSX1_8 ( .CLK(clk), .D(_0tx_clk_divider_10_0__2_), .Q(tx_clk_divider_2_));
DFFPOSX1 DFFPOSX1_9 ( .CLK(clk), .D(_0tx_clk_divider_10_0__3_), .Q(tx_clk_divider_3_));
INVX1 INVX1_1 ( .A(recv_state_0_), .Y(_abc_2284_new_n144_));
INVX1 INVX1_10 ( .A(tx_clk_divider_2_), .Y(_abc_2284_new_n162_));
INVX1 INVX1_100 ( .A(_abc_2284_new_n551_), .Y(_abc_2284_new_n591_));
INVX1 INVX1_101 ( .A(_abc_2284_new_n472_), .Y(_abc_2284_new_n606_));
INVX1 INVX1_102 ( .A(rx_bits_remaining_0_), .Y(_abc_2284_new_n611_));
INVX1 INVX1_103 ( .A(_abc_2284_new_n599_), .Y(_abc_2284_new_n616_));
INVX1 INVX1_104 ( .A(_abc_2284_new_n612_), .Y(_abc_2284_new_n619_));
INVX1 INVX1_105 ( .A(_abc_2284_new_n622_), .Y(_abc_2284_new_n628_));
INVX1 INVX1_106 ( .A(_abc_2284_new_n634_), .Y(_abc_2284_new_n635_));
INVX1 INVX1_107 ( .A(_abc_2284_new_n491_), .Y(_abc_2284_new_n639_));
INVX1 INVX1_108 ( .A(_abc_2284_new_n648_), .Y(_abc_2284_new_n653_));
INVX1 INVX1_109 ( .A(_abc_2284_new_n211_), .Y(_abc_2284_new_n657_));
INVX1 INVX1_11 ( .A(tx_clk_divider_3_), .Y(_abc_2284_new_n163_));
INVX1 INVX1_110 ( .A(_abc_2284_new_n208_), .Y(_abc_2284_new_n660_));
INVX1 INVX1_111 ( .A(_abc_2284_new_n204_), .Y(_abc_2284_new_n662_));
INVX1 INVX1_112 ( .A(_abc_2284_new_n196_), .Y(_abc_2284_new_n664_));
INVX1 INVX1_113 ( .A(_abc_2284_new_n187_), .Y(_abc_2284_new_n666_));
INVX1 INVX1_114 ( .A(_abc_2284_new_n184_), .Y(_abc_2284_new_n669_));
INVX1 INVX1_115 ( .A(_abc_2284_new_n182_), .Y(_abc_2284_new_n671_));
INVX1 INVX1_116 ( .A(rx_clk_divider_0_), .Y(_abc_2284_new_n674_));
INVX1 INVX1_117 ( .A(_abc_2284_new_n480_), .Y(_abc_2284_new_n675_));
INVX1 INVX1_118 ( .A(_abc_2284_new_n422_), .Y(_abc_2284_new_n677_));
INVX1 INVX1_119 ( .A(rx_clk_divider_2_), .Y(_abc_2284_new_n682_));
INVX1 INVX1_12 ( .A(tx_clk_divider_1_), .Y(_abc_2284_new_n165_));
INVX1 INVX1_120 ( .A(_abc_2284_new_n683_), .Y(_abc_2284_new_n688_));
INVX1 INVX1_121 ( .A(_abc_2284_new_n504_), .Y(_abc_2284_new_n694_));
INVX1 INVX1_122 ( .A(_abc_2284_new_n501_), .Y(_abc_2284_new_n696_));
INVX1 INVX1_123 ( .A(_abc_2284_new_n497_), .Y(_abc_2284_new_n700_));
INVX1 INVX1_124 ( .A(_abc_2284_new_n495_), .Y(_abc_2284_new_n706_));
INVX1 INVX1_125 ( .A(\rx_byte[1] ), .Y(_abc_2284_new_n710_));
INVX1 INVX1_126 ( .A(_abc_2284_new_n711_), .Y(_abc_2284_new_n712_));
INVX1 INVX1_127 ( .A(\rx_byte[2] ), .Y(_abc_2284_new_n715_));
INVX1 INVX1_128 ( .A(_abc_2284_new_n716_), .Y(_abc_2284_new_n717_));
INVX1 INVX1_129 ( .A(\rx_byte[3] ), .Y(_abc_2284_new_n720_));
INVX1 INVX1_13 ( .A(tx_clk_divider_0_), .Y(_abc_2284_new_n166_));
INVX1 INVX1_130 ( .A(_abc_2284_new_n721_), .Y(_abc_2284_new_n722_));
INVX1 INVX1_131 ( .A(\rx_byte[4] ), .Y(_abc_2284_new_n725_));
INVX1 INVX1_132 ( .A(_abc_2284_new_n726_), .Y(_abc_2284_new_n727_));
INVX1 INVX1_133 ( .A(\rx_byte[5] ), .Y(_abc_2284_new_n730_));
INVX1 INVX1_134 ( .A(_abc_2284_new_n731_), .Y(_abc_2284_new_n732_));
INVX1 INVX1_135 ( .A(\rx_byte[6] ), .Y(_abc_2284_new_n735_));
INVX1 INVX1_136 ( .A(_abc_2284_new_n736_), .Y(_abc_2284_new_n737_));
INVX1 INVX1_137 ( .A(\rx_byte[7] ), .Y(_abc_2284_new_n740_));
INVX1 INVX1_138 ( .A(_abc_2284_new_n741_), .Y(_abc_2284_new_n742_));
INVX1 INVX1_139 ( .A(_abc_2284_new_n744_), .Y(_abc_2284_new_n745_));
INVX1 INVX1_14 ( .A(tx_clk_divider_4_), .Y(_abc_2284_new_n169_));
INVX1 INVX1_15 ( .A(tx_clk_divider_5_), .Y(_abc_2284_new_n170_));
INVX1 INVX1_16 ( .A(tx_clk_divider_6_), .Y(_abc_2284_new_n172_));
INVX1 INVX1_17 ( .A(tx_clk_divider_7_), .Y(_abc_2284_new_n173_));
INVX1 INVX1_18 ( .A(_abc_2284_new_n178_), .Y(_abc_2284_new_n179_));
INVX1 INVX1_19 ( .A(_abc_2284_new_n177_), .Y(_abc_2284_new_n185_));
INVX1 INVX1_2 ( .A(recv_state_2_), .Y(_abc_2284_new_n145_));
INVX1 INVX1_20 ( .A(_abc_2284_new_n176_), .Y(_abc_2284_new_n192_));
INVX1 INVX1_21 ( .A(_abc_2284_new_n171_), .Y(_abc_2284_new_n200_));
INVX1 INVX1_22 ( .A(tx_countdown_0_), .Y(_abc_2284_new_n216_));
INVX1 INVX1_23 ( .A(tx_countdown_1_), .Y(_abc_2284_new_n217_));
INVX1 INVX1_24 ( .A(_abc_2284_new_n221_), .Y(_abc_2284_new_n222_));
INVX1 INVX1_25 ( .A(_abc_2284_new_n232_), .Y(_abc_2284_new_n233_));
INVX1 INVX1_26 ( .A(tx_countdown_2_), .Y(_abc_2284_new_n237_));
INVX1 INVX1_27 ( .A(tx_countdown_3_), .Y(_abc_2284_new_n240_));
INVX1 INVX1_28 ( .A(_abc_2284_new_n238_), .Y(_abc_2284_new_n241_));
INVX1 INVX1_29 ( .A(_abc_2284_new_n244_), .Y(_abc_2284_new_n245_));
INVX1 INVX1_3 ( .A(_abc_2284_new_n146_), .Y(_abc_2284_new_n147_));
INVX1 INVX1_30 ( .A(_abc_2284_new_n218_), .Y(_abc_2284_new_n249_));
INVX1 INVX1_31 ( .A(_abc_2284_new_n252_), .Y(_abc_2284_new_n253_));
INVX1 INVX1_32 ( .A(tx_countdown_4_), .Y(_abc_2284_new_n258_));
INVX1 INVX1_33 ( .A(_abc_2284_new_n261_), .Y(_abc_2284_new_n262_));
INVX1 INVX1_34 ( .A(tx_countdown_5_), .Y(_abc_2284_new_n264_));
INVX1 INVX1_35 ( .A(_abc_2284_new_n267_), .Y(_abc_2284_new_n268_));
INVX1 INVX1_36 ( .A(_abc_2284_new_n260_), .Y(_abc_2284_new_n271_));
INVX1 INVX1_37 ( .A(_abc_2284_new_n274_), .Y(_abc_2284_new_n275_));
INVX1 INVX1_38 ( .A(_abc_2284_new_n283_), .Y(_abc_2284_new_n284_));
INVX1 INVX1_39 ( .A(_abc_2284_new_n157_), .Y(_abc_2284_new_n289_));
INVX1 INVX1_4 ( .A(recv_state_1_), .Y(_abc_2284_new_n152_));
INVX1 INVX1_40 ( .A(_abc_2284_new_n290_), .Y(_abc_2284_new_n291_));
INVX1 INVX1_41 ( .A(transmit), .Y(_abc_2284_new_n295_));
INVX1 INVX1_42 ( .A(tx_bits_remaining_0_), .Y(_abc_2284_new_n355_));
INVX1 INVX1_43 ( .A(_abc_2284_new_n279_), .Y(_abc_2284_new_n357_));
INVX1 INVX1_44 ( .A(_abc_2284_new_n280_), .Y(_abc_2284_new_n363_));
INVX1 INVX1_45 ( .A(_abc_2284_new_n356_), .Y(_abc_2284_new_n366_));
INVX1 INVX1_46 ( .A(tx_bits_remaining_2_), .Y(_abc_2284_new_n372_));
INVX1 INVX1_47 ( .A(_abc_2284_new_n364_), .Y(_abc_2284_new_n376_));
INVX1 INVX1_48 ( .A(_abc_2284_new_n381_), .Y(_abc_2284_new_n382_));
INVX1 INVX1_49 ( .A(_abc_2284_new_n235_), .Y(_abc_2284_new_n385_));
INVX1 INVX1_5 ( .A(tx_state_1_), .Y(_abc_2284_new_n155_));
INVX1 INVX1_50 ( .A(_abc_2284_new_n293_), .Y(_abc_2284_new_n386_));
INVX1 INVX1_51 ( .A(_abc_2284_new_n224_), .Y(_abc_2284_new_n388_));
INVX1 INVX1_52 ( .A(_abc_2284_new_n255_), .Y(_abc_2284_new_n391_));
INVX1 INVX1_53 ( .A(_abc_2284_new_n247_), .Y(_abc_2284_new_n394_));
INVX1 INVX1_54 ( .A(_abc_2284_new_n282_), .Y(_abc_2284_new_n395_));
INVX1 INVX1_55 ( .A(_abc_2284_new_n277_), .Y(_abc_2284_new_n400_));
INVX1 INVX1_56 ( .A(_abc_2284_new_n270_), .Y(_abc_2284_new_n402_));
INVX1 INVX1_57 ( .A(_abc_2284_new_n404_), .Y(_abc_2284_new_n405_));
INVX1 INVX1_58 ( .A(_abc_2284_new_n409_), .Y(_abc_2284_new_n410_));
INVX1 INVX1_59 ( .A(tx_data_0_), .Y(_abc_2284_new_n412_));
INVX1 INVX1_6 ( .A(rst), .Y(_abc_2284_new_n156_));
INVX1 INVX1_60 ( .A(_abc_2284_new_n413_), .Y(_abc_2284_new_n414_));
INVX1 INVX1_61 ( .A(rx_clk_divider_10_), .Y(_abc_2284_new_n420_));
INVX1 INVX1_62 ( .A(rx_clk_divider_4_), .Y(_abc_2284_new_n424_));
INVX1 INVX1_63 ( .A(rx_clk_divider_5_), .Y(_abc_2284_new_n425_));
INVX1 INVX1_64 ( .A(_abc_2284_new_n426_), .Y(_abc_2284_new_n427_));
INVX1 INVX1_65 ( .A(rx_clk_divider_9_), .Y(_abc_2284_new_n433_));
INVX1 INVX1_66 ( .A(rx_clk_divider_8_), .Y(_abc_2284_new_n434_));
INVX1 INVX1_67 ( .A(_abc_2284_new_n428_), .Y(_abc_2284_new_n435_));
INVX1 INVX1_68 ( .A(_abc_2284_new_n429_), .Y(_abc_2284_new_n436_));
INVX1 INVX1_69 ( .A(_abc_2284_new_n442_), .Y(_abc_2284_new_n443_));
INVX1 INVX1_7 ( .A(tx_clk_divider_10_), .Y(_abc_2284_new_n159_));
INVX1 INVX1_70 ( .A(_abc_2284_new_n423_), .Y(_abc_2284_new_n445_));
INVX1 INVX1_71 ( .A(_abc_2284_new_n448_), .Y(_abc_2284_new_n449_));
INVX1 INVX1_72 ( .A(_abc_2284_new_n421_), .Y(_abc_2284_new_n450_));
INVX1 INVX1_73 ( .A(rx_clk_divider_1_), .Y(_abc_2284_new_n451_));
INVX1 INVX1_74 ( .A(rx_clk_divider_6_), .Y(_abc_2284_new_n454_));
INVX1 INVX1_75 ( .A(_abc_2284_new_n461_), .Y(_abc_2284_new_n462_));
INVX1 INVX1_76 ( .A(rx_countdown_0_), .Y(_abc_2284_new_n464_));
INVX1 INVX1_77 ( .A(_abc_2284_new_n467_), .Y(_abc_2284_new_n468_));
INVX1 INVX1_78 ( .A(rx), .Y(_abc_2284_new_n479_));
INVX1 INVX1_79 ( .A(_abc_2284_new_n465_), .Y(_abc_2284_new_n481_));
INVX1 INVX1_8 ( .A(tx_clk_divider_9_), .Y(_abc_2284_new_n160_));
INVX1 INVX1_80 ( .A(rx_countdown_1_), .Y(_abc_2284_new_n483_));
INVX1 INVX1_81 ( .A(_abc_2284_new_n487_), .Y(_abc_2284_new_n488_));
INVX1 INVX1_82 ( .A(rx_countdown_2_), .Y(_abc_2284_new_n511_));
INVX1 INVX1_83 ( .A(_abc_2284_new_n509_), .Y(_abc_2284_new_n512_));
INVX1 INVX1_84 ( .A(_abc_2284_new_n515_), .Y(_abc_2284_new_n516_));
INVX1 INVX1_85 ( .A(rx_countdown_4_), .Y(_abc_2284_new_n521_));
INVX1 INVX1_86 ( .A(rx_countdown_5_), .Y(_abc_2284_new_n525_));
INVX1 INVX1_87 ( .A(_abc_2284_new_n527_), .Y(_abc_2284_new_n528_));
INVX1 INVX1_88 ( .A(_abc_2284_new_n529_), .Y(_abc_2284_new_n530_));
INVX1 INVX1_89 ( .A(_abc_2284_new_n534_), .Y(_abc_2284_new_n535_));
INVX1 INVX1_9 ( .A(tx_clk_divider_8_), .Y(_abc_2284_new_n161_));
INVX1 INVX1_90 ( .A(_abc_2284_new_n540_), .Y(_abc_2284_new_n541_));
INVX1 INVX1_91 ( .A(rx_countdown_3_), .Y(_abc_2284_new_n542_));
INVX1 INVX1_92 ( .A(_abc_2284_new_n517_), .Y(_abc_2284_new_n548_));
INVX1 INVX1_93 ( .A(_abc_2284_new_n543_), .Y(_abc_2284_new_n556_));
INVX1 INVX1_94 ( .A(_abc_2284_new_n569_), .Y(_abc_2284_new_n571_));
INVX1 INVX1_95 ( .A(_abc_2284_new_n537_), .Y(_abc_2284_new_n575_));
INVX1 INVX1_96 ( .A(_abc_2284_new_n546_), .Y(_abc_2284_new_n578_));
INVX1 INVX1_97 ( .A(rx_bits_remaining_1_), .Y(_abc_2284_new_n582_));
INVX1 INVX1_98 ( .A(rx_bits_remaining_2_), .Y(_abc_2284_new_n584_));
INVX1 INVX1_99 ( .A(rx_bits_remaining_3_), .Y(_abc_2284_new_n585_));
OR2X2 OR2X2_1 ( .A(_abc_2284_new_n147_), .B(recv_state_1_), .Y(is_receiving));
OR2X2 OR2X2_10 ( .A(_abc_2284_new_n199_), .B(_abc_2284_new_n200_), .Y(_abc_2284_new_n201_));
OR2X2 OR2X2_100 ( .A(_abc_2284_new_n508_), .B(_abc_2284_new_n525_), .Y(_abc_2284_new_n536_));
OR2X2 OR2X2_101 ( .A(_abc_2284_new_n528_), .B(_abc_2284_new_n538_), .Y(_abc_2284_new_n539_));
OR2X2 OR2X2_102 ( .A(_abc_2284_new_n508_), .B(_abc_2284_new_n542_), .Y(_abc_2284_new_n543_));
OR2X2 OR2X2_103 ( .A(_abc_2284_new_n548_), .B(_abc_2284_new_n515_), .Y(_abc_2284_new_n549_));
OR2X2 OR2X2_104 ( .A(_abc_2284_new_n552_), .B(_abc_2284_new_n549_), .Y(_abc_2284_new_n553_));
OR2X2 OR2X2_105 ( .A(_abc_2284_new_n554_), .B(_abc_2284_new_n547_), .Y(_0rx_countdown_5_0__2_));
OR2X2 OR2X2_106 ( .A(_abc_2284_new_n556_), .B(_abc_2284_new_n540_), .Y(_abc_2284_new_n557_));
OR2X2 OR2X2_107 ( .A(_abc_2284_new_n558_), .B(_abc_2284_new_n487_), .Y(_0rx_countdown_5_0__3_));
OR2X2 OR2X2_108 ( .A(_abc_2284_new_n572_), .B(_abc_2284_new_n570_), .Y(_abc_2284_new_n573_));
OR2X2 OR2X2_109 ( .A(_abc_2284_new_n579_), .B(_abc_2284_new_n551_), .Y(_abc_2284_new_n580_));
OR2X2 OR2X2_11 ( .A(_abc_2284_new_n201_), .B(tx_clk_divider_6_), .Y(_abc_2284_new_n202_));
OR2X2 OR2X2_110 ( .A(_abc_2284_new_n579_), .B(_abc_2284_new_n588_), .Y(_abc_2284_new_n589_));
OR2X2 OR2X2_111 ( .A(_abc_2284_new_n480_), .B(_abc_2284_new_n593_), .Y(_abc_2284_new_n594_));
OR2X2 OR2X2_112 ( .A(_abc_2284_new_n592_), .B(_abc_2284_new_n594_), .Y(_abc_2284_new_n595_));
OR2X2 OR2X2_113 ( .A(_abc_2284_new_n595_), .B(_abc_2284_new_n590_), .Y(_abc_2284_new_n596_));
OR2X2 OR2X2_114 ( .A(_abc_2284_new_n596_), .B(_abc_2284_new_n581_), .Y(_0recv_state_2_0__0_));
OR2X2 OR2X2_115 ( .A(_abc_2284_new_n552_), .B(_abc_2284_new_n491_), .Y(_abc_2284_new_n599_));
OR2X2 OR2X2_116 ( .A(_abc_2284_new_n599_), .B(_abc_2284_new_n598_), .Y(_abc_2284_new_n600_));
OR2X2 OR2X2_117 ( .A(_abc_2284_new_n600_), .B(_abc_2284_new_n593_), .Y(_0recv_state_2_0__1_));
OR2X2 OR2X2_118 ( .A(_abc_2284_new_n603_), .B(_abc_2284_new_n604_), .Y(_abc_2284_new_n605_));
OR2X2 OR2X2_119 ( .A(_abc_2284_new_n608_), .B(_abc_2284_new_n486_), .Y(_abc_2284_new_n609_));
OR2X2 OR2X2_12 ( .A(_abc_2284_new_n193_), .B(_abc_2284_new_n172_), .Y(_abc_2284_new_n203_));
OR2X2 OR2X2_120 ( .A(_abc_2284_new_n609_), .B(_abc_2284_new_n605_), .Y(_0recv_state_2_0__2_));
OR2X2 OR2X2_121 ( .A(_abc_2284_new_n613_), .B(_abc_2284_new_n612_), .Y(_abc_2284_new_n614_));
OR2X2 OR2X2_122 ( .A(_abc_2284_new_n617_), .B(_abc_2284_new_n615_), .Y(_0rx_bits_remaining_3_0__0_));
OR2X2 OR2X2_123 ( .A(_abc_2284_new_n620_), .B(_abc_2284_new_n622_), .Y(_abc_2284_new_n623_));
OR2X2 OR2X2_124 ( .A(_abc_2284_new_n624_), .B(_abc_2284_new_n625_), .Y(_0rx_bits_remaining_3_0__1_));
OR2X2 OR2X2_125 ( .A(_abc_2284_new_n629_), .B(_abc_2284_new_n627_), .Y(_abc_2284_new_n630_));
OR2X2 OR2X2_126 ( .A(_abc_2284_new_n631_), .B(_abc_2284_new_n632_), .Y(_0rx_bits_remaining_3_0__2_));
OR2X2 OR2X2_127 ( .A(_abc_2284_new_n627_), .B(rx_bits_remaining_3_), .Y(_abc_2284_new_n636_));
OR2X2 OR2X2_128 ( .A(_abc_2284_new_n552_), .B(_abc_2284_new_n640_), .Y(_abc_2284_new_n641_));
OR2X2 OR2X2_129 ( .A(_abc_2284_new_n638_), .B(_abc_2284_new_n641_), .Y(_0rx_bits_remaining_3_0__3_));
OR2X2 OR2X2_13 ( .A(_abc_2284_new_n206_), .B(_abc_2284_new_n170_), .Y(_abc_2284_new_n207_));
OR2X2 OR2X2_130 ( .A(_abc_2284_new_n167_), .B(_abc_2284_new_n644_), .Y(_abc_2284_new_n645_));
OR2X2 OR2X2_131 ( .A(_abc_2284_new_n293_), .B(_abc_2284_new_n645_), .Y(_abc_2284_new_n646_));
OR2X2 OR2X2_132 ( .A(_abc_2284_new_n231_), .B(_abc_2284_new_n646_), .Y(_0tx_clk_divider_10_0__1_));
OR2X2 OR2X2_133 ( .A(_abc_2284_new_n648_), .B(_abc_2284_new_n649_), .Y(_abc_2284_new_n650_));
OR2X2 OR2X2_134 ( .A(_abc_2284_new_n293_), .B(_abc_2284_new_n650_), .Y(_abc_2284_new_n651_));
OR2X2 OR2X2_135 ( .A(_abc_2284_new_n231_), .B(_abc_2284_new_n651_), .Y(_0tx_clk_divider_10_0__2_));
OR2X2 OR2X2_136 ( .A(_abc_2284_new_n654_), .B(_abc_2284_new_n168_), .Y(_abc_2284_new_n655_));
OR2X2 OR2X2_137 ( .A(_abc_2284_new_n657_), .B(_abc_2284_new_n293_), .Y(_abc_2284_new_n658_));
OR2X2 OR2X2_138 ( .A(_abc_2284_new_n231_), .B(_abc_2284_new_n658_), .Y(_0tx_clk_divider_10_0__4_));
OR2X2 OR2X2_139 ( .A(_abc_2284_new_n666_), .B(_abc_2284_new_n293_), .Y(_abc_2284_new_n667_));
OR2X2 OR2X2_14 ( .A(_abc_2284_new_n199_), .B(tx_clk_divider_4_), .Y(_abc_2284_new_n209_));
OR2X2 OR2X2_140 ( .A(_abc_2284_new_n231_), .B(_abc_2284_new_n667_), .Y(_0tx_clk_divider_10_0__8_));
OR2X2 OR2X2_141 ( .A(_abc_2284_new_n230_), .B(_abc_2284_new_n293_), .Y(_abc_2284_new_n672_));
OR2X2 OR2X2_142 ( .A(_abc_2284_new_n672_), .B(_abc_2284_new_n671_), .Y(_0tx_clk_divider_10_0__10_));
OR2X2 OR2X2_143 ( .A(_abc_2284_new_n677_), .B(_abc_2284_new_n678_), .Y(_abc_2284_new_n679_));
OR2X2 OR2X2_144 ( .A(_abc_2284_new_n480_), .B(_abc_2284_new_n679_), .Y(_abc_2284_new_n680_));
OR2X2 OR2X2_145 ( .A(_abc_2284_new_n461_), .B(_abc_2284_new_n680_), .Y(_0rx_clk_divider_10_0__1_));
OR2X2 OR2X2_146 ( .A(_abc_2284_new_n683_), .B(_abc_2284_new_n684_), .Y(_abc_2284_new_n685_));
OR2X2 OR2X2_147 ( .A(_abc_2284_new_n480_), .B(_abc_2284_new_n685_), .Y(_abc_2284_new_n686_));
OR2X2 OR2X2_148 ( .A(_abc_2284_new_n461_), .B(_abc_2284_new_n686_), .Y(_0rx_clk_divider_10_0__2_));
OR2X2 OR2X2_149 ( .A(_abc_2284_new_n689_), .B(_abc_2284_new_n445_), .Y(_abc_2284_new_n690_));
OR2X2 OR2X2_15 ( .A(_abc_2284_new_n168_), .B(_abc_2284_new_n169_), .Y(_abc_2284_new_n210_));
OR2X2 OR2X2_150 ( .A(_abc_2284_new_n480_), .B(_abc_2284_new_n448_), .Y(_abc_2284_new_n692_));
OR2X2 OR2X2_151 ( .A(_abc_2284_new_n461_), .B(_abc_2284_new_n692_), .Y(_0rx_clk_divider_10_0__4_));
OR2X2 OR2X2_152 ( .A(_abc_2284_new_n442_), .B(_abc_2284_new_n437_), .Y(_abc_2284_new_n698_));
OR2X2 OR2X2_153 ( .A(_abc_2284_new_n700_), .B(_abc_2284_new_n480_), .Y(_abc_2284_new_n701_));
OR2X2 OR2X2_154 ( .A(_abc_2284_new_n461_), .B(_abc_2284_new_n701_), .Y(_0rx_clk_divider_10_0__8_));
OR2X2 OR2X2_155 ( .A(_abc_2284_new_n493_), .B(_abc_2284_new_n703_), .Y(_abc_2284_new_n704_));
OR2X2 OR2X2_156 ( .A(_abc_2284_new_n460_), .B(_abc_2284_new_n480_), .Y(_abc_2284_new_n707_));
OR2X2 OR2X2_157 ( .A(_abc_2284_new_n707_), .B(_abc_2284_new_n706_), .Y(_0rx_clk_divider_10_0__10_));
OR2X2 OR2X2_158 ( .A(_abc_2284_new_n547_), .B(\rx_byte[0] ), .Y(_abc_2284_new_n709_));
OR2X2 OR2X2_159 ( .A(_abc_2284_new_n547_), .B(\rx_byte[1] ), .Y(_abc_2284_new_n714_));
OR2X2 OR2X2_16 ( .A(_abc_2284_new_n218_), .B(_abc_2284_new_n219_), .Y(_abc_2284_new_n220_));
OR2X2 OR2X2_160 ( .A(_abc_2284_new_n547_), .B(\rx_byte[2] ), .Y(_abc_2284_new_n719_));
OR2X2 OR2X2_161 ( .A(_abc_2284_new_n547_), .B(\rx_byte[3] ), .Y(_abc_2284_new_n724_));
OR2X2 OR2X2_162 ( .A(_abc_2284_new_n547_), .B(\rx_byte[4] ), .Y(_abc_2284_new_n729_));
OR2X2 OR2X2_163 ( .A(_abc_2284_new_n547_), .B(\rx_byte[5] ), .Y(_abc_2284_new_n734_));
OR2X2 OR2X2_164 ( .A(_abc_2284_new_n547_), .B(\rx_byte[6] ), .Y(_abc_2284_new_n739_));
OR2X2 OR2X2_165 ( .A(_abc_2284_new_n547_), .B(\rx_byte[7] ), .Y(_abc_2284_new_n746_));
OR2X2 OR2X2_17 ( .A(_abc_2284_new_n215_), .B(_abc_2284_new_n217_), .Y(_abc_2284_new_n223_));
OR2X2 OR2X2_18 ( .A(_abc_2284_new_n231_), .B(_abc_2284_new_n216_), .Y(_abc_2284_new_n234_));
OR2X2 OR2X2_19 ( .A(_abc_2284_new_n238_), .B(tx_countdown_3_), .Y(_abc_2284_new_n239_));
OR2X2 OR2X2_2 ( .A(tx_state_1_), .B(tx_state_0_), .Y(is_transmitting));
OR2X2 OR2X2_20 ( .A(_abc_2284_new_n241_), .B(_abc_2284_new_n240_), .Y(_abc_2284_new_n242_));
OR2X2 OR2X2_21 ( .A(_abc_2284_new_n215_), .B(_abc_2284_new_n240_), .Y(_abc_2284_new_n246_));
OR2X2 OR2X2_22 ( .A(_abc_2284_new_n218_), .B(tx_countdown_2_), .Y(_abc_2284_new_n248_));
OR2X2 OR2X2_23 ( .A(_abc_2284_new_n249_), .B(_abc_2284_new_n237_), .Y(_abc_2284_new_n250_));
OR2X2 OR2X2_24 ( .A(_abc_2284_new_n215_), .B(_abc_2284_new_n237_), .Y(_abc_2284_new_n254_));
OR2X2 OR2X2_25 ( .A(_abc_2284_new_n263_), .B(_abc_2284_new_n265_), .Y(_abc_2284_new_n266_));
OR2X2 OR2X2_26 ( .A(_abc_2284_new_n215_), .B(_abc_2284_new_n264_), .Y(_abc_2284_new_n269_));
OR2X2 OR2X2_27 ( .A(_abc_2284_new_n272_), .B(_abc_2284_new_n261_), .Y(_abc_2284_new_n273_));
OR2X2 OR2X2_28 ( .A(_abc_2284_new_n215_), .B(_abc_2284_new_n258_), .Y(_abc_2284_new_n276_));
OR2X2 OR2X2_29 ( .A(tx_bits_remaining_1_), .B(tx_bits_remaining_0_), .Y(_abc_2284_new_n280_));
OR2X2 OR2X2_3 ( .A(_abc_2284_new_n180_), .B(_abc_2284_new_n181_), .Y(_abc_2284_new_n182_));
OR2X2 OR2X2_30 ( .A(tx_bits_remaining_3_), .B(tx_bits_remaining_2_), .Y(_abc_2284_new_n281_));
OR2X2 OR2X2_31 ( .A(_abc_2284_new_n280_), .B(_abc_2284_new_n281_), .Y(_abc_2284_new_n282_));
OR2X2 OR2X2_32 ( .A(_abc_2284_new_n285_), .B(_abc_2284_new_n286_), .Y(_abc_2284_new_n287_));
OR2X2 OR2X2_33 ( .A(_abc_2284_new_n296_), .B(_abc_2284_new_n290_), .Y(_abc_2284_new_n297_));
OR2X2 OR2X2_34 ( .A(_abc_2284_new_n298_), .B(_abc_2284_new_n294_), .Y(_abc_2284_new_n299_));
OR2X2 OR2X2_35 ( .A(_abc_2284_new_n288_), .B(_abc_2284_new_n299_), .Y(_0tx_data_7_0__0_));
OR2X2 OR2X2_36 ( .A(_abc_2284_new_n301_), .B(_abc_2284_new_n302_), .Y(_abc_2284_new_n303_));
OR2X2 OR2X2_37 ( .A(_abc_2284_new_n306_), .B(_abc_2284_new_n305_), .Y(_abc_2284_new_n307_));
OR2X2 OR2X2_38 ( .A(_abc_2284_new_n304_), .B(_abc_2284_new_n307_), .Y(_0tx_data_7_0__1_));
OR2X2 OR2X2_39 ( .A(_abc_2284_new_n309_), .B(_abc_2284_new_n310_), .Y(_abc_2284_new_n311_));
OR2X2 OR2X2_4 ( .A(_abc_2284_new_n177_), .B(_abc_2284_new_n160_), .Y(_abc_2284_new_n183_));
OR2X2 OR2X2_40 ( .A(_abc_2284_new_n314_), .B(_abc_2284_new_n313_), .Y(_abc_2284_new_n315_));
OR2X2 OR2X2_41 ( .A(_abc_2284_new_n312_), .B(_abc_2284_new_n315_), .Y(_0tx_data_7_0__2_));
OR2X2 OR2X2_42 ( .A(_abc_2284_new_n317_), .B(_abc_2284_new_n318_), .Y(_abc_2284_new_n319_));
OR2X2 OR2X2_43 ( .A(_abc_2284_new_n322_), .B(_abc_2284_new_n321_), .Y(_abc_2284_new_n323_));
OR2X2 OR2X2_44 ( .A(_abc_2284_new_n320_), .B(_abc_2284_new_n323_), .Y(_0tx_data_7_0__3_));
OR2X2 OR2X2_45 ( .A(_abc_2284_new_n325_), .B(_abc_2284_new_n326_), .Y(_abc_2284_new_n327_));
OR2X2 OR2X2_46 ( .A(_abc_2284_new_n330_), .B(_abc_2284_new_n329_), .Y(_abc_2284_new_n331_));
OR2X2 OR2X2_47 ( .A(_abc_2284_new_n328_), .B(_abc_2284_new_n331_), .Y(_0tx_data_7_0__4_));
OR2X2 OR2X2_48 ( .A(_abc_2284_new_n333_), .B(_abc_2284_new_n334_), .Y(_abc_2284_new_n335_));
OR2X2 OR2X2_49 ( .A(_abc_2284_new_n338_), .B(_abc_2284_new_n337_), .Y(_abc_2284_new_n339_));
OR2X2 OR2X2_5 ( .A(_abc_2284_new_n176_), .B(_abc_2284_new_n161_), .Y(_abc_2284_new_n186_));
OR2X2 OR2X2_50 ( .A(_abc_2284_new_n336_), .B(_abc_2284_new_n339_), .Y(_0tx_data_7_0__5_));
OR2X2 OR2X2_51 ( .A(_abc_2284_new_n283_), .B(tx_data_6_), .Y(_abc_2284_new_n341_));
OR2X2 OR2X2_52 ( .A(_abc_2284_new_n343_), .B(_abc_2284_new_n342_), .Y(_abc_2284_new_n344_));
OR2X2 OR2X2_53 ( .A(_abc_2284_new_n347_), .B(_abc_2284_new_n346_), .Y(_abc_2284_new_n348_));
OR2X2 OR2X2_54 ( .A(_abc_2284_new_n345_), .B(_abc_2284_new_n348_), .Y(_0tx_data_7_0__6_));
OR2X2 OR2X2_55 ( .A(_abc_2284_new_n343_), .B(_abc_2284_new_n297_), .Y(_abc_2284_new_n351_));
OR2X2 OR2X2_56 ( .A(_abc_2284_new_n352_), .B(_abc_2284_new_n350_), .Y(_0tx_data_7_0__7_));
OR2X2 OR2X2_57 ( .A(_abc_2284_new_n358_), .B(_abc_2284_new_n356_), .Y(_abc_2284_new_n359_));
OR2X2 OR2X2_58 ( .A(_abc_2284_new_n360_), .B(_abc_2284_new_n361_), .Y(_0tx_bits_remaining_3_0__0_));
OR2X2 OR2X2_59 ( .A(_abc_2284_new_n367_), .B(_abc_2284_new_n365_), .Y(_abc_2284_new_n368_));
OR2X2 OR2X2_6 ( .A(_abc_2284_new_n194_), .B(_abc_2284_new_n173_), .Y(_abc_2284_new_n195_));
OR2X2 OR2X2_60 ( .A(_abc_2284_new_n369_), .B(_abc_2284_new_n370_), .Y(_0tx_bits_remaining_3_0__1_));
OR2X2 OR2X2_61 ( .A(_abc_2284_new_n377_), .B(_abc_2284_new_n297_), .Y(_abc_2284_new_n378_));
OR2X2 OR2X2_62 ( .A(_abc_2284_new_n379_), .B(_abc_2284_new_n375_), .Y(_0tx_bits_remaining_3_0__2_));
OR2X2 OR2X2_63 ( .A(_abc_2284_new_n383_), .B(_abc_2284_new_n293_), .Y(_0tx_bits_remaining_3_0__3_));
OR2X2 OR2X2_64 ( .A(_abc_2284_new_n391_), .B(_abc_2284_new_n293_), .Y(_abc_2284_new_n392_));
OR2X2 OR2X2_65 ( .A(_abc_2284_new_n390_), .B(_abc_2284_new_n392_), .Y(_0tx_countdown_5_0__2_));
OR2X2 OR2X2_66 ( .A(_abc_2284_new_n397_), .B(_abc_2284_new_n394_), .Y(_abc_2284_new_n398_));
OR2X2 OR2X2_67 ( .A(_abc_2284_new_n406_), .B(_abc_2284_new_n293_), .Y(_0tx_state_1_0__0_));
OR2X2 OR2X2_68 ( .A(_abc_2284_new_n396_), .B(_abc_2284_new_n290_), .Y(_abc_2284_new_n408_));
OR2X2 OR2X2_69 ( .A(_abc_2284_new_n279_), .B(tx), .Y(_abc_2284_new_n415_));
OR2X2 OR2X2_7 ( .A(tx_clk_divider_2_), .B(tx_clk_divider_3_), .Y(_abc_2284_new_n197_));
OR2X2 OR2X2_70 ( .A(_abc_2284_new_n417_), .B(_abc_2284_new_n418_), .Y(_0tx_out_0_0_));
OR2X2 OR2X2_71 ( .A(rx_clk_divider_2_), .B(rx_clk_divider_3_), .Y(_abc_2284_new_n421_));
OR2X2 OR2X2_72 ( .A(rx_clk_divider_1_), .B(rx_clk_divider_0_), .Y(_abc_2284_new_n422_));
OR2X2 OR2X2_73 ( .A(_abc_2284_new_n421_), .B(_abc_2284_new_n422_), .Y(_abc_2284_new_n423_));
OR2X2 OR2X2_74 ( .A(_abc_2284_new_n423_), .B(_abc_2284_new_n427_), .Y(_abc_2284_new_n428_));
OR2X2 OR2X2_75 ( .A(rx_clk_divider_6_), .B(rx_clk_divider_7_), .Y(_abc_2284_new_n429_));
OR2X2 OR2X2_76 ( .A(_abc_2284_new_n428_), .B(_abc_2284_new_n429_), .Y(_abc_2284_new_n430_));
OR2X2 OR2X2_77 ( .A(_abc_2284_new_n430_), .B(rx_clk_divider_8_), .Y(_abc_2284_new_n431_));
OR2X2 OR2X2_78 ( .A(_abc_2284_new_n431_), .B(rx_clk_divider_9_), .Y(_abc_2284_new_n432_));
OR2X2 OR2X2_79 ( .A(_abc_2284_new_n438_), .B(_abc_2284_new_n433_), .Y(_abc_2284_new_n439_));
OR2X2 OR2X2_8 ( .A(tx_clk_divider_1_), .B(tx_clk_divider_0_), .Y(_abc_2284_new_n198_));
OR2X2 OR2X2_80 ( .A(_abc_2284_new_n428_), .B(rx_clk_divider_6_), .Y(_abc_2284_new_n441_));
OR2X2 OR2X2_81 ( .A(_abc_2284_new_n446_), .B(_abc_2284_new_n447_), .Y(_abc_2284_new_n448_));
OR2X2 OR2X2_82 ( .A(_abc_2284_new_n463_), .B(_abc_2284_new_n465_), .Y(_abc_2284_new_n466_));
OR2X2 OR2X2_83 ( .A(_abc_2284_new_n474_), .B(_abc_2284_new_n472_), .Y(_abc_2284_new_n475_));
OR2X2 OR2X2_84 ( .A(_abc_2284_new_n475_), .B(_abc_2284_new_n471_), .Y(_abc_2284_new_n476_));
OR2X2 OR2X2_85 ( .A(_abc_2284_new_n469_), .B(_abc_2284_new_n476_), .Y(_abc_2284_new_n477_));
OR2X2 OR2X2_86 ( .A(_abc_2284_new_n482_), .B(_abc_2284_new_n484_), .Y(_abc_2284_new_n485_));
OR2X2 OR2X2_87 ( .A(_abc_2284_new_n489_), .B(_abc_2284_new_n480_), .Y(_0rx_countdown_5_0__1_));
OR2X2 OR2X2_88 ( .A(_abc_2284_new_n494_), .B(_abc_2284_new_n492_), .Y(_abc_2284_new_n495_));
OR2X2 OR2X2_89 ( .A(_abc_2284_new_n437_), .B(_abc_2284_new_n434_), .Y(_abc_2284_new_n496_));
OR2X2 OR2X2_9 ( .A(_abc_2284_new_n197_), .B(_abc_2284_new_n198_), .Y(_abc_2284_new_n199_));
OR2X2 OR2X2_90 ( .A(_abc_2284_new_n435_), .B(_abc_2284_new_n454_), .Y(_abc_2284_new_n500_));
OR2X2 OR2X2_91 ( .A(_abc_2284_new_n446_), .B(_abc_2284_new_n425_), .Y(_abc_2284_new_n503_));
OR2X2 OR2X2_92 ( .A(_abc_2284_new_n509_), .B(rx_countdown_2_), .Y(_abc_2284_new_n510_));
OR2X2 OR2X2_93 ( .A(_abc_2284_new_n512_), .B(_abc_2284_new_n511_), .Y(_abc_2284_new_n513_));
OR2X2 OR2X2_94 ( .A(_abc_2284_new_n508_), .B(_abc_2284_new_n511_), .Y(_abc_2284_new_n517_));
OR2X2 OR2X2_95 ( .A(_abc_2284_new_n461_), .B(_abc_2284_new_n464_), .Y(_abc_2284_new_n519_));
OR2X2 OR2X2_96 ( .A(_abc_2284_new_n512_), .B(rx_countdown_2_), .Y(_abc_2284_new_n526_));
OR2X2 OR2X2_97 ( .A(_abc_2284_new_n526_), .B(rx_countdown_3_), .Y(_abc_2284_new_n527_));
OR2X2 OR2X2_98 ( .A(_abc_2284_new_n530_), .B(_abc_2284_new_n525_), .Y(_abc_2284_new_n531_));
OR2X2 OR2X2_99 ( .A(_abc_2284_new_n529_), .B(rx_countdown_5_), .Y(_abc_2284_new_n532_));


endmodule