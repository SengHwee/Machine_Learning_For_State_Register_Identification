module MEMORY_INTERFACE(clock, resetn, \rs1[0] , \rs1[1] , \rs1[2] , \rs1[3] , \rs1[4] , \rs1[5] , \rs1[6] , \rs1[7] , \rs1[8] , \rs1[9] , \rs1[10] , \rs1[11] , \rs1[12] , \rs1[13] , \rs1[14] , \rs1[15] , \rs1[16] , \rs1[17] , \rs1[18] , \rs1[19] , \rs1[20] , \rs1[21] , \rs1[22] , \rs1[23] , \rs1[24] , \rs1[25] , \rs1[26] , \rs1[27] , \rs1[28] , \rs1[29] , \rs1[30] , \rs1[31] , \rs2[0] , \rs2[1] , \rs2[2] , \rs2[3] , \rs2[4] , \rs2[5] , \rs2[6] , \rs2[7] , \rs2[8] , \rs2[9] , \rs2[10] , \rs2[11] , \rs2[12] , \rs2[13] , \rs2[14] , \rs2[15] , \rs2[16] , \rs2[17] , \rs2[18] , \rs2[19] , \rs2[20] , \rs2[21] , \rs2[22] , \rs2[23] , \rs2[24] , \rs2[25] , \rs2[26] , \rs2[27] , \rs2[28] , \rs2[29] , \rs2[30] , \rs2[31] , \Rdata_mem[0] , \Rdata_mem[1] , \Rdata_mem[2] , \Rdata_mem[3] , \Rdata_mem[4] , \Rdata_mem[5] , \Rdata_mem[6] , \Rdata_mem[7] , \Rdata_mem[8] , \Rdata_mem[9] , \Rdata_mem[10] , \Rdata_mem[11] , \Rdata_mem[12] , \Rdata_mem[13] , \Rdata_mem[14] , \Rdata_mem[15] , \Rdata_mem[16] , \Rdata_mem[17] , \Rdata_mem[18] , \Rdata_mem[19] , \Rdata_mem[20] , \Rdata_mem[21] , \Rdata_mem[22] , \Rdata_mem[23] , \Rdata_mem[24] , \Rdata_mem[25] , \Rdata_mem[26] , \Rdata_mem[27] , \Rdata_mem[28] , \Rdata_mem[29] , \Rdata_mem[30] , \Rdata_mem[31] , ARready, Rvalid, AWready, Wready, Bvalid, \imm[0] , \imm[1] , \imm[2] , \imm[3] , \imm[4] , \imm[5] , \imm[6] , \imm[7] , \imm[8] , \imm[9] , \imm[10] , \imm[11] , \imm[12] , \imm[13] , \imm[14] , \imm[15] , \imm[16] , \imm[17] , \imm[18] , \imm[19] , \imm[20] , \imm[21] , \imm[22] , \imm[23] , \imm[24] , \imm[25] , \imm[26] , \imm[27] , \imm[28] , \imm[29] , \imm[30] , \imm[31] , \W_R[0] , \W_R[1] , \wordsize[0] , \wordsize[1] , enable, \pc[0] , \pc[1] , \pc[2] , \pc[3] , \pc[4] , \pc[5] , \pc[6] , \pc[7] , \pc[8] , \pc[9] , \pc[10] , \pc[11] , \pc[12] , \pc[13] , \pc[14] , \pc[15] , \pc[16] , \pc[17] , \pc[18] , \pc[19] , \pc[20] , \pc[21] , \pc[22] , \pc[23] , \pc[24] , \pc[25] , \pc[26] , \pc[27] , \pc[28] , \pc[29] , \pc[30] , \pc[31] , signo, busy, done, align, \AWdata[0] , \AWdata[1] , \AWdata[2] , \AWdata[3] , \AWdata[4] , \AWdata[5] , \AWdata[6] , \AWdata[7] , \AWdata[8] , \AWdata[9] , \AWdata[10] , \AWdata[11] , \AWdata[12] , \AWdata[13] , \AWdata[14] , \AWdata[15] , \AWdata[16] , \AWdata[17] , \AWdata[18] , \AWdata[19] , \AWdata[20] , \AWdata[21] , \AWdata[22] , \AWdata[23] , \AWdata[24] , \AWdata[25] , \AWdata[26] , \AWdata[27] , \AWdata[28] , \AWdata[29] , \AWdata[30] , \AWdata[31] , \ARdata[0] , \ARdata[1] , \ARdata[2] , \ARdata[3] , \ARdata[4] , \ARdata[5] , \ARdata[6] , \ARdata[7] , \ARdata[8] , \ARdata[9] , \ARdata[10] , \ARdata[11] , \ARdata[12] , \ARdata[13] , \ARdata[14] , \ARdata[15] , \ARdata[16] , \ARdata[17] , \ARdata[18] , \ARdata[19] , \ARdata[20] , \ARdata[21] , \ARdata[22] , \ARdata[23] , \ARdata[24] , \ARdata[25] , \ARdata[26] , \ARdata[27] , \ARdata[28] , \ARdata[29] , \ARdata[30] , \ARdata[31] , \Wdata[0] , \Wdata[1] , \Wdata[2] , \Wdata[3] , \Wdata[4] , \Wdata[5] , \Wdata[6] , \Wdata[7] , \Wdata[8] , \Wdata[9] , \Wdata[10] , \Wdata[11] , \Wdata[12] , \Wdata[13] , \Wdata[14] , \Wdata[15] , \Wdata[16] , \Wdata[17] , \Wdata[18] , \Wdata[19] , \Wdata[20] , \Wdata[21] , \Wdata[22] , \Wdata[23] , \Wdata[24] , \Wdata[25] , \Wdata[26] , \Wdata[27] , \Wdata[28] , \Wdata[29] , \Wdata[30] , \Wdata[31] , \rd[0] , \rd[1] , \rd[2] , \rd[3] , \rd[4] , \rd[5] , \rd[6] , \rd[7] , \rd[8] , \rd[9] , \rd[10] , \rd[11] , \rd[12] , \rd[13] , \rd[14] , \rd[15] , \rd[16] , \rd[17] , \rd[18] , \rd[19] , \rd[20] , \rd[21] , \rd[22] , \rd[23] , \rd[24] , \rd[25] , \rd[26] , \rd[27] , \rd[28] , \rd[29] , \rd[30] , \rd[31] , \inst[0] , \inst[1] , \inst[2] , \inst[3] , \inst[4] , \inst[5] , \inst[6] , \inst[7] , \inst[8] , \inst[9] , \inst[10] , \inst[11] , \inst[12] , \inst[13] , \inst[14] , \inst[15] , \inst[16] , \inst[17] , \inst[18] , \inst[19] , \inst[20] , \inst[21] , \inst[22] , \inst[23] , \inst[24] , \inst[25] , \inst[26] , \inst[27] , \inst[28] , \inst[29] , \inst[30] , \inst[31] , ARvalid, RReady, AWvalid, Wvalid, \arprot[0] , \arprot[1] , \arprot[2] , \awprot[0] , \awprot[1] , \awprot[2] , Bready, \Wstrb[0] , \Wstrb[1] , \Wstrb[2] , \Wstrb[3] , rd_en);
  output \ARdata[0] ;
  output \ARdata[10] ;
  output \ARdata[11] ;
  output \ARdata[12] ;
  output \ARdata[13] ;
  output \ARdata[14] ;
  output \ARdata[15] ;
  output \ARdata[16] ;
  output \ARdata[17] ;
  output \ARdata[18] ;
  output \ARdata[19] ;
  output \ARdata[1] ;
  output \ARdata[20] ;
  output \ARdata[21] ;
  output \ARdata[22] ;
  output \ARdata[23] ;
  output \ARdata[24] ;
  output \ARdata[25] ;
  output \ARdata[26] ;
  output \ARdata[27] ;
  output \ARdata[28] ;
  output \ARdata[29] ;
  output \ARdata[2] ;
  output \ARdata[30] ;
  output \ARdata[31] ;
  output \ARdata[3] ;
  output \ARdata[4] ;
  output \ARdata[5] ;
  output \ARdata[6] ;
  output \ARdata[7] ;
  output \ARdata[8] ;
  output \ARdata[9] ;
  input ARready;
  output ARvalid;
  output \AWdata[0] ;
  output \AWdata[10] ;
  output \AWdata[11] ;
  output \AWdata[12] ;
  output \AWdata[13] ;
  output \AWdata[14] ;
  output \AWdata[15] ;
  output \AWdata[16] ;
  output \AWdata[17] ;
  output \AWdata[18] ;
  output \AWdata[19] ;
  output \AWdata[1] ;
  output \AWdata[20] ;
  output \AWdata[21] ;
  output \AWdata[22] ;
  output \AWdata[23] ;
  output \AWdata[24] ;
  output \AWdata[25] ;
  output \AWdata[26] ;
  output \AWdata[27] ;
  output \AWdata[28] ;
  output \AWdata[29] ;
  output \AWdata[2] ;
  output \AWdata[30] ;
  output \AWdata[31] ;
  output \AWdata[3] ;
  output \AWdata[4] ;
  output \AWdata[5] ;
  output \AWdata[6] ;
  output \AWdata[7] ;
  output \AWdata[8] ;
  output \AWdata[9] ;
  input AWready;
  output AWvalid;
  output Bready;
  input Bvalid;
  output RReady;
  input \Rdata_mem[0] ;
  input \Rdata_mem[10] ;
  input \Rdata_mem[11] ;
  input \Rdata_mem[12] ;
  input \Rdata_mem[13] ;
  input \Rdata_mem[14] ;
  input \Rdata_mem[15] ;
  input \Rdata_mem[16] ;
  input \Rdata_mem[17] ;
  input \Rdata_mem[18] ;
  input \Rdata_mem[19] ;
  input \Rdata_mem[1] ;
  input \Rdata_mem[20] ;
  input \Rdata_mem[21] ;
  input \Rdata_mem[22] ;
  input \Rdata_mem[23] ;
  input \Rdata_mem[24] ;
  input \Rdata_mem[25] ;
  input \Rdata_mem[26] ;
  input \Rdata_mem[27] ;
  input \Rdata_mem[28] ;
  input \Rdata_mem[29] ;
  input \Rdata_mem[2] ;
  input \Rdata_mem[30] ;
  input \Rdata_mem[31] ;
  input \Rdata_mem[3] ;
  input \Rdata_mem[4] ;
  input \Rdata_mem[5] ;
  input \Rdata_mem[6] ;
  input \Rdata_mem[7] ;
  input \Rdata_mem[8] ;
  input \Rdata_mem[9] ;
  input Rvalid;
  input \W_R[0] ;
  input \W_R[1] ;
  wire W_R_1_bF_buf0;
  wire W_R_1_bF_buf1;
  wire W_R_1_bF_buf2;
  wire W_R_1_bF_buf3;
  wire W_R_1_bF_buf4;
  wire W_R_1_bF_buf5;
  output \Wdata[0] ;
  output \Wdata[10] ;
  output \Wdata[11] ;
  output \Wdata[12] ;
  output \Wdata[13] ;
  output \Wdata[14] ;
  output \Wdata[15] ;
  output \Wdata[16] ;
  output \Wdata[17] ;
  output \Wdata[18] ;
  output \Wdata[19] ;
  output \Wdata[1] ;
  output \Wdata[20] ;
  output \Wdata[21] ;
  output \Wdata[22] ;
  output \Wdata[23] ;
  output \Wdata[24] ;
  output \Wdata[25] ;
  output \Wdata[26] ;
  output \Wdata[27] ;
  output \Wdata[28] ;
  output \Wdata[29] ;
  output \Wdata[2] ;
  output \Wdata[30] ;
  output \Wdata[31] ;
  output \Wdata[3] ;
  output \Wdata[4] ;
  output \Wdata[5] ;
  output \Wdata[6] ;
  output \Wdata[7] ;
  output \Wdata[8] ;
  output \Wdata[9] ;
  wire Wdata_0__FF_INPUT;
  wire Wdata_10__FF_INPUT;
  wire Wdata_11__FF_INPUT;
  wire Wdata_12__FF_INPUT;
  wire Wdata_13__FF_INPUT;
  wire Wdata_14__FF_INPUT;
  wire Wdata_15__FF_INPUT;
  wire Wdata_16__FF_INPUT;
  wire Wdata_17__FF_INPUT;
  wire Wdata_18__FF_INPUT;
  wire Wdata_19__FF_INPUT;
  wire Wdata_1__FF_INPUT;
  wire Wdata_20__FF_INPUT;
  wire Wdata_21__FF_INPUT;
  wire Wdata_22__FF_INPUT;
  wire Wdata_23__FF_INPUT;
  wire Wdata_24__FF_INPUT;
  wire Wdata_25__FF_INPUT;
  wire Wdata_26__FF_INPUT;
  wire Wdata_27__FF_INPUT;
  wire Wdata_28__FF_INPUT;
  wire Wdata_29__FF_INPUT;
  wire Wdata_2__FF_INPUT;
  wire Wdata_30__FF_INPUT;
  wire Wdata_31__FF_INPUT;
  wire Wdata_3__FF_INPUT;
  wire Wdata_4__FF_INPUT;
  wire Wdata_5__FF_INPUT;
  wire Wdata_6__FF_INPUT;
  wire Wdata_7__FF_INPUT;
  wire Wdata_8__FF_INPUT;
  wire Wdata_9__FF_INPUT;
  input Wready;
  output \Wstrb[0] ;
  output \Wstrb[1] ;
  output \Wstrb[2] ;
  output \Wstrb[3] ;
  wire Wstrb_0__FF_INPUT;
  wire Wstrb_1__FF_INPUT;
  wire Wstrb_2__FF_INPUT;
  wire Wstrb_3__FF_INPUT;
  output Wvalid;
  wire _abc_3815_n122;
  wire _abc_3815_n132;
  wire _abc_3815_n14;
  wire _abc_3815_n152;
  wire _abc_3815_n23;
  wire _abc_3815_n52;
  wire _abc_3815_n99;
  wire _abc_4513_n1000;
  wire _abc_4513_n1001;
  wire _abc_4513_n1002;
  wire _abc_4513_n1003;
  wire _abc_4513_n1004;
  wire _abc_4513_n1005;
  wire _abc_4513_n1006;
  wire _abc_4513_n1007;
  wire _abc_4513_n1008;
  wire _abc_4513_n1009;
  wire _abc_4513_n1010;
  wire _abc_4513_n1011;
  wire _abc_4513_n1012;
  wire _abc_4513_n1013;
  wire _abc_4513_n1014;
  wire _abc_4513_n1016;
  wire _abc_4513_n1017;
  wire _abc_4513_n1018;
  wire _abc_4513_n1019;
  wire _abc_4513_n1020;
  wire _abc_4513_n1021;
  wire _abc_4513_n1022;
  wire _abc_4513_n1023;
  wire _abc_4513_n1024;
  wire _abc_4513_n1025;
  wire _abc_4513_n1026;
  wire _abc_4513_n1027;
  wire _abc_4513_n1029;
  wire _abc_4513_n1030;
  wire _abc_4513_n1031;
  wire _abc_4513_n1032;
  wire _abc_4513_n1033;
  wire _abc_4513_n1034;
  wire _abc_4513_n1035;
  wire _abc_4513_n1036;
  wire _abc_4513_n1037;
  wire _abc_4513_n1038;
  wire _abc_4513_n1039;
  wire _abc_4513_n1040;
  wire _abc_4513_n1041;
  wire _abc_4513_n1042;
  wire _abc_4513_n1043;
  wire _abc_4513_n1044;
  wire _abc_4513_n1045;
  wire _abc_4513_n1046;
  wire _abc_4513_n1048;
  wire _abc_4513_n1049;
  wire _abc_4513_n1050;
  wire _abc_4513_n1051;
  wire _abc_4513_n1052;
  wire _abc_4513_n1053;
  wire _abc_4513_n1054;
  wire _abc_4513_n1055;
  wire _abc_4513_n1056;
  wire _abc_4513_n1057;
  wire _abc_4513_n1058;
  wire _abc_4513_n1059;
  wire _abc_4513_n1061;
  wire _abc_4513_n1062;
  wire _abc_4513_n1063;
  wire _abc_4513_n1064;
  wire _abc_4513_n1065;
  wire _abc_4513_n1066;
  wire _abc_4513_n1067;
  wire _abc_4513_n1068;
  wire _abc_4513_n1069;
  wire _abc_4513_n1070;
  wire _abc_4513_n1071;
  wire _abc_4513_n1072;
  wire _abc_4513_n1073;
  wire _abc_4513_n1074;
  wire _abc_4513_n1075;
  wire _abc_4513_n1077;
  wire _abc_4513_n1078;
  wire _abc_4513_n1079;
  wire _abc_4513_n1080;
  wire _abc_4513_n1081;
  wire _abc_4513_n1082;
  wire _abc_4513_n1083;
  wire _abc_4513_n1084;
  wire _abc_4513_n1085;
  wire _abc_4513_n1086;
  wire _abc_4513_n1087;
  wire _abc_4513_n1088;
  wire _abc_4513_n1090;
  wire _abc_4513_n1091;
  wire _abc_4513_n1092;
  wire _abc_4513_n1093;
  wire _abc_4513_n1094;
  wire _abc_4513_n1095;
  wire _abc_4513_n1096;
  wire _abc_4513_n1097;
  wire _abc_4513_n1098;
  wire _abc_4513_n1099;
  wire _abc_4513_n1100;
  wire _abc_4513_n1101;
  wire _abc_4513_n1102;
  wire _abc_4513_n1103;
  wire _abc_4513_n1104;
  wire _abc_4513_n1105;
  wire _abc_4513_n1106;
  wire _abc_4513_n1107;
  wire _abc_4513_n1109;
  wire _abc_4513_n1110;
  wire _abc_4513_n1111;
  wire _abc_4513_n1112;
  wire _abc_4513_n1113;
  wire _abc_4513_n1114;
  wire _abc_4513_n1115;
  wire _abc_4513_n1116;
  wire _abc_4513_n1117;
  wire _abc_4513_n1118;
  wire _abc_4513_n1119;
  wire _abc_4513_n1120;
  wire _abc_4513_n1122;
  wire _abc_4513_n1123;
  wire _abc_4513_n1124;
  wire _abc_4513_n1125;
  wire _abc_4513_n1126;
  wire _abc_4513_n1127;
  wire _abc_4513_n1128;
  wire _abc_4513_n1129;
  wire _abc_4513_n1130;
  wire _abc_4513_n1131;
  wire _abc_4513_n1132;
  wire _abc_4513_n1133;
  wire _abc_4513_n1134;
  wire _abc_4513_n1135;
  wire _abc_4513_n1136;
  wire _abc_4513_n1137;
  wire _abc_4513_n1139;
  wire _abc_4513_n1140;
  wire _abc_4513_n1141;
  wire _abc_4513_n1142;
  wire _abc_4513_n1143;
  wire _abc_4513_n1144;
  wire _abc_4513_n1145;
  wire _abc_4513_n1146;
  wire _abc_4513_n1147;
  wire _abc_4513_n1148;
  wire _abc_4513_n1149;
  wire _abc_4513_n1150;
  wire _abc_4513_n1152;
  wire _abc_4513_n1153;
  wire _abc_4513_n1154;
  wire _abc_4513_n1155;
  wire _abc_4513_n1156;
  wire _abc_4513_n1157;
  wire _abc_4513_n1158;
  wire _abc_4513_n1159;
  wire _abc_4513_n1160;
  wire _abc_4513_n1161;
  wire _abc_4513_n1162;
  wire _abc_4513_n1163;
  wire _abc_4513_n1164;
  wire _abc_4513_n1165;
  wire _abc_4513_n1166;
  wire _abc_4513_n1167;
  wire _abc_4513_n1168;
  wire _abc_4513_n1169;
  wire _abc_4513_n1170;
  wire _abc_4513_n1171;
  wire _abc_4513_n1172;
  wire _abc_4513_n1174;
  wire _abc_4513_n1175;
  wire _abc_4513_n1176;
  wire _abc_4513_n1177;
  wire _abc_4513_n1178;
  wire _abc_4513_n1179;
  wire _abc_4513_n1180;
  wire _abc_4513_n1181;
  wire _abc_4513_n1182;
  wire _abc_4513_n1183;
  wire _abc_4513_n1184;
  wire _abc_4513_n1185;
  wire _abc_4513_n1187;
  wire _abc_4513_n1188;
  wire _abc_4513_n1189;
  wire _abc_4513_n1190;
  wire _abc_4513_n1191;
  wire _abc_4513_n1192;
  wire _abc_4513_n1193;
  wire _abc_4513_n1194;
  wire _abc_4513_n1195;
  wire _abc_4513_n1196;
  wire _abc_4513_n1197;
  wire _abc_4513_n1198;
  wire _abc_4513_n1199;
  wire _abc_4513_n1200;
  wire _abc_4513_n1201;
  wire _abc_4513_n1202;
  wire _abc_4513_n1204;
  wire _abc_4513_n1205;
  wire _abc_4513_n1206;
  wire _abc_4513_n1207;
  wire _abc_4513_n1208;
  wire _abc_4513_n1209;
  wire _abc_4513_n1210;
  wire _abc_4513_n1211;
  wire _abc_4513_n1212;
  wire _abc_4513_n1213;
  wire _abc_4513_n1214;
  wire _abc_4513_n1215;
  wire _abc_4513_n1217;
  wire _abc_4513_n1218;
  wire _abc_4513_n1219;
  wire _abc_4513_n1220;
  wire _abc_4513_n1221;
  wire _abc_4513_n1222;
  wire _abc_4513_n1223;
  wire _abc_4513_n1224;
  wire _abc_4513_n1225;
  wire _abc_4513_n1226;
  wire _abc_4513_n1227;
  wire _abc_4513_n1228;
  wire _abc_4513_n1229;
  wire _abc_4513_n1230;
  wire _abc_4513_n1231;
  wire _abc_4513_n1232;
  wire _abc_4513_n1233;
  wire _abc_4513_n1234;
  wire _abc_4513_n1235;
  wire _abc_4513_n1237;
  wire _abc_4513_n1238;
  wire _abc_4513_n1239;
  wire _abc_4513_n1240;
  wire _abc_4513_n1241;
  wire _abc_4513_n1242;
  wire _abc_4513_n1243;
  wire _abc_4513_n1244;
  wire _abc_4513_n1245;
  wire _abc_4513_n1246;
  wire _abc_4513_n1247;
  wire _abc_4513_n1248;
  wire _abc_4513_n1250;
  wire _abc_4513_n1251;
  wire _abc_4513_n1252;
  wire _abc_4513_n1253;
  wire _abc_4513_n1254;
  wire _abc_4513_n1255;
  wire _abc_4513_n1256;
  wire _abc_4513_n1257;
  wire _abc_4513_n1258;
  wire _abc_4513_n1259;
  wire _abc_4513_n1260;
  wire _abc_4513_n1261;
  wire _abc_4513_n1262;
  wire _abc_4513_n1263;
  wire _abc_4513_n1264;
  wire _abc_4513_n1265;
  wire _abc_4513_n1267;
  wire _abc_4513_n1268;
  wire _abc_4513_n1269;
  wire _abc_4513_n1270;
  wire _abc_4513_n1271;
  wire _abc_4513_n1272;
  wire _abc_4513_n1273;
  wire _abc_4513_n1274;
  wire _abc_4513_n1275;
  wire _abc_4513_n1276;
  wire _abc_4513_n1277;
  wire _abc_4513_n1278;
  wire _abc_4513_n1280;
  wire _abc_4513_n1281;
  wire _abc_4513_n1282;
  wire _abc_4513_n1283;
  wire _abc_4513_n1284;
  wire _abc_4513_n1285;
  wire _abc_4513_n1286;
  wire _abc_4513_n1287;
  wire _abc_4513_n1288;
  wire _abc_4513_n1289;
  wire _abc_4513_n1290;
  wire _abc_4513_n1291;
  wire _abc_4513_n1292;
  wire _abc_4513_n1293;
  wire _abc_4513_n1294;
  wire _abc_4513_n1295;
  wire _abc_4513_n1296;
  wire _abc_4513_n1297;
  wire _abc_4513_n1298;
  wire _abc_4513_n1299;
  wire _abc_4513_n1300;
  wire _abc_4513_n1302;
  wire _abc_4513_n1303;
  wire _abc_4513_n1304;
  wire _abc_4513_n1305;
  wire _abc_4513_n1306;
  wire _abc_4513_n1307;
  wire _abc_4513_n1308;
  wire _abc_4513_n1309;
  wire _abc_4513_n1310;
  wire _abc_4513_n1311;
  wire _abc_4513_n1312;
  wire _abc_4513_n1313;
  wire _abc_4513_n1315;
  wire _abc_4513_n1316;
  wire _abc_4513_n1317;
  wire _abc_4513_n1318;
  wire _abc_4513_n1319;
  wire _abc_4513_n1320;
  wire _abc_4513_n1321;
  wire _abc_4513_n1322;
  wire _abc_4513_n1323;
  wire _abc_4513_n1324;
  wire _abc_4513_n1325;
  wire _abc_4513_n1326;
  wire _abc_4513_n1327;
  wire _abc_4513_n1328;
  wire _abc_4513_n1329;
  wire _abc_4513_n1330;
  wire _abc_4513_n1332;
  wire _abc_4513_n1333;
  wire _abc_4513_n1334;
  wire _abc_4513_n1335;
  wire _abc_4513_n1336;
  wire _abc_4513_n1337;
  wire _abc_4513_n1338;
  wire _abc_4513_n1339;
  wire _abc_4513_n1340;
  wire _abc_4513_n1341;
  wire _abc_4513_n1342;
  wire _abc_4513_n1343;
  wire _abc_4513_n1345;
  wire _abc_4513_n1346;
  wire _abc_4513_n1347;
  wire _abc_4513_n1348;
  wire _abc_4513_n1349;
  wire _abc_4513_n1350;
  wire _abc_4513_n1351;
  wire _abc_4513_n1352;
  wire _abc_4513_n1353;
  wire _abc_4513_n1354;
  wire _abc_4513_n1355;
  wire _abc_4513_n1356;
  wire _abc_4513_n1357;
  wire _abc_4513_n1358;
  wire _abc_4513_n1359;
  wire _abc_4513_n1360;
  wire _abc_4513_n1361;
  wire _abc_4513_n1362;
  wire _abc_4513_n1364;
  wire _abc_4513_n1365;
  wire _abc_4513_n1366;
  wire _abc_4513_n1367;
  wire _abc_4513_n1368;
  wire _abc_4513_n1369;
  wire _abc_4513_n1370;
  wire _abc_4513_n1371;
  wire _abc_4513_n1372;
  wire _abc_4513_n1373;
  wire _abc_4513_n1374;
  wire _abc_4513_n1375;
  wire _abc_4513_n1377;
  wire _abc_4513_n1378;
  wire _abc_4513_n1379;
  wire _abc_4513_n1380;
  wire _abc_4513_n1381;
  wire _abc_4513_n1382;
  wire _abc_4513_n1383;
  wire _abc_4513_n1384;
  wire _abc_4513_n1385;
  wire _abc_4513_n1386;
  wire _abc_4513_n1387;
  wire _abc_4513_n1388;
  wire _abc_4513_n1389;
  wire _abc_4513_n1390;
  wire _abc_4513_n1391;
  wire _abc_4513_n1392;
  wire _abc_4513_n1393;
  wire _abc_4513_n1394;
  wire _abc_4513_n1395;
  wire _abc_4513_n1396;
  wire _abc_4513_n1397;
  wire _abc_4513_n1398;
  wire _abc_4513_n1399;
  wire _abc_4513_n1400;
  wire _abc_4513_n1401;
  wire _abc_4513_n1402;
  wire _abc_4513_n1403;
  wire _abc_4513_n1404;
  wire _abc_4513_n1405;
  wire _abc_4513_n1406;
  wire _abc_4513_n1407;
  wire _abc_4513_n1408;
  wire _abc_4513_n1409;
  wire _abc_4513_n1410;
  wire _abc_4513_n1411;
  wire _abc_4513_n1412;
  wire _abc_4513_n1413;
  wire _abc_4513_n1414;
  wire _abc_4513_n1415;
  wire _abc_4513_n1416;
  wire _abc_4513_n1417;
  wire _abc_4513_n1419;
  wire _abc_4513_n1420;
  wire _abc_4513_n1421;
  wire _abc_4513_n1422;
  wire _abc_4513_n1423;
  wire _abc_4513_n1424;
  wire _abc_4513_n1425;
  wire _abc_4513_n1426;
  wire _abc_4513_n1427;
  wire _abc_4513_n1428;
  wire _abc_4513_n1429;
  wire _abc_4513_n1430;
  wire _abc_4513_n1431;
  wire _abc_4513_n1432;
  wire _abc_4513_n1435;
  wire _abc_4513_n1437;
  wire _abc_4513_n1439;
  wire _abc_4513_n1441;
  wire _abc_4513_n361;
  wire _abc_4513_n362_1;
  wire _abc_4513_n363_1;
  wire _abc_4513_n364;
  wire _abc_4513_n365;
  wire _abc_4513_n368;
  wire _abc_4513_n369;
  wire _abc_4513_n370_1;
  wire _abc_4513_n371_1;
  wire _abc_4513_n372;
  wire _abc_4513_n373;
  wire _abc_4513_n374_1;
  wire _abc_4513_n375_1;
  wire _abc_4513_n376;
  wire _abc_4513_n377_1;
  wire _abc_4513_n378_1;
  wire _abc_4513_n379;
  wire _abc_4513_n380_1;
  wire _abc_4513_n381_1;
  wire _abc_4513_n382;
  wire _abc_4513_n383_1;
  wire _abc_4513_n384_1;
  wire _abc_4513_n385;
  wire _abc_4513_n387_1;
  wire _abc_4513_n388;
  wire _abc_4513_n389_1;
  wire _abc_4513_n390_1;
  wire _abc_4513_n391;
  wire _abc_4513_n393_1;
  wire _abc_4513_n394;
  wire _abc_4513_n395_1;
  wire _abc_4513_n396_1;
  wire _abc_4513_n397;
  wire _abc_4513_n398_1;
  wire _abc_4513_n399_1;
  wire _abc_4513_n400;
  wire _abc_4513_n401_1;
  wire _abc_4513_n402_1;
  wire _abc_4513_n403;
  wire _abc_4513_n404_1;
  wire _abc_4513_n405_1;
  wire _abc_4513_n406;
  wire _abc_4513_n407_1;
  wire _abc_4513_n408_1;
  wire _abc_4513_n409;
  wire _abc_4513_n410_1;
  wire _abc_4513_n411_1;
  wire _abc_4513_n412;
  wire _abc_4513_n413_1;
  wire _abc_4513_n414_1;
  wire _abc_4513_n415;
  wire _abc_4513_n416_1;
  wire _abc_4513_n417_1;
  wire _abc_4513_n418;
  wire _abc_4513_n419_1;
  wire _abc_4513_n420_1;
  wire _abc_4513_n421;
  wire _abc_4513_n422_1;
  wire _abc_4513_n423;
  wire _abc_4513_n424;
  wire _abc_4513_n426;
  wire _abc_4513_n427_1;
  wire _abc_4513_n428;
  wire _abc_4513_n429;
  wire _abc_4513_n430;
  wire _abc_4513_n431;
  wire _abc_4513_n432;
  wire _abc_4513_n433;
  wire _abc_4513_n434;
  wire _abc_4513_n436;
  wire _abc_4513_n437;
  wire _abc_4513_n438_1;
  wire _abc_4513_n439;
  wire _abc_4513_n440;
  wire _abc_4513_n442;
  wire _abc_4513_n443;
  wire _abc_4513_n444;
  wire _abc_4513_n446_1;
  wire _abc_4513_n447;
  wire _abc_4513_n448;
  wire _abc_4513_n449;
  wire _abc_4513_n450;
  wire _abc_4513_n451;
  wire _abc_4513_n452;
  wire _abc_4513_n453;
  wire _abc_4513_n454_1;
  wire _abc_4513_n455;
  wire _abc_4513_n456;
  wire _abc_4513_n457;
  wire _abc_4513_n458;
  wire _abc_4513_n459;
  wire _abc_4513_n460;
  wire _abc_4513_n461;
  wire _abc_4513_n462_1;
  wire _abc_4513_n463;
  wire _abc_4513_n464;
  wire _abc_4513_n465;
  wire _abc_4513_n466;
  wire _abc_4513_n467;
  wire _abc_4513_n470_1;
  wire _abc_4513_n471;
  wire _abc_4513_n472;
  wire _abc_4513_n473;
  wire _abc_4513_n473_bF_buf0;
  wire _abc_4513_n473_bF_buf1;
  wire _abc_4513_n473_bF_buf2;
  wire _abc_4513_n473_bF_buf3;
  wire _abc_4513_n473_bF_buf4;
  wire _abc_4513_n473_bF_buf5;
  wire _abc_4513_n474;
  wire _abc_4513_n475;
  wire _abc_4513_n476;
  wire _abc_4513_n477;
  wire _abc_4513_n478_1;
  wire _abc_4513_n479;
  wire _abc_4513_n480;
  wire _abc_4513_n481;
  wire _abc_4513_n482;
  wire _abc_4513_n483;
  wire _abc_4513_n484;
  wire _abc_4513_n485;
  wire _abc_4513_n486_1;
  wire _abc_4513_n487;
  wire _abc_4513_n488;
  wire _abc_4513_n489;
  wire _abc_4513_n490;
  wire _abc_4513_n491;
  wire _abc_4513_n492;
  wire _abc_4513_n493;
  wire _abc_4513_n494_1;
  wire _abc_4513_n495_1;
  wire _abc_4513_n495_1_bF_buf0;
  wire _abc_4513_n495_1_bF_buf1;
  wire _abc_4513_n495_1_bF_buf2;
  wire _abc_4513_n495_1_bF_buf3;
  wire _abc_4513_n495_1_bF_buf4;
  wire _abc_4513_n495_1_bF_buf5;
  wire _abc_4513_n496;
  wire _abc_4513_n497;
  wire _abc_4513_n498;
  wire _abc_4513_n499;
  wire _abc_4513_n501;
  wire _abc_4513_n502;
  wire _abc_4513_n503;
  wire _abc_4513_n505;
  wire _abc_4513_n506;
  wire _abc_4513_n507_1;
  wire _abc_4513_n508;
  wire _abc_4513_n509;
  wire _abc_4513_n510_1;
  wire _abc_4513_n512;
  wire _abc_4513_n513_1;
  wire _abc_4513_n514;
  wire _abc_4513_n516_1;
  wire _abc_4513_n517;
  wire _abc_4513_n518;
  wire _abc_4513_n519_1;
  wire _abc_4513_n519_1_bF_buf0;
  wire _abc_4513_n519_1_bF_buf1;
  wire _abc_4513_n519_1_bF_buf2;
  wire _abc_4513_n519_1_bF_buf3;
  wire _abc_4513_n519_1_bF_buf4;
  wire _abc_4513_n520;
  wire _abc_4513_n521;
  wire _abc_4513_n521_bF_buf0;
  wire _abc_4513_n521_bF_buf1;
  wire _abc_4513_n521_bF_buf2;
  wire _abc_4513_n521_bF_buf3;
  wire _abc_4513_n521_bF_buf4;
  wire _abc_4513_n522_1;
  wire _abc_4513_n523;
  wire _abc_4513_n525_1;
  wire _abc_4513_n526;
  wire _abc_4513_n527;
  wire _abc_4513_n529;
  wire _abc_4513_n530;
  wire _abc_4513_n531;
  wire _abc_4513_n533_1;
  wire _abc_4513_n534;
  wire _abc_4513_n535_1;
  wire _abc_4513_n537_1;
  wire _abc_4513_n538;
  wire _abc_4513_n539_1;
  wire _abc_4513_n541_1;
  wire _abc_4513_n542;
  wire _abc_4513_n543_1;
  wire _abc_4513_n545_1;
  wire _abc_4513_n546;
  wire _abc_4513_n547_1;
  wire _abc_4513_n549_1;
  wire _abc_4513_n550;
  wire _abc_4513_n551_1;
  wire _abc_4513_n553_1;
  wire _abc_4513_n554;
  wire _abc_4513_n555_1;
  wire _abc_4513_n557_1;
  wire _abc_4513_n558;
  wire _abc_4513_n559_1;
  wire _abc_4513_n561_1;
  wire _abc_4513_n562;
  wire _abc_4513_n563_1;
  wire _abc_4513_n565_1;
  wire _abc_4513_n566_1;
  wire _abc_4513_n567_1;
  wire _abc_4513_n569_1;
  wire _abc_4513_n570;
  wire _abc_4513_n571;
  wire _abc_4513_n573;
  wire _abc_4513_n574_1;
  wire _abc_4513_n575_1;
  wire _abc_4513_n577_1;
  wire _abc_4513_n578;
  wire _abc_4513_n579;
  wire _abc_4513_n581;
  wire _abc_4513_n582;
  wire _abc_4513_n583_1;
  wire _abc_4513_n585_1;
  wire _abc_4513_n586_1;
  wire _abc_4513_n587;
  wire _abc_4513_n589;
  wire _abc_4513_n590;
  wire _abc_4513_n591;
  wire _abc_4513_n593;
  wire _abc_4513_n594_1;
  wire _abc_4513_n595_1;
  wire _abc_4513_n597_1;
  wire _abc_4513_n598;
  wire _abc_4513_n599;
  wire _abc_4513_n601;
  wire _abc_4513_n602_1;
  wire _abc_4513_n603_1;
  wire _abc_4513_n605_1;
  wire _abc_4513_n606;
  wire _abc_4513_n607;
  wire _abc_4513_n609;
  wire _abc_4513_n610;
  wire _abc_4513_n611;
  wire _abc_4513_n613_1;
  wire _abc_4513_n614_1;
  wire _abc_4513_n615_1;
  wire _abc_4513_n617;
  wire _abc_4513_n618;
  wire _abc_4513_n619;
  wire _abc_4513_n621;
  wire _abc_4513_n622_1;
  wire _abc_4513_n623_1;
  wire _abc_4513_n625_1;
  wire _abc_4513_n626;
  wire _abc_4513_n627;
  wire _abc_4513_n629;
  wire _abc_4513_n630;
  wire _abc_4513_n631;
  wire _abc_4513_n633;
  wire _abc_4513_n634;
  wire _abc_4513_n635;
  wire _abc_4513_n637_1;
  wire _abc_4513_n638_1;
  wire _abc_4513_n639_1;
  wire _abc_4513_n641;
  wire _abc_4513_n642;
  wire _abc_4513_n643;
  wire _abc_4513_n645_1;
  wire _abc_4513_n646_1;
  wire _abc_4513_n647_1;
  wire _abc_4513_n657_1;
  wire _abc_4513_n658_1;
  wire _abc_4513_n659_1;
  wire _abc_4513_n660_1;
  wire _abc_4513_n662;
  wire _abc_4513_n663;
  wire _abc_4513_n664;
  wire _abc_4513_n666_1;
  wire _abc_4513_n667_1;
  wire _abc_4513_n668_1;
  wire _abc_4513_n670;
  wire _abc_4513_n671;
  wire _abc_4513_n672;
  wire _abc_4513_n674;
  wire _abc_4513_n675;
  wire _abc_4513_n676;
  wire _abc_4513_n678;
  wire _abc_4513_n679;
  wire _abc_4513_n680_1;
  wire _abc_4513_n682_1;
  wire _abc_4513_n683_1;
  wire _abc_4513_n684;
  wire _abc_4513_n686;
  wire _abc_4513_n687;
  wire _abc_4513_n688_1;
  wire _abc_4513_n690_1;
  wire _abc_4513_n691_1;
  wire _abc_4513_n692;
  wire _abc_4513_n694;
  wire _abc_4513_n695;
  wire _abc_4513_n696;
  wire _abc_4513_n698;
  wire _abc_4513_n699_1;
  wire _abc_4513_n700_1;
  wire _abc_4513_n702_1;
  wire _abc_4513_n703;
  wire _abc_4513_n704;
  wire _abc_4513_n706;
  wire _abc_4513_n707;
  wire _abc_4513_n708_1;
  wire _abc_4513_n710_1;
  wire _abc_4513_n711_1;
  wire _abc_4513_n712;
  wire _abc_4513_n714;
  wire _abc_4513_n715;
  wire _abc_4513_n716;
  wire _abc_4513_n718;
  wire _abc_4513_n719;
  wire _abc_4513_n720;
  wire _abc_4513_n722;
  wire _abc_4513_n723;
  wire _abc_4513_n724;
  wire _abc_4513_n725;
  wire _abc_4513_n727_1;
  wire _abc_4513_n728_1;
  wire _abc_4513_n729_1;
  wire _abc_4513_n730;
  wire _abc_4513_n732;
  wire _abc_4513_n733;
  wire _abc_4513_n734;
  wire _abc_4513_n735_1;
  wire _abc_4513_n737_1;
  wire _abc_4513_n738_1;
  wire _abc_4513_n739;
  wire _abc_4513_n740;
  wire _abc_4513_n742;
  wire _abc_4513_n743;
  wire _abc_4513_n744;
  wire _abc_4513_n745_1;
  wire _abc_4513_n747_1;
  wire _abc_4513_n748_1;
  wire _abc_4513_n749;
  wire _abc_4513_n750;
  wire _abc_4513_n752;
  wire _abc_4513_n753_1;
  wire _abc_4513_n754_1;
  wire _abc_4513_n755_1;
  wire _abc_4513_n757;
  wire _abc_4513_n758;
  wire _abc_4513_n759;
  wire _abc_4513_n760;
  wire _abc_4513_n762;
  wire _abc_4513_n763;
  wire _abc_4513_n764;
  wire _abc_4513_n765;
  wire _abc_4513_n766_1;
  wire _abc_4513_n767_1;
  wire _abc_4513_n769_1;
  wire _abc_4513_n769_1_bF_buf0;
  wire _abc_4513_n769_1_bF_buf1;
  wire _abc_4513_n769_1_bF_buf2;
  wire _abc_4513_n769_1_bF_buf3;
  wire _abc_4513_n769_1_bF_buf4;
  wire _abc_4513_n770;
  wire _abc_4513_n771;
  wire _abc_4513_n771_bF_buf0;
  wire _abc_4513_n771_bF_buf1;
  wire _abc_4513_n771_bF_buf2;
  wire _abc_4513_n771_bF_buf3;
  wire _abc_4513_n771_bF_buf4;
  wire _abc_4513_n772;
  wire _abc_4513_n773;
  wire _abc_4513_n774_1;
  wire _abc_4513_n775_1;
  wire _abc_4513_n776_1;
  wire _abc_4513_n777_1;
  wire _abc_4513_n778;
  wire _abc_4513_n779;
  wire _abc_4513_n781;
  wire _abc_4513_n782;
  wire _abc_4513_n783;
  wire _abc_4513_n784;
  wire _abc_4513_n785;
  wire _abc_4513_n786_1;
  wire _abc_4513_n787_1;
  wire _abc_4513_n789_1;
  wire _abc_4513_n790;
  wire _abc_4513_n791;
  wire _abc_4513_n792;
  wire _abc_4513_n793;
  wire _abc_4513_n794_1;
  wire _abc_4513_n795_1;
  wire _abc_4513_n797_1;
  wire _abc_4513_n798;
  wire _abc_4513_n799;
  wire _abc_4513_n800;
  wire _abc_4513_n801;
  wire _abc_4513_n802;
  wire _abc_4513_n803;
  wire _abc_4513_n805;
  wire _abc_4513_n806;
  wire _abc_4513_n807;
  wire _abc_4513_n808;
  wire _abc_4513_n809;
  wire _abc_4513_n810;
  wire _abc_4513_n811_1;
  wire _abc_4513_n813_1;
  wire _abc_4513_n814_1;
  wire _abc_4513_n815;
  wire _abc_4513_n816;
  wire _abc_4513_n817;
  wire _abc_4513_n818;
  wire _abc_4513_n819_1;
  wire _abc_4513_n821_1;
  wire _abc_4513_n822_1;
  wire _abc_4513_n823;
  wire _abc_4513_n824;
  wire _abc_4513_n825;
  wire _abc_4513_n826;
  wire _abc_4513_n827;
  wire _abc_4513_n829;
  wire _abc_4513_n830;
  wire _abc_4513_n831;
  wire _abc_4513_n832;
  wire _abc_4513_n833_1;
  wire _abc_4513_n834_1;
  wire _abc_4513_n835_1;
  wire _abc_4513_n836_1;
  wire _abc_4513_n837;
  wire _abc_4513_n838;
  wire _abc_4513_n839;
  wire _abc_4513_n840;
  wire _abc_4513_n842_1;
  wire _abc_4513_n843_1;
  wire _abc_4513_n844_1;
  wire _abc_4513_n845;
  wire _abc_4513_n846;
  wire _abc_4513_n847;
  wire _abc_4513_n848;
  wire _abc_4513_n849;
  wire _abc_4513_n851;
  wire _abc_4513_n852;
  wire _abc_4513_n853;
  wire _abc_4513_n854;
  wire _abc_4513_n856_1;
  wire _abc_4513_n857_1;
  wire _abc_4513_n858_1;
  wire _abc_4513_n859_1;
  wire _abc_4513_n861;
  wire _abc_4513_n862;
  wire _abc_4513_n863;
  wire _abc_4513_n864;
  wire _abc_4513_n866_1;
  wire _abc_4513_n867_1;
  wire _abc_4513_n868_1;
  wire _abc_4513_n869_1;
  wire _abc_4513_n871;
  wire _abc_4513_n872;
  wire _abc_4513_n873;
  wire _abc_4513_n874;
  wire _abc_4513_n876;
  wire _abc_4513_n877;
  wire _abc_4513_n878_1;
  wire _abc_4513_n879_1;
  wire _abc_4513_n881_1;
  wire _abc_4513_n882;
  wire _abc_4513_n883;
  wire _abc_4513_n884;
  wire _abc_4513_n886_1;
  wire _abc_4513_n887_1;
  wire _abc_4513_n888_1;
  wire _abc_4513_n889;
  wire _abc_4513_n890;
  wire _abc_4513_n891;
  wire _abc_4513_n892;
  wire _abc_4513_n893;
  wire _abc_4513_n895;
  wire _abc_4513_n896_1;
  wire _abc_4513_n898;
  wire _abc_4513_n899_1;
  wire _abc_4513_n901;
  wire _abc_4513_n902_1;
  wire _abc_4513_n904_1;
  wire _abc_4513_n905;
  wire _abc_4513_n907;
  wire _abc_4513_n908;
  wire _abc_4513_n910;
  wire _abc_4513_n911;
  wire _abc_4513_n913;
  wire _abc_4513_n914;
  wire _abc_4513_n916;
  wire _abc_4513_n917;
  wire _abc_4513_n919;
  wire _abc_4513_n920;
  wire _abc_4513_n922;
  wire _abc_4513_n923;
  wire _abc_4513_n925;
  wire _abc_4513_n926;
  wire _abc_4513_n928;
  wire _abc_4513_n929;
  wire _abc_4513_n931;
  wire _abc_4513_n932;
  wire _abc_4513_n934;
  wire _abc_4513_n935;
  wire _abc_4513_n937;
  wire _abc_4513_n938;
  wire _abc_4513_n940;
  wire _abc_4513_n941;
  wire _abc_4513_n943;
  wire _abc_4513_n944;
  wire _abc_4513_n946;
  wire _abc_4513_n947;
  wire _abc_4513_n948;
  wire _abc_4513_n949;
  wire _abc_4513_n950;
  wire _abc_4513_n951;
  wire _abc_4513_n952;
  wire _abc_4513_n953;
  wire _abc_4513_n954;
  wire _abc_4513_n955;
  wire _abc_4513_n956;
  wire _abc_4513_n958;
  wire _abc_4513_n959;
  wire _abc_4513_n960;
  wire _abc_4513_n961;
  wire _abc_4513_n962;
  wire _abc_4513_n963;
  wire _abc_4513_n964;
  wire _abc_4513_n965;
  wire _abc_4513_n966;
  wire _abc_4513_n967;
  wire _abc_4513_n968;
  wire _abc_4513_n969;
  wire _abc_4513_n971;
  wire _abc_4513_n972;
  wire _abc_4513_n973;
  wire _abc_4513_n974;
  wire _abc_4513_n975;
  wire _abc_4513_n976;
  wire _abc_4513_n977;
  wire _abc_4513_n978;
  wire _abc_4513_n979;
  wire _abc_4513_n980;
  wire _abc_4513_n981;
  wire _abc_4513_n982;
  wire _abc_4513_n983;
  wire _abc_4513_n984;
  wire _abc_4513_n985;
  wire _abc_4513_n987;
  wire _abc_4513_n988;
  wire _abc_4513_n989;
  wire _abc_4513_n990;
  wire _abc_4513_n991;
  wire _abc_4513_n992;
  wire _abc_4513_n993;
  wire _abc_4513_n994;
  wire _abc_4513_n995;
  wire _abc_4513_n996;
  wire _abc_4513_n997;
  wire _abc_4513_n998;
  output align;
  output \arprot[0] ;
  output \arprot[1] ;
  output \arprot[2] ;
  output \awprot[0] ;
  output \awprot[1] ;
  output \awprot[2] ;
  output busy;
  input clock;
  wire clock_bF_buf0;
  wire clock_bF_buf1;
  wire clock_bF_buf2;
  wire clock_bF_buf3;
  wire clock_bF_buf4;
  wire clock_bF_buf5;
  wire clock_bF_buf6;
  wire clock_bF_buf7;
  output done;
  wire en_instr;
  input enable;
  input \imm[0] ;
  input \imm[10] ;
  input \imm[11] ;
  input \imm[12] ;
  input \imm[13] ;
  input \imm[14] ;
  input \imm[15] ;
  input \imm[16] ;
  input \imm[17] ;
  input \imm[18] ;
  input \imm[19] ;
  input \imm[1] ;
  input \imm[20] ;
  input \imm[21] ;
  input \imm[22] ;
  input \imm[23] ;
  input \imm[24] ;
  input \imm[25] ;
  input \imm[26] ;
  input \imm[27] ;
  input \imm[28] ;
  input \imm[29] ;
  input \imm[2] ;
  input \imm[30] ;
  input \imm[31] ;
  input \imm[3] ;
  input \imm[4] ;
  input \imm[5] ;
  input \imm[6] ;
  input \imm[7] ;
  input \imm[8] ;
  input \imm[9] ;
  output \inst[0] ;
  output \inst[10] ;
  output \inst[11] ;
  output \inst[12] ;
  output \inst[13] ;
  output \inst[14] ;
  output \inst[15] ;
  output \inst[16] ;
  output \inst[17] ;
  output \inst[18] ;
  output \inst[19] ;
  output \inst[1] ;
  output \inst[20] ;
  output \inst[21] ;
  output \inst[22] ;
  output \inst[23] ;
  output \inst[24] ;
  output \inst[25] ;
  output \inst[26] ;
  output \inst[27] ;
  output \inst[28] ;
  output \inst[29] ;
  output \inst[2] ;
  output \inst[30] ;
  output \inst[31] ;
  output \inst[3] ;
  output \inst[4] ;
  output \inst[5] ;
  output \inst[6] ;
  output \inst[7] ;
  output \inst[8] ;
  output \inst[9] ;
  wire inst_0__FF_INPUT;
  wire inst_10__FF_INPUT;
  wire inst_11__FF_INPUT;
  wire inst_12__FF_INPUT;
  wire inst_13__FF_INPUT;
  wire inst_14__FF_INPUT;
  wire inst_15__FF_INPUT;
  wire inst_16__FF_INPUT;
  wire inst_17__FF_INPUT;
  wire inst_18__FF_INPUT;
  wire inst_19__FF_INPUT;
  wire inst_1__FF_INPUT;
  wire inst_20__FF_INPUT;
  wire inst_21__FF_INPUT;
  wire inst_22__FF_INPUT;
  wire inst_23__FF_INPUT;
  wire inst_24__FF_INPUT;
  wire inst_25__FF_INPUT;
  wire inst_26__FF_INPUT;
  wire inst_27__FF_INPUT;
  wire inst_28__FF_INPUT;
  wire inst_29__FF_INPUT;
  wire inst_2__FF_INPUT;
  wire inst_30__FF_INPUT;
  wire inst_31__FF_INPUT;
  wire inst_3__FF_INPUT;
  wire inst_4__FF_INPUT;
  wire inst_5__FF_INPUT;
  wire inst_6__FF_INPUT;
  wire inst_7__FF_INPUT;
  wire inst_8__FF_INPUT;
  wire inst_9__FF_INPUT;
  input \pc[0] ;
  input \pc[10] ;
  input \pc[11] ;
  input \pc[12] ;
  input \pc[13] ;
  input \pc[14] ;
  input \pc[15] ;
  input \pc[16] ;
  input \pc[17] ;
  input \pc[18] ;
  input \pc[19] ;
  input \pc[1] ;
  input \pc[20] ;
  input \pc[21] ;
  input \pc[22] ;
  input \pc[23] ;
  input \pc[24] ;
  input \pc[25] ;
  input \pc[26] ;
  input \pc[27] ;
  input \pc[28] ;
  input \pc[29] ;
  input \pc[2] ;
  input \pc[30] ;
  input \pc[31] ;
  input \pc[3] ;
  input \pc[4] ;
  input \pc[5] ;
  input \pc[6] ;
  input \pc[7] ;
  input \pc[8] ;
  input \pc[9] ;
  output \rd[0] ;
  output \rd[10] ;
  output \rd[11] ;
  output \rd[12] ;
  output \rd[13] ;
  output \rd[14] ;
  output \rd[15] ;
  output \rd[16] ;
  output \rd[17] ;
  output \rd[18] ;
  output \rd[19] ;
  output \rd[1] ;
  output \rd[20] ;
  output \rd[21] ;
  output \rd[22] ;
  output \rd[23] ;
  output \rd[24] ;
  output \rd[25] ;
  output \rd[26] ;
  output \rd[27] ;
  output \rd[28] ;
  output \rd[29] ;
  output \rd[2] ;
  output \rd[30] ;
  output \rd[31] ;
  output \rd[3] ;
  output \rd[4] ;
  output \rd[5] ;
  output \rd[6] ;
  output \rd[7] ;
  output \rd[8] ;
  output \rd[9] ;
  output rd_en;
  input resetn;
  wire resetn_bF_buf0;
  wire resetn_bF_buf1;
  wire resetn_bF_buf2;
  wire resetn_bF_buf3;
  wire resetn_bF_buf4;
  wire resetn_bF_buf5;
  input \rs1[0] ;
  input \rs1[10] ;
  input \rs1[11] ;
  input \rs1[12] ;
  input \rs1[13] ;
  input \rs1[14] ;
  input \rs1[15] ;
  input \rs1[16] ;
  input \rs1[17] ;
  input \rs1[18] ;
  input \rs1[19] ;
  input \rs1[1] ;
  input \rs1[20] ;
  input \rs1[21] ;
  input \rs1[22] ;
  input \rs1[23] ;
  input \rs1[24] ;
  input \rs1[25] ;
  input \rs1[26] ;
  input \rs1[27] ;
  input \rs1[28] ;
  input \rs1[29] ;
  input \rs1[2] ;
  input \rs1[30] ;
  input \rs1[31] ;
  input \rs1[3] ;
  input \rs1[4] ;
  input \rs1[5] ;
  input \rs1[6] ;
  input \rs1[7] ;
  input \rs1[8] ;
  input \rs1[9] ;
  input \rs2[0] ;
  input \rs2[10] ;
  input \rs2[11] ;
  input \rs2[12] ;
  input \rs2[13] ;
  input \rs2[14] ;
  input \rs2[15] ;
  input \rs2[16] ;
  input \rs2[17] ;
  input \rs2[18] ;
  input \rs2[19] ;
  input \rs2[1] ;
  input \rs2[20] ;
  input \rs2[21] ;
  input \rs2[22] ;
  input \rs2[23] ;
  input \rs2[24] ;
  input \rs2[25] ;
  input \rs2[26] ;
  input \rs2[27] ;
  input \rs2[28] ;
  input \rs2[29] ;
  input \rs2[2] ;
  input \rs2[30] ;
  input \rs2[31] ;
  input \rs2[3] ;
  input \rs2[4] ;
  input \rs2[5] ;
  input \rs2[6] ;
  input \rs2[7] ;
  input \rs2[8] ;
  input \rs2[9] ;
  input signo;
  wire state_0_;
  wire state_1_;
  wire state_2_;
  wire state_3_;
  wire state_4_;
  wire state_5_;
  wire state_6_;
  input \wordsize[0] ;
  input \wordsize[1] ;
  AND2X2 AND2X2_1 ( .A(_abc_4513_n362_1), .B(enable), .Y(_abc_4513_n363_1) );
  AND2X2 AND2X2_10 ( .A(_abc_4513_n375_1), .B(resetn), .Y(_abc_4513_n376) );
  AND2X2 AND2X2_100 ( .A(_abc_4513_n521), .B(\inst[4] ), .Y(_abc_4513_n538) );
  AND2X2 AND2X2_101 ( .A(_abc_4513_n539_1), .B(resetn), .Y(inst_4__FF_INPUT) );
  AND2X2 AND2X2_102 ( .A(_abc_4513_n519_1), .B(\Rdata_mem[5] ), .Y(_abc_4513_n541_1) );
  AND2X2 AND2X2_103 ( .A(_abc_4513_n521), .B(\inst[5] ), .Y(_abc_4513_n542) );
  AND2X2 AND2X2_104 ( .A(_abc_4513_n543_1), .B(resetn), .Y(inst_5__FF_INPUT) );
  AND2X2 AND2X2_105 ( .A(_abc_4513_n519_1), .B(\Rdata_mem[6] ), .Y(_abc_4513_n545_1) );
  AND2X2 AND2X2_106 ( .A(_abc_4513_n521), .B(\inst[6] ), .Y(_abc_4513_n546) );
  AND2X2 AND2X2_107 ( .A(_abc_4513_n547_1), .B(resetn), .Y(inst_6__FF_INPUT) );
  AND2X2 AND2X2_108 ( .A(_abc_4513_n519_1), .B(\Rdata_mem[7] ), .Y(_abc_4513_n549_1) );
  AND2X2 AND2X2_109 ( .A(_abc_4513_n521), .B(\inst[7] ), .Y(_abc_4513_n550) );
  AND2X2 AND2X2_11 ( .A(_abc_4513_n372), .B(AWready), .Y(_abc_4513_n377_1) );
  AND2X2 AND2X2_110 ( .A(_abc_4513_n551_1), .B(resetn), .Y(inst_7__FF_INPUT) );
  AND2X2 AND2X2_111 ( .A(_abc_4513_n519_1), .B(\Rdata_mem[8] ), .Y(_abc_4513_n553_1) );
  AND2X2 AND2X2_112 ( .A(_abc_4513_n521), .B(\inst[8] ), .Y(_abc_4513_n554) );
  AND2X2 AND2X2_113 ( .A(_abc_4513_n555_1), .B(resetn), .Y(inst_8__FF_INPUT) );
  AND2X2 AND2X2_114 ( .A(_abc_4513_n519_1), .B(\Rdata_mem[9] ), .Y(_abc_4513_n557_1) );
  AND2X2 AND2X2_115 ( .A(_abc_4513_n521), .B(\inst[9] ), .Y(_abc_4513_n558) );
  AND2X2 AND2X2_116 ( .A(_abc_4513_n559_1), .B(resetn), .Y(inst_9__FF_INPUT) );
  AND2X2 AND2X2_117 ( .A(_abc_4513_n519_1), .B(\Rdata_mem[10] ), .Y(_abc_4513_n561_1) );
  AND2X2 AND2X2_118 ( .A(_abc_4513_n521), .B(\inst[10] ), .Y(_abc_4513_n562) );
  AND2X2 AND2X2_119 ( .A(_abc_4513_n563_1), .B(resetn), .Y(inst_10__FF_INPUT) );
  AND2X2 AND2X2_12 ( .A(resetn), .B(state_4_), .Y(_abc_4513_n378_1) );
  AND2X2 AND2X2_120 ( .A(_abc_4513_n519_1), .B(\Rdata_mem[11] ), .Y(_abc_4513_n565_1) );
  AND2X2 AND2X2_121 ( .A(_abc_4513_n521), .B(\inst[11] ), .Y(_abc_4513_n566_1) );
  AND2X2 AND2X2_122 ( .A(_abc_4513_n567_1), .B(resetn), .Y(inst_11__FF_INPUT) );
  AND2X2 AND2X2_123 ( .A(_abc_4513_n519_1), .B(\Rdata_mem[12] ), .Y(_abc_4513_n569_1) );
  AND2X2 AND2X2_124 ( .A(_abc_4513_n521), .B(\inst[12] ), .Y(_abc_4513_n570) );
  AND2X2 AND2X2_125 ( .A(_abc_4513_n571), .B(resetn), .Y(inst_12__FF_INPUT) );
  AND2X2 AND2X2_126 ( .A(_abc_4513_n519_1), .B(\Rdata_mem[13] ), .Y(_abc_4513_n573) );
  AND2X2 AND2X2_127 ( .A(_abc_4513_n521), .B(\inst[13] ), .Y(_abc_4513_n574_1) );
  AND2X2 AND2X2_128 ( .A(_abc_4513_n575_1), .B(resetn), .Y(inst_13__FF_INPUT) );
  AND2X2 AND2X2_129 ( .A(_abc_4513_n519_1), .B(\Rdata_mem[14] ), .Y(_abc_4513_n577_1) );
  AND2X2 AND2X2_13 ( .A(enable), .B(state_0_), .Y(_abc_4513_n380_1) );
  AND2X2 AND2X2_130 ( .A(_abc_4513_n521), .B(\inst[14] ), .Y(_abc_4513_n578) );
  AND2X2 AND2X2_131 ( .A(_abc_4513_n579), .B(resetn), .Y(inst_14__FF_INPUT) );
  AND2X2 AND2X2_132 ( .A(_abc_4513_n519_1), .B(\Rdata_mem[15] ), .Y(_abc_4513_n581) );
  AND2X2 AND2X2_133 ( .A(_abc_4513_n521), .B(\inst[15] ), .Y(_abc_4513_n582) );
  AND2X2 AND2X2_134 ( .A(_abc_4513_n583_1), .B(resetn), .Y(inst_15__FF_INPUT) );
  AND2X2 AND2X2_135 ( .A(_abc_4513_n519_1), .B(\Rdata_mem[16] ), .Y(_abc_4513_n585_1) );
  AND2X2 AND2X2_136 ( .A(_abc_4513_n521), .B(\inst[16] ), .Y(_abc_4513_n586_1) );
  AND2X2 AND2X2_137 ( .A(_abc_4513_n587), .B(resetn), .Y(inst_16__FF_INPUT) );
  AND2X2 AND2X2_138 ( .A(_abc_4513_n519_1), .B(\Rdata_mem[17] ), .Y(_abc_4513_n589) );
  AND2X2 AND2X2_139 ( .A(_abc_4513_n521), .B(\inst[17] ), .Y(_abc_4513_n590) );
  AND2X2 AND2X2_14 ( .A(_abc_4513_n379), .B(_abc_4513_n380_1), .Y(_abc_4513_n381_1) );
  AND2X2 AND2X2_140 ( .A(_abc_4513_n591), .B(resetn), .Y(inst_17__FF_INPUT) );
  AND2X2 AND2X2_141 ( .A(_abc_4513_n519_1), .B(\Rdata_mem[18] ), .Y(_abc_4513_n593) );
  AND2X2 AND2X2_142 ( .A(_abc_4513_n521), .B(\inst[18] ), .Y(_abc_4513_n594_1) );
  AND2X2 AND2X2_143 ( .A(_abc_4513_n595_1), .B(resetn), .Y(inst_18__FF_INPUT) );
  AND2X2 AND2X2_144 ( .A(_abc_4513_n519_1), .B(\Rdata_mem[19] ), .Y(_abc_4513_n597_1) );
  AND2X2 AND2X2_145 ( .A(_abc_4513_n521), .B(\inst[19] ), .Y(_abc_4513_n598) );
  AND2X2 AND2X2_146 ( .A(_abc_4513_n599), .B(resetn), .Y(inst_19__FF_INPUT) );
  AND2X2 AND2X2_147 ( .A(_abc_4513_n519_1), .B(\Rdata_mem[20] ), .Y(_abc_4513_n601) );
  AND2X2 AND2X2_148 ( .A(_abc_4513_n521), .B(\inst[20] ), .Y(_abc_4513_n602_1) );
  AND2X2 AND2X2_149 ( .A(_abc_4513_n603_1), .B(resetn), .Y(inst_20__FF_INPUT) );
  AND2X2 AND2X2_15 ( .A(_abc_4513_n381_1), .B(resetn), .Y(_abc_4513_n382) );
  AND2X2 AND2X2_150 ( .A(_abc_4513_n519_1), .B(\Rdata_mem[21] ), .Y(_abc_4513_n605_1) );
  AND2X2 AND2X2_151 ( .A(_abc_4513_n521), .B(\inst[21] ), .Y(_abc_4513_n606) );
  AND2X2 AND2X2_152 ( .A(_abc_4513_n607), .B(resetn), .Y(inst_21__FF_INPUT) );
  AND2X2 AND2X2_153 ( .A(_abc_4513_n519_1), .B(\Rdata_mem[22] ), .Y(_abc_4513_n609) );
  AND2X2 AND2X2_154 ( .A(_abc_4513_n521), .B(\inst[22] ), .Y(_abc_4513_n610) );
  AND2X2 AND2X2_155 ( .A(_abc_4513_n611), .B(resetn), .Y(inst_22__FF_INPUT) );
  AND2X2 AND2X2_156 ( .A(_abc_4513_n519_1), .B(\Rdata_mem[23] ), .Y(_abc_4513_n613_1) );
  AND2X2 AND2X2_157 ( .A(_abc_4513_n521), .B(\inst[23] ), .Y(_abc_4513_n614_1) );
  AND2X2 AND2X2_158 ( .A(_abc_4513_n615_1), .B(resetn), .Y(inst_23__FF_INPUT) );
  AND2X2 AND2X2_159 ( .A(_abc_4513_n519_1), .B(\Rdata_mem[24] ), .Y(_abc_4513_n617) );
  AND2X2 AND2X2_16 ( .A(_abc_4513_n382), .B(AWready), .Y(_abc_4513_n383_1) );
  AND2X2 AND2X2_160 ( .A(_abc_4513_n521), .B(\inst[24] ), .Y(_abc_4513_n618) );
  AND2X2 AND2X2_161 ( .A(_abc_4513_n619), .B(resetn), .Y(inst_24__FF_INPUT) );
  AND2X2 AND2X2_162 ( .A(_abc_4513_n519_1), .B(\Rdata_mem[25] ), .Y(_abc_4513_n621) );
  AND2X2 AND2X2_163 ( .A(_abc_4513_n521), .B(\inst[25] ), .Y(_abc_4513_n622_1) );
  AND2X2 AND2X2_164 ( .A(_abc_4513_n623_1), .B(resetn), .Y(inst_25__FF_INPUT) );
  AND2X2 AND2X2_165 ( .A(_abc_4513_n519_1), .B(\Rdata_mem[26] ), .Y(_abc_4513_n625_1) );
  AND2X2 AND2X2_166 ( .A(_abc_4513_n521), .B(\inst[26] ), .Y(_abc_4513_n626) );
  AND2X2 AND2X2_167 ( .A(_abc_4513_n627), .B(resetn), .Y(inst_26__FF_INPUT) );
  AND2X2 AND2X2_168 ( .A(_abc_4513_n519_1), .B(\Rdata_mem[27] ), .Y(_abc_4513_n629) );
  AND2X2 AND2X2_169 ( .A(_abc_4513_n521), .B(\inst[27] ), .Y(_abc_4513_n630) );
  AND2X2 AND2X2_17 ( .A(_abc_4513_n384_1), .B(_abc_4513_n377_1), .Y(_abc_4513_n385) );
  AND2X2 AND2X2_170 ( .A(_abc_4513_n631), .B(resetn), .Y(inst_27__FF_INPUT) );
  AND2X2 AND2X2_171 ( .A(_abc_4513_n519_1), .B(\Rdata_mem[28] ), .Y(_abc_4513_n633) );
  AND2X2 AND2X2_172 ( .A(_abc_4513_n521), .B(\inst[28] ), .Y(_abc_4513_n634) );
  AND2X2 AND2X2_173 ( .A(_abc_4513_n635), .B(resetn), .Y(inst_28__FF_INPUT) );
  AND2X2 AND2X2_174 ( .A(_abc_4513_n519_1), .B(\Rdata_mem[29] ), .Y(_abc_4513_n637_1) );
  AND2X2 AND2X2_175 ( .A(_abc_4513_n521), .B(\inst[29] ), .Y(_abc_4513_n638_1) );
  AND2X2 AND2X2_176 ( .A(_abc_4513_n639_1), .B(resetn), .Y(inst_29__FF_INPUT) );
  AND2X2 AND2X2_177 ( .A(_abc_4513_n519_1), .B(\Rdata_mem[30] ), .Y(_abc_4513_n641) );
  AND2X2 AND2X2_178 ( .A(_abc_4513_n521), .B(\inst[30] ), .Y(_abc_4513_n642) );
  AND2X2 AND2X2_179 ( .A(_abc_4513_n643), .B(resetn), .Y(inst_30__FF_INPUT) );
  AND2X2 AND2X2_18 ( .A(_abc_4513_n387_1), .B(state_5_), .Y(_abc_4513_n388) );
  AND2X2 AND2X2_180 ( .A(_abc_4513_n519_1), .B(\Rdata_mem[31] ), .Y(_abc_4513_n645_1) );
  AND2X2 AND2X2_181 ( .A(_abc_4513_n521), .B(\inst[31] ), .Y(_abc_4513_n646_1) );
  AND2X2 AND2X2_182 ( .A(_abc_4513_n647_1), .B(resetn), .Y(inst_31__FF_INPUT) );
  AND2X2 AND2X2_183 ( .A(_abc_4513_n473), .B(\rs2[0] ), .Y(Wdata_0__FF_INPUT) );
  AND2X2 AND2X2_184 ( .A(_abc_4513_n473), .B(\rs2[1] ), .Y(Wdata_1__FF_INPUT) );
  AND2X2 AND2X2_185 ( .A(_abc_4513_n473), .B(\rs2[2] ), .Y(Wdata_2__FF_INPUT) );
  AND2X2 AND2X2_186 ( .A(_abc_4513_n473), .B(\rs2[3] ), .Y(Wdata_3__FF_INPUT) );
  AND2X2 AND2X2_187 ( .A(_abc_4513_n473), .B(\rs2[4] ), .Y(Wdata_4__FF_INPUT) );
  AND2X2 AND2X2_188 ( .A(_abc_4513_n473), .B(\rs2[5] ), .Y(Wdata_5__FF_INPUT) );
  AND2X2 AND2X2_189 ( .A(_abc_4513_n473), .B(\rs2[6] ), .Y(Wdata_6__FF_INPUT) );
  AND2X2 AND2X2_19 ( .A(_abc_4513_n388), .B(resetn), .Y(_abc_4513_n389_1) );
  AND2X2 AND2X2_190 ( .A(_abc_4513_n473), .B(\rs2[7] ), .Y(Wdata_7__FF_INPUT) );
  AND2X2 AND2X2_191 ( .A(_abc_4513_n476), .B(\rs2[0] ), .Y(_abc_4513_n657_1) );
  AND2X2 AND2X2_192 ( .A(_abc_4513_n658_1), .B(\rs2[8] ), .Y(_abc_4513_n659_1) );
  AND2X2 AND2X2_193 ( .A(_abc_4513_n660_1), .B(_abc_4513_n473), .Y(Wdata_8__FF_INPUT) );
  AND2X2 AND2X2_194 ( .A(_abc_4513_n476), .B(\rs2[1] ), .Y(_abc_4513_n662) );
  AND2X2 AND2X2_195 ( .A(_abc_4513_n658_1), .B(\rs2[9] ), .Y(_abc_4513_n663) );
  AND2X2 AND2X2_196 ( .A(_abc_4513_n664), .B(_abc_4513_n473), .Y(Wdata_9__FF_INPUT) );
  AND2X2 AND2X2_197 ( .A(_abc_4513_n476), .B(\rs2[2] ), .Y(_abc_4513_n666_1) );
  AND2X2 AND2X2_198 ( .A(_abc_4513_n658_1), .B(\rs2[10] ), .Y(_abc_4513_n667_1) );
  AND2X2 AND2X2_199 ( .A(_abc_4513_n668_1), .B(_abc_4513_n473), .Y(Wdata_10__FF_INPUT) );
  AND2X2 AND2X2_2 ( .A(_abc_4513_n363_1), .B(state_0_), .Y(_abc_4513_n364) );
  AND2X2 AND2X2_20 ( .A(_abc_4513_n387_1), .B(ARready), .Y(_abc_4513_n390_1) );
  AND2X2 AND2X2_200 ( .A(_abc_4513_n476), .B(\rs2[3] ), .Y(_abc_4513_n670) );
  AND2X2 AND2X2_201 ( .A(_abc_4513_n658_1), .B(\rs2[11] ), .Y(_abc_4513_n671) );
  AND2X2 AND2X2_202 ( .A(_abc_4513_n672), .B(_abc_4513_n473), .Y(Wdata_11__FF_INPUT) );
  AND2X2 AND2X2_203 ( .A(_abc_4513_n476), .B(\rs2[4] ), .Y(_abc_4513_n674) );
  AND2X2 AND2X2_204 ( .A(_abc_4513_n658_1), .B(\rs2[12] ), .Y(_abc_4513_n675) );
  AND2X2 AND2X2_205 ( .A(_abc_4513_n676), .B(_abc_4513_n473), .Y(Wdata_12__FF_INPUT) );
  AND2X2 AND2X2_206 ( .A(_abc_4513_n476), .B(\rs2[5] ), .Y(_abc_4513_n678) );
  AND2X2 AND2X2_207 ( .A(_abc_4513_n658_1), .B(\rs2[13] ), .Y(_abc_4513_n679) );
  AND2X2 AND2X2_208 ( .A(_abc_4513_n680_1), .B(_abc_4513_n473), .Y(Wdata_13__FF_INPUT) );
  AND2X2 AND2X2_209 ( .A(_abc_4513_n476), .B(\rs2[6] ), .Y(_abc_4513_n682_1) );
  AND2X2 AND2X2_21 ( .A(ARvalid), .B(_abc_4513_n390_1), .Y(_abc_4513_n391) );
  AND2X2 AND2X2_210 ( .A(_abc_4513_n658_1), .B(\rs2[14] ), .Y(_abc_4513_n683_1) );
  AND2X2 AND2X2_211 ( .A(_abc_4513_n684), .B(_abc_4513_n473), .Y(Wdata_14__FF_INPUT) );
  AND2X2 AND2X2_212 ( .A(_abc_4513_n476), .B(\rs2[7] ), .Y(_abc_4513_n686) );
  AND2X2 AND2X2_213 ( .A(_abc_4513_n658_1), .B(\rs2[15] ), .Y(_abc_4513_n687) );
  AND2X2 AND2X2_214 ( .A(_abc_4513_n688_1), .B(_abc_4513_n473), .Y(Wdata_15__FF_INPUT) );
  AND2X2 AND2X2_215 ( .A(_abc_4513_n475), .B(\rs2[0] ), .Y(_abc_4513_n690_1) );
  AND2X2 AND2X2_216 ( .A(_abc_4513_n495_1), .B(\rs2[16] ), .Y(_abc_4513_n691_1) );
  AND2X2 AND2X2_217 ( .A(_abc_4513_n692), .B(_abc_4513_n473), .Y(Wdata_16__FF_INPUT) );
  AND2X2 AND2X2_218 ( .A(_abc_4513_n475), .B(\rs2[1] ), .Y(_abc_4513_n694) );
  AND2X2 AND2X2_219 ( .A(_abc_4513_n495_1), .B(\rs2[17] ), .Y(_abc_4513_n695) );
  AND2X2 AND2X2_22 ( .A(Wready), .B(Bvalid), .Y(_abc_4513_n393_1) );
  AND2X2 AND2X2_220 ( .A(_abc_4513_n696), .B(_abc_4513_n473), .Y(Wdata_17__FF_INPUT) );
  AND2X2 AND2X2_221 ( .A(_abc_4513_n475), .B(\rs2[2] ), .Y(_abc_4513_n698) );
  AND2X2 AND2X2_222 ( .A(_abc_4513_n495_1), .B(\rs2[18] ), .Y(_abc_4513_n699_1) );
  AND2X2 AND2X2_223 ( .A(_abc_4513_n700_1), .B(_abc_4513_n473), .Y(Wdata_18__FF_INPUT) );
  AND2X2 AND2X2_224 ( .A(_abc_4513_n475), .B(\rs2[3] ), .Y(_abc_4513_n702_1) );
  AND2X2 AND2X2_225 ( .A(_abc_4513_n495_1), .B(\rs2[19] ), .Y(_abc_4513_n703) );
  AND2X2 AND2X2_226 ( .A(_abc_4513_n704), .B(_abc_4513_n473), .Y(Wdata_19__FF_INPUT) );
  AND2X2 AND2X2_227 ( .A(_abc_4513_n475), .B(\rs2[4] ), .Y(_abc_4513_n706) );
  AND2X2 AND2X2_228 ( .A(_abc_4513_n495_1), .B(\rs2[20] ), .Y(_abc_4513_n707) );
  AND2X2 AND2X2_229 ( .A(_abc_4513_n708_1), .B(_abc_4513_n473), .Y(Wdata_20__FF_INPUT) );
  AND2X2 AND2X2_23 ( .A(_abc_4513_n394), .B(Wready), .Y(_abc_4513_n395_1) );
  AND2X2 AND2X2_230 ( .A(_abc_4513_n475), .B(\rs2[5] ), .Y(_abc_4513_n710_1) );
  AND2X2 AND2X2_231 ( .A(_abc_4513_n495_1), .B(\rs2[21] ), .Y(_abc_4513_n711_1) );
  AND2X2 AND2X2_232 ( .A(_abc_4513_n712), .B(_abc_4513_n473), .Y(Wdata_21__FF_INPUT) );
  AND2X2 AND2X2_233 ( .A(_abc_4513_n475), .B(\rs2[6] ), .Y(_abc_4513_n714) );
  AND2X2 AND2X2_234 ( .A(_abc_4513_n495_1), .B(\rs2[22] ), .Y(_abc_4513_n715) );
  AND2X2 AND2X2_235 ( .A(_abc_4513_n716), .B(_abc_4513_n473), .Y(Wdata_22__FF_INPUT) );
  AND2X2 AND2X2_236 ( .A(_abc_4513_n475), .B(\rs2[7] ), .Y(_abc_4513_n718) );
  AND2X2 AND2X2_237 ( .A(_abc_4513_n495_1), .B(\rs2[23] ), .Y(_abc_4513_n719) );
  AND2X2 AND2X2_238 ( .A(_abc_4513_n720), .B(_abc_4513_n473), .Y(Wdata_23__FF_INPUT) );
  AND2X2 AND2X2_239 ( .A(_abc_4513_n496), .B(\rs2[8] ), .Y(_abc_4513_n722) );
  AND2X2 AND2X2_24 ( .A(_abc_4513_n397), .B(AWready), .Y(_abc_4513_n398_1) );
  AND2X2 AND2X2_240 ( .A(_abc_4513_n495_1), .B(\rs2[24] ), .Y(_abc_4513_n724) );
  AND2X2 AND2X2_241 ( .A(_abc_4513_n725), .B(_abc_4513_n473), .Y(Wdata_24__FF_INPUT) );
  AND2X2 AND2X2_242 ( .A(_abc_4513_n496), .B(\rs2[9] ), .Y(_abc_4513_n727_1) );
  AND2X2 AND2X2_243 ( .A(_abc_4513_n495_1), .B(\rs2[25] ), .Y(_abc_4513_n729_1) );
  AND2X2 AND2X2_244 ( .A(_abc_4513_n730), .B(_abc_4513_n473), .Y(Wdata_25__FF_INPUT) );
  AND2X2 AND2X2_245 ( .A(_abc_4513_n496), .B(\rs2[10] ), .Y(_abc_4513_n732) );
  AND2X2 AND2X2_246 ( .A(_abc_4513_n495_1), .B(\rs2[26] ), .Y(_abc_4513_n734) );
  AND2X2 AND2X2_247 ( .A(_abc_4513_n735_1), .B(_abc_4513_n473), .Y(Wdata_26__FF_INPUT) );
  AND2X2 AND2X2_248 ( .A(_abc_4513_n496), .B(\rs2[11] ), .Y(_abc_4513_n737_1) );
  AND2X2 AND2X2_249 ( .A(_abc_4513_n495_1), .B(\rs2[27] ), .Y(_abc_4513_n739) );
  AND2X2 AND2X2_25 ( .A(_abc_4513_n396_1), .B(_abc_4513_n399_1), .Y(_abc_4513_n400) );
  AND2X2 AND2X2_250 ( .A(_abc_4513_n740), .B(_abc_4513_n473), .Y(Wdata_27__FF_INPUT) );
  AND2X2 AND2X2_251 ( .A(_abc_4513_n496), .B(\rs2[12] ), .Y(_abc_4513_n742) );
  AND2X2 AND2X2_252 ( .A(_abc_4513_n495_1), .B(\rs2[28] ), .Y(_abc_4513_n744) );
  AND2X2 AND2X2_253 ( .A(_abc_4513_n745_1), .B(_abc_4513_n473), .Y(Wdata_28__FF_INPUT) );
  AND2X2 AND2X2_254 ( .A(_abc_4513_n496), .B(\rs2[13] ), .Y(_abc_4513_n747_1) );
  AND2X2 AND2X2_255 ( .A(_abc_4513_n495_1), .B(\rs2[29] ), .Y(_abc_4513_n749) );
  AND2X2 AND2X2_256 ( .A(_abc_4513_n750), .B(_abc_4513_n473), .Y(Wdata_29__FF_INPUT) );
  AND2X2 AND2X2_257 ( .A(_abc_4513_n496), .B(\rs2[14] ), .Y(_abc_4513_n752) );
  AND2X2 AND2X2_258 ( .A(_abc_4513_n495_1), .B(\rs2[30] ), .Y(_abc_4513_n754_1) );
  AND2X2 AND2X2_259 ( .A(_abc_4513_n755_1), .B(_abc_4513_n473), .Y(Wdata_30__FF_INPUT) );
  AND2X2 AND2X2_26 ( .A(_abc_4513_n401_1), .B(resetn), .Y(_abc_4513_n402_1) );
  AND2X2 AND2X2_260 ( .A(_abc_4513_n496), .B(\rs2[15] ), .Y(_abc_4513_n757) );
  AND2X2 AND2X2_261 ( .A(_abc_4513_n495_1), .B(\rs2[31] ), .Y(_abc_4513_n759) );
  AND2X2 AND2X2_262 ( .A(_abc_4513_n760), .B(_abc_4513_n473), .Y(Wdata_31__FF_INPUT) );
  AND2X2 AND2X2_263 ( .A(_abc_4513_n493), .B(_abc_4513_n495_1), .Y(_abc_4513_n762) );
  AND2X2 AND2X2_264 ( .A(_abc_4513_n492), .B(_abc_4513_n496), .Y(_abc_4513_n763) );
  AND2X2 AND2X2_265 ( .A(_abc_4513_n769_1), .B(\W_R[0] ), .Y(_abc_4513_n770) );
  AND2X2 AND2X2_266 ( .A(_abc_4513_n471), .B(_abc_4513_n770), .Y(_abc_4513_n771) );
  AND2X2 AND2X2_267 ( .A(_abc_4513_n772), .B(\Rdata_mem[16] ), .Y(_abc_4513_n773) );
  AND2X2 AND2X2_268 ( .A(_abc_4513_n499), .B(\Rdata_mem[0] ), .Y(_abc_4513_n774_1) );
  AND2X2 AND2X2_269 ( .A(_abc_4513_n502), .B(\Rdata_mem[8] ), .Y(_abc_4513_n775_1) );
  AND2X2 AND2X2_27 ( .A(_abc_4513_n400), .B(_abc_4513_n402_1), .Y(_abc_4513_n403) );
  AND2X2 AND2X2_270 ( .A(_abc_4513_n513_1), .B(\Rdata_mem[24] ), .Y(_abc_4513_n776_1) );
  AND2X2 AND2X2_271 ( .A(_abc_4513_n779), .B(_abc_4513_n771), .Y(\rd[0] ) );
  AND2X2 AND2X2_272 ( .A(_abc_4513_n499), .B(\Rdata_mem[1] ), .Y(_abc_4513_n781) );
  AND2X2 AND2X2_273 ( .A(_abc_4513_n772), .B(\Rdata_mem[17] ), .Y(_abc_4513_n782) );
  AND2X2 AND2X2_274 ( .A(_abc_4513_n502), .B(\Rdata_mem[9] ), .Y(_abc_4513_n783) );
  AND2X2 AND2X2_275 ( .A(_abc_4513_n513_1), .B(\Rdata_mem[25] ), .Y(_abc_4513_n784) );
  AND2X2 AND2X2_276 ( .A(_abc_4513_n787_1), .B(_abc_4513_n771), .Y(\rd[1] ) );
  AND2X2 AND2X2_277 ( .A(_abc_4513_n772), .B(\Rdata_mem[18] ), .Y(_abc_4513_n789_1) );
  AND2X2 AND2X2_278 ( .A(_abc_4513_n499), .B(\Rdata_mem[2] ), .Y(_abc_4513_n790) );
  AND2X2 AND2X2_279 ( .A(_abc_4513_n513_1), .B(\Rdata_mem[26] ), .Y(_abc_4513_n791) );
  AND2X2 AND2X2_28 ( .A(_abc_4513_n403), .B(state_4_), .Y(_abc_4513_n404_1) );
  AND2X2 AND2X2_280 ( .A(_abc_4513_n502), .B(\Rdata_mem[10] ), .Y(_abc_4513_n792) );
  AND2X2 AND2X2_281 ( .A(_abc_4513_n795_1), .B(_abc_4513_n771), .Y(\rd[2] ) );
  AND2X2 AND2X2_282 ( .A(_abc_4513_n499), .B(\Rdata_mem[3] ), .Y(_abc_4513_n797_1) );
  AND2X2 AND2X2_283 ( .A(_abc_4513_n772), .B(\Rdata_mem[19] ), .Y(_abc_4513_n798) );
  AND2X2 AND2X2_284 ( .A(_abc_4513_n502), .B(\Rdata_mem[11] ), .Y(_abc_4513_n799) );
  AND2X2 AND2X2_285 ( .A(_abc_4513_n513_1), .B(\Rdata_mem[27] ), .Y(_abc_4513_n800) );
  AND2X2 AND2X2_286 ( .A(_abc_4513_n803), .B(_abc_4513_n771), .Y(\rd[3] ) );
  AND2X2 AND2X2_287 ( .A(_abc_4513_n772), .B(\Rdata_mem[20] ), .Y(_abc_4513_n805) );
  AND2X2 AND2X2_288 ( .A(_abc_4513_n499), .B(\Rdata_mem[4] ), .Y(_abc_4513_n806) );
  AND2X2 AND2X2_289 ( .A(_abc_4513_n502), .B(\Rdata_mem[12] ), .Y(_abc_4513_n807) );
  AND2X2 AND2X2_29 ( .A(_abc_4513_n405_1), .B(AWready), .Y(_abc_4513_n406) );
  AND2X2 AND2X2_290 ( .A(_abc_4513_n513_1), .B(\Rdata_mem[28] ), .Y(_abc_4513_n808) );
  AND2X2 AND2X2_291 ( .A(_abc_4513_n811_1), .B(_abc_4513_n771), .Y(\rd[4] ) );
  AND2X2 AND2X2_292 ( .A(_abc_4513_n499), .B(\Rdata_mem[5] ), .Y(_abc_4513_n813_1) );
  AND2X2 AND2X2_293 ( .A(_abc_4513_n772), .B(\Rdata_mem[21] ), .Y(_abc_4513_n814_1) );
  AND2X2 AND2X2_294 ( .A(_abc_4513_n502), .B(\Rdata_mem[13] ), .Y(_abc_4513_n815) );
  AND2X2 AND2X2_295 ( .A(_abc_4513_n513_1), .B(\Rdata_mem[29] ), .Y(_abc_4513_n816) );
  AND2X2 AND2X2_296 ( .A(_abc_4513_n819_1), .B(_abc_4513_n771), .Y(\rd[5] ) );
  AND2X2 AND2X2_297 ( .A(_abc_4513_n772), .B(\Rdata_mem[22] ), .Y(_abc_4513_n821_1) );
  AND2X2 AND2X2_298 ( .A(_abc_4513_n499), .B(\Rdata_mem[6] ), .Y(_abc_4513_n822_1) );
  AND2X2 AND2X2_299 ( .A(_abc_4513_n513_1), .B(\Rdata_mem[30] ), .Y(_abc_4513_n823) );
  AND2X2 AND2X2_3 ( .A(_abc_4513_n365), .B(resetn), .Y(ARvalid) );
  AND2X2 AND2X2_30 ( .A(_abc_4513_n407_1), .B(_abc_4513_n393_1), .Y(_abc_4513_n408_1) );
  AND2X2 AND2X2_300 ( .A(_abc_4513_n502), .B(\Rdata_mem[14] ), .Y(_abc_4513_n824) );
  AND2X2 AND2X2_301 ( .A(_abc_4513_n827), .B(_abc_4513_n771), .Y(\rd[6] ) );
  AND2X2 AND2X2_302 ( .A(_abc_4513_n508), .B(\Rdata_mem[23] ), .Y(_abc_4513_n829) );
  AND2X2 AND2X2_303 ( .A(_abc_4513_n512), .B(\Rdata_mem[31] ), .Y(_abc_4513_n830) );
  AND2X2 AND2X2_304 ( .A(_abc_4513_n493), .B(\Rdata_mem[7] ), .Y(_abc_4513_n832) );
  AND2X2 AND2X2_305 ( .A(_abc_4513_n501), .B(\Rdata_mem[15] ), .Y(_abc_4513_n833_1) );
  AND2X2 AND2X2_306 ( .A(_abc_4513_n835_1), .B(_abc_4513_n476), .Y(_abc_4513_n836_1) );
  AND2X2 AND2X2_307 ( .A(_abc_4513_n506), .B(\Rdata_mem[23] ), .Y(_abc_4513_n837) );
  AND2X2 AND2X2_308 ( .A(_abc_4513_n498), .B(\Rdata_mem[7] ), .Y(_abc_4513_n838) );
  AND2X2 AND2X2_309 ( .A(_abc_4513_n840), .B(_abc_4513_n771), .Y(\rd[7] ) );
  AND2X2 AND2X2_31 ( .A(Rvalid), .B(ARready), .Y(_abc_4513_n409) );
  AND2X2 AND2X2_310 ( .A(_abc_4513_n843_1), .B(signo), .Y(_abc_4513_n844_1) );
  AND2X2 AND2X2_311 ( .A(_abc_4513_n836_1), .B(_abc_4513_n844_1), .Y(_abc_4513_n845) );
  AND2X2 AND2X2_312 ( .A(_abc_4513_n506), .B(\Rdata_mem[24] ), .Y(_abc_4513_n846) );
  AND2X2 AND2X2_313 ( .A(_abc_4513_n498), .B(\Rdata_mem[8] ), .Y(_abc_4513_n847) );
  AND2X2 AND2X2_314 ( .A(_abc_4513_n849), .B(_abc_4513_n771), .Y(\rd[8] ) );
  AND2X2 AND2X2_315 ( .A(_abc_4513_n506), .B(\Rdata_mem[25] ), .Y(_abc_4513_n851) );
  AND2X2 AND2X2_316 ( .A(_abc_4513_n498), .B(\Rdata_mem[9] ), .Y(_abc_4513_n852) );
  AND2X2 AND2X2_317 ( .A(_abc_4513_n854), .B(_abc_4513_n771), .Y(\rd[9] ) );
  AND2X2 AND2X2_318 ( .A(_abc_4513_n506), .B(\Rdata_mem[26] ), .Y(_abc_4513_n856_1) );
  AND2X2 AND2X2_319 ( .A(_abc_4513_n498), .B(\Rdata_mem[10] ), .Y(_abc_4513_n857_1) );
  AND2X2 AND2X2_32 ( .A(_abc_4513_n364), .B(_abc_4513_n409), .Y(_abc_4513_n410_1) );
  AND2X2 AND2X2_320 ( .A(_abc_4513_n859_1), .B(_abc_4513_n771), .Y(\rd[10] ) );
  AND2X2 AND2X2_321 ( .A(_abc_4513_n506), .B(\Rdata_mem[27] ), .Y(_abc_4513_n861) );
  AND2X2 AND2X2_322 ( .A(_abc_4513_n498), .B(\Rdata_mem[11] ), .Y(_abc_4513_n862) );
  AND2X2 AND2X2_323 ( .A(_abc_4513_n864), .B(_abc_4513_n771), .Y(\rd[11] ) );
  AND2X2 AND2X2_324 ( .A(_abc_4513_n506), .B(\Rdata_mem[28] ), .Y(_abc_4513_n866_1) );
  AND2X2 AND2X2_325 ( .A(_abc_4513_n498), .B(\Rdata_mem[12] ), .Y(_abc_4513_n867_1) );
  AND2X2 AND2X2_326 ( .A(_abc_4513_n869_1), .B(_abc_4513_n771), .Y(\rd[12] ) );
  AND2X2 AND2X2_327 ( .A(_abc_4513_n506), .B(\Rdata_mem[29] ), .Y(_abc_4513_n871) );
  AND2X2 AND2X2_328 ( .A(_abc_4513_n498), .B(\Rdata_mem[13] ), .Y(_abc_4513_n872) );
  AND2X2 AND2X2_329 ( .A(_abc_4513_n874), .B(_abc_4513_n771), .Y(\rd[13] ) );
  AND2X2 AND2X2_33 ( .A(Rvalid), .B(state_5_), .Y(_abc_4513_n411_1) );
  AND2X2 AND2X2_330 ( .A(_abc_4513_n506), .B(\Rdata_mem[30] ), .Y(_abc_4513_n876) );
  AND2X2 AND2X2_331 ( .A(_abc_4513_n498), .B(\Rdata_mem[14] ), .Y(_abc_4513_n877) );
  AND2X2 AND2X2_332 ( .A(_abc_4513_n879_1), .B(_abc_4513_n771), .Y(\rd[14] ) );
  AND2X2 AND2X2_333 ( .A(_abc_4513_n498), .B(\Rdata_mem[15] ), .Y(_abc_4513_n881_1) );
  AND2X2 AND2X2_334 ( .A(_abc_4513_n506), .B(\Rdata_mem[31] ), .Y(_abc_4513_n882) );
  AND2X2 AND2X2_335 ( .A(_abc_4513_n884), .B(_abc_4513_n771), .Y(\rd[15] ) );
  AND2X2 AND2X2_336 ( .A(_abc_4513_n495_1), .B(\Rdata_mem[16] ), .Y(_abc_4513_n886_1) );
  AND2X2 AND2X2_337 ( .A(_abc_4513_n489), .B(\Rdata_mem[15] ), .Y(_abc_4513_n887_1) );
  AND2X2 AND2X2_338 ( .A(_abc_4513_n505), .B(\Rdata_mem[31] ), .Y(_abc_4513_n888_1) );
  AND2X2 AND2X2_339 ( .A(_abc_4513_n496), .B(signo), .Y(_abc_4513_n890) );
  AND2X2 AND2X2_34 ( .A(_abc_4513_n409), .B(state_2_), .Y(_abc_4513_n412) );
  AND2X2 AND2X2_340 ( .A(_abc_4513_n889), .B(_abc_4513_n890), .Y(_abc_4513_n891) );
  AND2X2 AND2X2_341 ( .A(_abc_4513_n893), .B(_abc_4513_n771), .Y(\rd[16] ) );
  AND2X2 AND2X2_342 ( .A(_abc_4513_n495_1), .B(\Rdata_mem[17] ), .Y(_abc_4513_n895) );
  AND2X2 AND2X2_343 ( .A(_abc_4513_n896_1), .B(_abc_4513_n771), .Y(\rd[17] ) );
  AND2X2 AND2X2_344 ( .A(_abc_4513_n495_1), .B(\Rdata_mem[18] ), .Y(_abc_4513_n898) );
  AND2X2 AND2X2_345 ( .A(_abc_4513_n899_1), .B(_abc_4513_n771), .Y(\rd[18] ) );
  AND2X2 AND2X2_346 ( .A(_abc_4513_n495_1), .B(\Rdata_mem[19] ), .Y(_abc_4513_n901) );
  AND2X2 AND2X2_347 ( .A(_abc_4513_n902_1), .B(_abc_4513_n771), .Y(\rd[19] ) );
  AND2X2 AND2X2_348 ( .A(_abc_4513_n495_1), .B(\Rdata_mem[20] ), .Y(_abc_4513_n904_1) );
  AND2X2 AND2X2_349 ( .A(_abc_4513_n905), .B(_abc_4513_n771), .Y(\rd[20] ) );
  AND2X2 AND2X2_35 ( .A(AWready), .B(Bvalid), .Y(_abc_4513_n414_1) );
  AND2X2 AND2X2_350 ( .A(_abc_4513_n495_1), .B(\Rdata_mem[21] ), .Y(_abc_4513_n907) );
  AND2X2 AND2X2_351 ( .A(_abc_4513_n908), .B(_abc_4513_n771), .Y(\rd[21] ) );
  AND2X2 AND2X2_352 ( .A(_abc_4513_n495_1), .B(\Rdata_mem[22] ), .Y(_abc_4513_n910) );
  AND2X2 AND2X2_353 ( .A(_abc_4513_n911), .B(_abc_4513_n771), .Y(\rd[22] ) );
  AND2X2 AND2X2_354 ( .A(_abc_4513_n495_1), .B(\Rdata_mem[23] ), .Y(_abc_4513_n913) );
  AND2X2 AND2X2_355 ( .A(_abc_4513_n914), .B(_abc_4513_n771), .Y(\rd[23] ) );
  AND2X2 AND2X2_356 ( .A(_abc_4513_n495_1), .B(\Rdata_mem[24] ), .Y(_abc_4513_n916) );
  AND2X2 AND2X2_357 ( .A(_abc_4513_n917), .B(_abc_4513_n771), .Y(\rd[24] ) );
  AND2X2 AND2X2_358 ( .A(_abc_4513_n495_1), .B(\Rdata_mem[25] ), .Y(_abc_4513_n919) );
  AND2X2 AND2X2_359 ( .A(_abc_4513_n920), .B(_abc_4513_n771), .Y(\rd[25] ) );
  AND2X2 AND2X2_36 ( .A(_abc_4513_n414_1), .B(state_6_), .Y(_abc_4513_n415) );
  AND2X2 AND2X2_360 ( .A(_abc_4513_n495_1), .B(\Rdata_mem[26] ), .Y(_abc_4513_n922) );
  AND2X2 AND2X2_361 ( .A(_abc_4513_n923), .B(_abc_4513_n771), .Y(\rd[26] ) );
  AND2X2 AND2X2_362 ( .A(_abc_4513_n495_1), .B(\Rdata_mem[27] ), .Y(_abc_4513_n925) );
  AND2X2 AND2X2_363 ( .A(_abc_4513_n926), .B(_abc_4513_n771), .Y(\rd[27] ) );
  AND2X2 AND2X2_364 ( .A(_abc_4513_n495_1), .B(\Rdata_mem[28] ), .Y(_abc_4513_n928) );
  AND2X2 AND2X2_365 ( .A(_abc_4513_n929), .B(_abc_4513_n771), .Y(\rd[28] ) );
  AND2X2 AND2X2_366 ( .A(_abc_4513_n495_1), .B(\Rdata_mem[29] ), .Y(_abc_4513_n931) );
  AND2X2 AND2X2_367 ( .A(_abc_4513_n932), .B(_abc_4513_n771), .Y(\rd[29] ) );
  AND2X2 AND2X2_368 ( .A(_abc_4513_n495_1), .B(\Rdata_mem[30] ), .Y(_abc_4513_n934) );
  AND2X2 AND2X2_369 ( .A(_abc_4513_n935), .B(_abc_4513_n771), .Y(\rd[30] ) );
  AND2X2 AND2X2_37 ( .A(Bvalid), .B(state_1_), .Y(_abc_4513_n417_1) );
  AND2X2 AND2X2_370 ( .A(_abc_4513_n495_1), .B(\Rdata_mem[31] ), .Y(_abc_4513_n937) );
  AND2X2 AND2X2_371 ( .A(_abc_4513_n938), .B(_abc_4513_n771), .Y(\rd[31] ) );
  AND2X2 AND2X2_372 ( .A(_abc_4513_n940), .B(_abc_4513_n941), .Y(\AWdata[0] ) );
  AND2X2 AND2X2_373 ( .A(_abc_4513_n943), .B(_abc_4513_n944), .Y(\AWdata[1] ) );
  AND2X2 AND2X2_374 ( .A(\imm[2] ), .B(\rs1[2] ), .Y(_abc_4513_n947) );
  AND2X2 AND2X2_375 ( .A(_abc_4513_n948), .B(_abc_4513_n949), .Y(_abc_4513_n950) );
  AND2X2 AND2X2_376 ( .A(_abc_4513_n946), .B(_abc_4513_n950), .Y(_abc_4513_n951) );
  AND2X2 AND2X2_377 ( .A(_abc_4513_n952), .B(_abc_4513_n953), .Y(_abc_4513_n954) );
  AND2X2 AND2X2_378 ( .A(_abc_4513_n955), .B(_abc_4513_n956), .Y(\AWdata[2] ) );
  AND2X2 AND2X2_379 ( .A(_abc_4513_n952), .B(_abc_4513_n948), .Y(_abc_4513_n958) );
  AND2X2 AND2X2_38 ( .A(_abc_4513_n419_1), .B(state_0_), .Y(_abc_4513_n420_1) );
  AND2X2 AND2X2_380 ( .A(\imm[3] ), .B(\rs1[3] ), .Y(_abc_4513_n961) );
  AND2X2 AND2X2_381 ( .A(_abc_4513_n962), .B(_abc_4513_n960), .Y(_abc_4513_n963) );
  AND2X2 AND2X2_382 ( .A(_abc_4513_n959), .B(_abc_4513_n964), .Y(_abc_4513_n965) );
  AND2X2 AND2X2_383 ( .A(_abc_4513_n958), .B(_abc_4513_n963), .Y(_abc_4513_n966) );
  AND2X2 AND2X2_384 ( .A(_abc_4513_n967), .B(_abc_4513_n769_1), .Y(_abc_4513_n968) );
  AND2X2 AND2X2_385 ( .A(\W_R[1] ), .B(\pc[3] ), .Y(_abc_4513_n969) );
  AND2X2 AND2X2_386 ( .A(_abc_4513_n950), .B(_abc_4513_n963), .Y(_abc_4513_n971) );
  AND2X2 AND2X2_387 ( .A(_abc_4513_n946), .B(_abc_4513_n971), .Y(_abc_4513_n972) );
  AND2X2 AND2X2_388 ( .A(_abc_4513_n960), .B(_abc_4513_n947), .Y(_abc_4513_n973) );
  AND2X2 AND2X2_389 ( .A(\imm[4] ), .B(\rs1[4] ), .Y(_abc_4513_n977) );
  AND2X2 AND2X2_39 ( .A(_abc_4513_n402_1), .B(_abc_4513_n428), .Y(_abc_4513_n429) );
  AND2X2 AND2X2_390 ( .A(_abc_4513_n978), .B(_abc_4513_n976), .Y(_abc_4513_n979) );
  AND2X2 AND2X2_391 ( .A(_abc_4513_n975), .B(_abc_4513_n979), .Y(_abc_4513_n980) );
  AND2X2 AND2X2_392 ( .A(_abc_4513_n981), .B(_abc_4513_n982), .Y(_abc_4513_n983) );
  AND2X2 AND2X2_393 ( .A(_abc_4513_n984), .B(_abc_4513_n985), .Y(\AWdata[4] ) );
  AND2X2 AND2X2_394 ( .A(_abc_4513_n981), .B(_abc_4513_n978), .Y(_abc_4513_n987) );
  AND2X2 AND2X2_395 ( .A(\imm[5] ), .B(\rs1[5] ), .Y(_abc_4513_n990) );
  AND2X2 AND2X2_396 ( .A(_abc_4513_n991), .B(_abc_4513_n989), .Y(_abc_4513_n992) );
  AND2X2 AND2X2_397 ( .A(_abc_4513_n993), .B(_abc_4513_n995), .Y(_abc_4513_n996) );
  AND2X2 AND2X2_398 ( .A(_abc_4513_n997), .B(_abc_4513_n998), .Y(\AWdata[5] ) );
  AND2X2 AND2X2_399 ( .A(\W_R[1] ), .B(\pc[6] ), .Y(_abc_4513_n1000) );
  AND2X2 AND2X2_4 ( .A(ARvalid), .B(_abc_4513_n361), .Y(_abc_3815_n14) );
  AND2X2 AND2X2_40 ( .A(_abc_4513_n394), .B(_abc_4513_n397), .Y(_abc_4513_n430) );
  AND2X2 AND2X2_400 ( .A(_abc_4513_n1001), .B(_abc_4513_n989), .Y(_abc_4513_n1002) );
  AND2X2 AND2X2_401 ( .A(_abc_4513_n979), .B(_abc_4513_n992), .Y(_abc_4513_n1003) );
  AND2X2 AND2X2_402 ( .A(_abc_4513_n975), .B(_abc_4513_n1003), .Y(_abc_4513_n1004) );
  AND2X2 AND2X2_403 ( .A(\imm[6] ), .B(\rs1[6] ), .Y(_abc_4513_n1006) );
  AND2X2 AND2X2_404 ( .A(_abc_4513_n1007), .B(_abc_4513_n1008), .Y(_abc_4513_n1009) );
  AND2X2 AND2X2_405 ( .A(_abc_4513_n1005), .B(_abc_4513_n1009), .Y(_abc_4513_n1011) );
  AND2X2 AND2X2_406 ( .A(_abc_4513_n1012), .B(_abc_4513_n1010), .Y(_abc_4513_n1013) );
  AND2X2 AND2X2_407 ( .A(_abc_4513_n1013), .B(_abc_4513_n769_1), .Y(_abc_4513_n1014) );
  AND2X2 AND2X2_408 ( .A(_abc_4513_n1012), .B(_abc_4513_n1007), .Y(_abc_4513_n1017) );
  AND2X2 AND2X2_409 ( .A(\imm[7] ), .B(\rs1[7] ), .Y(_abc_4513_n1019) );
  AND2X2 AND2X2_41 ( .A(_abc_4513_n382), .B(_abc_4513_n431), .Y(_abc_4513_n432) );
  AND2X2 AND2X2_410 ( .A(_abc_4513_n1020), .B(_abc_4513_n1018), .Y(_abc_4513_n1021) );
  AND2X2 AND2X2_411 ( .A(_abc_4513_n1025), .B(_abc_4513_n1023), .Y(_abc_4513_n1026) );
  AND2X2 AND2X2_412 ( .A(_abc_4513_n1027), .B(_abc_4513_n1016), .Y(\AWdata[7] ) );
  AND2X2 AND2X2_413 ( .A(\W_R[1] ), .B(\pc[8] ), .Y(_abc_4513_n1029) );
  AND2X2 AND2X2_414 ( .A(_abc_4513_n1009), .B(_abc_4513_n1021), .Y(_abc_4513_n1030) );
  AND2X2 AND2X2_415 ( .A(_abc_4513_n1003), .B(_abc_4513_n1030), .Y(_abc_4513_n1031) );
  AND2X2 AND2X2_416 ( .A(_abc_4513_n975), .B(_abc_4513_n1031), .Y(_abc_4513_n1032) );
  AND2X2 AND2X2_417 ( .A(_abc_4513_n1030), .B(_abc_4513_n1002), .Y(_abc_4513_n1033) );
  AND2X2 AND2X2_418 ( .A(_abc_4513_n1018), .B(_abc_4513_n1006), .Y(_abc_4513_n1034) );
  AND2X2 AND2X2_419 ( .A(\imm[8] ), .B(\rs1[8] ), .Y(_abc_4513_n1038) );
  AND2X2 AND2X2_42 ( .A(_abc_4513_n433), .B(_abc_4513_n398_1), .Y(_abc_4513_n434) );
  AND2X2 AND2X2_420 ( .A(_abc_4513_n1039), .B(_abc_4513_n1040), .Y(_abc_4513_n1041) );
  AND2X2 AND2X2_421 ( .A(_abc_4513_n1037), .B(_abc_4513_n1041), .Y(_abc_4513_n1043) );
  AND2X2 AND2X2_422 ( .A(_abc_4513_n1044), .B(_abc_4513_n1042), .Y(_abc_4513_n1045) );
  AND2X2 AND2X2_423 ( .A(_abc_4513_n1045), .B(_abc_4513_n769_1), .Y(_abc_4513_n1046) );
  AND2X2 AND2X2_424 ( .A(_abc_4513_n1044), .B(_abc_4513_n1039), .Y(_abc_4513_n1048) );
  AND2X2 AND2X2_425 ( .A(\imm[9] ), .B(\rs1[9] ), .Y(_abc_4513_n1051) );
  AND2X2 AND2X2_426 ( .A(_abc_4513_n1052), .B(_abc_4513_n1050), .Y(_abc_4513_n1053) );
  AND2X2 AND2X2_427 ( .A(_abc_4513_n1054), .B(_abc_4513_n1056), .Y(_abc_4513_n1057) );
  AND2X2 AND2X2_428 ( .A(_abc_4513_n1058), .B(_abc_4513_n1059), .Y(\AWdata[9] ) );
  AND2X2 AND2X2_429 ( .A(\W_R[1] ), .B(\pc[10] ), .Y(_abc_4513_n1061) );
  AND2X2 AND2X2_43 ( .A(_abc_4513_n393_1), .B(AWready), .Y(_abc_4513_n436) );
  AND2X2 AND2X2_430 ( .A(_abc_4513_n1062), .B(_abc_4513_n1050), .Y(_abc_4513_n1063) );
  AND2X2 AND2X2_431 ( .A(_abc_4513_n1041), .B(_abc_4513_n1053), .Y(_abc_4513_n1064) );
  AND2X2 AND2X2_432 ( .A(_abc_4513_n1037), .B(_abc_4513_n1064), .Y(_abc_4513_n1065) );
  AND2X2 AND2X2_433 ( .A(\imm[10] ), .B(\rs1[10] ), .Y(_abc_4513_n1067) );
  AND2X2 AND2X2_434 ( .A(_abc_4513_n1068), .B(_abc_4513_n1069), .Y(_abc_4513_n1070) );
  AND2X2 AND2X2_435 ( .A(_abc_4513_n1066), .B(_abc_4513_n1070), .Y(_abc_4513_n1072) );
  AND2X2 AND2X2_436 ( .A(_abc_4513_n1073), .B(_abc_4513_n1071), .Y(_abc_4513_n1074) );
  AND2X2 AND2X2_437 ( .A(_abc_4513_n1074), .B(_abc_4513_n769_1), .Y(_abc_4513_n1075) );
  AND2X2 AND2X2_438 ( .A(_abc_4513_n1073), .B(_abc_4513_n1068), .Y(_abc_4513_n1077) );
  AND2X2 AND2X2_439 ( .A(\imm[11] ), .B(\rs1[11] ), .Y(_abc_4513_n1079) );
  AND2X2 AND2X2_44 ( .A(_abc_4513_n437), .B(state_4_), .Y(_abc_4513_n438_1) );
  AND2X2 AND2X2_440 ( .A(_abc_4513_n1080), .B(_abc_4513_n1078), .Y(_abc_4513_n1081) );
  AND2X2 AND2X2_441 ( .A(_abc_4513_n1085), .B(_abc_4513_n1083), .Y(_abc_4513_n1086) );
  AND2X2 AND2X2_442 ( .A(_abc_4513_n1087), .B(_abc_4513_n1088), .Y(\AWdata[11] ) );
  AND2X2 AND2X2_443 ( .A(\W_R[1] ), .B(\pc[12] ), .Y(_abc_4513_n1090) );
  AND2X2 AND2X2_444 ( .A(_abc_4513_n1070), .B(_abc_4513_n1081), .Y(_abc_4513_n1091) );
  AND2X2 AND2X2_445 ( .A(_abc_4513_n1091), .B(_abc_4513_n1063), .Y(_abc_4513_n1092) );
  AND2X2 AND2X2_446 ( .A(_abc_4513_n1078), .B(_abc_4513_n1067), .Y(_abc_4513_n1093) );
  AND2X2 AND2X2_447 ( .A(_abc_4513_n1064), .B(_abc_4513_n1091), .Y(_abc_4513_n1096) );
  AND2X2 AND2X2_448 ( .A(_abc_4513_n1037), .B(_abc_4513_n1096), .Y(_abc_4513_n1097) );
  AND2X2 AND2X2_449 ( .A(\imm[12] ), .B(\rs1[12] ), .Y(_abc_4513_n1100) );
  AND2X2 AND2X2_45 ( .A(_abc_4513_n403), .B(_abc_4513_n438_1), .Y(_abc_4513_n439) );
  AND2X2 AND2X2_450 ( .A(_abc_4513_n1101), .B(_abc_4513_n1099), .Y(_abc_4513_n1102) );
  AND2X2 AND2X2_451 ( .A(_abc_4513_n1098), .B(_abc_4513_n1102), .Y(_abc_4513_n1104) );
  AND2X2 AND2X2_452 ( .A(_abc_4513_n1105), .B(_abc_4513_n1103), .Y(_abc_4513_n1106) );
  AND2X2 AND2X2_453 ( .A(_abc_4513_n1106), .B(_abc_4513_n769_1), .Y(_abc_4513_n1107) );
  AND2X2 AND2X2_454 ( .A(_abc_4513_n1105), .B(_abc_4513_n1101), .Y(_abc_4513_n1109) );
  AND2X2 AND2X2_455 ( .A(\imm[13] ), .B(\rs1[13] ), .Y(_abc_4513_n1112) );
  AND2X2 AND2X2_456 ( .A(_abc_4513_n1113), .B(_abc_4513_n1111), .Y(_abc_4513_n1114) );
  AND2X2 AND2X2_457 ( .A(_abc_4513_n1115), .B(_abc_4513_n1117), .Y(_abc_4513_n1118) );
  AND2X2 AND2X2_458 ( .A(_abc_4513_n1119), .B(_abc_4513_n1120), .Y(\AWdata[13] ) );
  AND2X2 AND2X2_459 ( .A(\W_R[1] ), .B(\pc[14] ), .Y(_abc_4513_n1122) );
  AND2X2 AND2X2_46 ( .A(_abc_4513_n382), .B(_abc_4513_n430), .Y(_abc_4513_n440) );
  AND2X2 AND2X2_460 ( .A(_abc_4513_n1123), .B(_abc_4513_n1113), .Y(_abc_4513_n1124) );
  AND2X2 AND2X2_461 ( .A(_abc_4513_n1102), .B(_abc_4513_n1114), .Y(_abc_4513_n1126) );
  AND2X2 AND2X2_462 ( .A(_abc_4513_n1098), .B(_abc_4513_n1126), .Y(_abc_4513_n1127) );
  AND2X2 AND2X2_463 ( .A(\imm[14] ), .B(\rs1[14] ), .Y(_abc_4513_n1129) );
  AND2X2 AND2X2_464 ( .A(_abc_4513_n1130), .B(_abc_4513_n1131), .Y(_abc_4513_n1132) );
  AND2X2 AND2X2_465 ( .A(_abc_4513_n1128), .B(_abc_4513_n1132), .Y(_abc_4513_n1134) );
  AND2X2 AND2X2_466 ( .A(_abc_4513_n1135), .B(_abc_4513_n1133), .Y(_abc_4513_n1136) );
  AND2X2 AND2X2_467 ( .A(_abc_4513_n1136), .B(_abc_4513_n769_1), .Y(_abc_4513_n1137) );
  AND2X2 AND2X2_468 ( .A(_abc_4513_n1135), .B(_abc_4513_n1130), .Y(_abc_4513_n1140) );
  AND2X2 AND2X2_469 ( .A(\imm[15] ), .B(\rs1[15] ), .Y(_abc_4513_n1142) );
  AND2X2 AND2X2_47 ( .A(resetn), .B(state_6_), .Y(_abc_4513_n442) );
  AND2X2 AND2X2_470 ( .A(_abc_4513_n1143), .B(_abc_4513_n1141), .Y(_abc_4513_n1144) );
  AND2X2 AND2X2_471 ( .A(_abc_4513_n1148), .B(_abc_4513_n1146), .Y(_abc_4513_n1149) );
  AND2X2 AND2X2_472 ( .A(_abc_4513_n1150), .B(_abc_4513_n1139), .Y(\AWdata[15] ) );
  AND2X2 AND2X2_473 ( .A(\W_R[1] ), .B(\pc[16] ), .Y(_abc_4513_n1152) );
  AND2X2 AND2X2_474 ( .A(_abc_4513_n1132), .B(_abc_4513_n1144), .Y(_abc_4513_n1153) );
  AND2X2 AND2X2_475 ( .A(_abc_4513_n1126), .B(_abc_4513_n1153), .Y(_abc_4513_n1154) );
  AND2X2 AND2X2_476 ( .A(_abc_4513_n1096), .B(_abc_4513_n1154), .Y(_abc_4513_n1155) );
  AND2X2 AND2X2_477 ( .A(_abc_4513_n1037), .B(_abc_4513_n1155), .Y(_abc_4513_n1156) );
  AND2X2 AND2X2_478 ( .A(_abc_4513_n1095), .B(_abc_4513_n1154), .Y(_abc_4513_n1157) );
  AND2X2 AND2X2_479 ( .A(_abc_4513_n1125), .B(_abc_4513_n1153), .Y(_abc_4513_n1158) );
  AND2X2 AND2X2_48 ( .A(_abc_4513_n442), .B(_abc_4513_n394), .Y(_abc_4513_n443) );
  AND2X2 AND2X2_480 ( .A(_abc_4513_n1141), .B(_abc_4513_n1129), .Y(_abc_4513_n1159) );
  AND2X2 AND2X2_481 ( .A(\imm[16] ), .B(\rs1[16] ), .Y(_abc_4513_n1164) );
  AND2X2 AND2X2_482 ( .A(_abc_4513_n1165), .B(_abc_4513_n1166), .Y(_abc_4513_n1167) );
  AND2X2 AND2X2_483 ( .A(_abc_4513_n1163), .B(_abc_4513_n1167), .Y(_abc_4513_n1169) );
  AND2X2 AND2X2_484 ( .A(_abc_4513_n1170), .B(_abc_4513_n1168), .Y(_abc_4513_n1171) );
  AND2X2 AND2X2_485 ( .A(_abc_4513_n1171), .B(_abc_4513_n769_1), .Y(_abc_4513_n1172) );
  AND2X2 AND2X2_486 ( .A(_abc_4513_n1170), .B(_abc_4513_n1165), .Y(_abc_4513_n1174) );
  AND2X2 AND2X2_487 ( .A(\imm[17] ), .B(\rs1[17] ), .Y(_abc_4513_n1176) );
  AND2X2 AND2X2_488 ( .A(_abc_4513_n1177), .B(_abc_4513_n1178), .Y(_abc_4513_n1179) );
  AND2X2 AND2X2_489 ( .A(_abc_4513_n1180), .B(_abc_4513_n1182), .Y(_abc_4513_n1183) );
  AND2X2 AND2X2_49 ( .A(_abc_4513_n433), .B(_abc_4513_n395_1), .Y(_abc_4513_n444) );
  AND2X2 AND2X2_490 ( .A(_abc_4513_n1184), .B(_abc_4513_n1185), .Y(\AWdata[17] ) );
  AND2X2 AND2X2_491 ( .A(\W_R[1] ), .B(\pc[18] ), .Y(_abc_4513_n1187) );
  AND2X2 AND2X2_492 ( .A(_abc_4513_n1188), .B(_abc_4513_n1177), .Y(_abc_4513_n1189) );
  AND2X2 AND2X2_493 ( .A(_abc_4513_n1167), .B(_abc_4513_n1179), .Y(_abc_4513_n1191) );
  AND2X2 AND2X2_494 ( .A(_abc_4513_n1163), .B(_abc_4513_n1191), .Y(_abc_4513_n1192) );
  AND2X2 AND2X2_495 ( .A(\imm[18] ), .B(\rs1[18] ), .Y(_abc_4513_n1194) );
  AND2X2 AND2X2_496 ( .A(_abc_4513_n1195), .B(_abc_4513_n1196), .Y(_abc_4513_n1197) );
  AND2X2 AND2X2_497 ( .A(_abc_4513_n1193), .B(_abc_4513_n1197), .Y(_abc_4513_n1199) );
  AND2X2 AND2X2_498 ( .A(_abc_4513_n1200), .B(_abc_4513_n1198), .Y(_abc_4513_n1201) );
  AND2X2 AND2X2_499 ( .A(_abc_4513_n1201), .B(_abc_4513_n769_1), .Y(_abc_4513_n1202) );
  AND2X2 AND2X2_5 ( .A(_abc_4513_n368), .B(AWready), .Y(_abc_4513_n369) );
  AND2X2 AND2X2_50 ( .A(_abc_4513_n365), .B(_abc_4513_n446_1), .Y(_abc_4513_n447) );
  AND2X2 AND2X2_500 ( .A(_abc_4513_n1200), .B(_abc_4513_n1195), .Y(_abc_4513_n1205) );
  AND2X2 AND2X2_501 ( .A(\imm[19] ), .B(\rs1[19] ), .Y(_abc_4513_n1206) );
  AND2X2 AND2X2_502 ( .A(_abc_4513_n1207), .B(_abc_4513_n1208), .Y(_abc_4513_n1209) );
  AND2X2 AND2X2_503 ( .A(_abc_4513_n1213), .B(_abc_4513_n1211), .Y(_abc_4513_n1214) );
  AND2X2 AND2X2_504 ( .A(_abc_4513_n1215), .B(_abc_4513_n1204), .Y(\AWdata[19] ) );
  AND2X2 AND2X2_505 ( .A(\W_R[1] ), .B(\pc[20] ), .Y(_abc_4513_n1217) );
  AND2X2 AND2X2_506 ( .A(_abc_4513_n1197), .B(_abc_4513_n1209), .Y(_abc_4513_n1218) );
  AND2X2 AND2X2_507 ( .A(_abc_4513_n1190), .B(_abc_4513_n1218), .Y(_abc_4513_n1219) );
  AND2X2 AND2X2_508 ( .A(_abc_4513_n1208), .B(_abc_4513_n1194), .Y(_abc_4513_n1220) );
  AND2X2 AND2X2_509 ( .A(_abc_4513_n1191), .B(_abc_4513_n1218), .Y(_abc_4513_n1223) );
  AND2X2 AND2X2_51 ( .A(_abc_4513_n449), .B(_abc_4513_n437), .Y(_abc_4513_n450) );
  AND2X2 AND2X2_510 ( .A(_abc_4513_n1163), .B(_abc_4513_n1223), .Y(_abc_4513_n1224) );
  AND2X2 AND2X2_511 ( .A(\imm[20] ), .B(\rs1[20] ), .Y(_abc_4513_n1226) );
  AND2X2 AND2X2_512 ( .A(_abc_4513_n1227), .B(_abc_4513_n1228), .Y(_abc_4513_n1229) );
  AND2X2 AND2X2_513 ( .A(_abc_4513_n1233), .B(_abc_4513_n1230), .Y(_abc_4513_n1234) );
  AND2X2 AND2X2_514 ( .A(_abc_4513_n1234), .B(_abc_4513_n769_1), .Y(_abc_4513_n1235) );
  AND2X2 AND2X2_515 ( .A(_abc_4513_n1233), .B(_abc_4513_n1227), .Y(_abc_4513_n1237) );
  AND2X2 AND2X2_516 ( .A(\imm[21] ), .B(\rs1[21] ), .Y(_abc_4513_n1238) );
  AND2X2 AND2X2_517 ( .A(_abc_4513_n1239), .B(_abc_4513_n1240), .Y(_abc_4513_n1241) );
  AND2X2 AND2X2_518 ( .A(_abc_4513_n1245), .B(_abc_4513_n1243), .Y(_abc_4513_n1246) );
  AND2X2 AND2X2_519 ( .A(_abc_4513_n1247), .B(_abc_4513_n1248), .Y(\AWdata[21] ) );
  AND2X2 AND2X2_52 ( .A(_abc_4513_n456), .B(_abc_4513_n453), .Y(_abc_4513_n457) );
  AND2X2 AND2X2_520 ( .A(\W_R[1] ), .B(\pc[22] ), .Y(_abc_4513_n1250) );
  AND2X2 AND2X2_521 ( .A(_abc_4513_n1251), .B(_abc_4513_n1239), .Y(_abc_4513_n1252) );
  AND2X2 AND2X2_522 ( .A(_abc_4513_n1229), .B(_abc_4513_n1241), .Y(_abc_4513_n1254) );
  AND2X2 AND2X2_523 ( .A(_abc_4513_n1225), .B(_abc_4513_n1254), .Y(_abc_4513_n1255) );
  AND2X2 AND2X2_524 ( .A(\imm[22] ), .B(\rs1[22] ), .Y(_abc_4513_n1257) );
  AND2X2 AND2X2_525 ( .A(_abc_4513_n1258), .B(_abc_4513_n1259), .Y(_abc_4513_n1260) );
  AND2X2 AND2X2_526 ( .A(_abc_4513_n1256), .B(_abc_4513_n1260), .Y(_abc_4513_n1262) );
  AND2X2 AND2X2_527 ( .A(_abc_4513_n1263), .B(_abc_4513_n1261), .Y(_abc_4513_n1264) );
  AND2X2 AND2X2_528 ( .A(_abc_4513_n1264), .B(_abc_4513_n769_1), .Y(_abc_4513_n1265) );
  AND2X2 AND2X2_529 ( .A(_abc_4513_n1263), .B(_abc_4513_n1258), .Y(_abc_4513_n1268) );
  AND2X2 AND2X2_53 ( .A(_abc_4513_n457), .B(_abc_4513_n451), .Y(_abc_4513_n458) );
  AND2X2 AND2X2_530 ( .A(\imm[23] ), .B(\rs1[23] ), .Y(_abc_4513_n1269) );
  AND2X2 AND2X2_531 ( .A(_abc_4513_n1270), .B(_abc_4513_n1271), .Y(_abc_4513_n1272) );
  AND2X2 AND2X2_532 ( .A(_abc_4513_n1276), .B(_abc_4513_n1274), .Y(_abc_4513_n1277) );
  AND2X2 AND2X2_533 ( .A(_abc_4513_n1278), .B(_abc_4513_n1267), .Y(\AWdata[23] ) );
  AND2X2 AND2X2_534 ( .A(\W_R[1] ), .B(\pc[24] ), .Y(_abc_4513_n1280) );
  AND2X2 AND2X2_535 ( .A(_abc_4513_n1260), .B(_abc_4513_n1272), .Y(_abc_4513_n1281) );
  AND2X2 AND2X2_536 ( .A(_abc_4513_n1254), .B(_abc_4513_n1281), .Y(_abc_4513_n1282) );
  AND2X2 AND2X2_537 ( .A(_abc_4513_n1223), .B(_abc_4513_n1282), .Y(_abc_4513_n1283) );
  AND2X2 AND2X2_538 ( .A(_abc_4513_n1163), .B(_abc_4513_n1283), .Y(_abc_4513_n1284) );
  AND2X2 AND2X2_539 ( .A(_abc_4513_n1222), .B(_abc_4513_n1282), .Y(_abc_4513_n1285) );
  AND2X2 AND2X2_54 ( .A(_abc_4513_n458), .B(_abc_4513_n448), .Y(_abc_4513_n459) );
  AND2X2 AND2X2_540 ( .A(_abc_4513_n1253), .B(_abc_4513_n1281), .Y(_abc_4513_n1286) );
  AND2X2 AND2X2_541 ( .A(_abc_4513_n1271), .B(_abc_4513_n1257), .Y(_abc_4513_n1287) );
  AND2X2 AND2X2_542 ( .A(\imm[24] ), .B(\rs1[24] ), .Y(_abc_4513_n1292) );
  AND2X2 AND2X2_543 ( .A(_abc_4513_n1293), .B(_abc_4513_n1294), .Y(_abc_4513_n1295) );
  AND2X2 AND2X2_544 ( .A(_abc_4513_n1291), .B(_abc_4513_n1295), .Y(_abc_4513_n1297) );
  AND2X2 AND2X2_545 ( .A(_abc_4513_n1298), .B(_abc_4513_n1296), .Y(_abc_4513_n1299) );
  AND2X2 AND2X2_546 ( .A(_abc_4513_n1299), .B(_abc_4513_n769_1), .Y(_abc_4513_n1300) );
  AND2X2 AND2X2_547 ( .A(_abc_4513_n1298), .B(_abc_4513_n1293), .Y(_abc_4513_n1302) );
  AND2X2 AND2X2_548 ( .A(\imm[25] ), .B(\rs1[25] ), .Y(_abc_4513_n1304) );
  AND2X2 AND2X2_549 ( .A(_abc_4513_n1305), .B(_abc_4513_n1306), .Y(_abc_4513_n1307) );
  AND2X2 AND2X2_55 ( .A(_abc_4513_n466), .B(resetn), .Y(_abc_4513_n467) );
  AND2X2 AND2X2_550 ( .A(_abc_4513_n1308), .B(_abc_4513_n1310), .Y(_abc_4513_n1311) );
  AND2X2 AND2X2_551 ( .A(_abc_4513_n1312), .B(_abc_4513_n1313), .Y(\AWdata[25] ) );
  AND2X2 AND2X2_552 ( .A(\W_R[1] ), .B(\pc[26] ), .Y(_abc_4513_n1315) );
  AND2X2 AND2X2_553 ( .A(_abc_4513_n1316), .B(_abc_4513_n1305), .Y(_abc_4513_n1317) );
  AND2X2 AND2X2_554 ( .A(_abc_4513_n1295), .B(_abc_4513_n1307), .Y(_abc_4513_n1319) );
  AND2X2 AND2X2_555 ( .A(_abc_4513_n1291), .B(_abc_4513_n1319), .Y(_abc_4513_n1320) );
  AND2X2 AND2X2_556 ( .A(\imm[26] ), .B(\rs1[26] ), .Y(_abc_4513_n1322) );
  AND2X2 AND2X2_557 ( .A(_abc_4513_n1323), .B(_abc_4513_n1324), .Y(_abc_4513_n1325) );
  AND2X2 AND2X2_558 ( .A(_abc_4513_n1321), .B(_abc_4513_n1325), .Y(_abc_4513_n1327) );
  AND2X2 AND2X2_559 ( .A(_abc_4513_n1328), .B(_abc_4513_n1326), .Y(_abc_4513_n1329) );
  AND2X2 AND2X2_56 ( .A(_abc_4513_n460), .B(_abc_4513_n467), .Y(busy) );
  AND2X2 AND2X2_560 ( .A(_abc_4513_n1329), .B(_abc_4513_n769_1), .Y(_abc_4513_n1330) );
  AND2X2 AND2X2_561 ( .A(_abc_4513_n1328), .B(_abc_4513_n1323), .Y(_abc_4513_n1333) );
  AND2X2 AND2X2_562 ( .A(\imm[27] ), .B(\rs1[27] ), .Y(_abc_4513_n1335) );
  AND2X2 AND2X2_563 ( .A(_abc_4513_n1336), .B(_abc_4513_n1334), .Y(_abc_4513_n1337) );
  AND2X2 AND2X2_564 ( .A(_abc_4513_n1341), .B(_abc_4513_n1339), .Y(_abc_4513_n1342) );
  AND2X2 AND2X2_565 ( .A(_abc_4513_n1343), .B(_abc_4513_n1332), .Y(\AWdata[27] ) );
  AND2X2 AND2X2_566 ( .A(\W_R[1] ), .B(\pc[28] ), .Y(_abc_4513_n1345) );
  AND2X2 AND2X2_567 ( .A(_abc_4513_n1325), .B(_abc_4513_n1337), .Y(_abc_4513_n1346) );
  AND2X2 AND2X2_568 ( .A(_abc_4513_n1319), .B(_abc_4513_n1346), .Y(_abc_4513_n1347) );
  AND2X2 AND2X2_569 ( .A(_abc_4513_n1291), .B(_abc_4513_n1347), .Y(_abc_4513_n1348) );
  AND2X2 AND2X2_57 ( .A(\wordsize[0] ), .B(\wordsize[1] ), .Y(_abc_4513_n470_1) );
  AND2X2 AND2X2_570 ( .A(_abc_4513_n1318), .B(_abc_4513_n1346), .Y(_abc_4513_n1349) );
  AND2X2 AND2X2_571 ( .A(_abc_4513_n1334), .B(_abc_4513_n1322), .Y(_abc_4513_n1350) );
  AND2X2 AND2X2_572 ( .A(\imm[28] ), .B(\rs1[28] ), .Y(_abc_4513_n1355) );
  AND2X2 AND2X2_573 ( .A(_abc_4513_n1356), .B(_abc_4513_n1354), .Y(_abc_4513_n1357) );
  AND2X2 AND2X2_574 ( .A(_abc_4513_n1353), .B(_abc_4513_n1357), .Y(_abc_4513_n1359) );
  AND2X2 AND2X2_575 ( .A(_abc_4513_n1360), .B(_abc_4513_n1358), .Y(_abc_4513_n1361) );
  AND2X2 AND2X2_576 ( .A(_abc_4513_n1361), .B(_abc_4513_n769_1), .Y(_abc_4513_n1362) );
  AND2X2 AND2X2_577 ( .A(_abc_4513_n1360), .B(_abc_4513_n1356), .Y(_abc_4513_n1364) );
  AND2X2 AND2X2_578 ( .A(\imm[29] ), .B(\rs1[29] ), .Y(_abc_4513_n1367) );
  AND2X2 AND2X2_579 ( .A(_abc_4513_n1368), .B(_abc_4513_n1366), .Y(_abc_4513_n1369) );
  AND2X2 AND2X2_58 ( .A(_abc_4513_n471), .B(resetn), .Y(_abc_4513_n472) );
  AND2X2 AND2X2_580 ( .A(_abc_4513_n1370), .B(_abc_4513_n1372), .Y(_abc_4513_n1373) );
  AND2X2 AND2X2_581 ( .A(_abc_4513_n1374), .B(_abc_4513_n1375), .Y(\AWdata[29] ) );
  AND2X2 AND2X2_582 ( .A(\W_R[1] ), .B(\pc[30] ), .Y(_abc_4513_n1377) );
  AND2X2 AND2X2_583 ( .A(_abc_4513_n1357), .B(_abc_4513_n1369), .Y(_abc_4513_n1378) );
  AND2X2 AND2X2_584 ( .A(_abc_4513_n1353), .B(_abc_4513_n1378), .Y(_abc_4513_n1379) );
  AND2X2 AND2X2_585 ( .A(_abc_4513_n1366), .B(_abc_4513_n1355), .Y(_abc_4513_n1380) );
  AND2X2 AND2X2_586 ( .A(\imm[30] ), .B(\rs1[30] ), .Y(_abc_4513_n1384) );
  AND2X2 AND2X2_587 ( .A(_abc_4513_n1385), .B(_abc_4513_n1383), .Y(_abc_4513_n1386) );
  AND2X2 AND2X2_588 ( .A(_abc_4513_n1388), .B(_abc_4513_n480), .Y(_abc_4513_n1389) );
  AND2X2 AND2X2_589 ( .A(_abc_4513_n1391), .B(_abc_4513_n1392), .Y(_abc_4513_n1393) );
  AND2X2 AND2X2_59 ( .A(_abc_4513_n472), .B(_abc_4513_n379), .Y(_abc_4513_n473) );
  AND2X2 AND2X2_590 ( .A(_abc_4513_n1395), .B(_abc_4513_n1396), .Y(_abc_4513_n1397) );
  AND2X2 AND2X2_591 ( .A(_abc_4513_n1399), .B(_abc_4513_n1400), .Y(_abc_4513_n1401) );
  AND2X2 AND2X2_592 ( .A(_abc_4513_n1403), .B(_abc_4513_n1404), .Y(_abc_4513_n1405) );
  AND2X2 AND2X2_593 ( .A(_abc_4513_n1407), .B(_abc_4513_n1408), .Y(_abc_4513_n1409) );
  AND2X2 AND2X2_594 ( .A(_abc_4513_n1411), .B(_abc_4513_n1412), .Y(_abc_4513_n1413) );
  AND2X2 AND2X2_595 ( .A(_abc_4513_n1415), .B(_abc_4513_n1387), .Y(_abc_4513_n1416) );
  AND2X2 AND2X2_596 ( .A(_abc_4513_n1416), .B(_abc_4513_n769_1), .Y(_abc_4513_n1417) );
  AND2X2 AND2X2_597 ( .A(_abc_4513_n1382), .B(_abc_4513_n1386), .Y(_abc_4513_n1419) );
  AND2X2 AND2X2_598 ( .A(_abc_4513_n1422), .B(_abc_4513_n1424), .Y(_abc_4513_n1425) );
  AND2X2 AND2X2_599 ( .A(_abc_4513_n1415), .B(_abc_4513_n1385), .Y(_abc_4513_n1428) );
  AND2X2 AND2X2_6 ( .A(_abc_4513_n369), .B(state_6_), .Y(_abc_4513_n370_1) );
  AND2X2 AND2X2_60 ( .A(_abc_4513_n474), .B(_abc_4513_n475), .Y(_abc_4513_n476) );
  AND2X2 AND2X2_600 ( .A(_abc_4513_n1429), .B(_abc_4513_n1427), .Y(_abc_4513_n1430) );
  AND2X2 AND2X2_601 ( .A(_abc_4513_n1431), .B(_abc_4513_n1432), .Y(\AWdata[31] ) );
  AND2X2 AND2X2_602 ( .A(_abc_4513_n518), .B(_abc_4513_n770), .Y(rd_en) );
  AND2X2 AND2X2_603 ( .A(_abc_4513_n1435), .B(resetn), .Y(Bready) );
  AND2X2 AND2X2_604 ( .A(_abc_4513_n1437), .B(resetn), .Y(Wvalid) );
  AND2X2 AND2X2_605 ( .A(_abc_4513_n1439), .B(resetn), .Y(AWvalid) );
  AND2X2 AND2X2_606 ( .A(_abc_4513_n1441), .B(_abc_4513_n516_1), .Y(RReady) );
  AND2X2 AND2X2_61 ( .A(\imm[0] ), .B(\rs1[0] ), .Y(_abc_4513_n477) );
  AND2X2 AND2X2_62 ( .A(\imm[1] ), .B(\rs1[1] ), .Y(_abc_4513_n479) );
  AND2X2 AND2X2_63 ( .A(_abc_4513_n480), .B(_abc_4513_n478_1), .Y(_abc_4513_n481) );
  AND2X2 AND2X2_64 ( .A(_abc_4513_n481), .B(_abc_4513_n477), .Y(_abc_4513_n482) );
  AND2X2 AND2X2_65 ( .A(_abc_4513_n484), .B(_abc_4513_n485), .Y(_abc_4513_n486_1) );
  AND2X2 AND2X2_66 ( .A(_abc_4513_n487), .B(_abc_4513_n483), .Y(_abc_4513_n488) );
  AND2X2 AND2X2_67 ( .A(_abc_4513_n483), .B(_abc_4513_n490), .Y(_abc_4513_n491) );
  AND2X2 AND2X2_68 ( .A(_abc_4513_n489), .B(_abc_4513_n492), .Y(_abc_4513_n493) );
  AND2X2 AND2X2_69 ( .A(_abc_4513_n493), .B(_abc_4513_n476), .Y(_abc_4513_n494_1) );
  AND2X2 AND2X2_7 ( .A(_abc_4513_n368), .B(state_1_), .Y(_abc_4513_n371_1) );
  AND2X2 AND2X2_70 ( .A(_abc_4513_n474), .B(\wordsize[1] ), .Y(_abc_4513_n495_1) );
  AND2X2 AND2X2_71 ( .A(_abc_4513_n475), .B(\wordsize[0] ), .Y(_abc_4513_n496) );
  AND2X2 AND2X2_72 ( .A(_abc_4513_n489), .B(_abc_4513_n496), .Y(_abc_4513_n497) );
  AND2X2 AND2X2_73 ( .A(_abc_4513_n499), .B(_abc_4513_n473), .Y(Wstrb_0__FF_INPUT) );
  AND2X2 AND2X2_74 ( .A(_abc_4513_n489), .B(_abc_4513_n491), .Y(_abc_4513_n501) );
  AND2X2 AND2X2_75 ( .A(_abc_4513_n501), .B(_abc_4513_n476), .Y(_abc_4513_n502) );
  AND2X2 AND2X2_76 ( .A(_abc_4513_n503), .B(_abc_4513_n473), .Y(Wstrb_1__FF_INPUT) );
  AND2X2 AND2X2_77 ( .A(_abc_4513_n505), .B(_abc_4513_n496), .Y(_abc_4513_n506) );
  AND2X2 AND2X2_78 ( .A(_abc_4513_n505), .B(_abc_4513_n492), .Y(_abc_4513_n508) );
  AND2X2 AND2X2_79 ( .A(_abc_4513_n508), .B(_abc_4513_n476), .Y(_abc_4513_n509) );
  AND2X2 AND2X2_8 ( .A(_abc_4513_n368), .B(Wready), .Y(_abc_4513_n372) );
  AND2X2 AND2X2_80 ( .A(_abc_4513_n510_1), .B(_abc_4513_n473), .Y(Wstrb_2__FF_INPUT) );
  AND2X2 AND2X2_81 ( .A(_abc_4513_n505), .B(_abc_4513_n491), .Y(_abc_4513_n512) );
  AND2X2 AND2X2_82 ( .A(_abc_4513_n512), .B(_abc_4513_n476), .Y(_abc_4513_n513_1) );
  AND2X2 AND2X2_83 ( .A(_abc_4513_n514), .B(_abc_4513_n473), .Y(Wstrb_3__FF_INPUT) );
  AND2X2 AND2X2_84 ( .A(_abc_4513_n462_1), .B(resetn), .Y(_abc_4513_n516_1) );
  AND2X2 AND2X2_85 ( .A(_abc_4513_n517), .B(_abc_4513_n516_1), .Y(_abc_4513_n518) );
  AND2X2 AND2X2_86 ( .A(_abc_4513_n518), .B(\W_R[1] ), .Y(_abc_4513_n519_1) );
  AND2X2 AND2X2_87 ( .A(_abc_4513_n519_1), .B(\Rdata_mem[0] ), .Y(_abc_4513_n520) );
  AND2X2 AND2X2_88 ( .A(_abc_4513_n521), .B(\inst[0] ), .Y(_abc_4513_n522_1) );
  AND2X2 AND2X2_89 ( .A(_abc_4513_n523), .B(resetn), .Y(inst_0__FF_INPUT) );
  AND2X2 AND2X2_9 ( .A(_abc_4513_n372), .B(state_3_), .Y(_abc_4513_n373) );
  AND2X2 AND2X2_90 ( .A(_abc_4513_n519_1), .B(\Rdata_mem[1] ), .Y(_abc_4513_n525_1) );
  AND2X2 AND2X2_91 ( .A(_abc_4513_n521), .B(\inst[1] ), .Y(_abc_4513_n526) );
  AND2X2 AND2X2_92 ( .A(_abc_4513_n527), .B(resetn), .Y(inst_1__FF_INPUT) );
  AND2X2 AND2X2_93 ( .A(_abc_4513_n519_1), .B(\Rdata_mem[2] ), .Y(_abc_4513_n529) );
  AND2X2 AND2X2_94 ( .A(_abc_4513_n521), .B(\inst[2] ), .Y(_abc_4513_n530) );
  AND2X2 AND2X2_95 ( .A(_abc_4513_n531), .B(resetn), .Y(inst_2__FF_INPUT) );
  AND2X2 AND2X2_96 ( .A(_abc_4513_n519_1), .B(\Rdata_mem[3] ), .Y(_abc_4513_n533_1) );
  AND2X2 AND2X2_97 ( .A(_abc_4513_n521), .B(\inst[3] ), .Y(_abc_4513_n534) );
  AND2X2 AND2X2_98 ( .A(_abc_4513_n535_1), .B(resetn), .Y(inst_3__FF_INPUT) );
  AND2X2 AND2X2_99 ( .A(_abc_4513_n519_1), .B(\Rdata_mem[4] ), .Y(_abc_4513_n537_1) );
  DFFPOSX1 DFFPOSX1_1 ( .CLK(clock), .D(_abc_3815_n99), .Q(state_0_) );
  DFFPOSX1 DFFPOSX1_10 ( .CLK(clock), .D(Wdata_2__FF_INPUT), .Q(\Wdata[2] ) );
  DFFPOSX1 DFFPOSX1_11 ( .CLK(clock), .D(Wdata_3__FF_INPUT), .Q(\Wdata[3] ) );
  DFFPOSX1 DFFPOSX1_12 ( .CLK(clock), .D(Wdata_4__FF_INPUT), .Q(\Wdata[4] ) );
  DFFPOSX1 DFFPOSX1_13 ( .CLK(clock), .D(Wdata_5__FF_INPUT), .Q(\Wdata[5] ) );
  DFFPOSX1 DFFPOSX1_14 ( .CLK(clock), .D(Wdata_6__FF_INPUT), .Q(\Wdata[6] ) );
  DFFPOSX1 DFFPOSX1_15 ( .CLK(clock), .D(Wdata_7__FF_INPUT), .Q(\Wdata[7] ) );
  DFFPOSX1 DFFPOSX1_16 ( .CLK(clock), .D(Wdata_8__FF_INPUT), .Q(\Wdata[8] ) );
  DFFPOSX1 DFFPOSX1_17 ( .CLK(clock), .D(Wdata_9__FF_INPUT), .Q(\Wdata[9] ) );
  DFFPOSX1 DFFPOSX1_18 ( .CLK(clock), .D(Wdata_10__FF_INPUT), .Q(\Wdata[10] ) );
  DFFPOSX1 DFFPOSX1_19 ( .CLK(clock), .D(Wdata_11__FF_INPUT), .Q(\Wdata[11] ) );
  DFFPOSX1 DFFPOSX1_2 ( .CLK(clock), .D(_abc_3815_n23), .Q(state_1_) );
  DFFPOSX1 DFFPOSX1_20 ( .CLK(clock), .D(Wdata_12__FF_INPUT), .Q(\Wdata[12] ) );
  DFFPOSX1 DFFPOSX1_21 ( .CLK(clock), .D(Wdata_13__FF_INPUT), .Q(\Wdata[13] ) );
  DFFPOSX1 DFFPOSX1_22 ( .CLK(clock), .D(Wdata_14__FF_INPUT), .Q(\Wdata[14] ) );
  DFFPOSX1 DFFPOSX1_23 ( .CLK(clock), .D(Wdata_15__FF_INPUT), .Q(\Wdata[15] ) );
  DFFPOSX1 DFFPOSX1_24 ( .CLK(clock), .D(Wdata_16__FF_INPUT), .Q(\Wdata[16] ) );
  DFFPOSX1 DFFPOSX1_25 ( .CLK(clock), .D(Wdata_17__FF_INPUT), .Q(\Wdata[17] ) );
  DFFPOSX1 DFFPOSX1_26 ( .CLK(clock), .D(Wdata_18__FF_INPUT), .Q(\Wdata[18] ) );
  DFFPOSX1 DFFPOSX1_27 ( .CLK(clock), .D(Wdata_19__FF_INPUT), .Q(\Wdata[19] ) );
  DFFPOSX1 DFFPOSX1_28 ( .CLK(clock), .D(Wdata_20__FF_INPUT), .Q(\Wdata[20] ) );
  DFFPOSX1 DFFPOSX1_29 ( .CLK(clock), .D(Wdata_21__FF_INPUT), .Q(\Wdata[21] ) );
  DFFPOSX1 DFFPOSX1_3 ( .CLK(clock), .D(_abc_3815_n14), .Q(state_2_) );
  DFFPOSX1 DFFPOSX1_30 ( .CLK(clock), .D(Wdata_22__FF_INPUT), .Q(\Wdata[22] ) );
  DFFPOSX1 DFFPOSX1_31 ( .CLK(clock), .D(Wdata_23__FF_INPUT), .Q(\Wdata[23] ) );
  DFFPOSX1 DFFPOSX1_32 ( .CLK(clock), .D(Wdata_24__FF_INPUT), .Q(\Wdata[24] ) );
  DFFPOSX1 DFFPOSX1_33 ( .CLK(clock), .D(Wdata_25__FF_INPUT), .Q(\Wdata[25] ) );
  DFFPOSX1 DFFPOSX1_34 ( .CLK(clock), .D(Wdata_26__FF_INPUT), .Q(\Wdata[26] ) );
  DFFPOSX1 DFFPOSX1_35 ( .CLK(clock), .D(Wdata_27__FF_INPUT), .Q(\Wdata[27] ) );
  DFFPOSX1 DFFPOSX1_36 ( .CLK(clock), .D(Wdata_28__FF_INPUT), .Q(\Wdata[28] ) );
  DFFPOSX1 DFFPOSX1_37 ( .CLK(clock), .D(Wdata_29__FF_INPUT), .Q(\Wdata[29] ) );
  DFFPOSX1 DFFPOSX1_38 ( .CLK(clock), .D(Wdata_30__FF_INPUT), .Q(\Wdata[30] ) );
  DFFPOSX1 DFFPOSX1_39 ( .CLK(clock), .D(Wdata_31__FF_INPUT), .Q(\Wdata[31] ) );
  DFFPOSX1 DFFPOSX1_4 ( .CLK(clock), .D(_abc_3815_n122), .Q(state_3_) );
  DFFPOSX1 DFFPOSX1_40 ( .CLK(clock), .D(inst_0__FF_INPUT), .Q(\inst[0] ) );
  DFFPOSX1 DFFPOSX1_41 ( .CLK(clock), .D(inst_1__FF_INPUT), .Q(\inst[1] ) );
  DFFPOSX1 DFFPOSX1_42 ( .CLK(clock), .D(inst_2__FF_INPUT), .Q(\inst[2] ) );
  DFFPOSX1 DFFPOSX1_43 ( .CLK(clock), .D(inst_3__FF_INPUT), .Q(\inst[3] ) );
  DFFPOSX1 DFFPOSX1_44 ( .CLK(clock), .D(inst_4__FF_INPUT), .Q(\inst[4] ) );
  DFFPOSX1 DFFPOSX1_45 ( .CLK(clock), .D(inst_5__FF_INPUT), .Q(\inst[5] ) );
  DFFPOSX1 DFFPOSX1_46 ( .CLK(clock), .D(inst_6__FF_INPUT), .Q(\inst[6] ) );
  DFFPOSX1 DFFPOSX1_47 ( .CLK(clock), .D(inst_7__FF_INPUT), .Q(\inst[7] ) );
  DFFPOSX1 DFFPOSX1_48 ( .CLK(clock), .D(inst_8__FF_INPUT), .Q(\inst[8] ) );
  DFFPOSX1 DFFPOSX1_49 ( .CLK(clock), .D(inst_9__FF_INPUT), .Q(\inst[9] ) );
  DFFPOSX1 DFFPOSX1_5 ( .CLK(clock), .D(_abc_3815_n132), .Q(state_4_) );
  DFFPOSX1 DFFPOSX1_50 ( .CLK(clock), .D(inst_10__FF_INPUT), .Q(\inst[10] ) );
  DFFPOSX1 DFFPOSX1_51 ( .CLK(clock), .D(inst_11__FF_INPUT), .Q(\inst[11] ) );
  DFFPOSX1 DFFPOSX1_52 ( .CLK(clock), .D(inst_12__FF_INPUT), .Q(\inst[12] ) );
  DFFPOSX1 DFFPOSX1_53 ( .CLK(clock), .D(inst_13__FF_INPUT), .Q(\inst[13] ) );
  DFFPOSX1 DFFPOSX1_54 ( .CLK(clock), .D(inst_14__FF_INPUT), .Q(\inst[14] ) );
  DFFPOSX1 DFFPOSX1_55 ( .CLK(clock), .D(inst_15__FF_INPUT), .Q(\inst[15] ) );
  DFFPOSX1 DFFPOSX1_56 ( .CLK(clock), .D(inst_16__FF_INPUT), .Q(\inst[16] ) );
  DFFPOSX1 DFFPOSX1_57 ( .CLK(clock), .D(inst_17__FF_INPUT), .Q(\inst[17] ) );
  DFFPOSX1 DFFPOSX1_58 ( .CLK(clock), .D(inst_18__FF_INPUT), .Q(\inst[18] ) );
  DFFPOSX1 DFFPOSX1_59 ( .CLK(clock), .D(inst_19__FF_INPUT), .Q(\inst[19] ) );
  DFFPOSX1 DFFPOSX1_6 ( .CLK(clock), .D(_abc_3815_n52), .Q(state_5_) );
  DFFPOSX1 DFFPOSX1_60 ( .CLK(clock), .D(inst_20__FF_INPUT), .Q(\inst[20] ) );
  DFFPOSX1 DFFPOSX1_61 ( .CLK(clock), .D(inst_21__FF_INPUT), .Q(\inst[21] ) );
  DFFPOSX1 DFFPOSX1_62 ( .CLK(clock), .D(inst_22__FF_INPUT), .Q(\inst[22] ) );
  DFFPOSX1 DFFPOSX1_63 ( .CLK(clock), .D(inst_23__FF_INPUT), .Q(\inst[23] ) );
  DFFPOSX1 DFFPOSX1_64 ( .CLK(clock), .D(inst_24__FF_INPUT), .Q(\inst[24] ) );
  DFFPOSX1 DFFPOSX1_65 ( .CLK(clock), .D(inst_25__FF_INPUT), .Q(\inst[25] ) );
  DFFPOSX1 DFFPOSX1_66 ( .CLK(clock), .D(inst_26__FF_INPUT), .Q(\inst[26] ) );
  DFFPOSX1 DFFPOSX1_67 ( .CLK(clock), .D(inst_27__FF_INPUT), .Q(\inst[27] ) );
  DFFPOSX1 DFFPOSX1_68 ( .CLK(clock), .D(inst_28__FF_INPUT), .Q(\inst[28] ) );
  DFFPOSX1 DFFPOSX1_69 ( .CLK(clock), .D(inst_29__FF_INPUT), .Q(\inst[29] ) );
  DFFPOSX1 DFFPOSX1_7 ( .CLK(clock), .D(_abc_3815_n152), .Q(state_6_) );
  DFFPOSX1 DFFPOSX1_70 ( .CLK(clock), .D(inst_30__FF_INPUT), .Q(\inst[30] ) );
  DFFPOSX1 DFFPOSX1_71 ( .CLK(clock), .D(inst_31__FF_INPUT), .Q(\inst[31] ) );
  DFFPOSX1 DFFPOSX1_72 ( .CLK(clock), .D(Wstrb_0__FF_INPUT), .Q(\Wstrb[0] ) );
  DFFPOSX1 DFFPOSX1_73 ( .CLK(clock), .D(Wstrb_1__FF_INPUT), .Q(\Wstrb[1] ) );
  DFFPOSX1 DFFPOSX1_74 ( .CLK(clock), .D(Wstrb_2__FF_INPUT), .Q(\Wstrb[2] ) );
  DFFPOSX1 DFFPOSX1_75 ( .CLK(clock), .D(Wstrb_3__FF_INPUT), .Q(\Wstrb[3] ) );
  DFFPOSX1 DFFPOSX1_8 ( .CLK(clock), .D(Wdata_0__FF_INPUT), .Q(\Wdata[0] ) );
  DFFPOSX1 DFFPOSX1_9 ( .CLK(clock), .D(Wdata_1__FF_INPUT), .Q(\Wdata[1] ) );
  INVX1 INVX1_1 ( .A(ARready), .Y(_abc_4513_n361) );
  INVX1 INVX1_10 ( .A(resetn), .Y(_abc_4513_n416_1) );
  INVX1 INVX1_100 ( .A(_abc_4513_n1337), .Y(_abc_4513_n1338) );
  INVX1 INVX1_101 ( .A(_abc_4513_n1333), .Y(_abc_4513_n1340) );
  INVX1 INVX1_102 ( .A(_abc_4513_n1355), .Y(_abc_4513_n1356) );
  INVX1 INVX1_103 ( .A(_abc_4513_n1359), .Y(_abc_4513_n1360) );
  INVX1 INVX1_104 ( .A(_abc_4513_n1364), .Y(_abc_4513_n1365) );
  INVX1 INVX1_105 ( .A(_abc_4513_n1367), .Y(_abc_4513_n1368) );
  INVX1 INVX1_106 ( .A(_abc_4513_n1369), .Y(_abc_4513_n1371) );
  INVX1 INVX1_107 ( .A(_abc_4513_n1384), .Y(_abc_4513_n1385) );
  INVX1 INVX1_108 ( .A(_abc_4513_n971), .Y(_abc_4513_n1390) );
  INVX1 INVX1_109 ( .A(_abc_4513_n974), .Y(_abc_4513_n1392) );
  INVX1 INVX1_11 ( .A(enable), .Y(_abc_4513_n419_1) );
  INVX1 INVX1_110 ( .A(_abc_4513_n1031), .Y(_abc_4513_n1394) );
  INVX1 INVX1_111 ( .A(_abc_4513_n1036), .Y(_abc_4513_n1396) );
  INVX1 INVX1_112 ( .A(_abc_4513_n1155), .Y(_abc_4513_n1398) );
  INVX1 INVX1_113 ( .A(_abc_4513_n1162), .Y(_abc_4513_n1400) );
  INVX1 INVX1_114 ( .A(_abc_4513_n1283), .Y(_abc_4513_n1402) );
  INVX1 INVX1_115 ( .A(_abc_4513_n1290), .Y(_abc_4513_n1404) );
  INVX1 INVX1_116 ( .A(_abc_4513_n1347), .Y(_abc_4513_n1406) );
  INVX1 INVX1_117 ( .A(_abc_4513_n1352), .Y(_abc_4513_n1408) );
  INVX1 INVX1_118 ( .A(_abc_4513_n1378), .Y(_abc_4513_n1410) );
  INVX1 INVX1_119 ( .A(_abc_4513_n1381), .Y(_abc_4513_n1412) );
  INVX1 INVX1_12 ( .A(state_3_), .Y(_abc_4513_n426) );
  INVX1 INVX1_120 ( .A(_abc_4513_n1386), .Y(_abc_4513_n1414) );
  INVX1 INVX1_121 ( .A(\imm[31] ), .Y(_abc_4513_n1421) );
  INVX1 INVX1_122 ( .A(\rs1[31] ), .Y(_abc_4513_n1423) );
  INVX1 INVX1_123 ( .A(_abc_4513_n1425), .Y(_abc_4513_n1426) );
  INVX1 INVX1_13 ( .A(_abc_4513_n427_1), .Y(_abc_4513_n428) );
  INVX1 INVX1_14 ( .A(_abc_4513_n430), .Y(_abc_4513_n431) );
  INVX1 INVX1_15 ( .A(_abc_4513_n436), .Y(_abc_4513_n437) );
  INVX1 INVX1_16 ( .A(_abc_4513_n409), .Y(_abc_4513_n446_1) );
  INVX1 INVX1_17 ( .A(_abc_4513_n447), .Y(_abc_4513_n448) );
  INVX1 INVX1_18 ( .A(_abc_4513_n450), .Y(_abc_4513_n451) );
  INVX1 INVX1_19 ( .A(state_6_), .Y(_abc_4513_n452) );
  INVX1 INVX1_2 ( .A(Bvalid), .Y(_abc_4513_n368) );
  INVX1 INVX1_20 ( .A(_abc_4513_n455), .Y(_abc_4513_n456) );
  INVX1 INVX1_21 ( .A(_abc_4513_n459), .Y(_abc_4513_n460) );
  INVX1 INVX1_22 ( .A(busy), .Y(done) );
  INVX1 INVX1_23 ( .A(_abc_4513_n470_1), .Y(_abc_4513_n471) );
  INVX1 INVX1_24 ( .A(\wordsize[0] ), .Y(_abc_4513_n474) );
  INVX1 INVX1_25 ( .A(_abc_4513_n479), .Y(_abc_4513_n480) );
  INVX1 INVX1_26 ( .A(_abc_4513_n477), .Y(_abc_4513_n483) );
  INVX1 INVX1_27 ( .A(\imm[1] ), .Y(_abc_4513_n484) );
  INVX1 INVX1_28 ( .A(\rs1[1] ), .Y(_abc_4513_n485) );
  INVX1 INVX1_29 ( .A(_abc_4513_n491), .Y(_abc_4513_n492) );
  INVX1 INVX1_3 ( .A(_abc_4513_n362_1), .Y(_abc_4513_n379) );
  INVX1 INVX1_30 ( .A(_abc_4513_n658_1), .Y(_abc_4513_n765) );
  INVX1 INVX1_31 ( .A(_abc_4513_n493), .Y(_abc_4513_n842_1) );
  INVX1 INVX1_32 ( .A(_abc_4513_n947), .Y(_abc_4513_n948) );
  INVX1 INVX1_33 ( .A(_abc_4513_n951), .Y(_abc_4513_n952) );
  INVX1 INVX1_34 ( .A(_abc_4513_n958), .Y(_abc_4513_n959) );
  INVX1 INVX1_35 ( .A(_abc_4513_n961), .Y(_abc_4513_n962) );
  INVX1 INVX1_36 ( .A(_abc_4513_n963), .Y(_abc_4513_n964) );
  INVX1 INVX1_37 ( .A(_abc_4513_n977), .Y(_abc_4513_n978) );
  INVX1 INVX1_38 ( .A(_abc_4513_n980), .Y(_abc_4513_n981) );
  INVX1 INVX1_39 ( .A(_abc_4513_n987), .Y(_abc_4513_n988) );
  INVX1 INVX1_4 ( .A(Rvalid), .Y(_abc_4513_n387_1) );
  INVX1 INVX1_40 ( .A(_abc_4513_n990), .Y(_abc_4513_n991) );
  INVX1 INVX1_41 ( .A(_abc_4513_n992), .Y(_abc_4513_n994) );
  INVX1 INVX1_42 ( .A(_abc_4513_n1006), .Y(_abc_4513_n1007) );
  INVX1 INVX1_43 ( .A(_abc_4513_n1011), .Y(_abc_4513_n1012) );
  INVX1 INVX1_44 ( .A(_abc_4513_n1019), .Y(_abc_4513_n1020) );
  INVX1 INVX1_45 ( .A(_abc_4513_n1021), .Y(_abc_4513_n1022) );
  INVX1 INVX1_46 ( .A(_abc_4513_n1017), .Y(_abc_4513_n1024) );
  INVX1 INVX1_47 ( .A(_abc_4513_n1038), .Y(_abc_4513_n1039) );
  INVX1 INVX1_48 ( .A(_abc_4513_n1043), .Y(_abc_4513_n1044) );
  INVX1 INVX1_49 ( .A(_abc_4513_n1048), .Y(_abc_4513_n1049) );
  INVX1 INVX1_5 ( .A(AWready), .Y(_abc_4513_n394) );
  INVX1 INVX1_50 ( .A(_abc_4513_n1051), .Y(_abc_4513_n1052) );
  INVX1 INVX1_51 ( .A(_abc_4513_n1053), .Y(_abc_4513_n1055) );
  INVX1 INVX1_52 ( .A(_abc_4513_n1067), .Y(_abc_4513_n1068) );
  INVX1 INVX1_53 ( .A(_abc_4513_n1072), .Y(_abc_4513_n1073) );
  INVX1 INVX1_54 ( .A(_abc_4513_n1079), .Y(_abc_4513_n1080) );
  INVX1 INVX1_55 ( .A(_abc_4513_n1081), .Y(_abc_4513_n1082) );
  INVX1 INVX1_56 ( .A(_abc_4513_n1077), .Y(_abc_4513_n1084) );
  INVX1 INVX1_57 ( .A(_abc_4513_n1100), .Y(_abc_4513_n1101) );
  INVX1 INVX1_58 ( .A(_abc_4513_n1104), .Y(_abc_4513_n1105) );
  INVX1 INVX1_59 ( .A(_abc_4513_n1109), .Y(_abc_4513_n1110) );
  INVX1 INVX1_6 ( .A(_abc_4513_n395_1), .Y(_abc_4513_n396_1) );
  INVX1 INVX1_60 ( .A(_abc_4513_n1112), .Y(_abc_4513_n1113) );
  INVX1 INVX1_61 ( .A(_abc_4513_n1114), .Y(_abc_4513_n1116) );
  INVX1 INVX1_62 ( .A(_abc_4513_n1124), .Y(_abc_4513_n1125) );
  INVX1 INVX1_63 ( .A(_abc_4513_n1129), .Y(_abc_4513_n1130) );
  INVX1 INVX1_64 ( .A(_abc_4513_n1134), .Y(_abc_4513_n1135) );
  INVX1 INVX1_65 ( .A(_abc_4513_n1142), .Y(_abc_4513_n1143) );
  INVX1 INVX1_66 ( .A(_abc_4513_n1144), .Y(_abc_4513_n1145) );
  INVX1 INVX1_67 ( .A(_abc_4513_n1140), .Y(_abc_4513_n1147) );
  INVX1 INVX1_68 ( .A(_abc_4513_n1164), .Y(_abc_4513_n1165) );
  INVX1 INVX1_69 ( .A(_abc_4513_n1169), .Y(_abc_4513_n1170) );
  INVX1 INVX1_7 ( .A(Wready), .Y(_abc_4513_n397) );
  INVX1 INVX1_70 ( .A(_abc_4513_n1174), .Y(_abc_4513_n1175) );
  INVX1 INVX1_71 ( .A(_abc_4513_n1176), .Y(_abc_4513_n1177) );
  INVX1 INVX1_72 ( .A(_abc_4513_n1179), .Y(_abc_4513_n1181) );
  INVX1 INVX1_73 ( .A(_abc_4513_n1189), .Y(_abc_4513_n1190) );
  INVX1 INVX1_74 ( .A(_abc_4513_n1194), .Y(_abc_4513_n1195) );
  INVX1 INVX1_75 ( .A(_abc_4513_n1199), .Y(_abc_4513_n1200) );
  INVX1 INVX1_76 ( .A(_abc_4513_n1206), .Y(_abc_4513_n1207) );
  INVX1 INVX1_77 ( .A(_abc_4513_n1209), .Y(_abc_4513_n1210) );
  INVX1 INVX1_78 ( .A(_abc_4513_n1205), .Y(_abc_4513_n1212) );
  INVX1 INVX1_79 ( .A(_abc_4513_n1226), .Y(_abc_4513_n1227) );
  INVX1 INVX1_8 ( .A(_abc_4513_n398_1), .Y(_abc_4513_n399_1) );
  INVX1 INVX1_80 ( .A(_abc_4513_n1225), .Y(_abc_4513_n1231) );
  INVX1 INVX1_81 ( .A(_abc_4513_n1229), .Y(_abc_4513_n1232) );
  INVX1 INVX1_82 ( .A(_abc_4513_n1238), .Y(_abc_4513_n1239) );
  INVX1 INVX1_83 ( .A(_abc_4513_n1241), .Y(_abc_4513_n1242) );
  INVX1 INVX1_84 ( .A(_abc_4513_n1237), .Y(_abc_4513_n1244) );
  INVX1 INVX1_85 ( .A(_abc_4513_n1252), .Y(_abc_4513_n1253) );
  INVX1 INVX1_86 ( .A(_abc_4513_n1257), .Y(_abc_4513_n1258) );
  INVX1 INVX1_87 ( .A(_abc_4513_n1262), .Y(_abc_4513_n1263) );
  INVX1 INVX1_88 ( .A(_abc_4513_n1269), .Y(_abc_4513_n1270) );
  INVX1 INVX1_89 ( .A(_abc_4513_n1272), .Y(_abc_4513_n1273) );
  INVX1 INVX1_9 ( .A(_abc_4513_n372), .Y(_abc_4513_n401_1) );
  INVX1 INVX1_90 ( .A(_abc_4513_n1268), .Y(_abc_4513_n1275) );
  INVX1 INVX1_91 ( .A(_abc_4513_n1292), .Y(_abc_4513_n1293) );
  INVX1 INVX1_92 ( .A(_abc_4513_n1297), .Y(_abc_4513_n1298) );
  INVX1 INVX1_93 ( .A(_abc_4513_n1302), .Y(_abc_4513_n1303) );
  INVX1 INVX1_94 ( .A(_abc_4513_n1304), .Y(_abc_4513_n1305) );
  INVX1 INVX1_95 ( .A(_abc_4513_n1307), .Y(_abc_4513_n1309) );
  INVX1 INVX1_96 ( .A(_abc_4513_n1317), .Y(_abc_4513_n1318) );
  INVX1 INVX1_97 ( .A(_abc_4513_n1322), .Y(_abc_4513_n1323) );
  INVX1 INVX1_98 ( .A(_abc_4513_n1327), .Y(_abc_4513_n1328) );
  INVX1 INVX1_99 ( .A(_abc_4513_n1335), .Y(_abc_4513_n1336) );
  INVX2 INVX2_1 ( .A(_abc_4513_n489), .Y(_abc_4513_n505) );
  INVX4 INVX4_1 ( .A(\wordsize[1] ), .Y(_abc_4513_n475) );
  INVX8 INVX8_1 ( .A(_abc_4513_n519_1), .Y(_abc_4513_n521) );
  INVX8 INVX8_2 ( .A(\W_R[1] ), .Y(_abc_4513_n769_1) );
  OR2X2 OR2X2_1 ( .A(\W_R[0] ), .B(\W_R[1] ), .Y(_abc_4513_n362_1) );
  OR2X2 OR2X2_10 ( .A(_abc_4513_n412), .B(_abc_4513_n411_1), .Y(_abc_4513_n413_1) );
  OR2X2 OR2X2_100 ( .A(_abc_4513_n674), .B(_abc_4513_n742), .Y(_abc_4513_n743) );
  OR2X2 OR2X2_101 ( .A(_abc_4513_n743), .B(_abc_4513_n744), .Y(_abc_4513_n745_1) );
  OR2X2 OR2X2_102 ( .A(_abc_4513_n678), .B(_abc_4513_n747_1), .Y(_abc_4513_n748_1) );
  OR2X2 OR2X2_103 ( .A(_abc_4513_n748_1), .B(_abc_4513_n749), .Y(_abc_4513_n750) );
  OR2X2 OR2X2_104 ( .A(_abc_4513_n682_1), .B(_abc_4513_n752), .Y(_abc_4513_n753_1) );
  OR2X2 OR2X2_105 ( .A(_abc_4513_n753_1), .B(_abc_4513_n754_1), .Y(_abc_4513_n755_1) );
  OR2X2 OR2X2_106 ( .A(_abc_4513_n686), .B(_abc_4513_n757), .Y(_abc_4513_n758) );
  OR2X2 OR2X2_107 ( .A(_abc_4513_n758), .B(_abc_4513_n759), .Y(_abc_4513_n760) );
  OR2X2 OR2X2_108 ( .A(_abc_4513_n419_1), .B(\W_R[1] ), .Y(_abc_4513_n764) );
  OR2X2 OR2X2_109 ( .A(_abc_4513_n765), .B(_abc_4513_n764), .Y(_abc_4513_n766_1) );
  OR2X2 OR2X2_11 ( .A(_abc_4513_n417_1), .B(_abc_4513_n416_1), .Y(_abc_4513_n418) );
  OR2X2 OR2X2_110 ( .A(_abc_4513_n766_1), .B(_abc_4513_n763), .Y(_abc_4513_n767_1) );
  OR2X2 OR2X2_111 ( .A(_abc_4513_n762), .B(_abc_4513_n767_1), .Y(align) );
  OR2X2 OR2X2_112 ( .A(_abc_4513_n509), .B(_abc_4513_n506), .Y(_abc_4513_n772) );
  OR2X2 OR2X2_113 ( .A(_abc_4513_n776_1), .B(_abc_4513_n775_1), .Y(_abc_4513_n777_1) );
  OR2X2 OR2X2_114 ( .A(_abc_4513_n777_1), .B(_abc_4513_n774_1), .Y(_abc_4513_n778) );
  OR2X2 OR2X2_115 ( .A(_abc_4513_n778), .B(_abc_4513_n773), .Y(_abc_4513_n779) );
  OR2X2 OR2X2_116 ( .A(_abc_4513_n784), .B(_abc_4513_n783), .Y(_abc_4513_n785) );
  OR2X2 OR2X2_117 ( .A(_abc_4513_n785), .B(_abc_4513_n782), .Y(_abc_4513_n786_1) );
  OR2X2 OR2X2_118 ( .A(_abc_4513_n786_1), .B(_abc_4513_n781), .Y(_abc_4513_n787_1) );
  OR2X2 OR2X2_119 ( .A(_abc_4513_n791), .B(_abc_4513_n792), .Y(_abc_4513_n793) );
  OR2X2 OR2X2_12 ( .A(_abc_4513_n418), .B(_abc_4513_n420_1), .Y(_abc_4513_n421) );
  OR2X2 OR2X2_120 ( .A(_abc_4513_n793), .B(_abc_4513_n790), .Y(_abc_4513_n794_1) );
  OR2X2 OR2X2_121 ( .A(_abc_4513_n794_1), .B(_abc_4513_n789_1), .Y(_abc_4513_n795_1) );
  OR2X2 OR2X2_122 ( .A(_abc_4513_n800), .B(_abc_4513_n799), .Y(_abc_4513_n801) );
  OR2X2 OR2X2_123 ( .A(_abc_4513_n801), .B(_abc_4513_n798), .Y(_abc_4513_n802) );
  OR2X2 OR2X2_124 ( .A(_abc_4513_n802), .B(_abc_4513_n797_1), .Y(_abc_4513_n803) );
  OR2X2 OR2X2_125 ( .A(_abc_4513_n808), .B(_abc_4513_n807), .Y(_abc_4513_n809) );
  OR2X2 OR2X2_126 ( .A(_abc_4513_n809), .B(_abc_4513_n806), .Y(_abc_4513_n810) );
  OR2X2 OR2X2_127 ( .A(_abc_4513_n810), .B(_abc_4513_n805), .Y(_abc_4513_n811_1) );
  OR2X2 OR2X2_128 ( .A(_abc_4513_n816), .B(_abc_4513_n815), .Y(_abc_4513_n817) );
  OR2X2 OR2X2_129 ( .A(_abc_4513_n817), .B(_abc_4513_n814_1), .Y(_abc_4513_n818) );
  OR2X2 OR2X2_13 ( .A(_abc_4513_n421), .B(_abc_4513_n415), .Y(_abc_4513_n422_1) );
  OR2X2 OR2X2_130 ( .A(_abc_4513_n818), .B(_abc_4513_n813_1), .Y(_abc_4513_n819_1) );
  OR2X2 OR2X2_131 ( .A(_abc_4513_n823), .B(_abc_4513_n824), .Y(_abc_4513_n825) );
  OR2X2 OR2X2_132 ( .A(_abc_4513_n825), .B(_abc_4513_n822_1), .Y(_abc_4513_n826) );
  OR2X2 OR2X2_133 ( .A(_abc_4513_n826), .B(_abc_4513_n821_1), .Y(_abc_4513_n827) );
  OR2X2 OR2X2_134 ( .A(_abc_4513_n829), .B(_abc_4513_n830), .Y(_abc_4513_n831) );
  OR2X2 OR2X2_135 ( .A(_abc_4513_n832), .B(_abc_4513_n833_1), .Y(_abc_4513_n834_1) );
  OR2X2 OR2X2_136 ( .A(_abc_4513_n831), .B(_abc_4513_n834_1), .Y(_abc_4513_n835_1) );
  OR2X2 OR2X2_137 ( .A(_abc_4513_n838), .B(_abc_4513_n837), .Y(_abc_4513_n839) );
  OR2X2 OR2X2_138 ( .A(_abc_4513_n836_1), .B(_abc_4513_n839), .Y(_abc_4513_n840) );
  OR2X2 OR2X2_139 ( .A(_abc_4513_n842_1), .B(\Rdata_mem[7] ), .Y(_abc_4513_n843_1) );
  OR2X2 OR2X2_14 ( .A(_abc_4513_n422_1), .B(_abc_4513_n413_1), .Y(_abc_4513_n423) );
  OR2X2 OR2X2_140 ( .A(_abc_4513_n847), .B(_abc_4513_n846), .Y(_abc_4513_n848) );
  OR2X2 OR2X2_141 ( .A(_abc_4513_n845), .B(_abc_4513_n848), .Y(_abc_4513_n849) );
  OR2X2 OR2X2_142 ( .A(_abc_4513_n852), .B(_abc_4513_n851), .Y(_abc_4513_n853) );
  OR2X2 OR2X2_143 ( .A(_abc_4513_n845), .B(_abc_4513_n853), .Y(_abc_4513_n854) );
  OR2X2 OR2X2_144 ( .A(_abc_4513_n857_1), .B(_abc_4513_n856_1), .Y(_abc_4513_n858_1) );
  OR2X2 OR2X2_145 ( .A(_abc_4513_n845), .B(_abc_4513_n858_1), .Y(_abc_4513_n859_1) );
  OR2X2 OR2X2_146 ( .A(_abc_4513_n862), .B(_abc_4513_n861), .Y(_abc_4513_n863) );
  OR2X2 OR2X2_147 ( .A(_abc_4513_n845), .B(_abc_4513_n863), .Y(_abc_4513_n864) );
  OR2X2 OR2X2_148 ( .A(_abc_4513_n867_1), .B(_abc_4513_n866_1), .Y(_abc_4513_n868_1) );
  OR2X2 OR2X2_149 ( .A(_abc_4513_n845), .B(_abc_4513_n868_1), .Y(_abc_4513_n869_1) );
  OR2X2 OR2X2_15 ( .A(_abc_4513_n423), .B(_abc_4513_n410_1), .Y(_abc_4513_n424) );
  OR2X2 OR2X2_150 ( .A(_abc_4513_n872), .B(_abc_4513_n871), .Y(_abc_4513_n873) );
  OR2X2 OR2X2_151 ( .A(_abc_4513_n845), .B(_abc_4513_n873), .Y(_abc_4513_n874) );
  OR2X2 OR2X2_152 ( .A(_abc_4513_n877), .B(_abc_4513_n876), .Y(_abc_4513_n878_1) );
  OR2X2 OR2X2_153 ( .A(_abc_4513_n845), .B(_abc_4513_n878_1), .Y(_abc_4513_n879_1) );
  OR2X2 OR2X2_154 ( .A(_abc_4513_n881_1), .B(_abc_4513_n882), .Y(_abc_4513_n883) );
  OR2X2 OR2X2_155 ( .A(_abc_4513_n845), .B(_abc_4513_n883), .Y(_abc_4513_n884) );
  OR2X2 OR2X2_156 ( .A(_abc_4513_n888_1), .B(_abc_4513_n887_1), .Y(_abc_4513_n889) );
  OR2X2 OR2X2_157 ( .A(_abc_4513_n845), .B(_abc_4513_n891), .Y(_abc_4513_n892) );
  OR2X2 OR2X2_158 ( .A(_abc_4513_n892), .B(_abc_4513_n886_1), .Y(_abc_4513_n893) );
  OR2X2 OR2X2_159 ( .A(_abc_4513_n892), .B(_abc_4513_n895), .Y(_abc_4513_n896_1) );
  OR2X2 OR2X2_16 ( .A(_abc_4513_n408_1), .B(_abc_4513_n424), .Y(_abc_3815_n99) );
  OR2X2 OR2X2_160 ( .A(_abc_4513_n892), .B(_abc_4513_n898), .Y(_abc_4513_n899_1) );
  OR2X2 OR2X2_161 ( .A(_abc_4513_n892), .B(_abc_4513_n901), .Y(_abc_4513_n902_1) );
  OR2X2 OR2X2_162 ( .A(_abc_4513_n892), .B(_abc_4513_n904_1), .Y(_abc_4513_n905) );
  OR2X2 OR2X2_163 ( .A(_abc_4513_n892), .B(_abc_4513_n907), .Y(_abc_4513_n908) );
  OR2X2 OR2X2_164 ( .A(_abc_4513_n892), .B(_abc_4513_n910), .Y(_abc_4513_n911) );
  OR2X2 OR2X2_165 ( .A(_abc_4513_n892), .B(_abc_4513_n913), .Y(_abc_4513_n914) );
  OR2X2 OR2X2_166 ( .A(_abc_4513_n892), .B(_abc_4513_n916), .Y(_abc_4513_n917) );
  OR2X2 OR2X2_167 ( .A(_abc_4513_n892), .B(_abc_4513_n919), .Y(_abc_4513_n920) );
  OR2X2 OR2X2_168 ( .A(_abc_4513_n892), .B(_abc_4513_n922), .Y(_abc_4513_n923) );
  OR2X2 OR2X2_169 ( .A(_abc_4513_n892), .B(_abc_4513_n925), .Y(_abc_4513_n926) );
  OR2X2 OR2X2_17 ( .A(_abc_4513_n393_1), .B(_abc_4513_n426), .Y(_abc_4513_n427_1) );
  OR2X2 OR2X2_170 ( .A(_abc_4513_n892), .B(_abc_4513_n928), .Y(_abc_4513_n929) );
  OR2X2 OR2X2_171 ( .A(_abc_4513_n892), .B(_abc_4513_n931), .Y(_abc_4513_n932) );
  OR2X2 OR2X2_172 ( .A(_abc_4513_n892), .B(_abc_4513_n934), .Y(_abc_4513_n935) );
  OR2X2 OR2X2_173 ( .A(_abc_4513_n892), .B(_abc_4513_n937), .Y(_abc_4513_n938) );
  OR2X2 OR2X2_174 ( .A(_abc_4513_n491), .B(\W_R[1] ), .Y(_abc_4513_n940) );
  OR2X2 OR2X2_175 ( .A(_abc_4513_n769_1), .B(\pc[0] ), .Y(_abc_4513_n941) );
  OR2X2 OR2X2_176 ( .A(_abc_4513_n505), .B(\W_R[1] ), .Y(_abc_4513_n943) );
  OR2X2 OR2X2_177 ( .A(_abc_4513_n769_1), .B(\pc[1] ), .Y(_abc_4513_n944) );
  OR2X2 OR2X2_178 ( .A(_abc_4513_n482), .B(_abc_4513_n479), .Y(_abc_4513_n946) );
  OR2X2 OR2X2_179 ( .A(\imm[2] ), .B(\rs1[2] ), .Y(_abc_4513_n949) );
  OR2X2 OR2X2_18 ( .A(_abc_4513_n432), .B(_abc_4513_n378_1), .Y(_abc_4513_n433) );
  OR2X2 OR2X2_180 ( .A(_abc_4513_n946), .B(_abc_4513_n950), .Y(_abc_4513_n953) );
  OR2X2 OR2X2_181 ( .A(_abc_4513_n954), .B(\W_R[1] ), .Y(_abc_4513_n955) );
  OR2X2 OR2X2_182 ( .A(_abc_4513_n769_1), .B(\pc[2] ), .Y(_abc_4513_n956) );
  OR2X2 OR2X2_183 ( .A(\imm[3] ), .B(\rs1[3] ), .Y(_abc_4513_n960) );
  OR2X2 OR2X2_184 ( .A(_abc_4513_n965), .B(_abc_4513_n966), .Y(_abc_4513_n967) );
  OR2X2 OR2X2_185 ( .A(_abc_4513_n968), .B(_abc_4513_n969), .Y(\AWdata[3] ) );
  OR2X2 OR2X2_186 ( .A(_abc_4513_n973), .B(_abc_4513_n961), .Y(_abc_4513_n974) );
  OR2X2 OR2X2_187 ( .A(_abc_4513_n972), .B(_abc_4513_n974), .Y(_abc_4513_n975) );
  OR2X2 OR2X2_188 ( .A(\imm[4] ), .B(\rs1[4] ), .Y(_abc_4513_n976) );
  OR2X2 OR2X2_189 ( .A(_abc_4513_n975), .B(_abc_4513_n979), .Y(_abc_4513_n982) );
  OR2X2 OR2X2_19 ( .A(_abc_4513_n434), .B(_abc_4513_n429), .Y(_abc_3815_n122) );
  OR2X2 OR2X2_190 ( .A(_abc_4513_n983), .B(\W_R[1] ), .Y(_abc_4513_n984) );
  OR2X2 OR2X2_191 ( .A(_abc_4513_n769_1), .B(\pc[4] ), .Y(_abc_4513_n985) );
  OR2X2 OR2X2_192 ( .A(\imm[5] ), .B(\rs1[5] ), .Y(_abc_4513_n989) );
  OR2X2 OR2X2_193 ( .A(_abc_4513_n988), .B(_abc_4513_n992), .Y(_abc_4513_n993) );
  OR2X2 OR2X2_194 ( .A(_abc_4513_n987), .B(_abc_4513_n994), .Y(_abc_4513_n995) );
  OR2X2 OR2X2_195 ( .A(_abc_4513_n996), .B(\W_R[1] ), .Y(_abc_4513_n997) );
  OR2X2 OR2X2_196 ( .A(_abc_4513_n769_1), .B(\pc[5] ), .Y(_abc_4513_n998) );
  OR2X2 OR2X2_197 ( .A(_abc_4513_n977), .B(_abc_4513_n990), .Y(_abc_4513_n1001) );
  OR2X2 OR2X2_198 ( .A(_abc_4513_n1004), .B(_abc_4513_n1002), .Y(_abc_4513_n1005) );
  OR2X2 OR2X2_199 ( .A(\imm[6] ), .B(\rs1[6] ), .Y(_abc_4513_n1008) );
  OR2X2 OR2X2_2 ( .A(_abc_4513_n364), .B(state_2_), .Y(_abc_4513_n365) );
  OR2X2 OR2X2_20 ( .A(_abc_4513_n439), .B(_abc_4513_n440), .Y(_abc_3815_n132) );
  OR2X2 OR2X2_200 ( .A(_abc_4513_n1005), .B(_abc_4513_n1009), .Y(_abc_4513_n1010) );
  OR2X2 OR2X2_201 ( .A(_abc_4513_n1014), .B(_abc_4513_n1000), .Y(\AWdata[6] ) );
  OR2X2 OR2X2_202 ( .A(_abc_4513_n769_1), .B(\pc[7] ), .Y(_abc_4513_n1016) );
  OR2X2 OR2X2_203 ( .A(\imm[7] ), .B(\rs1[7] ), .Y(_abc_4513_n1018) );
  OR2X2 OR2X2_204 ( .A(_abc_4513_n1017), .B(_abc_4513_n1022), .Y(_abc_4513_n1023) );
  OR2X2 OR2X2_205 ( .A(_abc_4513_n1024), .B(_abc_4513_n1021), .Y(_abc_4513_n1025) );
  OR2X2 OR2X2_206 ( .A(_abc_4513_n1026), .B(\W_R[1] ), .Y(_abc_4513_n1027) );
  OR2X2 OR2X2_207 ( .A(_abc_4513_n1034), .B(_abc_4513_n1019), .Y(_abc_4513_n1035) );
  OR2X2 OR2X2_208 ( .A(_abc_4513_n1033), .B(_abc_4513_n1035), .Y(_abc_4513_n1036) );
  OR2X2 OR2X2_209 ( .A(_abc_4513_n1032), .B(_abc_4513_n1036), .Y(_abc_4513_n1037) );
  OR2X2 OR2X2_21 ( .A(_abc_4513_n444), .B(_abc_4513_n443), .Y(_abc_3815_n152) );
  OR2X2 OR2X2_210 ( .A(\imm[8] ), .B(\rs1[8] ), .Y(_abc_4513_n1040) );
  OR2X2 OR2X2_211 ( .A(_abc_4513_n1037), .B(_abc_4513_n1041), .Y(_abc_4513_n1042) );
  OR2X2 OR2X2_212 ( .A(_abc_4513_n1046), .B(_abc_4513_n1029), .Y(\AWdata[8] ) );
  OR2X2 OR2X2_213 ( .A(\imm[9] ), .B(\rs1[9] ), .Y(_abc_4513_n1050) );
  OR2X2 OR2X2_214 ( .A(_abc_4513_n1049), .B(_abc_4513_n1053), .Y(_abc_4513_n1054) );
  OR2X2 OR2X2_215 ( .A(_abc_4513_n1048), .B(_abc_4513_n1055), .Y(_abc_4513_n1056) );
  OR2X2 OR2X2_216 ( .A(_abc_4513_n1057), .B(\W_R[1] ), .Y(_abc_4513_n1058) );
  OR2X2 OR2X2_217 ( .A(_abc_4513_n769_1), .B(\pc[9] ), .Y(_abc_4513_n1059) );
  OR2X2 OR2X2_218 ( .A(_abc_4513_n1038), .B(_abc_4513_n1051), .Y(_abc_4513_n1062) );
  OR2X2 OR2X2_219 ( .A(_abc_4513_n1065), .B(_abc_4513_n1063), .Y(_abc_4513_n1066) );
  OR2X2 OR2X2_22 ( .A(_abc_4513_n381_1), .B(state_4_), .Y(_abc_4513_n449) );
  OR2X2 OR2X2_220 ( .A(\imm[10] ), .B(\rs1[10] ), .Y(_abc_4513_n1069) );
  OR2X2 OR2X2_221 ( .A(_abc_4513_n1066), .B(_abc_4513_n1070), .Y(_abc_4513_n1071) );
  OR2X2 OR2X2_222 ( .A(_abc_4513_n1075), .B(_abc_4513_n1061), .Y(\AWdata[10] ) );
  OR2X2 OR2X2_223 ( .A(\imm[11] ), .B(\rs1[11] ), .Y(_abc_4513_n1078) );
  OR2X2 OR2X2_224 ( .A(_abc_4513_n1077), .B(_abc_4513_n1082), .Y(_abc_4513_n1083) );
  OR2X2 OR2X2_225 ( .A(_abc_4513_n1084), .B(_abc_4513_n1081), .Y(_abc_4513_n1085) );
  OR2X2 OR2X2_226 ( .A(_abc_4513_n1086), .B(\W_R[1] ), .Y(_abc_4513_n1087) );
  OR2X2 OR2X2_227 ( .A(_abc_4513_n769_1), .B(\pc[11] ), .Y(_abc_4513_n1088) );
  OR2X2 OR2X2_228 ( .A(_abc_4513_n1093), .B(_abc_4513_n1079), .Y(_abc_4513_n1094) );
  OR2X2 OR2X2_229 ( .A(_abc_4513_n1092), .B(_abc_4513_n1094), .Y(_abc_4513_n1095) );
  OR2X2 OR2X2_23 ( .A(_abc_4513_n414_1), .B(_abc_4513_n452), .Y(_abc_4513_n453) );
  OR2X2 OR2X2_230 ( .A(_abc_4513_n1097), .B(_abc_4513_n1095), .Y(_abc_4513_n1098) );
  OR2X2 OR2X2_231 ( .A(\imm[12] ), .B(\rs1[12] ), .Y(_abc_4513_n1099) );
  OR2X2 OR2X2_232 ( .A(_abc_4513_n1098), .B(_abc_4513_n1102), .Y(_abc_4513_n1103) );
  OR2X2 OR2X2_233 ( .A(_abc_4513_n1107), .B(_abc_4513_n1090), .Y(\AWdata[12] ) );
  OR2X2 OR2X2_234 ( .A(\imm[13] ), .B(\rs1[13] ), .Y(_abc_4513_n1111) );
  OR2X2 OR2X2_235 ( .A(_abc_4513_n1110), .B(_abc_4513_n1114), .Y(_abc_4513_n1115) );
  OR2X2 OR2X2_236 ( .A(_abc_4513_n1109), .B(_abc_4513_n1116), .Y(_abc_4513_n1117) );
  OR2X2 OR2X2_237 ( .A(_abc_4513_n1118), .B(\W_R[1] ), .Y(_abc_4513_n1119) );
  OR2X2 OR2X2_238 ( .A(_abc_4513_n769_1), .B(\pc[13] ), .Y(_abc_4513_n1120) );
  OR2X2 OR2X2_239 ( .A(_abc_4513_n1116), .B(_abc_4513_n1101), .Y(_abc_4513_n1123) );
  OR2X2 OR2X2_24 ( .A(_abc_4513_n371_1), .B(_abc_4513_n388), .Y(_abc_4513_n454_1) );
  OR2X2 OR2X2_240 ( .A(_abc_4513_n1127), .B(_abc_4513_n1125), .Y(_abc_4513_n1128) );
  OR2X2 OR2X2_241 ( .A(\imm[14] ), .B(\rs1[14] ), .Y(_abc_4513_n1131) );
  OR2X2 OR2X2_242 ( .A(_abc_4513_n1128), .B(_abc_4513_n1132), .Y(_abc_4513_n1133) );
  OR2X2 OR2X2_243 ( .A(_abc_4513_n1137), .B(_abc_4513_n1122), .Y(\AWdata[14] ) );
  OR2X2 OR2X2_244 ( .A(_abc_4513_n769_1), .B(\pc[15] ), .Y(_abc_4513_n1139) );
  OR2X2 OR2X2_245 ( .A(\imm[15] ), .B(\rs1[15] ), .Y(_abc_4513_n1141) );
  OR2X2 OR2X2_246 ( .A(_abc_4513_n1140), .B(_abc_4513_n1145), .Y(_abc_4513_n1146) );
  OR2X2 OR2X2_247 ( .A(_abc_4513_n1147), .B(_abc_4513_n1144), .Y(_abc_4513_n1148) );
  OR2X2 OR2X2_248 ( .A(_abc_4513_n1149), .B(\W_R[1] ), .Y(_abc_4513_n1150) );
  OR2X2 OR2X2_249 ( .A(_abc_4513_n1159), .B(_abc_4513_n1142), .Y(_abc_4513_n1160) );
  OR2X2 OR2X2_25 ( .A(_abc_4513_n454_1), .B(_abc_4513_n428), .Y(_abc_4513_n455) );
  OR2X2 OR2X2_250 ( .A(_abc_4513_n1158), .B(_abc_4513_n1160), .Y(_abc_4513_n1161) );
  OR2X2 OR2X2_251 ( .A(_abc_4513_n1161), .B(_abc_4513_n1157), .Y(_abc_4513_n1162) );
  OR2X2 OR2X2_252 ( .A(_abc_4513_n1156), .B(_abc_4513_n1162), .Y(_abc_4513_n1163) );
  OR2X2 OR2X2_253 ( .A(\imm[16] ), .B(\rs1[16] ), .Y(_abc_4513_n1166) );
  OR2X2 OR2X2_254 ( .A(_abc_4513_n1163), .B(_abc_4513_n1167), .Y(_abc_4513_n1168) );
  OR2X2 OR2X2_255 ( .A(_abc_4513_n1172), .B(_abc_4513_n1152), .Y(\AWdata[16] ) );
  OR2X2 OR2X2_256 ( .A(\imm[17] ), .B(\rs1[17] ), .Y(_abc_4513_n1178) );
  OR2X2 OR2X2_257 ( .A(_abc_4513_n1175), .B(_abc_4513_n1179), .Y(_abc_4513_n1180) );
  OR2X2 OR2X2_258 ( .A(_abc_4513_n1174), .B(_abc_4513_n1181), .Y(_abc_4513_n1182) );
  OR2X2 OR2X2_259 ( .A(_abc_4513_n1183), .B(\W_R[1] ), .Y(_abc_4513_n1184) );
  OR2X2 OR2X2_26 ( .A(state_2_), .B(state_5_), .Y(_abc_4513_n461) );
  OR2X2 OR2X2_260 ( .A(_abc_4513_n769_1), .B(\pc[17] ), .Y(_abc_4513_n1185) );
  OR2X2 OR2X2_261 ( .A(_abc_4513_n1181), .B(_abc_4513_n1165), .Y(_abc_4513_n1188) );
  OR2X2 OR2X2_262 ( .A(_abc_4513_n1192), .B(_abc_4513_n1190), .Y(_abc_4513_n1193) );
  OR2X2 OR2X2_263 ( .A(\imm[18] ), .B(\rs1[18] ), .Y(_abc_4513_n1196) );
  OR2X2 OR2X2_264 ( .A(_abc_4513_n1193), .B(_abc_4513_n1197), .Y(_abc_4513_n1198) );
  OR2X2 OR2X2_265 ( .A(_abc_4513_n1202), .B(_abc_4513_n1187), .Y(\AWdata[18] ) );
  OR2X2 OR2X2_266 ( .A(_abc_4513_n769_1), .B(\pc[19] ), .Y(_abc_4513_n1204) );
  OR2X2 OR2X2_267 ( .A(\imm[19] ), .B(\rs1[19] ), .Y(_abc_4513_n1208) );
  OR2X2 OR2X2_268 ( .A(_abc_4513_n1205), .B(_abc_4513_n1210), .Y(_abc_4513_n1211) );
  OR2X2 OR2X2_269 ( .A(_abc_4513_n1212), .B(_abc_4513_n1209), .Y(_abc_4513_n1213) );
  OR2X2 OR2X2_27 ( .A(_abc_4513_n461), .B(state_0_), .Y(_abc_4513_n462_1) );
  OR2X2 OR2X2_270 ( .A(_abc_4513_n1214), .B(\W_R[1] ), .Y(_abc_4513_n1215) );
  OR2X2 OR2X2_271 ( .A(_abc_4513_n1220), .B(_abc_4513_n1206), .Y(_abc_4513_n1221) );
  OR2X2 OR2X2_272 ( .A(_abc_4513_n1219), .B(_abc_4513_n1221), .Y(_abc_4513_n1222) );
  OR2X2 OR2X2_273 ( .A(_abc_4513_n1224), .B(_abc_4513_n1222), .Y(_abc_4513_n1225) );
  OR2X2 OR2X2_274 ( .A(\imm[20] ), .B(\rs1[20] ), .Y(_abc_4513_n1228) );
  OR2X2 OR2X2_275 ( .A(_abc_4513_n1225), .B(_abc_4513_n1229), .Y(_abc_4513_n1230) );
  OR2X2 OR2X2_276 ( .A(_abc_4513_n1231), .B(_abc_4513_n1232), .Y(_abc_4513_n1233) );
  OR2X2 OR2X2_277 ( .A(_abc_4513_n1235), .B(_abc_4513_n1217), .Y(\AWdata[20] ) );
  OR2X2 OR2X2_278 ( .A(\imm[21] ), .B(\rs1[21] ), .Y(_abc_4513_n1240) );
  OR2X2 OR2X2_279 ( .A(_abc_4513_n1237), .B(_abc_4513_n1242), .Y(_abc_4513_n1243) );
  OR2X2 OR2X2_28 ( .A(state_4_), .B(state_3_), .Y(_abc_4513_n463) );
  OR2X2 OR2X2_280 ( .A(_abc_4513_n1244), .B(_abc_4513_n1241), .Y(_abc_4513_n1245) );
  OR2X2 OR2X2_281 ( .A(_abc_4513_n1246), .B(\W_R[1] ), .Y(_abc_4513_n1247) );
  OR2X2 OR2X2_282 ( .A(_abc_4513_n769_1), .B(\pc[21] ), .Y(_abc_4513_n1248) );
  OR2X2 OR2X2_283 ( .A(_abc_4513_n1242), .B(_abc_4513_n1227), .Y(_abc_4513_n1251) );
  OR2X2 OR2X2_284 ( .A(_abc_4513_n1255), .B(_abc_4513_n1253), .Y(_abc_4513_n1256) );
  OR2X2 OR2X2_285 ( .A(\imm[22] ), .B(\rs1[22] ), .Y(_abc_4513_n1259) );
  OR2X2 OR2X2_286 ( .A(_abc_4513_n1256), .B(_abc_4513_n1260), .Y(_abc_4513_n1261) );
  OR2X2 OR2X2_287 ( .A(_abc_4513_n1265), .B(_abc_4513_n1250), .Y(\AWdata[22] ) );
  OR2X2 OR2X2_288 ( .A(_abc_4513_n769_1), .B(\pc[23] ), .Y(_abc_4513_n1267) );
  OR2X2 OR2X2_289 ( .A(\imm[23] ), .B(\rs1[23] ), .Y(_abc_4513_n1271) );
  OR2X2 OR2X2_29 ( .A(state_6_), .B(state_1_), .Y(_abc_4513_n464) );
  OR2X2 OR2X2_290 ( .A(_abc_4513_n1268), .B(_abc_4513_n1273), .Y(_abc_4513_n1274) );
  OR2X2 OR2X2_291 ( .A(_abc_4513_n1275), .B(_abc_4513_n1272), .Y(_abc_4513_n1276) );
  OR2X2 OR2X2_292 ( .A(_abc_4513_n1277), .B(\W_R[1] ), .Y(_abc_4513_n1278) );
  OR2X2 OR2X2_293 ( .A(_abc_4513_n1287), .B(_abc_4513_n1269), .Y(_abc_4513_n1288) );
  OR2X2 OR2X2_294 ( .A(_abc_4513_n1286), .B(_abc_4513_n1288), .Y(_abc_4513_n1289) );
  OR2X2 OR2X2_295 ( .A(_abc_4513_n1285), .B(_abc_4513_n1289), .Y(_abc_4513_n1290) );
  OR2X2 OR2X2_296 ( .A(_abc_4513_n1284), .B(_abc_4513_n1290), .Y(_abc_4513_n1291) );
  OR2X2 OR2X2_297 ( .A(\imm[24] ), .B(\rs1[24] ), .Y(_abc_4513_n1294) );
  OR2X2 OR2X2_298 ( .A(_abc_4513_n1291), .B(_abc_4513_n1295), .Y(_abc_4513_n1296) );
  OR2X2 OR2X2_299 ( .A(_abc_4513_n1300), .B(_abc_4513_n1280), .Y(\AWdata[24] ) );
  OR2X2 OR2X2_3 ( .A(_abc_4513_n373), .B(_abc_4513_n371_1), .Y(_abc_4513_n374_1) );
  OR2X2 OR2X2_30 ( .A(_abc_4513_n463), .B(_abc_4513_n464), .Y(_abc_4513_n465) );
  OR2X2 OR2X2_300 ( .A(\imm[25] ), .B(\rs1[25] ), .Y(_abc_4513_n1306) );
  OR2X2 OR2X2_301 ( .A(_abc_4513_n1303), .B(_abc_4513_n1307), .Y(_abc_4513_n1308) );
  OR2X2 OR2X2_302 ( .A(_abc_4513_n1302), .B(_abc_4513_n1309), .Y(_abc_4513_n1310) );
  OR2X2 OR2X2_303 ( .A(_abc_4513_n1311), .B(\W_R[1] ), .Y(_abc_4513_n1312) );
  OR2X2 OR2X2_304 ( .A(_abc_4513_n769_1), .B(\pc[25] ), .Y(_abc_4513_n1313) );
  OR2X2 OR2X2_305 ( .A(_abc_4513_n1309), .B(_abc_4513_n1293), .Y(_abc_4513_n1316) );
  OR2X2 OR2X2_306 ( .A(_abc_4513_n1320), .B(_abc_4513_n1318), .Y(_abc_4513_n1321) );
  OR2X2 OR2X2_307 ( .A(\imm[26] ), .B(\rs1[26] ), .Y(_abc_4513_n1324) );
  OR2X2 OR2X2_308 ( .A(_abc_4513_n1321), .B(_abc_4513_n1325), .Y(_abc_4513_n1326) );
  OR2X2 OR2X2_309 ( .A(_abc_4513_n1330), .B(_abc_4513_n1315), .Y(\AWdata[26] ) );
  OR2X2 OR2X2_31 ( .A(_abc_4513_n465), .B(_abc_4513_n462_1), .Y(_abc_4513_n466) );
  OR2X2 OR2X2_310 ( .A(_abc_4513_n769_1), .B(\pc[27] ), .Y(_abc_4513_n1332) );
  OR2X2 OR2X2_311 ( .A(\imm[27] ), .B(\rs1[27] ), .Y(_abc_4513_n1334) );
  OR2X2 OR2X2_312 ( .A(_abc_4513_n1333), .B(_abc_4513_n1338), .Y(_abc_4513_n1339) );
  OR2X2 OR2X2_313 ( .A(_abc_4513_n1340), .B(_abc_4513_n1337), .Y(_abc_4513_n1341) );
  OR2X2 OR2X2_314 ( .A(_abc_4513_n1342), .B(\W_R[1] ), .Y(_abc_4513_n1343) );
  OR2X2 OR2X2_315 ( .A(_abc_4513_n1350), .B(_abc_4513_n1335), .Y(_abc_4513_n1351) );
  OR2X2 OR2X2_316 ( .A(_abc_4513_n1349), .B(_abc_4513_n1351), .Y(_abc_4513_n1352) );
  OR2X2 OR2X2_317 ( .A(_abc_4513_n1348), .B(_abc_4513_n1352), .Y(_abc_4513_n1353) );
  OR2X2 OR2X2_318 ( .A(\imm[28] ), .B(\rs1[28] ), .Y(_abc_4513_n1354) );
  OR2X2 OR2X2_319 ( .A(_abc_4513_n1353), .B(_abc_4513_n1357), .Y(_abc_4513_n1358) );
  OR2X2 OR2X2_32 ( .A(\imm[1] ), .B(\rs1[1] ), .Y(_abc_4513_n478_1) );
  OR2X2 OR2X2_320 ( .A(_abc_4513_n1362), .B(_abc_4513_n1345), .Y(\AWdata[28] ) );
  OR2X2 OR2X2_321 ( .A(\imm[29] ), .B(\rs1[29] ), .Y(_abc_4513_n1366) );
  OR2X2 OR2X2_322 ( .A(_abc_4513_n1365), .B(_abc_4513_n1369), .Y(_abc_4513_n1370) );
  OR2X2 OR2X2_323 ( .A(_abc_4513_n1364), .B(_abc_4513_n1371), .Y(_abc_4513_n1372) );
  OR2X2 OR2X2_324 ( .A(_abc_4513_n1373), .B(\W_R[1] ), .Y(_abc_4513_n1374) );
  OR2X2 OR2X2_325 ( .A(_abc_4513_n769_1), .B(\pc[29] ), .Y(_abc_4513_n1375) );
  OR2X2 OR2X2_326 ( .A(_abc_4513_n1380), .B(_abc_4513_n1367), .Y(_abc_4513_n1381) );
  OR2X2 OR2X2_327 ( .A(_abc_4513_n1379), .B(_abc_4513_n1381), .Y(_abc_4513_n1382) );
  OR2X2 OR2X2_328 ( .A(\imm[30] ), .B(\rs1[30] ), .Y(_abc_4513_n1383) );
  OR2X2 OR2X2_329 ( .A(_abc_4513_n1382), .B(_abc_4513_n1386), .Y(_abc_4513_n1387) );
  OR2X2 OR2X2_33 ( .A(_abc_4513_n486_1), .B(_abc_4513_n479), .Y(_abc_4513_n487) );
  OR2X2 OR2X2_330 ( .A(_abc_4513_n487), .B(_abc_4513_n483), .Y(_abc_4513_n1388) );
  OR2X2 OR2X2_331 ( .A(_abc_4513_n1389), .B(_abc_4513_n1390), .Y(_abc_4513_n1391) );
  OR2X2 OR2X2_332 ( .A(_abc_4513_n1393), .B(_abc_4513_n1394), .Y(_abc_4513_n1395) );
  OR2X2 OR2X2_333 ( .A(_abc_4513_n1397), .B(_abc_4513_n1398), .Y(_abc_4513_n1399) );
  OR2X2 OR2X2_334 ( .A(_abc_4513_n1401), .B(_abc_4513_n1402), .Y(_abc_4513_n1403) );
  OR2X2 OR2X2_335 ( .A(_abc_4513_n1405), .B(_abc_4513_n1406), .Y(_abc_4513_n1407) );
  OR2X2 OR2X2_336 ( .A(_abc_4513_n1409), .B(_abc_4513_n1410), .Y(_abc_4513_n1411) );
  OR2X2 OR2X2_337 ( .A(_abc_4513_n1413), .B(_abc_4513_n1414), .Y(_abc_4513_n1415) );
  OR2X2 OR2X2_338 ( .A(_abc_4513_n1417), .B(_abc_4513_n1377), .Y(\AWdata[30] ) );
  OR2X2 OR2X2_339 ( .A(_abc_4513_n1419), .B(_abc_4513_n1384), .Y(_abc_4513_n1420) );
  OR2X2 OR2X2_34 ( .A(_abc_4513_n488), .B(_abc_4513_n482), .Y(_abc_4513_n489) );
  OR2X2 OR2X2_340 ( .A(_abc_4513_n1421), .B(\rs1[31] ), .Y(_abc_4513_n1422) );
  OR2X2 OR2X2_341 ( .A(_abc_4513_n1423), .B(\imm[31] ), .Y(_abc_4513_n1424) );
  OR2X2 OR2X2_342 ( .A(_abc_4513_n1420), .B(_abc_4513_n1426), .Y(_abc_4513_n1427) );
  OR2X2 OR2X2_343 ( .A(_abc_4513_n1428), .B(_abc_4513_n1425), .Y(_abc_4513_n1429) );
  OR2X2 OR2X2_344 ( .A(_abc_4513_n1430), .B(\W_R[1] ), .Y(_abc_4513_n1431) );
  OR2X2 OR2X2_345 ( .A(_abc_4513_n769_1), .B(\pc[31] ), .Y(_abc_4513_n1432) );
  OR2X2 OR2X2_346 ( .A(_abc_4513_n381_1), .B(_abc_4513_n465), .Y(_abc_4513_n1435) );
  OR2X2 OR2X2_347 ( .A(_abc_4513_n381_1), .B(_abc_4513_n463), .Y(_abc_4513_n1437) );
  OR2X2 OR2X2_348 ( .A(_abc_4513_n449), .B(state_6_), .Y(_abc_4513_n1439) );
  OR2X2 OR2X2_349 ( .A(_abc_4513_n364), .B(_abc_4513_n461), .Y(_abc_4513_n1441) );
  OR2X2 OR2X2_35 ( .A(\imm[0] ), .B(\rs1[0] ), .Y(_abc_4513_n490) );
  OR2X2 OR2X2_36 ( .A(_abc_4513_n497), .B(_abc_4513_n495_1), .Y(_abc_4513_n498) );
  OR2X2 OR2X2_37 ( .A(_abc_4513_n498), .B(_abc_4513_n494_1), .Y(_abc_4513_n499) );
  OR2X2 OR2X2_38 ( .A(_abc_4513_n498), .B(_abc_4513_n502), .Y(_abc_4513_n503) );
  OR2X2 OR2X2_39 ( .A(_abc_4513_n506), .B(_abc_4513_n495_1), .Y(_abc_4513_n507_1) );
  OR2X2 OR2X2_4 ( .A(_abc_4513_n374_1), .B(_abc_4513_n370_1), .Y(_abc_4513_n375_1) );
  OR2X2 OR2X2_40 ( .A(_abc_4513_n507_1), .B(_abc_4513_n509), .Y(_abc_4513_n510_1) );
  OR2X2 OR2X2_41 ( .A(_abc_4513_n507_1), .B(_abc_4513_n513_1), .Y(_abc_4513_n514) );
  OR2X2 OR2X2_42 ( .A(_abc_4513_n410_1), .B(_abc_4513_n413_1), .Y(_abc_4513_n517) );
  OR2X2 OR2X2_43 ( .A(_abc_4513_n522_1), .B(_abc_4513_n520), .Y(_abc_4513_n523) );
  OR2X2 OR2X2_44 ( .A(_abc_4513_n526), .B(_abc_4513_n525_1), .Y(_abc_4513_n527) );
  OR2X2 OR2X2_45 ( .A(_abc_4513_n530), .B(_abc_4513_n529), .Y(_abc_4513_n531) );
  OR2X2 OR2X2_46 ( .A(_abc_4513_n534), .B(_abc_4513_n533_1), .Y(_abc_4513_n535_1) );
  OR2X2 OR2X2_47 ( .A(_abc_4513_n538), .B(_abc_4513_n537_1), .Y(_abc_4513_n539_1) );
  OR2X2 OR2X2_48 ( .A(_abc_4513_n542), .B(_abc_4513_n541_1), .Y(_abc_4513_n543_1) );
  OR2X2 OR2X2_49 ( .A(_abc_4513_n546), .B(_abc_4513_n545_1), .Y(_abc_4513_n547_1) );
  OR2X2 OR2X2_5 ( .A(_abc_4513_n383_1), .B(_abc_4513_n378_1), .Y(_abc_4513_n384_1) );
  OR2X2 OR2X2_50 ( .A(_abc_4513_n550), .B(_abc_4513_n549_1), .Y(_abc_4513_n551_1) );
  OR2X2 OR2X2_51 ( .A(_abc_4513_n554), .B(_abc_4513_n553_1), .Y(_abc_4513_n555_1) );
  OR2X2 OR2X2_52 ( .A(_abc_4513_n558), .B(_abc_4513_n557_1), .Y(_abc_4513_n559_1) );
  OR2X2 OR2X2_53 ( .A(_abc_4513_n562), .B(_abc_4513_n561_1), .Y(_abc_4513_n563_1) );
  OR2X2 OR2X2_54 ( .A(_abc_4513_n566_1), .B(_abc_4513_n565_1), .Y(_abc_4513_n567_1) );
  OR2X2 OR2X2_55 ( .A(_abc_4513_n570), .B(_abc_4513_n569_1), .Y(_abc_4513_n571) );
  OR2X2 OR2X2_56 ( .A(_abc_4513_n574_1), .B(_abc_4513_n573), .Y(_abc_4513_n575_1) );
  OR2X2 OR2X2_57 ( .A(_abc_4513_n578), .B(_abc_4513_n577_1), .Y(_abc_4513_n579) );
  OR2X2 OR2X2_58 ( .A(_abc_4513_n582), .B(_abc_4513_n581), .Y(_abc_4513_n583_1) );
  OR2X2 OR2X2_59 ( .A(_abc_4513_n586_1), .B(_abc_4513_n585_1), .Y(_abc_4513_n587) );
  OR2X2 OR2X2_6 ( .A(_abc_4513_n385), .B(_abc_4513_n376), .Y(_abc_3815_n23) );
  OR2X2 OR2X2_60 ( .A(_abc_4513_n590), .B(_abc_4513_n589), .Y(_abc_4513_n591) );
  OR2X2 OR2X2_61 ( .A(_abc_4513_n594_1), .B(_abc_4513_n593), .Y(_abc_4513_n595_1) );
  OR2X2 OR2X2_62 ( .A(_abc_4513_n598), .B(_abc_4513_n597_1), .Y(_abc_4513_n599) );
  OR2X2 OR2X2_63 ( .A(_abc_4513_n602_1), .B(_abc_4513_n601), .Y(_abc_4513_n603_1) );
  OR2X2 OR2X2_64 ( .A(_abc_4513_n606), .B(_abc_4513_n605_1), .Y(_abc_4513_n607) );
  OR2X2 OR2X2_65 ( .A(_abc_4513_n610), .B(_abc_4513_n609), .Y(_abc_4513_n611) );
  OR2X2 OR2X2_66 ( .A(_abc_4513_n614_1), .B(_abc_4513_n613_1), .Y(_abc_4513_n615_1) );
  OR2X2 OR2X2_67 ( .A(_abc_4513_n618), .B(_abc_4513_n617), .Y(_abc_4513_n619) );
  OR2X2 OR2X2_68 ( .A(_abc_4513_n622_1), .B(_abc_4513_n621), .Y(_abc_4513_n623_1) );
  OR2X2 OR2X2_69 ( .A(_abc_4513_n626), .B(_abc_4513_n625_1), .Y(_abc_4513_n627) );
  OR2X2 OR2X2_7 ( .A(_abc_4513_n391), .B(_abc_4513_n389_1), .Y(_abc_3815_n52) );
  OR2X2 OR2X2_70 ( .A(_abc_4513_n630), .B(_abc_4513_n629), .Y(_abc_4513_n631) );
  OR2X2 OR2X2_71 ( .A(_abc_4513_n634), .B(_abc_4513_n633), .Y(_abc_4513_n635) );
  OR2X2 OR2X2_72 ( .A(_abc_4513_n638_1), .B(_abc_4513_n637_1), .Y(_abc_4513_n639_1) );
  OR2X2 OR2X2_73 ( .A(_abc_4513_n642), .B(_abc_4513_n641), .Y(_abc_4513_n643) );
  OR2X2 OR2X2_74 ( .A(_abc_4513_n646_1), .B(_abc_4513_n645_1), .Y(_abc_4513_n647_1) );
  OR2X2 OR2X2_75 ( .A(_abc_4513_n495_1), .B(_abc_4513_n496), .Y(_abc_4513_n658_1) );
  OR2X2 OR2X2_76 ( .A(_abc_4513_n659_1), .B(_abc_4513_n657_1), .Y(_abc_4513_n660_1) );
  OR2X2 OR2X2_77 ( .A(_abc_4513_n663), .B(_abc_4513_n662), .Y(_abc_4513_n664) );
  OR2X2 OR2X2_78 ( .A(_abc_4513_n667_1), .B(_abc_4513_n666_1), .Y(_abc_4513_n668_1) );
  OR2X2 OR2X2_79 ( .A(_abc_4513_n671), .B(_abc_4513_n670), .Y(_abc_4513_n672) );
  OR2X2 OR2X2_8 ( .A(_abc_4513_n404_1), .B(_abc_4513_n381_1), .Y(_abc_4513_n405_1) );
  OR2X2 OR2X2_80 ( .A(_abc_4513_n675), .B(_abc_4513_n674), .Y(_abc_4513_n676) );
  OR2X2 OR2X2_81 ( .A(_abc_4513_n679), .B(_abc_4513_n678), .Y(_abc_4513_n680_1) );
  OR2X2 OR2X2_82 ( .A(_abc_4513_n683_1), .B(_abc_4513_n682_1), .Y(_abc_4513_n684) );
  OR2X2 OR2X2_83 ( .A(_abc_4513_n687), .B(_abc_4513_n686), .Y(_abc_4513_n688_1) );
  OR2X2 OR2X2_84 ( .A(_abc_4513_n691_1), .B(_abc_4513_n690_1), .Y(_abc_4513_n692) );
  OR2X2 OR2X2_85 ( .A(_abc_4513_n695), .B(_abc_4513_n694), .Y(_abc_4513_n696) );
  OR2X2 OR2X2_86 ( .A(_abc_4513_n699_1), .B(_abc_4513_n698), .Y(_abc_4513_n700_1) );
  OR2X2 OR2X2_87 ( .A(_abc_4513_n703), .B(_abc_4513_n702_1), .Y(_abc_4513_n704) );
  OR2X2 OR2X2_88 ( .A(_abc_4513_n707), .B(_abc_4513_n706), .Y(_abc_4513_n708_1) );
  OR2X2 OR2X2_89 ( .A(_abc_4513_n711_1), .B(_abc_4513_n710_1), .Y(_abc_4513_n712) );
  OR2X2 OR2X2_9 ( .A(_abc_4513_n406), .B(state_3_), .Y(_abc_4513_n407_1) );
  OR2X2 OR2X2_90 ( .A(_abc_4513_n715), .B(_abc_4513_n714), .Y(_abc_4513_n716) );
  OR2X2 OR2X2_91 ( .A(_abc_4513_n719), .B(_abc_4513_n718), .Y(_abc_4513_n720) );
  OR2X2 OR2X2_92 ( .A(_abc_4513_n657_1), .B(_abc_4513_n722), .Y(_abc_4513_n723) );
  OR2X2 OR2X2_93 ( .A(_abc_4513_n723), .B(_abc_4513_n724), .Y(_abc_4513_n725) );
  OR2X2 OR2X2_94 ( .A(_abc_4513_n662), .B(_abc_4513_n727_1), .Y(_abc_4513_n728_1) );
  OR2X2 OR2X2_95 ( .A(_abc_4513_n728_1), .B(_abc_4513_n729_1), .Y(_abc_4513_n730) );
  OR2X2 OR2X2_96 ( .A(_abc_4513_n666_1), .B(_abc_4513_n732), .Y(_abc_4513_n733) );
  OR2X2 OR2X2_97 ( .A(_abc_4513_n733), .B(_abc_4513_n734), .Y(_abc_4513_n735_1) );
  OR2X2 OR2X2_98 ( .A(_abc_4513_n670), .B(_abc_4513_n737_1), .Y(_abc_4513_n738_1) );
  OR2X2 OR2X2_99 ( .A(_abc_4513_n738_1), .B(_abc_4513_n739), .Y(_abc_4513_n740) );
endmodule
