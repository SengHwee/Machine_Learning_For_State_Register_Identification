module altor32_lite(clk_i, rst_i, intr_i, nmi_i, enable_i, \mem_dat_i[0] , \mem_dat_i[1] , \mem_dat_i[2] , \mem_dat_i[3] , \mem_dat_i[4] , \mem_dat_i[5] , \mem_dat_i[6] , \mem_dat_i[7] , \mem_dat_i[8] , \mem_dat_i[9] , \mem_dat_i[10] , \mem_dat_i[11] , \mem_dat_i[12] , \mem_dat_i[13] , \mem_dat_i[14] , \mem_dat_i[15] , \mem_dat_i[16] , \mem_dat_i[17] , \mem_dat_i[18] , \mem_dat_i[19] , \mem_dat_i[20] , \mem_dat_i[21] , \mem_dat_i[22] , \mem_dat_i[23] , \mem_dat_i[24] , \mem_dat_i[25] , \mem_dat_i[26] , \mem_dat_i[27] , \mem_dat_i[28] , \mem_dat_i[29] , \mem_dat_i[30] , \mem_dat_i[31] , mem_stall_i, mem_ack_i, fault_o, break_o, \mem_addr_o[0] , \mem_addr_o[1] , \mem_addr_o[2] , \mem_addr_o[3] , \mem_addr_o[4] , \mem_addr_o[5] , \mem_addr_o[6] , \mem_addr_o[7] , \mem_addr_o[8] , \mem_addr_o[9] , \mem_addr_o[10] , \mem_addr_o[11] , \mem_addr_o[12] , \mem_addr_o[13] , \mem_addr_o[14] , \mem_addr_o[15] , \mem_addr_o[16] , \mem_addr_o[17] , \mem_addr_o[18] , \mem_addr_o[19] , \mem_addr_o[20] , \mem_addr_o[21] , \mem_addr_o[22] , \mem_addr_o[23] , \mem_addr_o[24] , \mem_addr_o[25] , \mem_addr_o[26] , \mem_addr_o[27] , \mem_addr_o[28] , \mem_addr_o[29] , \mem_addr_o[30] , \mem_addr_o[31] , \mem_dat_o[0] , \mem_dat_o[1] , \mem_dat_o[2] , \mem_dat_o[3] , \mem_dat_o[4] , \mem_dat_o[5] , \mem_dat_o[6] , \mem_dat_o[7] , \mem_dat_o[8] , \mem_dat_o[9] , \mem_dat_o[10] , \mem_dat_o[11] , \mem_dat_o[12] , \mem_dat_o[13] , \mem_dat_o[14] , \mem_dat_o[15] , \mem_dat_o[16] , \mem_dat_o[17] , \mem_dat_o[18] , \mem_dat_o[19] , \mem_dat_o[20] , \mem_dat_o[21] , \mem_dat_o[22] , \mem_dat_o[23] , \mem_dat_o[24] , \mem_dat_o[25] , \mem_dat_o[26] , \mem_dat_o[27] , \mem_dat_o[28] , \mem_dat_o[29] , \mem_dat_o[30] , \mem_dat_o[31] , \mem_cti_o[0] , \mem_cti_o[1] , \mem_cti_o[2] , mem_cyc_o, mem_stb_o, mem_we_o, \mem_sel_o[0] , \mem_sel_o[1] , \mem_sel_o[2] , \mem_sel_o[3] );

wire REGFILE_SIM_reg_bank__0reg_r10_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__9_; 
wire REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2099_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2100_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2101_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2102_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2103_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2104_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2105_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2106_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2108_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2109_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2111_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2112_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2114_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2115_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2117_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2118_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2120_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2121_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2123_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2124_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2126_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2127_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2129_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2130_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2132_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2133_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2135_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2136_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2138_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2139_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2141_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2142_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2144_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2145_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2147_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2148_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2150_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2151_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2153_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2154_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2156_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2157_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2159_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2160_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2162_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2163_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2165_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2166_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2168_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2169_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2171_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2172_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2174_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2175_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2177_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2178_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2180_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2181_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2183_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2184_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2186_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2187_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2189_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2190_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2192_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2193_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2195_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2196_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2198_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2199_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2201_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2202_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2203_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2204_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2205_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2207_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2209_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2211_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2213_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2215_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2217_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2219_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2221_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2223_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2225_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2227_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2229_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2231_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2233_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2235_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2237_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2239_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2241_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2243_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2245_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2247_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2249_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2251_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2253_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2255_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2257_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2259_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2261_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2263_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2265_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2267_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2269_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2270_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2271_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2272_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2274_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2276_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2278_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2280_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2282_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2284_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2286_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2288_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2290_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2292_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2294_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2296_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2298_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2300_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2302_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2304_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2306_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2308_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2310_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2312_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2314_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2316_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2318_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2320_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2322_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2324_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2326_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2328_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2330_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2332_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2334_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2336_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2337_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2338_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2339_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2341_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2343_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2345_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2347_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2349_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2351_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2353_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2355_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2357_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2359_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2361_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2363_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2365_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2367_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2369_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2371_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2373_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2375_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2377_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2379_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2381_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2383_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2385_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2387_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2389_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2391_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2393_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2395_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2397_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2399_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2401_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2403_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2404_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2405_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2406_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2407_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2409_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2411_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2413_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2415_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2417_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2419_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2421_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2423_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2425_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2427_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2429_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2431_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2433_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2435_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2437_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2439_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2441_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2443_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2445_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2447_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2449_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2451_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2453_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2455_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2457_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2459_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2461_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2463_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2465_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2467_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2469_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2471_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2472_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2473_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2475_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2477_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2479_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2481_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2483_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2485_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2487_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2489_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2491_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2493_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2495_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2497_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2499_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2501_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2503_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2505_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2507_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2509_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2511_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2513_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2515_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2517_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2519_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2521_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2523_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2525_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2527_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2529_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2531_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2533_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2535_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2537_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2538_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2539_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2541_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2543_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2545_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2547_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2549_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2551_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2553_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2555_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2557_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2559_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2561_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2563_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2565_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2567_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2569_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2571_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2573_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2575_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2577_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2579_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2581_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2583_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2585_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2587_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2589_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2591_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2593_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2595_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2597_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2599_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2601_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2603_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2604_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2606_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2608_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2610_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2612_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2614_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2616_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2618_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2620_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2622_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2624_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2626_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2628_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2630_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2632_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2634_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2636_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2638_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2640_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2642_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2644_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2646_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2648_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2650_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2652_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2654_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2656_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2658_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2660_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2662_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2664_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2666_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2668_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2669_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2670_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2671_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2673_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2675_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2677_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2679_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2681_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2683_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2685_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2687_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2689_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2691_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2693_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2695_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2697_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2699_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2701_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2703_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2705_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2707_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2709_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2711_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2713_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2715_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2717_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2719_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2721_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2723_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2725_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2727_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2729_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2731_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2733_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2735_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2736_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2737_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2739_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2741_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2743_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2745_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2747_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2749_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2751_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2753_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2755_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2757_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2759_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2761_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2763_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2765_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2767_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2769_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2771_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2773_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2775_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2777_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2779_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2781_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2783_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2785_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2787_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2789_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2791_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2793_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2795_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2797_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2799_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2801_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2802_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2803_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2805_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2807_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2809_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2811_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2813_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2815_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2817_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2819_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2821_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2823_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2825_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2827_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2829_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2831_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2833_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2835_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2837_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2839_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2841_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2843_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2845_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2847_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2849_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2851_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2853_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2855_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2857_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2859_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2861_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2863_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2865_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2867_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2868_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2870_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2872_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2874_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2876_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2878_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2880_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2882_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2884_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2886_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2888_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2890_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2892_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2894_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2896_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2898_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2900_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2902_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2904_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2906_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2908_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2910_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2912_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2914_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2916_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2918_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2920_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2922_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2924_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2926_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2928_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2930_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2932_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2933_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2934_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2935_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2936_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2938_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2940_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2942_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2944_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2946_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2948_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2950_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2952_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2954_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2956_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2958_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2960_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2962_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2964_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2966_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2968_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2970_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2972_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2974_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2976_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2978_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2980_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2982_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2984_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2986_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2988_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2990_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2992_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2994_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2996_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n2998_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3000_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3001_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3002_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3004_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3006_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3008_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3010_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3012_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3014_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3016_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3018_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3020_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3022_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3024_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3026_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3028_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3030_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3032_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3034_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3036_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3038_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3040_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3042_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3044_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3046_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3048_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3050_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3052_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3054_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3056_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3058_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3060_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3062_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3064_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3066_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3067_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3068_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3070_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3072_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3074_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3076_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3078_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3080_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3082_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3084_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3086_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3088_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3090_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3092_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3094_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3096_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3098_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3100_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3102_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3104_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3106_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3108_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3110_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3112_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3114_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3116_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3118_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3120_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3122_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3124_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3126_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3128_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3130_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3132_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3133_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3135_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3137_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3139_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3141_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3143_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3145_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3147_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3149_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3151_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3153_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3155_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3157_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3159_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3161_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3163_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3165_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3167_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3169_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3171_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3173_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3175_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3177_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3179_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3181_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3183_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3185_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3187_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3189_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3191_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3193_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3195_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3197_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3198_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3199_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3200_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3202_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3204_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3206_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3208_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3210_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3212_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3214_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3216_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3218_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3220_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3222_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3224_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3226_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3228_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3230_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3232_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3234_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3236_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3238_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3240_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3242_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3244_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3246_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3248_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3250_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3252_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3254_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3256_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3258_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3260_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3262_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3264_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3265_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3267_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3269_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3271_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3273_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3275_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3277_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3279_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3281_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3283_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3285_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3287_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3289_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3291_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3293_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3295_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3297_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3299_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3301_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3303_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3305_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3307_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3309_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3311_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3313_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3315_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3317_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3319_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3321_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3323_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3325_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3327_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3329_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3330_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3332_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3334_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3336_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3338_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3340_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3342_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3344_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3346_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3348_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3350_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3352_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3354_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3356_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3358_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3360_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3362_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3364_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3366_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3368_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3370_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3372_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3374_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3376_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3378_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3380_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3382_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3384_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3386_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3388_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3390_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3392_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3394_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3395_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3396_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3398_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3400_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3402_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3404_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3406_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3408_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3410_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3412_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3414_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3416_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3418_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3420_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3422_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3424_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3426_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3428_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3430_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3432_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3434_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3436_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3438_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3440_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3442_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3444_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3446_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3448_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3450_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3452_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3454_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3456_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3458_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3460_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3461_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3463_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3465_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3467_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3469_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3471_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3473_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3475_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3477_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3479_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3481_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3483_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3485_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3487_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3489_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3491_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3493_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3495_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3497_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3499_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3501_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3503_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3505_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3507_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3509_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3511_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3513_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3515_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3517_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3519_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3521_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3523_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3525_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3526_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3528_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3530_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3532_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3534_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3536_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3538_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3540_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3542_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3544_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3546_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3548_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3550_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3552_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3554_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3556_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3558_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3560_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3562_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3564_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3566_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3568_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3570_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3572_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3574_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3576_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3578_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3580_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3582_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3584_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3586_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3588_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3590_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3591_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3592_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3594_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3596_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3598_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3600_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3602_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3604_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3606_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3608_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3610_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3612_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3614_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3616_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3618_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3620_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3622_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3624_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3626_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3628_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3630_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3632_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3634_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3636_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3638_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3640_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3642_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3644_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3646_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3648_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3650_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3652_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3654_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3656_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3657_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3659_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3661_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3663_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3665_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3667_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3669_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3671_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3673_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3675_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3677_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3679_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3681_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3683_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3685_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3687_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3689_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3691_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3693_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3695_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3697_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3699_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3701_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3703_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3705_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3707_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3709_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3711_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3713_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3715_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3717_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3719_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3721_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3722_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3724_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3726_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3728_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3730_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3732_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3734_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3736_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3738_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3740_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3742_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3744_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3746_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3748_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3750_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3752_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3754_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3756_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3758_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3760_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3762_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3764_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3766_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3768_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3770_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3772_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3774_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3776_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3778_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3780_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3782_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3784_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3786_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3787_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3789_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3791_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3793_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3795_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3797_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3799_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3801_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3803_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3805_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3807_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3809_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3811_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3813_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3815_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3817_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3819_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3821_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3823_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3825_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3827_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3829_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3831_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3833_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3835_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3837_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3839_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3841_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3843_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3845_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3847_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3849_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3851_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3852_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3854_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3856_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3858_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3860_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3862_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3864_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3866_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3868_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3870_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3872_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3874_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3876_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3878_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3880_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3882_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3884_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3886_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3888_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3890_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3892_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3894_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3896_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3898_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3900_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3902_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3904_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3906_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3908_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3910_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3912_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3914_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3916_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3917_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3919_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3921_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3923_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3925_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3927_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3929_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3931_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3933_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3935_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3937_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3939_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3941_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3943_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3945_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3947_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3949_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3951_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3953_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3955_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3957_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3959_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3961_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3963_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3965_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3967_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3969_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3971_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3973_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3975_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3977_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3979_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3981_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3982_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3984_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3986_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3988_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3990_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3992_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3994_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3996_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n3998_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4000_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4002_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4004_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4006_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4008_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4010_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4012_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4014_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4016_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4018_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4020_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4022_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4024_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4026_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4028_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4030_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4032_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4034_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4036_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4038_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4040_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4042_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4044_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4046_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4047_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4049_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4051_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4053_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4055_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4057_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4059_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4061_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4063_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4065_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4067_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4069_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4071_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4073_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4075_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4077_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4079_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4081_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4083_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4085_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4087_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4089_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4091_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4093_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4095_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4097_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4099_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4101_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4103_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4105_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4107_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4109_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4111_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4112_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4114_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4116_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4118_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4120_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4122_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4124_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4126_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4128_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4130_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4132_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4134_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4136_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4138_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4140_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4142_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4144_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4146_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4148_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4150_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4152_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4154_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4156_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4158_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4160_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4162_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4164_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4166_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4168_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4170_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4172_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4174_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4176_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4177_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4178_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4179_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4180_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4181_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4182_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4183_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4184_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4185_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4186_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4187_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4188_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4189_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4190_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4191_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4192_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4193_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4194_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4195_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4196_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4197_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4198_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4199_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4200_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4201_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4202_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4203_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4204_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4205_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4206_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4207_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4208_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4209_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4210_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4211_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4212_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4213_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4214_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4215_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4216_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4217_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4218_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4219_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4220_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4221_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4222_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4223_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4224_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4225_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4226_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4227_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4228_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4229_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4230_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4231_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4232_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4233_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4234_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4235_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4236_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4237_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4238_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4239_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4240_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4241_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4242_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4243_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4244_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4245_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4246_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4247_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4248_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4249_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4250_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4251_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4252_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4253_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4254_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4256_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4257_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4258_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4259_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4260_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4261_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4262_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4263_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4264_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4265_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4266_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4267_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4268_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4269_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4270_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4271_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4272_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4273_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4274_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4275_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4276_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4277_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4278_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4279_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4280_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4281_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4282_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4283_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4284_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4285_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4286_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4288_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4289_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4290_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4291_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4292_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4293_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4294_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4295_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4296_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4297_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4298_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4299_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4300_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4301_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4302_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4303_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4304_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4305_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4306_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4307_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4308_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4309_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4310_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4311_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4312_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4313_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4314_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4315_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4316_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4317_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4318_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4320_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4321_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4322_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4323_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4324_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4325_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4326_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4327_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4328_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4329_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4330_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4331_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4332_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4333_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4334_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4335_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4336_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4337_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4338_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4339_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4340_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4341_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4342_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4343_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4344_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4345_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4346_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4347_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4348_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4349_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4350_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4352_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4353_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4354_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4355_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4356_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4357_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4358_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4359_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4360_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4361_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4362_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4363_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4364_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4365_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4366_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4367_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4368_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4369_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4370_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4371_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4372_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4373_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4374_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4375_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4376_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4377_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4378_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4379_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4380_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4381_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4382_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4384_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4385_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4386_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4387_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4388_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4389_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4390_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4391_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4392_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4393_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4394_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4395_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4396_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4397_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4398_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4399_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4400_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4401_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4402_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4403_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4404_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4405_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4406_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4407_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4408_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4409_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4410_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4411_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4412_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4413_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4414_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4416_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4417_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4418_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4419_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4420_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4421_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4422_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4423_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4424_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4425_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4426_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4427_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4428_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4429_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4430_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4431_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4432_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4433_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4434_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4435_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4436_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4437_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4438_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4439_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4440_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4441_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4442_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4443_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4444_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4445_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4446_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4448_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4449_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4450_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4451_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4452_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4453_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4454_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4455_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4456_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4457_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4458_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4459_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4460_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4461_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4462_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4463_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4464_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4465_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4466_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4467_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4468_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4469_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4470_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4471_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4472_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4473_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4474_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4475_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4476_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4477_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4478_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4480_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4481_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4482_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4483_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4484_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4485_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4486_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4487_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4488_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4489_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4490_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4491_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4492_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4493_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4494_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4495_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4496_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4497_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4498_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4499_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4500_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4501_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4502_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4503_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4504_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4505_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4506_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4507_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4508_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4509_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4510_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4512_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4513_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4514_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4515_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4516_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4517_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4518_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4519_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4520_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4521_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4522_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4523_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4524_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4525_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4526_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4527_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4528_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4529_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4530_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4531_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4532_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4533_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4534_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4535_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4536_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4537_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4538_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4539_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4540_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4541_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4542_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4544_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4545_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4546_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4547_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4548_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4549_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4550_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4551_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4552_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4553_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4554_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4555_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4556_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4557_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4558_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4559_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4560_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4561_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4562_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4563_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4564_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4565_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4566_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4567_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4568_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4569_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4570_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4571_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4572_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4573_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4574_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4576_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4577_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4578_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4579_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4580_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4581_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4582_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4583_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4584_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4585_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4586_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4587_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4588_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4589_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4590_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4591_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4592_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4593_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4594_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4595_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4596_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4597_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4598_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4599_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4600_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4601_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4602_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4603_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4604_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4605_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4606_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4608_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4609_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4610_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4611_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4612_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4613_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4614_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4615_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4616_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4617_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4618_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4619_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4620_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4621_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4622_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4623_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4624_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4625_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4626_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4627_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4628_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4629_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4630_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4631_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4632_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4633_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4634_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4635_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4636_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4637_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4638_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4640_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4641_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4642_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4643_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4644_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4645_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4646_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4647_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4648_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4649_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4650_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4651_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4652_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4653_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4654_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4655_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4656_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4657_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4658_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4659_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4660_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4661_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4662_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4663_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4664_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4665_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4666_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4667_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4668_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4669_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4670_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4672_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4673_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4674_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4675_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4676_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4677_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4678_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4679_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4680_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4681_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4682_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4683_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4684_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4685_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4686_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4687_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4688_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4689_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4690_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4691_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4692_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4693_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4694_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4695_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4696_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4697_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4698_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4699_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4700_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4701_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4702_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4704_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4705_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4706_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4707_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4708_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4709_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4710_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4711_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4712_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4713_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4714_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4715_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4716_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4717_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4718_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4719_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4720_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4721_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4722_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4723_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4724_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4725_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4726_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4727_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4728_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4729_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4730_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4731_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4732_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4733_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4734_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4736_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4737_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4738_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4739_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4740_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4741_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4742_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4743_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4744_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4745_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4746_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4747_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4748_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4749_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4750_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4751_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4752_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4753_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4754_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4755_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4756_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4757_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4758_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4759_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4760_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4761_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4762_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4763_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4764_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4765_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4766_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4768_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4769_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4770_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4771_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4772_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4773_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4774_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4775_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4776_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4777_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4778_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4779_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4780_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4781_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4782_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4783_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4784_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4785_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4786_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4787_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4788_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4789_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4790_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4791_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4792_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4793_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4794_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4795_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4796_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4797_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4798_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4800_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4801_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4802_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4803_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4804_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4805_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4806_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4807_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4808_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4809_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4810_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4811_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4812_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4813_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4814_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4815_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4816_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4817_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4818_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4819_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4820_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4821_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4822_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4823_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4824_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4825_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4826_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4827_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4828_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4829_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4830_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4832_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4833_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4834_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4835_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4836_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4837_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4838_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4839_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4840_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4841_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4842_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4843_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4844_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4845_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4846_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4847_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4848_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4849_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4850_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4851_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4852_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4853_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4854_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4855_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4856_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4857_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4858_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4859_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4860_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4861_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4862_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4864_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4865_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4866_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4867_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4868_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4869_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4870_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4871_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4872_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4873_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4874_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4875_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4876_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4877_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4878_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4879_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4880_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4881_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4882_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4883_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4884_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4885_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4886_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4887_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4888_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4889_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4890_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4891_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4892_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4893_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4894_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4896_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4897_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4898_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4899_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4900_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4901_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4902_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4903_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4904_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4905_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4906_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4907_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4908_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4909_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4910_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4911_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4912_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4913_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4914_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4915_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4916_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4917_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4918_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4919_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4920_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4921_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4922_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4923_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4924_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4925_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4926_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4928_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4929_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4930_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4931_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4932_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4933_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4934_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4935_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4936_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4937_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4938_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4939_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4940_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4941_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4942_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4943_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4944_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4945_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4946_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4947_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4948_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4949_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4950_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4951_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4952_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4953_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4954_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4955_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4956_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4957_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4958_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4960_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4961_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4962_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4963_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4964_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4965_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4966_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4967_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4968_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4969_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4970_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4971_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4972_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4973_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4974_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4975_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4976_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4977_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4978_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4979_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4980_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4981_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4982_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4983_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4984_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4985_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4986_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4987_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4988_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4989_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4990_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4992_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4993_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4994_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4995_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4996_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4997_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4998_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n4999_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5000_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5001_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5002_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5003_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5004_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5005_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5006_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5007_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5008_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5009_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5010_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5011_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5012_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5013_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5014_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5015_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5016_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5017_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5018_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5019_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5020_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5021_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5022_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5024_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5025_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5026_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5027_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5028_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5029_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5030_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5031_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5032_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5033_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5034_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5035_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5036_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5037_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5038_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5039_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5040_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5041_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5042_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5043_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5044_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5045_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5046_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5047_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5048_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5049_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5050_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5051_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5052_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5053_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5054_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5056_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5057_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5058_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5059_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5060_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5061_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5062_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5063_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5064_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5065_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5066_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5067_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5068_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5069_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5070_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5071_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5072_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5073_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5074_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5075_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5076_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5077_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5078_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5079_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5080_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5081_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5082_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5083_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5084_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5085_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5086_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5088_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5089_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5090_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5091_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5092_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5093_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5094_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5095_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5096_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5097_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5098_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5099_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5100_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5101_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5102_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5103_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5104_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5105_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5106_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5107_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5108_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5109_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5110_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5111_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5112_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5113_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5114_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5115_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5116_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5117_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5118_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5120_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5121_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5122_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5123_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5124_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5125_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5126_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5127_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5128_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5129_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5130_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5131_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5132_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5133_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5134_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5135_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5136_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5137_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5138_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5139_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5140_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5141_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5142_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5143_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5144_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5145_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5146_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5147_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5148_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5149_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5150_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5152_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5153_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5154_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5155_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5156_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5157_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5158_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5159_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5160_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5161_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5162_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5163_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5164_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5165_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5166_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5167_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5168_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5169_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5170_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5171_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5172_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5173_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5174_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5175_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5176_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5177_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5178_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5179_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5180_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5181_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5182_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5184_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5185_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5186_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5187_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5188_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5189_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5190_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5191_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5192_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5193_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5194_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5195_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5196_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5197_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5198_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5199_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5200_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5201_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5202_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5203_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5204_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5205_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5206_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5207_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5208_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5209_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5210_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5211_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5212_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5213_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5214_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5216_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5217_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5218_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5219_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5220_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5221_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5222_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5223_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5224_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5225_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5226_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5227_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5228_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5229_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5230_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5231_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5232_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5233_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5234_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5235_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5236_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5237_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5238_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5239_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5240_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5241_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5242_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5243_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5244_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5245_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5246_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5248_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5249_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5250_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5251_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5252_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5253_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5254_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5255_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5256_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5257_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5258_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5259_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5260_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5261_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5262_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5263_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5264_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5265_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5266_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5267_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5268_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5269_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5270_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5271_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5272_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5273_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5274_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5275_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5276_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5277_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5278_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5279_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5280_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5281_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5282_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5283_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5284_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5285_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5286_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5287_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5288_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5289_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5290_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5291_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5292_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5293_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5294_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5295_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5296_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5297_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5298_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5299_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5300_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5301_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5302_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5303_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5304_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5305_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5306_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5307_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5308_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5309_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5310_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5311_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5312_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5313_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5314_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5315_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5316_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5317_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5318_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5319_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5320_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5321_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5322_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5323_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5324_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5325_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5326_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5328_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5329_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5330_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5331_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5332_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5333_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5334_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5335_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5336_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5337_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5338_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5339_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5340_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5341_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5342_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5343_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5344_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5345_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5346_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5347_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5348_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5349_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5350_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5351_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5352_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5353_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5354_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5355_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5356_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5357_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5358_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5360_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5361_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5362_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5363_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5364_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5365_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5366_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5367_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5368_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5369_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5370_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5371_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5372_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5373_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5374_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5375_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5376_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5377_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5378_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5379_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5380_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5381_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5382_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5383_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5384_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5385_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5386_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5387_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5388_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5389_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5390_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5392_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5393_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5394_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5395_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5396_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5397_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5398_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5399_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5400_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5401_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5402_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5403_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5404_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5405_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5406_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5407_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5408_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5409_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5410_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5411_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5412_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5413_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5414_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5415_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5416_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5417_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5418_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5419_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5420_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5421_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5422_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5424_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5425_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5426_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5427_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5428_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5429_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5430_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5431_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5432_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5433_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5434_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5435_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5436_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5437_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5438_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5439_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5440_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5441_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5442_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5443_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5444_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5445_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5446_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5447_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5448_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5449_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5450_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5451_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5452_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5453_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5454_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5456_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5457_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5458_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5459_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5460_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5461_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5462_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5463_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5464_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5465_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5466_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5467_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5468_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5469_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5470_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5471_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5472_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5473_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5474_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5475_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5476_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5477_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5478_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5479_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5480_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5481_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5482_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5483_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5484_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5485_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5486_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5488_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5489_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5490_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5491_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5492_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5493_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5494_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5495_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5496_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5497_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5498_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5499_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5500_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5501_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5502_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5503_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5504_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5505_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5506_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5507_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5508_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5509_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5510_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5511_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5512_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5513_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5514_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5515_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5516_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5517_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5518_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5520_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5521_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5522_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5523_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5524_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5525_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5526_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5527_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5528_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5529_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5530_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5531_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5532_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5533_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5534_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5535_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5536_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5537_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5538_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5539_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5540_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5541_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5542_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5543_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5544_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5545_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5546_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5547_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5548_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5549_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5550_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5552_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5553_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5554_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5555_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5556_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5557_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5558_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5559_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5560_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5561_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5562_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5563_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5564_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5565_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5566_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5567_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5568_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5569_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5570_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5571_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5572_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5573_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5574_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5575_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5576_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5577_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5578_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5579_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5580_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5581_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5582_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5584_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5585_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5586_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5587_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5588_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5589_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5590_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5591_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5592_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5593_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5594_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5595_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5596_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5597_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5598_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5599_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5600_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5601_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5602_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5603_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5604_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5605_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5606_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5607_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5608_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5609_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5610_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5611_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5612_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5613_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5614_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5616_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5617_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5618_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5619_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5620_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5621_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5622_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5623_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5624_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5625_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5626_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5627_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5628_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5629_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5630_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5631_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5632_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5633_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5634_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5635_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5636_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5637_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5638_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5639_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5640_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5641_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5642_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5643_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5644_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5645_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5646_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5648_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5649_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5650_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5651_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5652_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5653_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5654_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5655_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5656_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5657_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5658_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5659_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5660_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5661_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5662_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5663_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5664_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5665_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5666_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5667_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5668_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5669_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5670_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5671_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5672_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5673_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5674_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5675_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5676_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5677_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5678_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5680_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5681_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5682_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5683_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5684_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5685_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5686_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5687_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5688_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5689_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5690_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5691_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5692_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5693_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5694_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5695_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5696_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5697_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5698_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5699_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5700_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5701_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5702_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5703_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5704_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5705_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5706_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5707_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5708_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5709_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5710_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5712_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5713_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5714_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5715_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5716_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5717_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5718_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5719_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5720_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5721_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5722_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5723_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5724_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5725_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5726_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5727_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5728_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5729_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5730_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5731_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5732_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5733_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5734_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5735_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5736_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5737_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5738_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5739_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5740_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5741_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5742_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5744_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5745_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5746_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5747_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5748_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5749_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5750_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5751_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5752_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5753_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5754_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5755_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5756_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5757_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5758_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5759_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5760_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5761_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5762_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5763_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5764_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5765_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5766_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5767_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5768_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5769_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5770_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5771_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5772_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5773_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5774_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5776_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5777_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5778_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5779_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5780_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5781_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5782_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5783_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5784_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5785_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5786_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5787_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5788_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5789_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5790_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5791_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5792_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5793_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5794_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5795_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5796_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5797_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5798_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5799_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5800_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5801_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5802_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5803_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5804_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5805_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5806_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5808_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5809_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5810_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5811_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5812_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5813_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5814_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5815_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5816_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5817_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5818_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5819_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5820_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5821_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5822_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5823_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5824_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5825_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5826_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5827_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5828_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5829_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5830_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5831_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5832_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5833_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5834_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5835_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5836_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5837_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5838_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5840_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5841_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5842_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5843_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5844_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5845_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5846_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5847_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5848_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5849_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5850_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5851_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5852_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5853_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5854_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5855_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5856_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5857_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5858_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5859_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5860_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5861_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5862_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5863_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5864_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5865_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5866_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5867_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5868_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5869_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5870_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5872_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5873_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5874_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5875_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5876_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5877_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5878_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5879_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5880_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5881_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5882_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5883_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5884_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5885_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5886_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5887_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5888_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5889_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5890_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5891_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5892_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5893_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5894_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5895_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5896_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5897_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5898_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5899_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5900_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5901_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5902_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5904_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5905_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5906_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5907_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5908_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5909_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5910_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5911_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5912_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5913_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5914_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5915_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5916_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5917_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5918_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5919_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5920_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5921_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5922_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5923_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5924_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5925_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5926_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5927_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5928_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5929_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5930_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5931_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5932_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5933_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5934_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5936_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5937_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5938_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5939_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5940_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5941_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5942_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5943_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5944_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5945_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5946_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5947_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5948_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5949_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5950_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5951_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5952_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5953_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5954_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5955_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5956_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5957_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5958_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5959_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5960_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5961_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5962_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5963_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5964_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5965_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5966_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5968_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5969_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5970_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5971_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5972_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5973_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5974_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5975_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5976_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5977_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5978_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5979_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5980_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5981_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5982_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5983_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5984_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5985_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5986_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5987_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5988_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5989_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5990_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5991_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5992_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5993_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5994_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5995_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5996_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5997_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n5998_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6000_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6001_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6002_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6003_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6004_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6005_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6006_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6007_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6008_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6009_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6010_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6011_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6012_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6013_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6014_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6015_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6016_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6017_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6018_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6019_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6020_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6021_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6022_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6023_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6024_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6025_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6026_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6027_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6028_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6029_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6030_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6032_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6033_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6034_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6035_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6036_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6037_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6038_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6039_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6040_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6041_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6042_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6043_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6044_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6045_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6046_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6047_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6048_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6049_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6050_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6051_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6052_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6053_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6054_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6055_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6056_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6057_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6058_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6059_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6060_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6061_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6062_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6064_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6065_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6066_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6067_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6068_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6069_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6070_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6071_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6072_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6073_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6074_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6075_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6076_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6077_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6078_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6079_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6080_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6081_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6082_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6083_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6084_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6085_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6086_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6087_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6088_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6089_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6090_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6091_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6092_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6093_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6094_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6096_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6097_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6098_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6099_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6100_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6101_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6102_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6103_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6104_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6105_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6106_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6107_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6108_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6109_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6110_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6111_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6112_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6113_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6114_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6115_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6116_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6117_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6118_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6119_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6120_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6121_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6122_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6123_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6124_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6125_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6126_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6128_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6129_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6130_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6131_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6132_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6133_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6134_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6135_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6136_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6137_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6138_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6139_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6140_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6141_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6142_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6143_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6144_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6145_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6146_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6147_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6148_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6149_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6150_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6151_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6152_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6153_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6154_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6155_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6156_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6157_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6158_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6160_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6161_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6162_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6163_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6164_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6165_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6166_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6167_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6168_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6169_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6170_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6171_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6172_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6173_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6174_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6175_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6176_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6177_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6178_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6179_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6180_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6181_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6182_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6183_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6184_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6185_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6186_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6187_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6188_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6189_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6190_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6192_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6193_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6194_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6195_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6196_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6197_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6198_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6199_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6200_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6201_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6202_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6203_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6204_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6205_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6206_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6207_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6208_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6209_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6210_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6211_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6212_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6213_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6214_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6215_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6216_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6217_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6218_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6219_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6220_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6221_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6222_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6224_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6225_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6226_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6227_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6228_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6229_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6230_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6231_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6232_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6233_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6234_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6235_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6236_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6237_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6238_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6239_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6240_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6241_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6242_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6243_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6244_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6245_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6246_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6247_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6248_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6249_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6250_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6251_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6252_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6253_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6254_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6256_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6257_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6258_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6259_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6260_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6261_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6262_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6263_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6264_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6265_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6266_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6267_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6268_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6269_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6270_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6271_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6272_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6273_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6274_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6275_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6276_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6277_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6278_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6279_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6280_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6281_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6282_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6283_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6284_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6285_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6286_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6288_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6289_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6290_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6291_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6292_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6293_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6294_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6295_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6296_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6297_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6298_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6299_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6300_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6301_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6302_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6303_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6304_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6305_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6306_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6307_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6308_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6309_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6310_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6311_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6312_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6313_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6314_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6315_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6316_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6317_; 
wire REGFILE_SIM_reg_bank__abc_34451_new_n6318_; 
wire REGFILE_SIM_reg_bank_ra_i_0_; 
wire REGFILE_SIM_reg_bank_ra_i_1_; 
wire REGFILE_SIM_reg_bank_ra_i_2_; 
wire REGFILE_SIM_reg_bank_ra_i_3_; 
wire REGFILE_SIM_reg_bank_ra_i_4_; 
wire REGFILE_SIM_reg_bank_rb_i_0_; 
wire REGFILE_SIM_reg_bank_rb_i_1_; 
wire REGFILE_SIM_reg_bank_rb_i_2_; 
wire REGFILE_SIM_reg_bank_rb_i_3_; 
wire REGFILE_SIM_reg_bank_rb_i_4_; 
wire REGFILE_SIM_reg_bank_rd_i_0_; 
wire REGFILE_SIM_reg_bank_rd_i_1_; 
wire REGFILE_SIM_reg_bank_rd_i_2_; 
wire REGFILE_SIM_reg_bank_rd_i_3_; 
wire REGFILE_SIM_reg_bank_rd_i_4_; 
wire REGFILE_SIM_reg_bank_reg_r10_0_; 
wire REGFILE_SIM_reg_bank_reg_r10_10_; 
wire REGFILE_SIM_reg_bank_reg_r10_11_; 
wire REGFILE_SIM_reg_bank_reg_r10_12_; 
wire REGFILE_SIM_reg_bank_reg_r10_13_; 
wire REGFILE_SIM_reg_bank_reg_r10_14_; 
wire REGFILE_SIM_reg_bank_reg_r10_15_; 
wire REGFILE_SIM_reg_bank_reg_r10_16_; 
wire REGFILE_SIM_reg_bank_reg_r10_17_; 
wire REGFILE_SIM_reg_bank_reg_r10_18_; 
wire REGFILE_SIM_reg_bank_reg_r10_19_; 
wire REGFILE_SIM_reg_bank_reg_r10_1_; 
wire REGFILE_SIM_reg_bank_reg_r10_20_; 
wire REGFILE_SIM_reg_bank_reg_r10_21_; 
wire REGFILE_SIM_reg_bank_reg_r10_22_; 
wire REGFILE_SIM_reg_bank_reg_r10_23_; 
wire REGFILE_SIM_reg_bank_reg_r10_24_; 
wire REGFILE_SIM_reg_bank_reg_r10_25_; 
wire REGFILE_SIM_reg_bank_reg_r10_26_; 
wire REGFILE_SIM_reg_bank_reg_r10_27_; 
wire REGFILE_SIM_reg_bank_reg_r10_28_; 
wire REGFILE_SIM_reg_bank_reg_r10_29_; 
wire REGFILE_SIM_reg_bank_reg_r10_2_; 
wire REGFILE_SIM_reg_bank_reg_r10_30_; 
wire REGFILE_SIM_reg_bank_reg_r10_31_; 
wire REGFILE_SIM_reg_bank_reg_r10_3_; 
wire REGFILE_SIM_reg_bank_reg_r10_4_; 
wire REGFILE_SIM_reg_bank_reg_r10_5_; 
wire REGFILE_SIM_reg_bank_reg_r10_6_; 
wire REGFILE_SIM_reg_bank_reg_r10_7_; 
wire REGFILE_SIM_reg_bank_reg_r10_8_; 
wire REGFILE_SIM_reg_bank_reg_r10_9_; 
wire REGFILE_SIM_reg_bank_reg_r11_0_; 
wire REGFILE_SIM_reg_bank_reg_r11_10_; 
wire REGFILE_SIM_reg_bank_reg_r11_11_; 
wire REGFILE_SIM_reg_bank_reg_r11_12_; 
wire REGFILE_SIM_reg_bank_reg_r11_13_; 
wire REGFILE_SIM_reg_bank_reg_r11_14_; 
wire REGFILE_SIM_reg_bank_reg_r11_15_; 
wire REGFILE_SIM_reg_bank_reg_r11_16_; 
wire REGFILE_SIM_reg_bank_reg_r11_17_; 
wire REGFILE_SIM_reg_bank_reg_r11_18_; 
wire REGFILE_SIM_reg_bank_reg_r11_19_; 
wire REGFILE_SIM_reg_bank_reg_r11_1_; 
wire REGFILE_SIM_reg_bank_reg_r11_20_; 
wire REGFILE_SIM_reg_bank_reg_r11_21_; 
wire REGFILE_SIM_reg_bank_reg_r11_22_; 
wire REGFILE_SIM_reg_bank_reg_r11_23_; 
wire REGFILE_SIM_reg_bank_reg_r11_24_; 
wire REGFILE_SIM_reg_bank_reg_r11_25_; 
wire REGFILE_SIM_reg_bank_reg_r11_26_; 
wire REGFILE_SIM_reg_bank_reg_r11_27_; 
wire REGFILE_SIM_reg_bank_reg_r11_28_; 
wire REGFILE_SIM_reg_bank_reg_r11_29_; 
wire REGFILE_SIM_reg_bank_reg_r11_2_; 
wire REGFILE_SIM_reg_bank_reg_r11_30_; 
wire REGFILE_SIM_reg_bank_reg_r11_31_; 
wire REGFILE_SIM_reg_bank_reg_r11_3_; 
wire REGFILE_SIM_reg_bank_reg_r11_4_; 
wire REGFILE_SIM_reg_bank_reg_r11_5_; 
wire REGFILE_SIM_reg_bank_reg_r11_6_; 
wire REGFILE_SIM_reg_bank_reg_r11_7_; 
wire REGFILE_SIM_reg_bank_reg_r11_8_; 
wire REGFILE_SIM_reg_bank_reg_r11_9_; 
wire REGFILE_SIM_reg_bank_reg_r12_0_; 
wire REGFILE_SIM_reg_bank_reg_r12_10_; 
wire REGFILE_SIM_reg_bank_reg_r12_11_; 
wire REGFILE_SIM_reg_bank_reg_r12_12_; 
wire REGFILE_SIM_reg_bank_reg_r12_13_; 
wire REGFILE_SIM_reg_bank_reg_r12_14_; 
wire REGFILE_SIM_reg_bank_reg_r12_15_; 
wire REGFILE_SIM_reg_bank_reg_r12_16_; 
wire REGFILE_SIM_reg_bank_reg_r12_17_; 
wire REGFILE_SIM_reg_bank_reg_r12_18_; 
wire REGFILE_SIM_reg_bank_reg_r12_19_; 
wire REGFILE_SIM_reg_bank_reg_r12_1_; 
wire REGFILE_SIM_reg_bank_reg_r12_20_; 
wire REGFILE_SIM_reg_bank_reg_r12_21_; 
wire REGFILE_SIM_reg_bank_reg_r12_22_; 
wire REGFILE_SIM_reg_bank_reg_r12_23_; 
wire REGFILE_SIM_reg_bank_reg_r12_24_; 
wire REGFILE_SIM_reg_bank_reg_r12_25_; 
wire REGFILE_SIM_reg_bank_reg_r12_26_; 
wire REGFILE_SIM_reg_bank_reg_r12_27_; 
wire REGFILE_SIM_reg_bank_reg_r12_28_; 
wire REGFILE_SIM_reg_bank_reg_r12_29_; 
wire REGFILE_SIM_reg_bank_reg_r12_2_; 
wire REGFILE_SIM_reg_bank_reg_r12_30_; 
wire REGFILE_SIM_reg_bank_reg_r12_31_; 
wire REGFILE_SIM_reg_bank_reg_r12_3_; 
wire REGFILE_SIM_reg_bank_reg_r12_4_; 
wire REGFILE_SIM_reg_bank_reg_r12_5_; 
wire REGFILE_SIM_reg_bank_reg_r12_6_; 
wire REGFILE_SIM_reg_bank_reg_r12_7_; 
wire REGFILE_SIM_reg_bank_reg_r12_8_; 
wire REGFILE_SIM_reg_bank_reg_r12_9_; 
wire REGFILE_SIM_reg_bank_reg_r13_0_; 
wire REGFILE_SIM_reg_bank_reg_r13_10_; 
wire REGFILE_SIM_reg_bank_reg_r13_11_; 
wire REGFILE_SIM_reg_bank_reg_r13_12_; 
wire REGFILE_SIM_reg_bank_reg_r13_13_; 
wire REGFILE_SIM_reg_bank_reg_r13_14_; 
wire REGFILE_SIM_reg_bank_reg_r13_15_; 
wire REGFILE_SIM_reg_bank_reg_r13_16_; 
wire REGFILE_SIM_reg_bank_reg_r13_17_; 
wire REGFILE_SIM_reg_bank_reg_r13_18_; 
wire REGFILE_SIM_reg_bank_reg_r13_19_; 
wire REGFILE_SIM_reg_bank_reg_r13_1_; 
wire REGFILE_SIM_reg_bank_reg_r13_20_; 
wire REGFILE_SIM_reg_bank_reg_r13_21_; 
wire REGFILE_SIM_reg_bank_reg_r13_22_; 
wire REGFILE_SIM_reg_bank_reg_r13_23_; 
wire REGFILE_SIM_reg_bank_reg_r13_24_; 
wire REGFILE_SIM_reg_bank_reg_r13_25_; 
wire REGFILE_SIM_reg_bank_reg_r13_26_; 
wire REGFILE_SIM_reg_bank_reg_r13_27_; 
wire REGFILE_SIM_reg_bank_reg_r13_28_; 
wire REGFILE_SIM_reg_bank_reg_r13_29_; 
wire REGFILE_SIM_reg_bank_reg_r13_2_; 
wire REGFILE_SIM_reg_bank_reg_r13_30_; 
wire REGFILE_SIM_reg_bank_reg_r13_31_; 
wire REGFILE_SIM_reg_bank_reg_r13_3_; 
wire REGFILE_SIM_reg_bank_reg_r13_4_; 
wire REGFILE_SIM_reg_bank_reg_r13_5_; 
wire REGFILE_SIM_reg_bank_reg_r13_6_; 
wire REGFILE_SIM_reg_bank_reg_r13_7_; 
wire REGFILE_SIM_reg_bank_reg_r13_8_; 
wire REGFILE_SIM_reg_bank_reg_r13_9_; 
wire REGFILE_SIM_reg_bank_reg_r14_0_; 
wire REGFILE_SIM_reg_bank_reg_r14_10_; 
wire REGFILE_SIM_reg_bank_reg_r14_11_; 
wire REGFILE_SIM_reg_bank_reg_r14_12_; 
wire REGFILE_SIM_reg_bank_reg_r14_13_; 
wire REGFILE_SIM_reg_bank_reg_r14_14_; 
wire REGFILE_SIM_reg_bank_reg_r14_15_; 
wire REGFILE_SIM_reg_bank_reg_r14_16_; 
wire REGFILE_SIM_reg_bank_reg_r14_17_; 
wire REGFILE_SIM_reg_bank_reg_r14_18_; 
wire REGFILE_SIM_reg_bank_reg_r14_19_; 
wire REGFILE_SIM_reg_bank_reg_r14_1_; 
wire REGFILE_SIM_reg_bank_reg_r14_20_; 
wire REGFILE_SIM_reg_bank_reg_r14_21_; 
wire REGFILE_SIM_reg_bank_reg_r14_22_; 
wire REGFILE_SIM_reg_bank_reg_r14_23_; 
wire REGFILE_SIM_reg_bank_reg_r14_24_; 
wire REGFILE_SIM_reg_bank_reg_r14_25_; 
wire REGFILE_SIM_reg_bank_reg_r14_26_; 
wire REGFILE_SIM_reg_bank_reg_r14_27_; 
wire REGFILE_SIM_reg_bank_reg_r14_28_; 
wire REGFILE_SIM_reg_bank_reg_r14_29_; 
wire REGFILE_SIM_reg_bank_reg_r14_2_; 
wire REGFILE_SIM_reg_bank_reg_r14_30_; 
wire REGFILE_SIM_reg_bank_reg_r14_31_; 
wire REGFILE_SIM_reg_bank_reg_r14_3_; 
wire REGFILE_SIM_reg_bank_reg_r14_4_; 
wire REGFILE_SIM_reg_bank_reg_r14_5_; 
wire REGFILE_SIM_reg_bank_reg_r14_6_; 
wire REGFILE_SIM_reg_bank_reg_r14_7_; 
wire REGFILE_SIM_reg_bank_reg_r14_8_; 
wire REGFILE_SIM_reg_bank_reg_r14_9_; 
wire REGFILE_SIM_reg_bank_reg_r15_0_; 
wire REGFILE_SIM_reg_bank_reg_r15_10_; 
wire REGFILE_SIM_reg_bank_reg_r15_11_; 
wire REGFILE_SIM_reg_bank_reg_r15_12_; 
wire REGFILE_SIM_reg_bank_reg_r15_13_; 
wire REGFILE_SIM_reg_bank_reg_r15_14_; 
wire REGFILE_SIM_reg_bank_reg_r15_15_; 
wire REGFILE_SIM_reg_bank_reg_r15_16_; 
wire REGFILE_SIM_reg_bank_reg_r15_17_; 
wire REGFILE_SIM_reg_bank_reg_r15_18_; 
wire REGFILE_SIM_reg_bank_reg_r15_19_; 
wire REGFILE_SIM_reg_bank_reg_r15_1_; 
wire REGFILE_SIM_reg_bank_reg_r15_20_; 
wire REGFILE_SIM_reg_bank_reg_r15_21_; 
wire REGFILE_SIM_reg_bank_reg_r15_22_; 
wire REGFILE_SIM_reg_bank_reg_r15_23_; 
wire REGFILE_SIM_reg_bank_reg_r15_24_; 
wire REGFILE_SIM_reg_bank_reg_r15_25_; 
wire REGFILE_SIM_reg_bank_reg_r15_26_; 
wire REGFILE_SIM_reg_bank_reg_r15_27_; 
wire REGFILE_SIM_reg_bank_reg_r15_28_; 
wire REGFILE_SIM_reg_bank_reg_r15_29_; 
wire REGFILE_SIM_reg_bank_reg_r15_2_; 
wire REGFILE_SIM_reg_bank_reg_r15_30_; 
wire REGFILE_SIM_reg_bank_reg_r15_31_; 
wire REGFILE_SIM_reg_bank_reg_r15_3_; 
wire REGFILE_SIM_reg_bank_reg_r15_4_; 
wire REGFILE_SIM_reg_bank_reg_r15_5_; 
wire REGFILE_SIM_reg_bank_reg_r15_6_; 
wire REGFILE_SIM_reg_bank_reg_r15_7_; 
wire REGFILE_SIM_reg_bank_reg_r15_8_; 
wire REGFILE_SIM_reg_bank_reg_r15_9_; 
wire REGFILE_SIM_reg_bank_reg_r16_0_; 
wire REGFILE_SIM_reg_bank_reg_r16_10_; 
wire REGFILE_SIM_reg_bank_reg_r16_11_; 
wire REGFILE_SIM_reg_bank_reg_r16_12_; 
wire REGFILE_SIM_reg_bank_reg_r16_13_; 
wire REGFILE_SIM_reg_bank_reg_r16_14_; 
wire REGFILE_SIM_reg_bank_reg_r16_15_; 
wire REGFILE_SIM_reg_bank_reg_r16_16_; 
wire REGFILE_SIM_reg_bank_reg_r16_17_; 
wire REGFILE_SIM_reg_bank_reg_r16_18_; 
wire REGFILE_SIM_reg_bank_reg_r16_19_; 
wire REGFILE_SIM_reg_bank_reg_r16_1_; 
wire REGFILE_SIM_reg_bank_reg_r16_20_; 
wire REGFILE_SIM_reg_bank_reg_r16_21_; 
wire REGFILE_SIM_reg_bank_reg_r16_22_; 
wire REGFILE_SIM_reg_bank_reg_r16_23_; 
wire REGFILE_SIM_reg_bank_reg_r16_24_; 
wire REGFILE_SIM_reg_bank_reg_r16_25_; 
wire REGFILE_SIM_reg_bank_reg_r16_26_; 
wire REGFILE_SIM_reg_bank_reg_r16_27_; 
wire REGFILE_SIM_reg_bank_reg_r16_28_; 
wire REGFILE_SIM_reg_bank_reg_r16_29_; 
wire REGFILE_SIM_reg_bank_reg_r16_2_; 
wire REGFILE_SIM_reg_bank_reg_r16_30_; 
wire REGFILE_SIM_reg_bank_reg_r16_31_; 
wire REGFILE_SIM_reg_bank_reg_r16_3_; 
wire REGFILE_SIM_reg_bank_reg_r16_4_; 
wire REGFILE_SIM_reg_bank_reg_r16_5_; 
wire REGFILE_SIM_reg_bank_reg_r16_6_; 
wire REGFILE_SIM_reg_bank_reg_r16_7_; 
wire REGFILE_SIM_reg_bank_reg_r16_8_; 
wire REGFILE_SIM_reg_bank_reg_r16_9_; 
wire REGFILE_SIM_reg_bank_reg_r17_0_; 
wire REGFILE_SIM_reg_bank_reg_r17_10_; 
wire REGFILE_SIM_reg_bank_reg_r17_11_; 
wire REGFILE_SIM_reg_bank_reg_r17_12_; 
wire REGFILE_SIM_reg_bank_reg_r17_13_; 
wire REGFILE_SIM_reg_bank_reg_r17_14_; 
wire REGFILE_SIM_reg_bank_reg_r17_15_; 
wire REGFILE_SIM_reg_bank_reg_r17_16_; 
wire REGFILE_SIM_reg_bank_reg_r17_17_; 
wire REGFILE_SIM_reg_bank_reg_r17_18_; 
wire REGFILE_SIM_reg_bank_reg_r17_19_; 
wire REGFILE_SIM_reg_bank_reg_r17_1_; 
wire REGFILE_SIM_reg_bank_reg_r17_20_; 
wire REGFILE_SIM_reg_bank_reg_r17_21_; 
wire REGFILE_SIM_reg_bank_reg_r17_22_; 
wire REGFILE_SIM_reg_bank_reg_r17_23_; 
wire REGFILE_SIM_reg_bank_reg_r17_24_; 
wire REGFILE_SIM_reg_bank_reg_r17_25_; 
wire REGFILE_SIM_reg_bank_reg_r17_26_; 
wire REGFILE_SIM_reg_bank_reg_r17_27_; 
wire REGFILE_SIM_reg_bank_reg_r17_28_; 
wire REGFILE_SIM_reg_bank_reg_r17_29_; 
wire REGFILE_SIM_reg_bank_reg_r17_2_; 
wire REGFILE_SIM_reg_bank_reg_r17_30_; 
wire REGFILE_SIM_reg_bank_reg_r17_31_; 
wire REGFILE_SIM_reg_bank_reg_r17_3_; 
wire REGFILE_SIM_reg_bank_reg_r17_4_; 
wire REGFILE_SIM_reg_bank_reg_r17_5_; 
wire REGFILE_SIM_reg_bank_reg_r17_6_; 
wire REGFILE_SIM_reg_bank_reg_r17_7_; 
wire REGFILE_SIM_reg_bank_reg_r17_8_; 
wire REGFILE_SIM_reg_bank_reg_r17_9_; 
wire REGFILE_SIM_reg_bank_reg_r18_0_; 
wire REGFILE_SIM_reg_bank_reg_r18_10_; 
wire REGFILE_SIM_reg_bank_reg_r18_11_; 
wire REGFILE_SIM_reg_bank_reg_r18_12_; 
wire REGFILE_SIM_reg_bank_reg_r18_13_; 
wire REGFILE_SIM_reg_bank_reg_r18_14_; 
wire REGFILE_SIM_reg_bank_reg_r18_15_; 
wire REGFILE_SIM_reg_bank_reg_r18_16_; 
wire REGFILE_SIM_reg_bank_reg_r18_17_; 
wire REGFILE_SIM_reg_bank_reg_r18_18_; 
wire REGFILE_SIM_reg_bank_reg_r18_19_; 
wire REGFILE_SIM_reg_bank_reg_r18_1_; 
wire REGFILE_SIM_reg_bank_reg_r18_20_; 
wire REGFILE_SIM_reg_bank_reg_r18_21_; 
wire REGFILE_SIM_reg_bank_reg_r18_22_; 
wire REGFILE_SIM_reg_bank_reg_r18_23_; 
wire REGFILE_SIM_reg_bank_reg_r18_24_; 
wire REGFILE_SIM_reg_bank_reg_r18_25_; 
wire REGFILE_SIM_reg_bank_reg_r18_26_; 
wire REGFILE_SIM_reg_bank_reg_r18_27_; 
wire REGFILE_SIM_reg_bank_reg_r18_28_; 
wire REGFILE_SIM_reg_bank_reg_r18_29_; 
wire REGFILE_SIM_reg_bank_reg_r18_2_; 
wire REGFILE_SIM_reg_bank_reg_r18_30_; 
wire REGFILE_SIM_reg_bank_reg_r18_31_; 
wire REGFILE_SIM_reg_bank_reg_r18_3_; 
wire REGFILE_SIM_reg_bank_reg_r18_4_; 
wire REGFILE_SIM_reg_bank_reg_r18_5_; 
wire REGFILE_SIM_reg_bank_reg_r18_6_; 
wire REGFILE_SIM_reg_bank_reg_r18_7_; 
wire REGFILE_SIM_reg_bank_reg_r18_8_; 
wire REGFILE_SIM_reg_bank_reg_r18_9_; 
wire REGFILE_SIM_reg_bank_reg_r19_0_; 
wire REGFILE_SIM_reg_bank_reg_r19_10_; 
wire REGFILE_SIM_reg_bank_reg_r19_11_; 
wire REGFILE_SIM_reg_bank_reg_r19_12_; 
wire REGFILE_SIM_reg_bank_reg_r19_13_; 
wire REGFILE_SIM_reg_bank_reg_r19_14_; 
wire REGFILE_SIM_reg_bank_reg_r19_15_; 
wire REGFILE_SIM_reg_bank_reg_r19_16_; 
wire REGFILE_SIM_reg_bank_reg_r19_17_; 
wire REGFILE_SIM_reg_bank_reg_r19_18_; 
wire REGFILE_SIM_reg_bank_reg_r19_19_; 
wire REGFILE_SIM_reg_bank_reg_r19_1_; 
wire REGFILE_SIM_reg_bank_reg_r19_20_; 
wire REGFILE_SIM_reg_bank_reg_r19_21_; 
wire REGFILE_SIM_reg_bank_reg_r19_22_; 
wire REGFILE_SIM_reg_bank_reg_r19_23_; 
wire REGFILE_SIM_reg_bank_reg_r19_24_; 
wire REGFILE_SIM_reg_bank_reg_r19_25_; 
wire REGFILE_SIM_reg_bank_reg_r19_26_; 
wire REGFILE_SIM_reg_bank_reg_r19_27_; 
wire REGFILE_SIM_reg_bank_reg_r19_28_; 
wire REGFILE_SIM_reg_bank_reg_r19_29_; 
wire REGFILE_SIM_reg_bank_reg_r19_2_; 
wire REGFILE_SIM_reg_bank_reg_r19_30_; 
wire REGFILE_SIM_reg_bank_reg_r19_31_; 
wire REGFILE_SIM_reg_bank_reg_r19_3_; 
wire REGFILE_SIM_reg_bank_reg_r19_4_; 
wire REGFILE_SIM_reg_bank_reg_r19_5_; 
wire REGFILE_SIM_reg_bank_reg_r19_6_; 
wire REGFILE_SIM_reg_bank_reg_r19_7_; 
wire REGFILE_SIM_reg_bank_reg_r19_8_; 
wire REGFILE_SIM_reg_bank_reg_r19_9_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_0_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_10_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_11_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_12_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_13_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_14_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_15_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_16_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_17_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_18_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_19_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_1_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_20_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_21_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_22_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_23_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_24_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_25_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_26_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_27_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_28_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_29_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_2_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_30_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_31_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_3_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_4_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_5_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_6_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_7_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_8_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_9_; 
wire REGFILE_SIM_reg_bank_reg_r20_0_; 
wire REGFILE_SIM_reg_bank_reg_r20_10_; 
wire REGFILE_SIM_reg_bank_reg_r20_11_; 
wire REGFILE_SIM_reg_bank_reg_r20_12_; 
wire REGFILE_SIM_reg_bank_reg_r20_13_; 
wire REGFILE_SIM_reg_bank_reg_r20_14_; 
wire REGFILE_SIM_reg_bank_reg_r20_15_; 
wire REGFILE_SIM_reg_bank_reg_r20_16_; 
wire REGFILE_SIM_reg_bank_reg_r20_17_; 
wire REGFILE_SIM_reg_bank_reg_r20_18_; 
wire REGFILE_SIM_reg_bank_reg_r20_19_; 
wire REGFILE_SIM_reg_bank_reg_r20_1_; 
wire REGFILE_SIM_reg_bank_reg_r20_20_; 
wire REGFILE_SIM_reg_bank_reg_r20_21_; 
wire REGFILE_SIM_reg_bank_reg_r20_22_; 
wire REGFILE_SIM_reg_bank_reg_r20_23_; 
wire REGFILE_SIM_reg_bank_reg_r20_24_; 
wire REGFILE_SIM_reg_bank_reg_r20_25_; 
wire REGFILE_SIM_reg_bank_reg_r20_26_; 
wire REGFILE_SIM_reg_bank_reg_r20_27_; 
wire REGFILE_SIM_reg_bank_reg_r20_28_; 
wire REGFILE_SIM_reg_bank_reg_r20_29_; 
wire REGFILE_SIM_reg_bank_reg_r20_2_; 
wire REGFILE_SIM_reg_bank_reg_r20_30_; 
wire REGFILE_SIM_reg_bank_reg_r20_31_; 
wire REGFILE_SIM_reg_bank_reg_r20_3_; 
wire REGFILE_SIM_reg_bank_reg_r20_4_; 
wire REGFILE_SIM_reg_bank_reg_r20_5_; 
wire REGFILE_SIM_reg_bank_reg_r20_6_; 
wire REGFILE_SIM_reg_bank_reg_r20_7_; 
wire REGFILE_SIM_reg_bank_reg_r20_8_; 
wire REGFILE_SIM_reg_bank_reg_r20_9_; 
wire REGFILE_SIM_reg_bank_reg_r21_0_; 
wire REGFILE_SIM_reg_bank_reg_r21_10_; 
wire REGFILE_SIM_reg_bank_reg_r21_11_; 
wire REGFILE_SIM_reg_bank_reg_r21_12_; 
wire REGFILE_SIM_reg_bank_reg_r21_13_; 
wire REGFILE_SIM_reg_bank_reg_r21_14_; 
wire REGFILE_SIM_reg_bank_reg_r21_15_; 
wire REGFILE_SIM_reg_bank_reg_r21_16_; 
wire REGFILE_SIM_reg_bank_reg_r21_17_; 
wire REGFILE_SIM_reg_bank_reg_r21_18_; 
wire REGFILE_SIM_reg_bank_reg_r21_19_; 
wire REGFILE_SIM_reg_bank_reg_r21_1_; 
wire REGFILE_SIM_reg_bank_reg_r21_20_; 
wire REGFILE_SIM_reg_bank_reg_r21_21_; 
wire REGFILE_SIM_reg_bank_reg_r21_22_; 
wire REGFILE_SIM_reg_bank_reg_r21_23_; 
wire REGFILE_SIM_reg_bank_reg_r21_24_; 
wire REGFILE_SIM_reg_bank_reg_r21_25_; 
wire REGFILE_SIM_reg_bank_reg_r21_26_; 
wire REGFILE_SIM_reg_bank_reg_r21_27_; 
wire REGFILE_SIM_reg_bank_reg_r21_28_; 
wire REGFILE_SIM_reg_bank_reg_r21_29_; 
wire REGFILE_SIM_reg_bank_reg_r21_2_; 
wire REGFILE_SIM_reg_bank_reg_r21_30_; 
wire REGFILE_SIM_reg_bank_reg_r21_31_; 
wire REGFILE_SIM_reg_bank_reg_r21_3_; 
wire REGFILE_SIM_reg_bank_reg_r21_4_; 
wire REGFILE_SIM_reg_bank_reg_r21_5_; 
wire REGFILE_SIM_reg_bank_reg_r21_6_; 
wire REGFILE_SIM_reg_bank_reg_r21_7_; 
wire REGFILE_SIM_reg_bank_reg_r21_8_; 
wire REGFILE_SIM_reg_bank_reg_r21_9_; 
wire REGFILE_SIM_reg_bank_reg_r22_0_; 
wire REGFILE_SIM_reg_bank_reg_r22_10_; 
wire REGFILE_SIM_reg_bank_reg_r22_11_; 
wire REGFILE_SIM_reg_bank_reg_r22_12_; 
wire REGFILE_SIM_reg_bank_reg_r22_13_; 
wire REGFILE_SIM_reg_bank_reg_r22_14_; 
wire REGFILE_SIM_reg_bank_reg_r22_15_; 
wire REGFILE_SIM_reg_bank_reg_r22_16_; 
wire REGFILE_SIM_reg_bank_reg_r22_17_; 
wire REGFILE_SIM_reg_bank_reg_r22_18_; 
wire REGFILE_SIM_reg_bank_reg_r22_19_; 
wire REGFILE_SIM_reg_bank_reg_r22_1_; 
wire REGFILE_SIM_reg_bank_reg_r22_20_; 
wire REGFILE_SIM_reg_bank_reg_r22_21_; 
wire REGFILE_SIM_reg_bank_reg_r22_22_; 
wire REGFILE_SIM_reg_bank_reg_r22_23_; 
wire REGFILE_SIM_reg_bank_reg_r22_24_; 
wire REGFILE_SIM_reg_bank_reg_r22_25_; 
wire REGFILE_SIM_reg_bank_reg_r22_26_; 
wire REGFILE_SIM_reg_bank_reg_r22_27_; 
wire REGFILE_SIM_reg_bank_reg_r22_28_; 
wire REGFILE_SIM_reg_bank_reg_r22_29_; 
wire REGFILE_SIM_reg_bank_reg_r22_2_; 
wire REGFILE_SIM_reg_bank_reg_r22_30_; 
wire REGFILE_SIM_reg_bank_reg_r22_31_; 
wire REGFILE_SIM_reg_bank_reg_r22_3_; 
wire REGFILE_SIM_reg_bank_reg_r22_4_; 
wire REGFILE_SIM_reg_bank_reg_r22_5_; 
wire REGFILE_SIM_reg_bank_reg_r22_6_; 
wire REGFILE_SIM_reg_bank_reg_r22_7_; 
wire REGFILE_SIM_reg_bank_reg_r22_8_; 
wire REGFILE_SIM_reg_bank_reg_r22_9_; 
wire REGFILE_SIM_reg_bank_reg_r23_0_; 
wire REGFILE_SIM_reg_bank_reg_r23_10_; 
wire REGFILE_SIM_reg_bank_reg_r23_11_; 
wire REGFILE_SIM_reg_bank_reg_r23_12_; 
wire REGFILE_SIM_reg_bank_reg_r23_13_; 
wire REGFILE_SIM_reg_bank_reg_r23_14_; 
wire REGFILE_SIM_reg_bank_reg_r23_15_; 
wire REGFILE_SIM_reg_bank_reg_r23_16_; 
wire REGFILE_SIM_reg_bank_reg_r23_17_; 
wire REGFILE_SIM_reg_bank_reg_r23_18_; 
wire REGFILE_SIM_reg_bank_reg_r23_19_; 
wire REGFILE_SIM_reg_bank_reg_r23_1_; 
wire REGFILE_SIM_reg_bank_reg_r23_20_; 
wire REGFILE_SIM_reg_bank_reg_r23_21_; 
wire REGFILE_SIM_reg_bank_reg_r23_22_; 
wire REGFILE_SIM_reg_bank_reg_r23_23_; 
wire REGFILE_SIM_reg_bank_reg_r23_24_; 
wire REGFILE_SIM_reg_bank_reg_r23_25_; 
wire REGFILE_SIM_reg_bank_reg_r23_26_; 
wire REGFILE_SIM_reg_bank_reg_r23_27_; 
wire REGFILE_SIM_reg_bank_reg_r23_28_; 
wire REGFILE_SIM_reg_bank_reg_r23_29_; 
wire REGFILE_SIM_reg_bank_reg_r23_2_; 
wire REGFILE_SIM_reg_bank_reg_r23_30_; 
wire REGFILE_SIM_reg_bank_reg_r23_31_; 
wire REGFILE_SIM_reg_bank_reg_r23_3_; 
wire REGFILE_SIM_reg_bank_reg_r23_4_; 
wire REGFILE_SIM_reg_bank_reg_r23_5_; 
wire REGFILE_SIM_reg_bank_reg_r23_6_; 
wire REGFILE_SIM_reg_bank_reg_r23_7_; 
wire REGFILE_SIM_reg_bank_reg_r23_8_; 
wire REGFILE_SIM_reg_bank_reg_r23_9_; 
wire REGFILE_SIM_reg_bank_reg_r24_0_; 
wire REGFILE_SIM_reg_bank_reg_r24_10_; 
wire REGFILE_SIM_reg_bank_reg_r24_11_; 
wire REGFILE_SIM_reg_bank_reg_r24_12_; 
wire REGFILE_SIM_reg_bank_reg_r24_13_; 
wire REGFILE_SIM_reg_bank_reg_r24_14_; 
wire REGFILE_SIM_reg_bank_reg_r24_15_; 
wire REGFILE_SIM_reg_bank_reg_r24_16_; 
wire REGFILE_SIM_reg_bank_reg_r24_17_; 
wire REGFILE_SIM_reg_bank_reg_r24_18_; 
wire REGFILE_SIM_reg_bank_reg_r24_19_; 
wire REGFILE_SIM_reg_bank_reg_r24_1_; 
wire REGFILE_SIM_reg_bank_reg_r24_20_; 
wire REGFILE_SIM_reg_bank_reg_r24_21_; 
wire REGFILE_SIM_reg_bank_reg_r24_22_; 
wire REGFILE_SIM_reg_bank_reg_r24_23_; 
wire REGFILE_SIM_reg_bank_reg_r24_24_; 
wire REGFILE_SIM_reg_bank_reg_r24_25_; 
wire REGFILE_SIM_reg_bank_reg_r24_26_; 
wire REGFILE_SIM_reg_bank_reg_r24_27_; 
wire REGFILE_SIM_reg_bank_reg_r24_28_; 
wire REGFILE_SIM_reg_bank_reg_r24_29_; 
wire REGFILE_SIM_reg_bank_reg_r24_2_; 
wire REGFILE_SIM_reg_bank_reg_r24_30_; 
wire REGFILE_SIM_reg_bank_reg_r24_31_; 
wire REGFILE_SIM_reg_bank_reg_r24_3_; 
wire REGFILE_SIM_reg_bank_reg_r24_4_; 
wire REGFILE_SIM_reg_bank_reg_r24_5_; 
wire REGFILE_SIM_reg_bank_reg_r24_6_; 
wire REGFILE_SIM_reg_bank_reg_r24_7_; 
wire REGFILE_SIM_reg_bank_reg_r24_8_; 
wire REGFILE_SIM_reg_bank_reg_r24_9_; 
wire REGFILE_SIM_reg_bank_reg_r25_0_; 
wire REGFILE_SIM_reg_bank_reg_r25_10_; 
wire REGFILE_SIM_reg_bank_reg_r25_11_; 
wire REGFILE_SIM_reg_bank_reg_r25_12_; 
wire REGFILE_SIM_reg_bank_reg_r25_13_; 
wire REGFILE_SIM_reg_bank_reg_r25_14_; 
wire REGFILE_SIM_reg_bank_reg_r25_15_; 
wire REGFILE_SIM_reg_bank_reg_r25_16_; 
wire REGFILE_SIM_reg_bank_reg_r25_17_; 
wire REGFILE_SIM_reg_bank_reg_r25_18_; 
wire REGFILE_SIM_reg_bank_reg_r25_19_; 
wire REGFILE_SIM_reg_bank_reg_r25_1_; 
wire REGFILE_SIM_reg_bank_reg_r25_20_; 
wire REGFILE_SIM_reg_bank_reg_r25_21_; 
wire REGFILE_SIM_reg_bank_reg_r25_22_; 
wire REGFILE_SIM_reg_bank_reg_r25_23_; 
wire REGFILE_SIM_reg_bank_reg_r25_24_; 
wire REGFILE_SIM_reg_bank_reg_r25_25_; 
wire REGFILE_SIM_reg_bank_reg_r25_26_; 
wire REGFILE_SIM_reg_bank_reg_r25_27_; 
wire REGFILE_SIM_reg_bank_reg_r25_28_; 
wire REGFILE_SIM_reg_bank_reg_r25_29_; 
wire REGFILE_SIM_reg_bank_reg_r25_2_; 
wire REGFILE_SIM_reg_bank_reg_r25_30_; 
wire REGFILE_SIM_reg_bank_reg_r25_31_; 
wire REGFILE_SIM_reg_bank_reg_r25_3_; 
wire REGFILE_SIM_reg_bank_reg_r25_4_; 
wire REGFILE_SIM_reg_bank_reg_r25_5_; 
wire REGFILE_SIM_reg_bank_reg_r25_6_; 
wire REGFILE_SIM_reg_bank_reg_r25_7_; 
wire REGFILE_SIM_reg_bank_reg_r25_8_; 
wire REGFILE_SIM_reg_bank_reg_r25_9_; 
wire REGFILE_SIM_reg_bank_reg_r26_0_; 
wire REGFILE_SIM_reg_bank_reg_r26_10_; 
wire REGFILE_SIM_reg_bank_reg_r26_11_; 
wire REGFILE_SIM_reg_bank_reg_r26_12_; 
wire REGFILE_SIM_reg_bank_reg_r26_13_; 
wire REGFILE_SIM_reg_bank_reg_r26_14_; 
wire REGFILE_SIM_reg_bank_reg_r26_15_; 
wire REGFILE_SIM_reg_bank_reg_r26_16_; 
wire REGFILE_SIM_reg_bank_reg_r26_17_; 
wire REGFILE_SIM_reg_bank_reg_r26_18_; 
wire REGFILE_SIM_reg_bank_reg_r26_19_; 
wire REGFILE_SIM_reg_bank_reg_r26_1_; 
wire REGFILE_SIM_reg_bank_reg_r26_20_; 
wire REGFILE_SIM_reg_bank_reg_r26_21_; 
wire REGFILE_SIM_reg_bank_reg_r26_22_; 
wire REGFILE_SIM_reg_bank_reg_r26_23_; 
wire REGFILE_SIM_reg_bank_reg_r26_24_; 
wire REGFILE_SIM_reg_bank_reg_r26_25_; 
wire REGFILE_SIM_reg_bank_reg_r26_26_; 
wire REGFILE_SIM_reg_bank_reg_r26_27_; 
wire REGFILE_SIM_reg_bank_reg_r26_28_; 
wire REGFILE_SIM_reg_bank_reg_r26_29_; 
wire REGFILE_SIM_reg_bank_reg_r26_2_; 
wire REGFILE_SIM_reg_bank_reg_r26_30_; 
wire REGFILE_SIM_reg_bank_reg_r26_31_; 
wire REGFILE_SIM_reg_bank_reg_r26_3_; 
wire REGFILE_SIM_reg_bank_reg_r26_4_; 
wire REGFILE_SIM_reg_bank_reg_r26_5_; 
wire REGFILE_SIM_reg_bank_reg_r26_6_; 
wire REGFILE_SIM_reg_bank_reg_r26_7_; 
wire REGFILE_SIM_reg_bank_reg_r26_8_; 
wire REGFILE_SIM_reg_bank_reg_r26_9_; 
wire REGFILE_SIM_reg_bank_reg_r27_0_; 
wire REGFILE_SIM_reg_bank_reg_r27_10_; 
wire REGFILE_SIM_reg_bank_reg_r27_11_; 
wire REGFILE_SIM_reg_bank_reg_r27_12_; 
wire REGFILE_SIM_reg_bank_reg_r27_13_; 
wire REGFILE_SIM_reg_bank_reg_r27_14_; 
wire REGFILE_SIM_reg_bank_reg_r27_15_; 
wire REGFILE_SIM_reg_bank_reg_r27_16_; 
wire REGFILE_SIM_reg_bank_reg_r27_17_; 
wire REGFILE_SIM_reg_bank_reg_r27_18_; 
wire REGFILE_SIM_reg_bank_reg_r27_19_; 
wire REGFILE_SIM_reg_bank_reg_r27_1_; 
wire REGFILE_SIM_reg_bank_reg_r27_20_; 
wire REGFILE_SIM_reg_bank_reg_r27_21_; 
wire REGFILE_SIM_reg_bank_reg_r27_22_; 
wire REGFILE_SIM_reg_bank_reg_r27_23_; 
wire REGFILE_SIM_reg_bank_reg_r27_24_; 
wire REGFILE_SIM_reg_bank_reg_r27_25_; 
wire REGFILE_SIM_reg_bank_reg_r27_26_; 
wire REGFILE_SIM_reg_bank_reg_r27_27_; 
wire REGFILE_SIM_reg_bank_reg_r27_28_; 
wire REGFILE_SIM_reg_bank_reg_r27_29_; 
wire REGFILE_SIM_reg_bank_reg_r27_2_; 
wire REGFILE_SIM_reg_bank_reg_r27_30_; 
wire REGFILE_SIM_reg_bank_reg_r27_31_; 
wire REGFILE_SIM_reg_bank_reg_r27_3_; 
wire REGFILE_SIM_reg_bank_reg_r27_4_; 
wire REGFILE_SIM_reg_bank_reg_r27_5_; 
wire REGFILE_SIM_reg_bank_reg_r27_6_; 
wire REGFILE_SIM_reg_bank_reg_r27_7_; 
wire REGFILE_SIM_reg_bank_reg_r27_8_; 
wire REGFILE_SIM_reg_bank_reg_r27_9_; 
wire REGFILE_SIM_reg_bank_reg_r28_0_; 
wire REGFILE_SIM_reg_bank_reg_r28_10_; 
wire REGFILE_SIM_reg_bank_reg_r28_11_; 
wire REGFILE_SIM_reg_bank_reg_r28_12_; 
wire REGFILE_SIM_reg_bank_reg_r28_13_; 
wire REGFILE_SIM_reg_bank_reg_r28_14_; 
wire REGFILE_SIM_reg_bank_reg_r28_15_; 
wire REGFILE_SIM_reg_bank_reg_r28_16_; 
wire REGFILE_SIM_reg_bank_reg_r28_17_; 
wire REGFILE_SIM_reg_bank_reg_r28_18_; 
wire REGFILE_SIM_reg_bank_reg_r28_19_; 
wire REGFILE_SIM_reg_bank_reg_r28_1_; 
wire REGFILE_SIM_reg_bank_reg_r28_20_; 
wire REGFILE_SIM_reg_bank_reg_r28_21_; 
wire REGFILE_SIM_reg_bank_reg_r28_22_; 
wire REGFILE_SIM_reg_bank_reg_r28_23_; 
wire REGFILE_SIM_reg_bank_reg_r28_24_; 
wire REGFILE_SIM_reg_bank_reg_r28_25_; 
wire REGFILE_SIM_reg_bank_reg_r28_26_; 
wire REGFILE_SIM_reg_bank_reg_r28_27_; 
wire REGFILE_SIM_reg_bank_reg_r28_28_; 
wire REGFILE_SIM_reg_bank_reg_r28_29_; 
wire REGFILE_SIM_reg_bank_reg_r28_2_; 
wire REGFILE_SIM_reg_bank_reg_r28_30_; 
wire REGFILE_SIM_reg_bank_reg_r28_31_; 
wire REGFILE_SIM_reg_bank_reg_r28_3_; 
wire REGFILE_SIM_reg_bank_reg_r28_4_; 
wire REGFILE_SIM_reg_bank_reg_r28_5_; 
wire REGFILE_SIM_reg_bank_reg_r28_6_; 
wire REGFILE_SIM_reg_bank_reg_r28_7_; 
wire REGFILE_SIM_reg_bank_reg_r28_8_; 
wire REGFILE_SIM_reg_bank_reg_r28_9_; 
wire REGFILE_SIM_reg_bank_reg_r29_0_; 
wire REGFILE_SIM_reg_bank_reg_r29_10_; 
wire REGFILE_SIM_reg_bank_reg_r29_11_; 
wire REGFILE_SIM_reg_bank_reg_r29_12_; 
wire REGFILE_SIM_reg_bank_reg_r29_13_; 
wire REGFILE_SIM_reg_bank_reg_r29_14_; 
wire REGFILE_SIM_reg_bank_reg_r29_15_; 
wire REGFILE_SIM_reg_bank_reg_r29_16_; 
wire REGFILE_SIM_reg_bank_reg_r29_17_; 
wire REGFILE_SIM_reg_bank_reg_r29_18_; 
wire REGFILE_SIM_reg_bank_reg_r29_19_; 
wire REGFILE_SIM_reg_bank_reg_r29_1_; 
wire REGFILE_SIM_reg_bank_reg_r29_20_; 
wire REGFILE_SIM_reg_bank_reg_r29_21_; 
wire REGFILE_SIM_reg_bank_reg_r29_22_; 
wire REGFILE_SIM_reg_bank_reg_r29_23_; 
wire REGFILE_SIM_reg_bank_reg_r29_24_; 
wire REGFILE_SIM_reg_bank_reg_r29_25_; 
wire REGFILE_SIM_reg_bank_reg_r29_26_; 
wire REGFILE_SIM_reg_bank_reg_r29_27_; 
wire REGFILE_SIM_reg_bank_reg_r29_28_; 
wire REGFILE_SIM_reg_bank_reg_r29_29_; 
wire REGFILE_SIM_reg_bank_reg_r29_2_; 
wire REGFILE_SIM_reg_bank_reg_r29_30_; 
wire REGFILE_SIM_reg_bank_reg_r29_31_; 
wire REGFILE_SIM_reg_bank_reg_r29_3_; 
wire REGFILE_SIM_reg_bank_reg_r29_4_; 
wire REGFILE_SIM_reg_bank_reg_r29_5_; 
wire REGFILE_SIM_reg_bank_reg_r29_6_; 
wire REGFILE_SIM_reg_bank_reg_r29_7_; 
wire REGFILE_SIM_reg_bank_reg_r29_8_; 
wire REGFILE_SIM_reg_bank_reg_r29_9_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_0_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_10_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_11_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_12_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_13_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_14_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_15_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_16_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_17_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_18_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_19_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_1_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_20_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_21_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_22_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_23_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_24_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_25_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_26_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_27_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_28_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_29_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_2_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_30_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_31_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_3_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_4_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_5_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_6_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_7_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_8_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_9_; 
wire REGFILE_SIM_reg_bank_reg_r30_0_; 
wire REGFILE_SIM_reg_bank_reg_r30_10_; 
wire REGFILE_SIM_reg_bank_reg_r30_11_; 
wire REGFILE_SIM_reg_bank_reg_r30_12_; 
wire REGFILE_SIM_reg_bank_reg_r30_13_; 
wire REGFILE_SIM_reg_bank_reg_r30_14_; 
wire REGFILE_SIM_reg_bank_reg_r30_15_; 
wire REGFILE_SIM_reg_bank_reg_r30_16_; 
wire REGFILE_SIM_reg_bank_reg_r30_17_; 
wire REGFILE_SIM_reg_bank_reg_r30_18_; 
wire REGFILE_SIM_reg_bank_reg_r30_19_; 
wire REGFILE_SIM_reg_bank_reg_r30_1_; 
wire REGFILE_SIM_reg_bank_reg_r30_20_; 
wire REGFILE_SIM_reg_bank_reg_r30_21_; 
wire REGFILE_SIM_reg_bank_reg_r30_22_; 
wire REGFILE_SIM_reg_bank_reg_r30_23_; 
wire REGFILE_SIM_reg_bank_reg_r30_24_; 
wire REGFILE_SIM_reg_bank_reg_r30_25_; 
wire REGFILE_SIM_reg_bank_reg_r30_26_; 
wire REGFILE_SIM_reg_bank_reg_r30_27_; 
wire REGFILE_SIM_reg_bank_reg_r30_28_; 
wire REGFILE_SIM_reg_bank_reg_r30_29_; 
wire REGFILE_SIM_reg_bank_reg_r30_2_; 
wire REGFILE_SIM_reg_bank_reg_r30_30_; 
wire REGFILE_SIM_reg_bank_reg_r30_31_; 
wire REGFILE_SIM_reg_bank_reg_r30_3_; 
wire REGFILE_SIM_reg_bank_reg_r30_4_; 
wire REGFILE_SIM_reg_bank_reg_r30_5_; 
wire REGFILE_SIM_reg_bank_reg_r30_6_; 
wire REGFILE_SIM_reg_bank_reg_r30_7_; 
wire REGFILE_SIM_reg_bank_reg_r30_8_; 
wire REGFILE_SIM_reg_bank_reg_r30_9_; 
wire REGFILE_SIM_reg_bank_reg_r31_0_; 
wire REGFILE_SIM_reg_bank_reg_r31_10_; 
wire REGFILE_SIM_reg_bank_reg_r31_11_; 
wire REGFILE_SIM_reg_bank_reg_r31_12_; 
wire REGFILE_SIM_reg_bank_reg_r31_13_; 
wire REGFILE_SIM_reg_bank_reg_r31_14_; 
wire REGFILE_SIM_reg_bank_reg_r31_15_; 
wire REGFILE_SIM_reg_bank_reg_r31_16_; 
wire REGFILE_SIM_reg_bank_reg_r31_17_; 
wire REGFILE_SIM_reg_bank_reg_r31_18_; 
wire REGFILE_SIM_reg_bank_reg_r31_19_; 
wire REGFILE_SIM_reg_bank_reg_r31_1_; 
wire REGFILE_SIM_reg_bank_reg_r31_20_; 
wire REGFILE_SIM_reg_bank_reg_r31_21_; 
wire REGFILE_SIM_reg_bank_reg_r31_22_; 
wire REGFILE_SIM_reg_bank_reg_r31_23_; 
wire REGFILE_SIM_reg_bank_reg_r31_24_; 
wire REGFILE_SIM_reg_bank_reg_r31_25_; 
wire REGFILE_SIM_reg_bank_reg_r31_26_; 
wire REGFILE_SIM_reg_bank_reg_r31_27_; 
wire REGFILE_SIM_reg_bank_reg_r31_28_; 
wire REGFILE_SIM_reg_bank_reg_r31_29_; 
wire REGFILE_SIM_reg_bank_reg_r31_2_; 
wire REGFILE_SIM_reg_bank_reg_r31_30_; 
wire REGFILE_SIM_reg_bank_reg_r31_31_; 
wire REGFILE_SIM_reg_bank_reg_r31_3_; 
wire REGFILE_SIM_reg_bank_reg_r31_4_; 
wire REGFILE_SIM_reg_bank_reg_r31_5_; 
wire REGFILE_SIM_reg_bank_reg_r31_6_; 
wire REGFILE_SIM_reg_bank_reg_r31_7_; 
wire REGFILE_SIM_reg_bank_reg_r31_8_; 
wire REGFILE_SIM_reg_bank_reg_r31_9_; 
wire REGFILE_SIM_reg_bank_reg_r3_0_; 
wire REGFILE_SIM_reg_bank_reg_r3_10_; 
wire REGFILE_SIM_reg_bank_reg_r3_11_; 
wire REGFILE_SIM_reg_bank_reg_r3_12_; 
wire REGFILE_SIM_reg_bank_reg_r3_13_; 
wire REGFILE_SIM_reg_bank_reg_r3_14_; 
wire REGFILE_SIM_reg_bank_reg_r3_15_; 
wire REGFILE_SIM_reg_bank_reg_r3_16_; 
wire REGFILE_SIM_reg_bank_reg_r3_17_; 
wire REGFILE_SIM_reg_bank_reg_r3_18_; 
wire REGFILE_SIM_reg_bank_reg_r3_19_; 
wire REGFILE_SIM_reg_bank_reg_r3_1_; 
wire REGFILE_SIM_reg_bank_reg_r3_20_; 
wire REGFILE_SIM_reg_bank_reg_r3_21_; 
wire REGFILE_SIM_reg_bank_reg_r3_22_; 
wire REGFILE_SIM_reg_bank_reg_r3_23_; 
wire REGFILE_SIM_reg_bank_reg_r3_24_; 
wire REGFILE_SIM_reg_bank_reg_r3_25_; 
wire REGFILE_SIM_reg_bank_reg_r3_26_; 
wire REGFILE_SIM_reg_bank_reg_r3_27_; 
wire REGFILE_SIM_reg_bank_reg_r3_28_; 
wire REGFILE_SIM_reg_bank_reg_r3_29_; 
wire REGFILE_SIM_reg_bank_reg_r3_2_; 
wire REGFILE_SIM_reg_bank_reg_r3_30_; 
wire REGFILE_SIM_reg_bank_reg_r3_31_; 
wire REGFILE_SIM_reg_bank_reg_r3_3_; 
wire REGFILE_SIM_reg_bank_reg_r3_4_; 
wire REGFILE_SIM_reg_bank_reg_r3_5_; 
wire REGFILE_SIM_reg_bank_reg_r3_6_; 
wire REGFILE_SIM_reg_bank_reg_r3_7_; 
wire REGFILE_SIM_reg_bank_reg_r3_8_; 
wire REGFILE_SIM_reg_bank_reg_r3_9_; 
wire REGFILE_SIM_reg_bank_reg_r4_0_; 
wire REGFILE_SIM_reg_bank_reg_r4_10_; 
wire REGFILE_SIM_reg_bank_reg_r4_11_; 
wire REGFILE_SIM_reg_bank_reg_r4_12_; 
wire REGFILE_SIM_reg_bank_reg_r4_13_; 
wire REGFILE_SIM_reg_bank_reg_r4_14_; 
wire REGFILE_SIM_reg_bank_reg_r4_15_; 
wire REGFILE_SIM_reg_bank_reg_r4_16_; 
wire REGFILE_SIM_reg_bank_reg_r4_17_; 
wire REGFILE_SIM_reg_bank_reg_r4_18_; 
wire REGFILE_SIM_reg_bank_reg_r4_19_; 
wire REGFILE_SIM_reg_bank_reg_r4_1_; 
wire REGFILE_SIM_reg_bank_reg_r4_20_; 
wire REGFILE_SIM_reg_bank_reg_r4_21_; 
wire REGFILE_SIM_reg_bank_reg_r4_22_; 
wire REGFILE_SIM_reg_bank_reg_r4_23_; 
wire REGFILE_SIM_reg_bank_reg_r4_24_; 
wire REGFILE_SIM_reg_bank_reg_r4_25_; 
wire REGFILE_SIM_reg_bank_reg_r4_26_; 
wire REGFILE_SIM_reg_bank_reg_r4_27_; 
wire REGFILE_SIM_reg_bank_reg_r4_28_; 
wire REGFILE_SIM_reg_bank_reg_r4_29_; 
wire REGFILE_SIM_reg_bank_reg_r4_2_; 
wire REGFILE_SIM_reg_bank_reg_r4_30_; 
wire REGFILE_SIM_reg_bank_reg_r4_31_; 
wire REGFILE_SIM_reg_bank_reg_r4_3_; 
wire REGFILE_SIM_reg_bank_reg_r4_4_; 
wire REGFILE_SIM_reg_bank_reg_r4_5_; 
wire REGFILE_SIM_reg_bank_reg_r4_6_; 
wire REGFILE_SIM_reg_bank_reg_r4_7_; 
wire REGFILE_SIM_reg_bank_reg_r4_8_; 
wire REGFILE_SIM_reg_bank_reg_r4_9_; 
wire REGFILE_SIM_reg_bank_reg_r5_0_; 
wire REGFILE_SIM_reg_bank_reg_r5_10_; 
wire REGFILE_SIM_reg_bank_reg_r5_11_; 
wire REGFILE_SIM_reg_bank_reg_r5_12_; 
wire REGFILE_SIM_reg_bank_reg_r5_13_; 
wire REGFILE_SIM_reg_bank_reg_r5_14_; 
wire REGFILE_SIM_reg_bank_reg_r5_15_; 
wire REGFILE_SIM_reg_bank_reg_r5_16_; 
wire REGFILE_SIM_reg_bank_reg_r5_17_; 
wire REGFILE_SIM_reg_bank_reg_r5_18_; 
wire REGFILE_SIM_reg_bank_reg_r5_19_; 
wire REGFILE_SIM_reg_bank_reg_r5_1_; 
wire REGFILE_SIM_reg_bank_reg_r5_20_; 
wire REGFILE_SIM_reg_bank_reg_r5_21_; 
wire REGFILE_SIM_reg_bank_reg_r5_22_; 
wire REGFILE_SIM_reg_bank_reg_r5_23_; 
wire REGFILE_SIM_reg_bank_reg_r5_24_; 
wire REGFILE_SIM_reg_bank_reg_r5_25_; 
wire REGFILE_SIM_reg_bank_reg_r5_26_; 
wire REGFILE_SIM_reg_bank_reg_r5_27_; 
wire REGFILE_SIM_reg_bank_reg_r5_28_; 
wire REGFILE_SIM_reg_bank_reg_r5_29_; 
wire REGFILE_SIM_reg_bank_reg_r5_2_; 
wire REGFILE_SIM_reg_bank_reg_r5_30_; 
wire REGFILE_SIM_reg_bank_reg_r5_31_; 
wire REGFILE_SIM_reg_bank_reg_r5_3_; 
wire REGFILE_SIM_reg_bank_reg_r5_4_; 
wire REGFILE_SIM_reg_bank_reg_r5_5_; 
wire REGFILE_SIM_reg_bank_reg_r5_6_; 
wire REGFILE_SIM_reg_bank_reg_r5_7_; 
wire REGFILE_SIM_reg_bank_reg_r5_8_; 
wire REGFILE_SIM_reg_bank_reg_r5_9_; 
wire REGFILE_SIM_reg_bank_reg_r6_0_; 
wire REGFILE_SIM_reg_bank_reg_r6_10_; 
wire REGFILE_SIM_reg_bank_reg_r6_11_; 
wire REGFILE_SIM_reg_bank_reg_r6_12_; 
wire REGFILE_SIM_reg_bank_reg_r6_13_; 
wire REGFILE_SIM_reg_bank_reg_r6_14_; 
wire REGFILE_SIM_reg_bank_reg_r6_15_; 
wire REGFILE_SIM_reg_bank_reg_r6_16_; 
wire REGFILE_SIM_reg_bank_reg_r6_17_; 
wire REGFILE_SIM_reg_bank_reg_r6_18_; 
wire REGFILE_SIM_reg_bank_reg_r6_19_; 
wire REGFILE_SIM_reg_bank_reg_r6_1_; 
wire REGFILE_SIM_reg_bank_reg_r6_20_; 
wire REGFILE_SIM_reg_bank_reg_r6_21_; 
wire REGFILE_SIM_reg_bank_reg_r6_22_; 
wire REGFILE_SIM_reg_bank_reg_r6_23_; 
wire REGFILE_SIM_reg_bank_reg_r6_24_; 
wire REGFILE_SIM_reg_bank_reg_r6_25_; 
wire REGFILE_SIM_reg_bank_reg_r6_26_; 
wire REGFILE_SIM_reg_bank_reg_r6_27_; 
wire REGFILE_SIM_reg_bank_reg_r6_28_; 
wire REGFILE_SIM_reg_bank_reg_r6_29_; 
wire REGFILE_SIM_reg_bank_reg_r6_2_; 
wire REGFILE_SIM_reg_bank_reg_r6_30_; 
wire REGFILE_SIM_reg_bank_reg_r6_31_; 
wire REGFILE_SIM_reg_bank_reg_r6_3_; 
wire REGFILE_SIM_reg_bank_reg_r6_4_; 
wire REGFILE_SIM_reg_bank_reg_r6_5_; 
wire REGFILE_SIM_reg_bank_reg_r6_6_; 
wire REGFILE_SIM_reg_bank_reg_r6_7_; 
wire REGFILE_SIM_reg_bank_reg_r6_8_; 
wire REGFILE_SIM_reg_bank_reg_r6_9_; 
wire REGFILE_SIM_reg_bank_reg_r7_0_; 
wire REGFILE_SIM_reg_bank_reg_r7_10_; 
wire REGFILE_SIM_reg_bank_reg_r7_11_; 
wire REGFILE_SIM_reg_bank_reg_r7_12_; 
wire REGFILE_SIM_reg_bank_reg_r7_13_; 
wire REGFILE_SIM_reg_bank_reg_r7_14_; 
wire REGFILE_SIM_reg_bank_reg_r7_15_; 
wire REGFILE_SIM_reg_bank_reg_r7_16_; 
wire REGFILE_SIM_reg_bank_reg_r7_17_; 
wire REGFILE_SIM_reg_bank_reg_r7_18_; 
wire REGFILE_SIM_reg_bank_reg_r7_19_; 
wire REGFILE_SIM_reg_bank_reg_r7_1_; 
wire REGFILE_SIM_reg_bank_reg_r7_20_; 
wire REGFILE_SIM_reg_bank_reg_r7_21_; 
wire REGFILE_SIM_reg_bank_reg_r7_22_; 
wire REGFILE_SIM_reg_bank_reg_r7_23_; 
wire REGFILE_SIM_reg_bank_reg_r7_24_; 
wire REGFILE_SIM_reg_bank_reg_r7_25_; 
wire REGFILE_SIM_reg_bank_reg_r7_26_; 
wire REGFILE_SIM_reg_bank_reg_r7_27_; 
wire REGFILE_SIM_reg_bank_reg_r7_28_; 
wire REGFILE_SIM_reg_bank_reg_r7_29_; 
wire REGFILE_SIM_reg_bank_reg_r7_2_; 
wire REGFILE_SIM_reg_bank_reg_r7_30_; 
wire REGFILE_SIM_reg_bank_reg_r7_31_; 
wire REGFILE_SIM_reg_bank_reg_r7_3_; 
wire REGFILE_SIM_reg_bank_reg_r7_4_; 
wire REGFILE_SIM_reg_bank_reg_r7_5_; 
wire REGFILE_SIM_reg_bank_reg_r7_6_; 
wire REGFILE_SIM_reg_bank_reg_r7_7_; 
wire REGFILE_SIM_reg_bank_reg_r7_8_; 
wire REGFILE_SIM_reg_bank_reg_r7_9_; 
wire REGFILE_SIM_reg_bank_reg_r8_0_; 
wire REGFILE_SIM_reg_bank_reg_r8_10_; 
wire REGFILE_SIM_reg_bank_reg_r8_11_; 
wire REGFILE_SIM_reg_bank_reg_r8_12_; 
wire REGFILE_SIM_reg_bank_reg_r8_13_; 
wire REGFILE_SIM_reg_bank_reg_r8_14_; 
wire REGFILE_SIM_reg_bank_reg_r8_15_; 
wire REGFILE_SIM_reg_bank_reg_r8_16_; 
wire REGFILE_SIM_reg_bank_reg_r8_17_; 
wire REGFILE_SIM_reg_bank_reg_r8_18_; 
wire REGFILE_SIM_reg_bank_reg_r8_19_; 
wire REGFILE_SIM_reg_bank_reg_r8_1_; 
wire REGFILE_SIM_reg_bank_reg_r8_20_; 
wire REGFILE_SIM_reg_bank_reg_r8_21_; 
wire REGFILE_SIM_reg_bank_reg_r8_22_; 
wire REGFILE_SIM_reg_bank_reg_r8_23_; 
wire REGFILE_SIM_reg_bank_reg_r8_24_; 
wire REGFILE_SIM_reg_bank_reg_r8_25_; 
wire REGFILE_SIM_reg_bank_reg_r8_26_; 
wire REGFILE_SIM_reg_bank_reg_r8_27_; 
wire REGFILE_SIM_reg_bank_reg_r8_28_; 
wire REGFILE_SIM_reg_bank_reg_r8_29_; 
wire REGFILE_SIM_reg_bank_reg_r8_2_; 
wire REGFILE_SIM_reg_bank_reg_r8_30_; 
wire REGFILE_SIM_reg_bank_reg_r8_31_; 
wire REGFILE_SIM_reg_bank_reg_r8_3_; 
wire REGFILE_SIM_reg_bank_reg_r8_4_; 
wire REGFILE_SIM_reg_bank_reg_r8_5_; 
wire REGFILE_SIM_reg_bank_reg_r8_6_; 
wire REGFILE_SIM_reg_bank_reg_r8_7_; 
wire REGFILE_SIM_reg_bank_reg_r8_8_; 
wire REGFILE_SIM_reg_bank_reg_r8_9_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_0_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_10_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_11_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_12_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_13_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_14_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_15_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_16_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_17_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_18_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_19_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_1_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_20_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_21_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_22_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_23_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_24_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_25_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_26_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_27_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_28_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_29_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_2_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_30_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_31_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_3_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_4_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_5_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_6_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_7_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_8_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_9_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_0_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_10_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_11_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_12_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_13_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_14_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_15_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_16_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_17_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_18_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_19_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_1_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_20_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_21_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_22_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_23_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_24_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_25_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_26_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_27_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_28_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_29_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_2_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_30_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_31_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_3_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_4_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_5_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_6_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_7_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_8_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_9_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_0_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_10_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_11_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_12_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_13_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_14_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_15_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_16_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_17_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_18_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_19_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_1_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_20_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_21_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_22_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_23_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_24_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_25_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_26_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_27_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_28_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_29_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_2_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_30_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_31_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_3_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_4_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_5_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_6_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_7_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_8_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_9_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_0_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_10_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_11_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_12_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_13_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_14_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_15_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_16_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_17_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_18_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_19_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_1_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_20_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_21_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_22_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_23_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_24_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_25_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_26_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_27_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_28_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_29_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_2_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_30_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_31_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_3_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_4_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_5_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_6_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_7_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_8_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_9_; 
wire REGFILE_SIM_reg_bank_wr_i; 
wire _0epc_q_31_0__0_; 
wire _0epc_q_31_0__10_; 
wire _0epc_q_31_0__11_; 
wire _0epc_q_31_0__12_; 
wire _0epc_q_31_0__13_; 
wire _0epc_q_31_0__14_; 
wire _0epc_q_31_0__15_; 
wire _0epc_q_31_0__16_; 
wire _0epc_q_31_0__17_; 
wire _0epc_q_31_0__18_; 
wire _0epc_q_31_0__19_; 
wire _0epc_q_31_0__1_; 
wire _0epc_q_31_0__20_; 
wire _0epc_q_31_0__21_; 
wire _0epc_q_31_0__22_; 
wire _0epc_q_31_0__23_; 
wire _0epc_q_31_0__24_; 
wire _0epc_q_31_0__25_; 
wire _0epc_q_31_0__26_; 
wire _0epc_q_31_0__27_; 
wire _0epc_q_31_0__28_; 
wire _0epc_q_31_0__29_; 
wire _0epc_q_31_0__2_; 
wire _0epc_q_31_0__30_; 
wire _0epc_q_31_0__31_; 
wire _0epc_q_31_0__3_; 
wire _0epc_q_31_0__4_; 
wire _0epc_q_31_0__5_; 
wire _0epc_q_31_0__6_; 
wire _0epc_q_31_0__7_; 
wire _0epc_q_31_0__8_; 
wire _0epc_q_31_0__9_; 
wire _0esr_q_31_0__10_; 
wire _0esr_q_31_0__2_; 
wire _0esr_q_31_0__9_; 
wire _0ex_rd_q_4_0__0_; 
wire _0ex_rd_q_4_0__1_; 
wire _0ex_rd_q_4_0__2_; 
wire _0ex_rd_q_4_0__3_; 
wire _0ex_rd_q_4_0__4_; 
wire _0fault_o_0_0_; 
wire _0mem_addr_o_31_0__0_; 
wire _0mem_addr_o_31_0__10_; 
wire _0mem_addr_o_31_0__11_; 
wire _0mem_addr_o_31_0__12_; 
wire _0mem_addr_o_31_0__13_; 
wire _0mem_addr_o_31_0__14_; 
wire _0mem_addr_o_31_0__15_; 
wire _0mem_addr_o_31_0__16_; 
wire _0mem_addr_o_31_0__17_; 
wire _0mem_addr_o_31_0__18_; 
wire _0mem_addr_o_31_0__19_; 
wire _0mem_addr_o_31_0__1_; 
wire _0mem_addr_o_31_0__20_; 
wire _0mem_addr_o_31_0__21_; 
wire _0mem_addr_o_31_0__22_; 
wire _0mem_addr_o_31_0__23_; 
wire _0mem_addr_o_31_0__24_; 
wire _0mem_addr_o_31_0__25_; 
wire _0mem_addr_o_31_0__26_; 
wire _0mem_addr_o_31_0__27_; 
wire _0mem_addr_o_31_0__28_; 
wire _0mem_addr_o_31_0__29_; 
wire _0mem_addr_o_31_0__2_; 
wire _0mem_addr_o_31_0__30_; 
wire _0mem_addr_o_31_0__31_; 
wire _0mem_addr_o_31_0__3_; 
wire _0mem_addr_o_31_0__4_; 
wire _0mem_addr_o_31_0__5_; 
wire _0mem_addr_o_31_0__6_; 
wire _0mem_addr_o_31_0__7_; 
wire _0mem_addr_o_31_0__8_; 
wire _0mem_addr_o_31_0__9_; 
wire _0mem_cyc_o_0_0_; 
wire _0mem_dat_o_31_0__0_; 
wire _0mem_dat_o_31_0__10_; 
wire _0mem_dat_o_31_0__11_; 
wire _0mem_dat_o_31_0__12_; 
wire _0mem_dat_o_31_0__13_; 
wire _0mem_dat_o_31_0__14_; 
wire _0mem_dat_o_31_0__15_; 
wire _0mem_dat_o_31_0__16_; 
wire _0mem_dat_o_31_0__17_; 
wire _0mem_dat_o_31_0__18_; 
wire _0mem_dat_o_31_0__19_; 
wire _0mem_dat_o_31_0__1_; 
wire _0mem_dat_o_31_0__20_; 
wire _0mem_dat_o_31_0__21_; 
wire _0mem_dat_o_31_0__22_; 
wire _0mem_dat_o_31_0__23_; 
wire _0mem_dat_o_31_0__24_; 
wire _0mem_dat_o_31_0__25_; 
wire _0mem_dat_o_31_0__26_; 
wire _0mem_dat_o_31_0__27_; 
wire _0mem_dat_o_31_0__28_; 
wire _0mem_dat_o_31_0__29_; 
wire _0mem_dat_o_31_0__2_; 
wire _0mem_dat_o_31_0__30_; 
wire _0mem_dat_o_31_0__31_; 
wire _0mem_dat_o_31_0__3_; 
wire _0mem_dat_o_31_0__4_; 
wire _0mem_dat_o_31_0__5_; 
wire _0mem_dat_o_31_0__6_; 
wire _0mem_dat_o_31_0__7_; 
wire _0mem_dat_o_31_0__8_; 
wire _0mem_dat_o_31_0__9_; 
wire _0mem_offset_q_1_0__0_; 
wire _0mem_offset_q_1_0__1_; 
wire _0mem_sel_o_3_0__0_; 
wire _0mem_sel_o_3_0__1_; 
wire _0mem_sel_o_3_0__2_; 
wire _0mem_sel_o_3_0__3_; 
wire _0mem_stb_o_0_0_; 
wire _0mem_we_o_0_0_; 
wire _0nmi_q_0_0_; 
wire _0opcode_q_31_0__0_; 
wire _0opcode_q_31_0__10_; 
wire _0opcode_q_31_0__11_; 
wire _0opcode_q_31_0__12_; 
wire _0opcode_q_31_0__13_; 
wire _0opcode_q_31_0__14_; 
wire _0opcode_q_31_0__15_; 
wire _0opcode_q_31_0__16_; 
wire _0opcode_q_31_0__17_; 
wire _0opcode_q_31_0__18_; 
wire _0opcode_q_31_0__19_; 
wire _0opcode_q_31_0__1_; 
wire _0opcode_q_31_0__20_; 
wire _0opcode_q_31_0__21_; 
wire _0opcode_q_31_0__22_; 
wire _0opcode_q_31_0__23_; 
wire _0opcode_q_31_0__24_; 
wire _0opcode_q_31_0__25_; 
wire _0opcode_q_31_0__26_; 
wire _0opcode_q_31_0__27_; 
wire _0opcode_q_31_0__28_; 
wire _0opcode_q_31_0__29_; 
wire _0opcode_q_31_0__2_; 
wire _0opcode_q_31_0__30_; 
wire _0opcode_q_31_0__31_; 
wire _0opcode_q_31_0__3_; 
wire _0opcode_q_31_0__4_; 
wire _0opcode_q_31_0__5_; 
wire _0opcode_q_31_0__6_; 
wire _0opcode_q_31_0__7_; 
wire _0opcode_q_31_0__8_; 
wire _0opcode_q_31_0__9_; 
wire _0pc_q_31_0__0_; 
wire _0pc_q_31_0__10_; 
wire _0pc_q_31_0__11_; 
wire _0pc_q_31_0__12_; 
wire _0pc_q_31_0__13_; 
wire _0pc_q_31_0__14_; 
wire _0pc_q_31_0__15_; 
wire _0pc_q_31_0__16_; 
wire _0pc_q_31_0__17_; 
wire _0pc_q_31_0__18_; 
wire _0pc_q_31_0__19_; 
wire _0pc_q_31_0__1_; 
wire _0pc_q_31_0__20_; 
wire _0pc_q_31_0__21_; 
wire _0pc_q_31_0__22_; 
wire _0pc_q_31_0__23_; 
wire _0pc_q_31_0__24_; 
wire _0pc_q_31_0__25_; 
wire _0pc_q_31_0__26_; 
wire _0pc_q_31_0__27_; 
wire _0pc_q_31_0__28_; 
wire _0pc_q_31_0__29_; 
wire _0pc_q_31_0__2_; 
wire _0pc_q_31_0__30_; 
wire _0pc_q_31_0__31_; 
wire _0pc_q_31_0__3_; 
wire _0pc_q_31_0__4_; 
wire _0pc_q_31_0__5_; 
wire _0pc_q_31_0__6_; 
wire _0pc_q_31_0__7_; 
wire _0pc_q_31_0__8_; 
wire _0pc_q_31_0__9_; 
wire _0sr_q_31_0__10_; 
wire _0sr_q_31_0__2_; 
wire _0sr_q_31_0__9_; 
wire _abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2382; 
wire _abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2420; 
wire _abc_27663_auto_fsm_map_cc_170_map_fsm_2376_1_; 
wire _abc_27663_auto_fsm_map_cc_170_map_fsm_2376_2_; 
wire _abc_27663_auto_fsm_map_cc_170_map_fsm_2376_3_; 
wire _abc_27663_auto_fsm_map_cc_170_map_fsm_2376_4_; 
wire _abc_40298_auto_rtlil_cc_1942_NotGate_33938; 
wire _abc_40298_new_n1000_; 
wire _abc_40298_new_n1001_; 
wire _abc_40298_new_n1002_; 
wire _abc_40298_new_n1003_; 
wire _abc_40298_new_n1004_; 
wire _abc_40298_new_n1005_; 
wire _abc_40298_new_n1006_; 
wire _abc_40298_new_n1007_; 
wire _abc_40298_new_n1008_; 
wire _abc_40298_new_n1009_; 
wire _abc_40298_new_n1010_; 
wire _abc_40298_new_n1011_; 
wire _abc_40298_new_n1012_; 
wire _abc_40298_new_n1013_; 
wire _abc_40298_new_n1014_; 
wire _abc_40298_new_n1015_; 
wire _abc_40298_new_n1016_; 
wire _abc_40298_new_n1017_; 
wire _abc_40298_new_n1018_; 
wire _abc_40298_new_n1019_; 
wire _abc_40298_new_n1020_; 
wire _abc_40298_new_n1021_; 
wire _abc_40298_new_n1022_; 
wire _abc_40298_new_n1023_; 
wire _abc_40298_new_n1024_; 
wire _abc_40298_new_n1025_; 
wire _abc_40298_new_n1026_; 
wire _abc_40298_new_n1027_; 
wire _abc_40298_new_n1028_; 
wire _abc_40298_new_n1029_; 
wire _abc_40298_new_n1030_; 
wire _abc_40298_new_n1031_; 
wire _abc_40298_new_n1032_; 
wire _abc_40298_new_n1033_; 
wire _abc_40298_new_n1034_; 
wire _abc_40298_new_n1035_; 
wire _abc_40298_new_n1036_; 
wire _abc_40298_new_n1037_; 
wire _abc_40298_new_n1038_; 
wire _abc_40298_new_n1039_; 
wire _abc_40298_new_n1040_; 
wire _abc_40298_new_n1041_; 
wire _abc_40298_new_n1042_; 
wire _abc_40298_new_n1043_; 
wire _abc_40298_new_n1044_; 
wire _abc_40298_new_n1045_; 
wire _abc_40298_new_n1046_; 
wire _abc_40298_new_n1047_; 
wire _abc_40298_new_n1048_; 
wire _abc_40298_new_n1049_; 
wire _abc_40298_new_n1050_; 
wire _abc_40298_new_n1051_; 
wire _abc_40298_new_n1052_; 
wire _abc_40298_new_n1053_; 
wire _abc_40298_new_n1054_; 
wire _abc_40298_new_n1055_; 
wire _abc_40298_new_n1056_; 
wire _abc_40298_new_n1057_; 
wire _abc_40298_new_n1058_; 
wire _abc_40298_new_n1059_; 
wire _abc_40298_new_n1060_; 
wire _abc_40298_new_n1061_; 
wire _abc_40298_new_n1062_; 
wire _abc_40298_new_n1063_; 
wire _abc_40298_new_n1064_; 
wire _abc_40298_new_n1065_; 
wire _abc_40298_new_n1066_; 
wire _abc_40298_new_n1067_; 
wire _abc_40298_new_n1068_; 
wire _abc_40298_new_n1069_; 
wire _abc_40298_new_n1070_; 
wire _abc_40298_new_n1071_; 
wire _abc_40298_new_n1072_; 
wire _abc_40298_new_n1073_; 
wire _abc_40298_new_n1074_; 
wire _abc_40298_new_n1075_; 
wire _abc_40298_new_n1076_; 
wire _abc_40298_new_n1077_; 
wire _abc_40298_new_n1078_; 
wire _abc_40298_new_n1079_; 
wire _abc_40298_new_n1080_; 
wire _abc_40298_new_n1081_; 
wire _abc_40298_new_n1082_; 
wire _abc_40298_new_n1083_; 
wire _abc_40298_new_n1084_; 
wire _abc_40298_new_n1085_; 
wire _abc_40298_new_n1086_; 
wire _abc_40298_new_n1087_; 
wire _abc_40298_new_n1089_; 
wire _abc_40298_new_n1090_; 
wire _abc_40298_new_n1091_; 
wire _abc_40298_new_n1092_; 
wire _abc_40298_new_n1093_; 
wire _abc_40298_new_n1094_; 
wire _abc_40298_new_n1095_; 
wire _abc_40298_new_n1096_; 
wire _abc_40298_new_n1097_; 
wire _abc_40298_new_n1098_; 
wire _abc_40298_new_n1099_; 
wire _abc_40298_new_n1100_; 
wire _abc_40298_new_n1101_; 
wire _abc_40298_new_n1102_; 
wire _abc_40298_new_n1103_; 
wire _abc_40298_new_n1104_; 
wire _abc_40298_new_n1105_; 
wire _abc_40298_new_n1106_; 
wire _abc_40298_new_n1107_; 
wire _abc_40298_new_n1108_; 
wire _abc_40298_new_n1109_; 
wire _abc_40298_new_n1110_; 
wire _abc_40298_new_n1111_; 
wire _abc_40298_new_n1112_; 
wire _abc_40298_new_n1113_; 
wire _abc_40298_new_n1114_; 
wire _abc_40298_new_n1115_; 
wire _abc_40298_new_n1116_; 
wire _abc_40298_new_n1117_; 
wire _abc_40298_new_n1118_; 
wire _abc_40298_new_n1119_; 
wire _abc_40298_new_n1120_; 
wire _abc_40298_new_n1121_; 
wire _abc_40298_new_n1122_; 
wire _abc_40298_new_n1123_; 
wire _abc_40298_new_n1124_; 
wire _abc_40298_new_n1125_; 
wire _abc_40298_new_n1126_; 
wire _abc_40298_new_n1127_; 
wire _abc_40298_new_n1128_; 
wire _abc_40298_new_n1129_; 
wire _abc_40298_new_n1130_; 
wire _abc_40298_new_n1131_; 
wire _abc_40298_new_n1132_; 
wire _abc_40298_new_n1133_; 
wire _abc_40298_new_n1134_; 
wire _abc_40298_new_n1135_; 
wire _abc_40298_new_n1136_; 
wire _abc_40298_new_n1137_; 
wire _abc_40298_new_n1138_; 
wire _abc_40298_new_n1139_; 
wire _abc_40298_new_n1140_; 
wire _abc_40298_new_n1141_; 
wire _abc_40298_new_n1142_; 
wire _abc_40298_new_n1143_; 
wire _abc_40298_new_n1145_; 
wire _abc_40298_new_n1146_; 
wire _abc_40298_new_n1147_; 
wire _abc_40298_new_n1148_; 
wire _abc_40298_new_n1149_; 
wire _abc_40298_new_n1150_; 
wire _abc_40298_new_n1151_; 
wire _abc_40298_new_n1152_; 
wire _abc_40298_new_n1153_; 
wire _abc_40298_new_n1154_; 
wire _abc_40298_new_n1155_; 
wire _abc_40298_new_n1156_; 
wire _abc_40298_new_n1157_; 
wire _abc_40298_new_n1159_; 
wire _abc_40298_new_n1160_; 
wire _abc_40298_new_n1161_; 
wire _abc_40298_new_n1163_; 
wire _abc_40298_new_n1164_; 
wire _abc_40298_new_n1166_; 
wire _abc_40298_new_n1167_; 
wire _abc_40298_new_n1168_; 
wire _abc_40298_new_n1169_; 
wire _abc_40298_new_n1170_; 
wire _abc_40298_new_n1171_; 
wire _abc_40298_new_n1173_; 
wire _abc_40298_new_n1174_; 
wire _abc_40298_new_n1175_; 
wire _abc_40298_new_n1176_; 
wire _abc_40298_new_n1177_; 
wire _abc_40298_new_n1178_; 
wire _abc_40298_new_n1179_; 
wire _abc_40298_new_n1180_; 
wire _abc_40298_new_n1181_; 
wire _abc_40298_new_n1182_; 
wire _abc_40298_new_n1183_; 
wire _abc_40298_new_n1184_; 
wire _abc_40298_new_n1185_; 
wire _abc_40298_new_n1186_; 
wire _abc_40298_new_n1187_; 
wire _abc_40298_new_n1188_; 
wire _abc_40298_new_n1189_; 
wire _abc_40298_new_n1190_; 
wire _abc_40298_new_n1191_; 
wire _abc_40298_new_n1192_; 
wire _abc_40298_new_n1193_; 
wire _abc_40298_new_n1194_; 
wire _abc_40298_new_n1196_; 
wire _abc_40298_new_n1197_; 
wire _abc_40298_new_n1198_; 
wire _abc_40298_new_n1199_; 
wire _abc_40298_new_n1200_; 
wire _abc_40298_new_n1201_; 
wire _abc_40298_new_n1202_; 
wire _abc_40298_new_n1203_; 
wire _abc_40298_new_n1204_; 
wire _abc_40298_new_n1205_; 
wire _abc_40298_new_n1206_; 
wire _abc_40298_new_n1208_; 
wire _abc_40298_new_n1209_; 
wire _abc_40298_new_n1210_; 
wire _abc_40298_new_n1211_; 
wire _abc_40298_new_n1212_; 
wire _abc_40298_new_n1213_; 
wire _abc_40298_new_n1214_; 
wire _abc_40298_new_n1215_; 
wire _abc_40298_new_n1216_; 
wire _abc_40298_new_n1217_; 
wire _abc_40298_new_n1218_; 
wire _abc_40298_new_n1219_; 
wire _abc_40298_new_n1220_; 
wire _abc_40298_new_n1221_; 
wire _abc_40298_new_n1222_; 
wire _abc_40298_new_n1223_; 
wire _abc_40298_new_n1224_; 
wire _abc_40298_new_n1225_; 
wire _abc_40298_new_n1226_; 
wire _abc_40298_new_n1227_; 
wire _abc_40298_new_n1229_; 
wire _abc_40298_new_n1230_; 
wire _abc_40298_new_n1231_; 
wire _abc_40298_new_n1232_; 
wire _abc_40298_new_n1233_; 
wire _abc_40298_new_n1234_; 
wire _abc_40298_new_n1235_; 
wire _abc_40298_new_n1236_; 
wire _abc_40298_new_n1237_; 
wire _abc_40298_new_n1238_; 
wire _abc_40298_new_n1239_; 
wire _abc_40298_new_n1240_; 
wire _abc_40298_new_n1241_; 
wire _abc_40298_new_n1242_; 
wire _abc_40298_new_n1243_; 
wire _abc_40298_new_n1244_; 
wire _abc_40298_new_n1245_; 
wire _abc_40298_new_n1246_; 
wire _abc_40298_new_n1247_; 
wire _abc_40298_new_n1248_; 
wire _abc_40298_new_n1249_; 
wire _abc_40298_new_n1250_; 
wire _abc_40298_new_n1252_; 
wire _abc_40298_new_n1253_; 
wire _abc_40298_new_n1254_; 
wire _abc_40298_new_n1255_; 
wire _abc_40298_new_n1256_; 
wire _abc_40298_new_n1257_; 
wire _abc_40298_new_n1258_; 
wire _abc_40298_new_n1259_; 
wire _abc_40298_new_n1260_; 
wire _abc_40298_new_n1261_; 
wire _abc_40298_new_n1262_; 
wire _abc_40298_new_n1263_; 
wire _abc_40298_new_n1264_; 
wire _abc_40298_new_n1265_; 
wire _abc_40298_new_n1266_; 
wire _abc_40298_new_n1267_; 
wire _abc_40298_new_n1268_; 
wire _abc_40298_new_n1269_; 
wire _abc_40298_new_n1270_; 
wire _abc_40298_new_n1271_; 
wire _abc_40298_new_n1272_; 
wire _abc_40298_new_n1273_; 
wire _abc_40298_new_n1274_; 
wire _abc_40298_new_n1275_; 
wire _abc_40298_new_n1276_; 
wire _abc_40298_new_n1278_; 
wire _abc_40298_new_n1279_; 
wire _abc_40298_new_n1280_; 
wire _abc_40298_new_n1281_; 
wire _abc_40298_new_n1282_; 
wire _abc_40298_new_n1283_; 
wire _abc_40298_new_n1284_; 
wire _abc_40298_new_n1285_; 
wire _abc_40298_new_n1286_; 
wire _abc_40298_new_n1287_; 
wire _abc_40298_new_n1288_; 
wire _abc_40298_new_n1289_; 
wire _abc_40298_new_n1290_; 
wire _abc_40298_new_n1291_; 
wire _abc_40298_new_n1292_; 
wire _abc_40298_new_n1293_; 
wire _abc_40298_new_n1294_; 
wire _abc_40298_new_n1295_; 
wire _abc_40298_new_n1296_; 
wire _abc_40298_new_n1297_; 
wire _abc_40298_new_n1298_; 
wire _abc_40298_new_n1299_; 
wire _abc_40298_new_n1300_; 
wire _abc_40298_new_n1302_; 
wire _abc_40298_new_n1303_; 
wire _abc_40298_new_n1304_; 
wire _abc_40298_new_n1305_; 
wire _abc_40298_new_n1306_; 
wire _abc_40298_new_n1307_; 
wire _abc_40298_new_n1308_; 
wire _abc_40298_new_n1309_; 
wire _abc_40298_new_n1310_; 
wire _abc_40298_new_n1311_; 
wire _abc_40298_new_n1312_; 
wire _abc_40298_new_n1313_; 
wire _abc_40298_new_n1314_; 
wire _abc_40298_new_n1315_; 
wire _abc_40298_new_n1316_; 
wire _abc_40298_new_n1317_; 
wire _abc_40298_new_n1318_; 
wire _abc_40298_new_n1319_; 
wire _abc_40298_new_n1320_; 
wire _abc_40298_new_n1321_; 
wire _abc_40298_new_n1322_; 
wire _abc_40298_new_n1323_; 
wire _abc_40298_new_n1324_; 
wire _abc_40298_new_n1325_; 
wire _abc_40298_new_n1326_; 
wire _abc_40298_new_n1327_; 
wire _abc_40298_new_n1328_; 
wire _abc_40298_new_n1329_; 
wire _abc_40298_new_n1331_; 
wire _abc_40298_new_n1332_; 
wire _abc_40298_new_n1333_; 
wire _abc_40298_new_n1334_; 
wire _abc_40298_new_n1335_; 
wire _abc_40298_new_n1336_; 
wire _abc_40298_new_n1337_; 
wire _abc_40298_new_n1338_; 
wire _abc_40298_new_n1339_; 
wire _abc_40298_new_n1340_; 
wire _abc_40298_new_n1341_; 
wire _abc_40298_new_n1342_; 
wire _abc_40298_new_n1343_; 
wire _abc_40298_new_n1344_; 
wire _abc_40298_new_n1345_; 
wire _abc_40298_new_n1346_; 
wire _abc_40298_new_n1347_; 
wire _abc_40298_new_n1348_; 
wire _abc_40298_new_n1349_; 
wire _abc_40298_new_n1350_; 
wire _abc_40298_new_n1351_; 
wire _abc_40298_new_n1352_; 
wire _abc_40298_new_n1353_; 
wire _abc_40298_new_n1354_; 
wire _abc_40298_new_n1355_; 
wire _abc_40298_new_n1356_; 
wire _abc_40298_new_n1357_; 
wire _abc_40298_new_n1358_; 
wire _abc_40298_new_n1359_; 
wire _abc_40298_new_n1360_; 
wire _abc_40298_new_n1362_; 
wire _abc_40298_new_n1363_; 
wire _abc_40298_new_n1364_; 
wire _abc_40298_new_n1365_; 
wire _abc_40298_new_n1366_; 
wire _abc_40298_new_n1367_; 
wire _abc_40298_new_n1368_; 
wire _abc_40298_new_n1369_; 
wire _abc_40298_new_n1370_; 
wire _abc_40298_new_n1371_; 
wire _abc_40298_new_n1372_; 
wire _abc_40298_new_n1373_; 
wire _abc_40298_new_n1374_; 
wire _abc_40298_new_n1375_; 
wire _abc_40298_new_n1376_; 
wire _abc_40298_new_n1377_; 
wire _abc_40298_new_n1378_; 
wire _abc_40298_new_n1379_; 
wire _abc_40298_new_n1380_; 
wire _abc_40298_new_n1381_; 
wire _abc_40298_new_n1382_; 
wire _abc_40298_new_n1383_; 
wire _abc_40298_new_n1384_; 
wire _abc_40298_new_n1385_; 
wire _abc_40298_new_n1386_; 
wire _abc_40298_new_n1387_; 
wire _abc_40298_new_n1388_; 
wire _abc_40298_new_n1389_; 
wire _abc_40298_new_n1391_; 
wire _abc_40298_new_n1392_; 
wire _abc_40298_new_n1393_; 
wire _abc_40298_new_n1394_; 
wire _abc_40298_new_n1395_; 
wire _abc_40298_new_n1396_; 
wire _abc_40298_new_n1397_; 
wire _abc_40298_new_n1398_; 
wire _abc_40298_new_n1399_; 
wire _abc_40298_new_n1400_; 
wire _abc_40298_new_n1401_; 
wire _abc_40298_new_n1402_; 
wire _abc_40298_new_n1403_; 
wire _abc_40298_new_n1404_; 
wire _abc_40298_new_n1405_; 
wire _abc_40298_new_n1406_; 
wire _abc_40298_new_n1407_; 
wire _abc_40298_new_n1408_; 
wire _abc_40298_new_n1409_; 
wire _abc_40298_new_n1410_; 
wire _abc_40298_new_n1411_; 
wire _abc_40298_new_n1412_; 
wire _abc_40298_new_n1414_; 
wire _abc_40298_new_n1415_; 
wire _abc_40298_new_n1416_; 
wire _abc_40298_new_n1417_; 
wire _abc_40298_new_n1418_; 
wire _abc_40298_new_n1419_; 
wire _abc_40298_new_n1420_; 
wire _abc_40298_new_n1421_; 
wire _abc_40298_new_n1422_; 
wire _abc_40298_new_n1423_; 
wire _abc_40298_new_n1424_; 
wire _abc_40298_new_n1425_; 
wire _abc_40298_new_n1426_; 
wire _abc_40298_new_n1427_; 
wire _abc_40298_new_n1428_; 
wire _abc_40298_new_n1429_; 
wire _abc_40298_new_n1430_; 
wire _abc_40298_new_n1431_; 
wire _abc_40298_new_n1432_; 
wire _abc_40298_new_n1433_; 
wire _abc_40298_new_n1434_; 
wire _abc_40298_new_n1435_; 
wire _abc_40298_new_n1436_; 
wire _abc_40298_new_n1437_; 
wire _abc_40298_new_n1438_; 
wire _abc_40298_new_n1439_; 
wire _abc_40298_new_n1440_; 
wire _abc_40298_new_n1441_; 
wire _abc_40298_new_n1442_; 
wire _abc_40298_new_n1443_; 
wire _abc_40298_new_n1444_; 
wire _abc_40298_new_n1446_; 
wire _abc_40298_new_n1447_; 
wire _abc_40298_new_n1448_; 
wire _abc_40298_new_n1449_; 
wire _abc_40298_new_n1450_; 
wire _abc_40298_new_n1451_; 
wire _abc_40298_new_n1452_; 
wire _abc_40298_new_n1453_; 
wire _abc_40298_new_n1454_; 
wire _abc_40298_new_n1455_; 
wire _abc_40298_new_n1456_; 
wire _abc_40298_new_n1457_; 
wire _abc_40298_new_n1458_; 
wire _abc_40298_new_n1459_; 
wire _abc_40298_new_n1460_; 
wire _abc_40298_new_n1461_; 
wire _abc_40298_new_n1462_; 
wire _abc_40298_new_n1463_; 
wire _abc_40298_new_n1464_; 
wire _abc_40298_new_n1465_; 
wire _abc_40298_new_n1466_; 
wire _abc_40298_new_n1467_; 
wire _abc_40298_new_n1468_; 
wire _abc_40298_new_n1469_; 
wire _abc_40298_new_n1470_; 
wire _abc_40298_new_n1471_; 
wire _abc_40298_new_n1473_; 
wire _abc_40298_new_n1474_; 
wire _abc_40298_new_n1475_; 
wire _abc_40298_new_n1476_; 
wire _abc_40298_new_n1477_; 
wire _abc_40298_new_n1478_; 
wire _abc_40298_new_n1479_; 
wire _abc_40298_new_n1480_; 
wire _abc_40298_new_n1481_; 
wire _abc_40298_new_n1482_; 
wire _abc_40298_new_n1483_; 
wire _abc_40298_new_n1484_; 
wire _abc_40298_new_n1485_; 
wire _abc_40298_new_n1486_; 
wire _abc_40298_new_n1487_; 
wire _abc_40298_new_n1488_; 
wire _abc_40298_new_n1489_; 
wire _abc_40298_new_n1490_; 
wire _abc_40298_new_n1491_; 
wire _abc_40298_new_n1492_; 
wire _abc_40298_new_n1493_; 
wire _abc_40298_new_n1494_; 
wire _abc_40298_new_n1495_; 
wire _abc_40298_new_n1496_; 
wire _abc_40298_new_n1497_; 
wire _abc_40298_new_n1498_; 
wire _abc_40298_new_n1499_; 
wire _abc_40298_new_n1500_; 
wire _abc_40298_new_n1501_; 
wire _abc_40298_new_n1502_; 
wire _abc_40298_new_n1503_; 
wire _abc_40298_new_n1504_; 
wire _abc_40298_new_n1505_; 
wire _abc_40298_new_n1506_; 
wire _abc_40298_new_n1507_; 
wire _abc_40298_new_n1509_; 
wire _abc_40298_new_n1510_; 
wire _abc_40298_new_n1511_; 
wire _abc_40298_new_n1512_; 
wire _abc_40298_new_n1513_; 
wire _abc_40298_new_n1514_; 
wire _abc_40298_new_n1515_; 
wire _abc_40298_new_n1516_; 
wire _abc_40298_new_n1517_; 
wire _abc_40298_new_n1518_; 
wire _abc_40298_new_n1519_; 
wire _abc_40298_new_n1520_; 
wire _abc_40298_new_n1521_; 
wire _abc_40298_new_n1522_; 
wire _abc_40298_new_n1523_; 
wire _abc_40298_new_n1524_; 
wire _abc_40298_new_n1525_; 
wire _abc_40298_new_n1526_; 
wire _abc_40298_new_n1527_; 
wire _abc_40298_new_n1528_; 
wire _abc_40298_new_n1529_; 
wire _abc_40298_new_n1530_; 
wire _abc_40298_new_n1532_; 
wire _abc_40298_new_n1533_; 
wire _abc_40298_new_n1534_; 
wire _abc_40298_new_n1535_; 
wire _abc_40298_new_n1536_; 
wire _abc_40298_new_n1537_; 
wire _abc_40298_new_n1538_; 
wire _abc_40298_new_n1539_; 
wire _abc_40298_new_n1540_; 
wire _abc_40298_new_n1541_; 
wire _abc_40298_new_n1542_; 
wire _abc_40298_new_n1543_; 
wire _abc_40298_new_n1544_; 
wire _abc_40298_new_n1545_; 
wire _abc_40298_new_n1546_; 
wire _abc_40298_new_n1547_; 
wire _abc_40298_new_n1548_; 
wire _abc_40298_new_n1549_; 
wire _abc_40298_new_n1550_; 
wire _abc_40298_new_n1551_; 
wire _abc_40298_new_n1552_; 
wire _abc_40298_new_n1553_; 
wire _abc_40298_new_n1554_; 
wire _abc_40298_new_n1555_; 
wire _abc_40298_new_n1556_; 
wire _abc_40298_new_n1557_; 
wire _abc_40298_new_n1558_; 
wire _abc_40298_new_n1559_; 
wire _abc_40298_new_n1561_; 
wire _abc_40298_new_n1562_; 
wire _abc_40298_new_n1563_; 
wire _abc_40298_new_n1564_; 
wire _abc_40298_new_n1565_; 
wire _abc_40298_new_n1566_; 
wire _abc_40298_new_n1567_; 
wire _abc_40298_new_n1568_; 
wire _abc_40298_new_n1569_; 
wire _abc_40298_new_n1570_; 
wire _abc_40298_new_n1571_; 
wire _abc_40298_new_n1572_; 
wire _abc_40298_new_n1573_; 
wire _abc_40298_new_n1574_; 
wire _abc_40298_new_n1575_; 
wire _abc_40298_new_n1576_; 
wire _abc_40298_new_n1577_; 
wire _abc_40298_new_n1578_; 
wire _abc_40298_new_n1579_; 
wire _abc_40298_new_n1580_; 
wire _abc_40298_new_n1581_; 
wire _abc_40298_new_n1582_; 
wire _abc_40298_new_n1583_; 
wire _abc_40298_new_n1584_; 
wire _abc_40298_new_n1585_; 
wire _abc_40298_new_n1587_; 
wire _abc_40298_new_n1588_; 
wire _abc_40298_new_n1589_; 
wire _abc_40298_new_n1590_; 
wire _abc_40298_new_n1591_; 
wire _abc_40298_new_n1592_; 
wire _abc_40298_new_n1593_; 
wire _abc_40298_new_n1594_; 
wire _abc_40298_new_n1595_; 
wire _abc_40298_new_n1596_; 
wire _abc_40298_new_n1597_; 
wire _abc_40298_new_n1598_; 
wire _abc_40298_new_n1599_; 
wire _abc_40298_new_n1600_; 
wire _abc_40298_new_n1601_; 
wire _abc_40298_new_n1602_; 
wire _abc_40298_new_n1603_; 
wire _abc_40298_new_n1604_; 
wire _abc_40298_new_n1605_; 
wire _abc_40298_new_n1606_; 
wire _abc_40298_new_n1607_; 
wire _abc_40298_new_n1608_; 
wire _abc_40298_new_n1609_; 
wire _abc_40298_new_n1610_; 
wire _abc_40298_new_n1611_; 
wire _abc_40298_new_n1612_; 
wire _abc_40298_new_n1613_; 
wire _abc_40298_new_n1614_; 
wire _abc_40298_new_n1615_; 
wire _abc_40298_new_n1616_; 
wire _abc_40298_new_n1617_; 
wire _abc_40298_new_n1618_; 
wire _abc_40298_new_n1620_; 
wire _abc_40298_new_n1621_; 
wire _abc_40298_new_n1622_; 
wire _abc_40298_new_n1623_; 
wire _abc_40298_new_n1624_; 
wire _abc_40298_new_n1625_; 
wire _abc_40298_new_n1626_; 
wire _abc_40298_new_n1627_; 
wire _abc_40298_new_n1628_; 
wire _abc_40298_new_n1629_; 
wire _abc_40298_new_n1630_; 
wire _abc_40298_new_n1631_; 
wire _abc_40298_new_n1632_; 
wire _abc_40298_new_n1633_; 
wire _abc_40298_new_n1634_; 
wire _abc_40298_new_n1635_; 
wire _abc_40298_new_n1636_; 
wire _abc_40298_new_n1637_; 
wire _abc_40298_new_n1638_; 
wire _abc_40298_new_n1639_; 
wire _abc_40298_new_n1640_; 
wire _abc_40298_new_n1641_; 
wire _abc_40298_new_n1642_; 
wire _abc_40298_new_n1644_; 
wire _abc_40298_new_n1645_; 
wire _abc_40298_new_n1646_; 
wire _abc_40298_new_n1647_; 
wire _abc_40298_new_n1648_; 
wire _abc_40298_new_n1649_; 
wire _abc_40298_new_n1650_; 
wire _abc_40298_new_n1651_; 
wire _abc_40298_new_n1652_; 
wire _abc_40298_new_n1653_; 
wire _abc_40298_new_n1654_; 
wire _abc_40298_new_n1655_; 
wire _abc_40298_new_n1656_; 
wire _abc_40298_new_n1657_; 
wire _abc_40298_new_n1658_; 
wire _abc_40298_new_n1659_; 
wire _abc_40298_new_n1660_; 
wire _abc_40298_new_n1661_; 
wire _abc_40298_new_n1662_; 
wire _abc_40298_new_n1663_; 
wire _abc_40298_new_n1664_; 
wire _abc_40298_new_n1665_; 
wire _abc_40298_new_n1666_; 
wire _abc_40298_new_n1667_; 
wire _abc_40298_new_n1668_; 
wire _abc_40298_new_n1669_; 
wire _abc_40298_new_n1670_; 
wire _abc_40298_new_n1671_; 
wire _abc_40298_new_n1672_; 
wire _abc_40298_new_n1674_; 
wire _abc_40298_new_n1675_; 
wire _abc_40298_new_n1676_; 
wire _abc_40298_new_n1677_; 
wire _abc_40298_new_n1678_; 
wire _abc_40298_new_n1679_; 
wire _abc_40298_new_n1680_; 
wire _abc_40298_new_n1681_; 
wire _abc_40298_new_n1682_; 
wire _abc_40298_new_n1683_; 
wire _abc_40298_new_n1684_; 
wire _abc_40298_new_n1685_; 
wire _abc_40298_new_n1686_; 
wire _abc_40298_new_n1687_; 
wire _abc_40298_new_n1688_; 
wire _abc_40298_new_n1689_; 
wire _abc_40298_new_n1690_; 
wire _abc_40298_new_n1691_; 
wire _abc_40298_new_n1692_; 
wire _abc_40298_new_n1693_; 
wire _abc_40298_new_n1694_; 
wire _abc_40298_new_n1695_; 
wire _abc_40298_new_n1697_; 
wire _abc_40298_new_n1698_; 
wire _abc_40298_new_n1699_; 
wire _abc_40298_new_n1700_; 
wire _abc_40298_new_n1701_; 
wire _abc_40298_new_n1702_; 
wire _abc_40298_new_n1703_; 
wire _abc_40298_new_n1704_; 
wire _abc_40298_new_n1705_; 
wire _abc_40298_new_n1706_; 
wire _abc_40298_new_n1707_; 
wire _abc_40298_new_n1708_; 
wire _abc_40298_new_n1709_; 
wire _abc_40298_new_n1710_; 
wire _abc_40298_new_n1711_; 
wire _abc_40298_new_n1712_; 
wire _abc_40298_new_n1713_; 
wire _abc_40298_new_n1714_; 
wire _abc_40298_new_n1715_; 
wire _abc_40298_new_n1716_; 
wire _abc_40298_new_n1717_; 
wire _abc_40298_new_n1718_; 
wire _abc_40298_new_n1719_; 
wire _abc_40298_new_n1720_; 
wire _abc_40298_new_n1721_; 
wire _abc_40298_new_n1722_; 
wire _abc_40298_new_n1723_; 
wire _abc_40298_new_n1724_; 
wire _abc_40298_new_n1726_; 
wire _abc_40298_new_n1727_; 
wire _abc_40298_new_n1728_; 
wire _abc_40298_new_n1729_; 
wire _abc_40298_new_n1730_; 
wire _abc_40298_new_n1731_; 
wire _abc_40298_new_n1732_; 
wire _abc_40298_new_n1733_; 
wire _abc_40298_new_n1734_; 
wire _abc_40298_new_n1735_; 
wire _abc_40298_new_n1736_; 
wire _abc_40298_new_n1737_; 
wire _abc_40298_new_n1738_; 
wire _abc_40298_new_n1739_; 
wire _abc_40298_new_n1740_; 
wire _abc_40298_new_n1741_; 
wire _abc_40298_new_n1742_; 
wire _abc_40298_new_n1743_; 
wire _abc_40298_new_n1744_; 
wire _abc_40298_new_n1745_; 
wire _abc_40298_new_n1746_; 
wire _abc_40298_new_n1747_; 
wire _abc_40298_new_n1748_; 
wire _abc_40298_new_n1749_; 
wire _abc_40298_new_n1750_; 
wire _abc_40298_new_n1751_; 
wire _abc_40298_new_n1753_; 
wire _abc_40298_new_n1754_; 
wire _abc_40298_new_n1755_; 
wire _abc_40298_new_n1756_; 
wire _abc_40298_new_n1757_; 
wire _abc_40298_new_n1758_; 
wire _abc_40298_new_n1759_; 
wire _abc_40298_new_n1760_; 
wire _abc_40298_new_n1761_; 
wire _abc_40298_new_n1762_; 
wire _abc_40298_new_n1763_; 
wire _abc_40298_new_n1764_; 
wire _abc_40298_new_n1765_; 
wire _abc_40298_new_n1766_; 
wire _abc_40298_new_n1767_; 
wire _abc_40298_new_n1768_; 
wire _abc_40298_new_n1769_; 
wire _abc_40298_new_n1770_; 
wire _abc_40298_new_n1771_; 
wire _abc_40298_new_n1772_; 
wire _abc_40298_new_n1773_; 
wire _abc_40298_new_n1774_; 
wire _abc_40298_new_n1775_; 
wire _abc_40298_new_n1776_; 
wire _abc_40298_new_n1777_; 
wire _abc_40298_new_n1778_; 
wire _abc_40298_new_n1779_; 
wire _abc_40298_new_n1780_; 
wire _abc_40298_new_n1782_; 
wire _abc_40298_new_n1783_; 
wire _abc_40298_new_n1784_; 
wire _abc_40298_new_n1785_; 
wire _abc_40298_new_n1786_; 
wire _abc_40298_new_n1787_; 
wire _abc_40298_new_n1788_; 
wire _abc_40298_new_n1789_; 
wire _abc_40298_new_n1790_; 
wire _abc_40298_new_n1791_; 
wire _abc_40298_new_n1792_; 
wire _abc_40298_new_n1793_; 
wire _abc_40298_new_n1794_; 
wire _abc_40298_new_n1795_; 
wire _abc_40298_new_n1796_; 
wire _abc_40298_new_n1797_; 
wire _abc_40298_new_n1798_; 
wire _abc_40298_new_n1799_; 
wire _abc_40298_new_n1800_; 
wire _abc_40298_new_n1801_; 
wire _abc_40298_new_n1802_; 
wire _abc_40298_new_n1803_; 
wire _abc_40298_new_n1805_; 
wire _abc_40298_new_n1806_; 
wire _abc_40298_new_n1807_; 
wire _abc_40298_new_n1808_; 
wire _abc_40298_new_n1809_; 
wire _abc_40298_new_n1810_; 
wire _abc_40298_new_n1811_; 
wire _abc_40298_new_n1812_; 
wire _abc_40298_new_n1813_; 
wire _abc_40298_new_n1814_; 
wire _abc_40298_new_n1815_; 
wire _abc_40298_new_n1816_; 
wire _abc_40298_new_n1817_; 
wire _abc_40298_new_n1818_; 
wire _abc_40298_new_n1819_; 
wire _abc_40298_new_n1820_; 
wire _abc_40298_new_n1821_; 
wire _abc_40298_new_n1822_; 
wire _abc_40298_new_n1823_; 
wire _abc_40298_new_n1824_; 
wire _abc_40298_new_n1825_; 
wire _abc_40298_new_n1826_; 
wire _abc_40298_new_n1827_; 
wire _abc_40298_new_n1828_; 
wire _abc_40298_new_n1829_; 
wire _abc_40298_new_n1830_; 
wire _abc_40298_new_n1831_; 
wire _abc_40298_new_n1832_; 
wire _abc_40298_new_n1833_; 
wire _abc_40298_new_n1834_; 
wire _abc_40298_new_n1835_; 
wire _abc_40298_new_n1836_; 
wire _abc_40298_new_n1837_; 
wire _abc_40298_new_n1838_; 
wire _abc_40298_new_n1839_; 
wire _abc_40298_new_n1841_; 
wire _abc_40298_new_n1842_; 
wire _abc_40298_new_n1843_; 
wire _abc_40298_new_n1844_; 
wire _abc_40298_new_n1845_; 
wire _abc_40298_new_n1846_; 
wire _abc_40298_new_n1847_; 
wire _abc_40298_new_n1848_; 
wire _abc_40298_new_n1849_; 
wire _abc_40298_new_n1850_; 
wire _abc_40298_new_n1851_; 
wire _abc_40298_new_n1852_; 
wire _abc_40298_new_n1853_; 
wire _abc_40298_new_n1854_; 
wire _abc_40298_new_n1855_; 
wire _abc_40298_new_n1856_; 
wire _abc_40298_new_n1857_; 
wire _abc_40298_new_n1858_; 
wire _abc_40298_new_n1859_; 
wire _abc_40298_new_n1860_; 
wire _abc_40298_new_n1862_; 
wire _abc_40298_new_n1863_; 
wire _abc_40298_new_n1864_; 
wire _abc_40298_new_n1865_; 
wire _abc_40298_new_n1866_; 
wire _abc_40298_new_n1867_; 
wire _abc_40298_new_n1868_; 
wire _abc_40298_new_n1869_; 
wire _abc_40298_new_n1870_; 
wire _abc_40298_new_n1871_; 
wire _abc_40298_new_n1872_; 
wire _abc_40298_new_n1873_; 
wire _abc_40298_new_n1874_; 
wire _abc_40298_new_n1875_; 
wire _abc_40298_new_n1876_; 
wire _abc_40298_new_n1877_; 
wire _abc_40298_new_n1878_; 
wire _abc_40298_new_n1879_; 
wire _abc_40298_new_n1880_; 
wire _abc_40298_new_n1881_; 
wire _abc_40298_new_n1882_; 
wire _abc_40298_new_n1883_; 
wire _abc_40298_new_n1884_; 
wire _abc_40298_new_n1885_; 
wire _abc_40298_new_n1886_; 
wire _abc_40298_new_n1887_; 
wire _abc_40298_new_n1888_; 
wire _abc_40298_new_n1889_; 
wire _abc_40298_new_n1891_; 
wire _abc_40298_new_n1892_; 
wire _abc_40298_new_n1893_; 
wire _abc_40298_new_n1894_; 
wire _abc_40298_new_n1895_; 
wire _abc_40298_new_n1896_; 
wire _abc_40298_new_n1897_; 
wire _abc_40298_new_n1898_; 
wire _abc_40298_new_n1899_; 
wire _abc_40298_new_n1900_; 
wire _abc_40298_new_n1901_; 
wire _abc_40298_new_n1902_; 
wire _abc_40298_new_n1903_; 
wire _abc_40298_new_n1904_; 
wire _abc_40298_new_n1905_; 
wire _abc_40298_new_n1906_; 
wire _abc_40298_new_n1907_; 
wire _abc_40298_new_n1908_; 
wire _abc_40298_new_n1909_; 
wire _abc_40298_new_n1911_; 
wire _abc_40298_new_n1912_; 
wire _abc_40298_new_n1913_; 
wire _abc_40298_new_n1914_; 
wire _abc_40298_new_n1915_; 
wire _abc_40298_new_n1916_; 
wire _abc_40298_new_n1917_; 
wire _abc_40298_new_n1918_; 
wire _abc_40298_new_n1919_; 
wire _abc_40298_new_n1920_; 
wire _abc_40298_new_n1921_; 
wire _abc_40298_new_n1922_; 
wire _abc_40298_new_n1923_; 
wire _abc_40298_new_n1924_; 
wire _abc_40298_new_n1925_; 
wire _abc_40298_new_n1926_; 
wire _abc_40298_new_n1927_; 
wire _abc_40298_new_n1928_; 
wire _abc_40298_new_n1929_; 
wire _abc_40298_new_n1930_; 
wire _abc_40298_new_n1931_; 
wire _abc_40298_new_n1932_; 
wire _abc_40298_new_n1933_; 
wire _abc_40298_new_n1934_; 
wire _abc_40298_new_n1935_; 
wire _abc_40298_new_n1936_; 
wire _abc_40298_new_n1937_; 
wire _abc_40298_new_n1938_; 
wire _abc_40298_new_n1939_; 
wire _abc_40298_new_n1941_; 
wire _abc_40298_new_n1942_; 
wire _abc_40298_new_n1943_; 
wire _abc_40298_new_n1944_; 
wire _abc_40298_new_n1945_; 
wire _abc_40298_new_n1946_; 
wire _abc_40298_new_n1947_; 
wire _abc_40298_new_n1948_; 
wire _abc_40298_new_n1949_; 
wire _abc_40298_new_n1950_; 
wire _abc_40298_new_n1951_; 
wire _abc_40298_new_n1952_; 
wire _abc_40298_new_n1953_; 
wire _abc_40298_new_n1954_; 
wire _abc_40298_new_n1955_; 
wire _abc_40298_new_n1956_; 
wire _abc_40298_new_n1957_; 
wire _abc_40298_new_n1958_; 
wire _abc_40298_new_n1960_; 
wire _abc_40298_new_n1961_; 
wire _abc_40298_new_n1962_; 
wire _abc_40298_new_n1963_; 
wire _abc_40298_new_n1964_; 
wire _abc_40298_new_n1965_; 
wire _abc_40298_new_n1966_; 
wire _abc_40298_new_n1967_; 
wire _abc_40298_new_n1968_; 
wire _abc_40298_new_n1969_; 
wire _abc_40298_new_n1970_; 
wire _abc_40298_new_n1971_; 
wire _abc_40298_new_n1972_; 
wire _abc_40298_new_n1973_; 
wire _abc_40298_new_n1974_; 
wire _abc_40298_new_n1975_; 
wire _abc_40298_new_n1976_; 
wire _abc_40298_new_n1977_; 
wire _abc_40298_new_n1978_; 
wire _abc_40298_new_n1979_; 
wire _abc_40298_new_n1980_; 
wire _abc_40298_new_n1981_; 
wire _abc_40298_new_n1982_; 
wire _abc_40298_new_n1983_; 
wire _abc_40298_new_n1984_; 
wire _abc_40298_new_n1985_; 
wire _abc_40298_new_n1986_; 
wire _abc_40298_new_n1987_; 
wire _abc_40298_new_n1989_; 
wire _abc_40298_new_n1990_; 
wire _abc_40298_new_n1991_; 
wire _abc_40298_new_n1992_; 
wire _abc_40298_new_n1993_; 
wire _abc_40298_new_n1994_; 
wire _abc_40298_new_n1995_; 
wire _abc_40298_new_n1996_; 
wire _abc_40298_new_n1997_; 
wire _abc_40298_new_n1998_; 
wire _abc_40298_new_n1999_; 
wire _abc_40298_new_n2000_; 
wire _abc_40298_new_n2001_; 
wire _abc_40298_new_n2002_; 
wire _abc_40298_new_n2003_; 
wire _abc_40298_new_n2004_; 
wire _abc_40298_new_n2005_; 
wire _abc_40298_new_n2006_; 
wire _abc_40298_new_n2007_; 
wire _abc_40298_new_n2008_; 
wire _abc_40298_new_n2009_; 
wire _abc_40298_new_n2010_; 
wire _abc_40298_new_n2011_; 
wire _abc_40298_new_n2012_; 
wire _abc_40298_new_n2014_; 
wire _abc_40298_new_n2015_; 
wire _abc_40298_new_n2016_; 
wire _abc_40298_new_n2018_; 
wire _abc_40298_new_n2019_; 
wire _abc_40298_new_n2021_; 
wire _abc_40298_new_n2022_; 
wire _abc_40298_new_n2024_; 
wire _abc_40298_new_n2025_; 
wire _abc_40298_new_n2026_; 
wire _abc_40298_new_n2028_; 
wire _abc_40298_new_n2029_; 
wire _abc_40298_new_n2031_; 
wire _abc_40298_new_n2032_; 
wire _abc_40298_new_n2034_; 
wire _abc_40298_new_n2035_; 
wire _abc_40298_new_n2037_; 
wire _abc_40298_new_n2038_; 
wire _abc_40298_new_n2040_; 
wire _abc_40298_new_n2041_; 
wire _abc_40298_new_n2043_; 
wire _abc_40298_new_n2044_; 
wire _abc_40298_new_n2045_; 
wire _abc_40298_new_n2046_; 
wire _abc_40298_new_n2047_; 
wire _abc_40298_new_n2049_; 
wire _abc_40298_new_n2050_; 
wire _abc_40298_new_n2051_; 
wire _abc_40298_new_n2052_; 
wire _abc_40298_new_n2054_; 
wire _abc_40298_new_n2055_; 
wire _abc_40298_new_n2056_; 
wire _abc_40298_new_n2058_; 
wire _abc_40298_new_n2059_; 
wire _abc_40298_new_n2061_; 
wire _abc_40298_new_n2062_; 
wire _abc_40298_new_n2064_; 
wire _abc_40298_new_n2065_; 
wire _abc_40298_new_n2067_; 
wire _abc_40298_new_n2068_; 
wire _abc_40298_new_n2070_; 
wire _abc_40298_new_n2071_; 
wire _abc_40298_new_n2073_; 
wire _abc_40298_new_n2074_; 
wire _abc_40298_new_n2076_; 
wire _abc_40298_new_n2077_; 
wire _abc_40298_new_n2079_; 
wire _abc_40298_new_n2080_; 
wire _abc_40298_new_n2082_; 
wire _abc_40298_new_n2083_; 
wire _abc_40298_new_n2085_; 
wire _abc_40298_new_n2086_; 
wire _abc_40298_new_n2088_; 
wire _abc_40298_new_n2089_; 
wire _abc_40298_new_n2091_; 
wire _abc_40298_new_n2092_; 
wire _abc_40298_new_n2094_; 
wire _abc_40298_new_n2095_; 
wire _abc_40298_new_n2097_; 
wire _abc_40298_new_n2098_; 
wire _abc_40298_new_n2100_; 
wire _abc_40298_new_n2101_; 
wire _abc_40298_new_n2103_; 
wire _abc_40298_new_n2104_; 
wire _abc_40298_new_n2106_; 
wire _abc_40298_new_n2107_; 
wire _abc_40298_new_n2109_; 
wire _abc_40298_new_n2110_; 
wire _abc_40298_new_n2112_; 
wire _abc_40298_new_n2113_; 
wire _abc_40298_new_n2115_; 
wire _abc_40298_new_n2116_; 
wire _abc_40298_new_n2117_; 
wire _abc_40298_new_n2119_; 
wire _abc_40298_new_n2120_; 
wire _abc_40298_new_n2121_; 
wire _abc_40298_new_n2122_; 
wire _abc_40298_new_n2123_; 
wire _abc_40298_new_n2124_; 
wire _abc_40298_new_n2125_; 
wire _abc_40298_new_n2126_; 
wire _abc_40298_new_n2127_; 
wire _abc_40298_new_n2128_; 
wire _abc_40298_new_n2129_; 
wire _abc_40298_new_n2130_; 
wire _abc_40298_new_n2132_; 
wire _abc_40298_new_n2134_; 
wire _abc_40298_new_n2137_; 
wire _abc_40298_new_n2139_; 
wire _abc_40298_new_n2140_; 
wire _abc_40298_new_n2141_; 
wire _abc_40298_new_n2142_; 
wire _abc_40298_new_n2143_; 
wire _abc_40298_new_n2144_; 
wire _abc_40298_new_n2145_; 
wire _abc_40298_new_n2146_; 
wire _abc_40298_new_n2147_; 
wire _abc_40298_new_n2148_; 
wire _abc_40298_new_n2149_; 
wire _abc_40298_new_n2150_; 
wire _abc_40298_new_n2151_; 
wire _abc_40298_new_n2153_; 
wire _abc_40298_new_n2159_; 
wire _abc_40298_new_n2160_; 
wire _abc_40298_new_n2161_; 
wire _abc_40298_new_n2162_; 
wire _abc_40298_new_n2163_; 
wire _abc_40298_new_n2164_; 
wire _abc_40298_new_n2165_; 
wire _abc_40298_new_n2166_; 
wire _abc_40298_new_n2167_; 
wire _abc_40298_new_n2168_; 
wire _abc_40298_new_n2169_; 
wire _abc_40298_new_n2170_; 
wire _abc_40298_new_n2171_; 
wire _abc_40298_new_n2172_; 
wire _abc_40298_new_n2173_; 
wire _abc_40298_new_n2174_; 
wire _abc_40298_new_n2175_; 
wire _abc_40298_new_n2176_; 
wire _abc_40298_new_n2178_; 
wire _abc_40298_new_n2180_; 
wire _abc_40298_new_n2182_; 
wire _abc_40298_new_n2184_; 
wire _abc_40298_new_n2186_; 
wire _abc_40298_new_n2188_; 
wire _abc_40298_new_n2190_; 
wire _abc_40298_new_n2191_; 
wire _abc_40298_new_n2193_; 
wire _abc_40298_new_n2194_; 
wire _abc_40298_new_n2196_; 
wire _abc_40298_new_n2197_; 
wire _abc_40298_new_n2198_; 
wire _abc_40298_new_n2199_; 
wire _abc_40298_new_n2200_; 
wire _abc_40298_new_n2202_; 
wire _abc_40298_new_n2203_; 
wire _abc_40298_new_n2204_; 
wire _abc_40298_new_n2205_; 
wire _abc_40298_new_n2206_; 
wire _abc_40298_new_n2207_; 
wire _abc_40298_new_n2208_; 
wire _abc_40298_new_n2209_; 
wire _abc_40298_new_n2211_; 
wire _abc_40298_new_n2212_; 
wire _abc_40298_new_n2213_; 
wire _abc_40298_new_n2214_; 
wire _abc_40298_new_n2216_; 
wire _abc_40298_new_n2217_; 
wire _abc_40298_new_n2218_; 
wire _abc_40298_new_n2219_; 
wire _abc_40298_new_n2221_; 
wire _abc_40298_new_n2222_; 
wire _abc_40298_new_n2223_; 
wire _abc_40298_new_n2224_; 
wire _abc_40298_new_n2226_; 
wire _abc_40298_new_n2227_; 
wire _abc_40298_new_n2228_; 
wire _abc_40298_new_n2229_; 
wire _abc_40298_new_n2231_; 
wire _abc_40298_new_n2232_; 
wire _abc_40298_new_n2233_; 
wire _abc_40298_new_n2234_; 
wire _abc_40298_new_n2236_; 
wire _abc_40298_new_n2237_; 
wire _abc_40298_new_n2238_; 
wire _abc_40298_new_n2239_; 
wire _abc_40298_new_n2241_; 
wire _abc_40298_new_n2242_; 
wire _abc_40298_new_n2243_; 
wire _abc_40298_new_n2244_; 
wire _abc_40298_new_n2246_; 
wire _abc_40298_new_n2247_; 
wire _abc_40298_new_n2248_; 
wire _abc_40298_new_n2250_; 
wire _abc_40298_new_n2251_; 
wire _abc_40298_new_n2252_; 
wire _abc_40298_new_n2254_; 
wire _abc_40298_new_n2255_; 
wire _abc_40298_new_n2256_; 
wire _abc_40298_new_n2258_; 
wire _abc_40298_new_n2259_; 
wire _abc_40298_new_n2260_; 
wire _abc_40298_new_n2261_; 
wire _abc_40298_new_n2263_; 
wire _abc_40298_new_n2264_; 
wire _abc_40298_new_n2265_; 
wire _abc_40298_new_n2266_; 
wire _abc_40298_new_n2268_; 
wire _abc_40298_new_n2269_; 
wire _abc_40298_new_n2270_; 
wire _abc_40298_new_n2272_; 
wire _abc_40298_new_n2273_; 
wire _abc_40298_new_n2274_; 
wire _abc_40298_new_n2276_; 
wire _abc_40298_new_n2277_; 
wire _abc_40298_new_n2278_; 
wire _abc_40298_new_n2280_; 
wire _abc_40298_new_n2281_; 
wire _abc_40298_new_n2282_; 
wire _abc_40298_new_n2283_; 
wire _abc_40298_new_n2284_; 
wire _abc_40298_new_n2285_; 
wire _abc_40298_new_n2286_; 
wire _abc_40298_new_n2287_; 
wire _abc_40298_new_n2288_; 
wire _abc_40298_new_n2289_; 
wire _abc_40298_new_n2290_; 
wire _abc_40298_new_n2292_; 
wire _abc_40298_new_n2293_; 
wire _abc_40298_new_n2294_; 
wire _abc_40298_new_n2295_; 
wire _abc_40298_new_n2296_; 
wire _abc_40298_new_n2297_; 
wire _abc_40298_new_n2299_; 
wire _abc_40298_new_n2300_; 
wire _abc_40298_new_n2301_; 
wire _abc_40298_new_n2302_; 
wire _abc_40298_new_n2303_; 
wire _abc_40298_new_n2304_; 
wire _abc_40298_new_n2305_; 
wire _abc_40298_new_n2307_; 
wire _abc_40298_new_n2308_; 
wire _abc_40298_new_n2309_; 
wire _abc_40298_new_n2310_; 
wire _abc_40298_new_n2311_; 
wire _abc_40298_new_n2312_; 
wire _abc_40298_new_n2314_; 
wire _abc_40298_new_n2315_; 
wire _abc_40298_new_n2316_; 
wire _abc_40298_new_n2317_; 
wire _abc_40298_new_n2318_; 
wire _abc_40298_new_n2319_; 
wire _abc_40298_new_n2321_; 
wire _abc_40298_new_n2322_; 
wire _abc_40298_new_n2323_; 
wire _abc_40298_new_n2324_; 
wire _abc_40298_new_n2325_; 
wire _abc_40298_new_n2327_; 
wire _abc_40298_new_n2328_; 
wire _abc_40298_new_n2329_; 
wire _abc_40298_new_n2330_; 
wire _abc_40298_new_n2331_; 
wire _abc_40298_new_n2332_; 
wire _abc_40298_new_n2334_; 
wire _abc_40298_new_n2335_; 
wire _abc_40298_new_n2336_; 
wire _abc_40298_new_n2337_; 
wire _abc_40298_new_n2338_; 
wire _abc_40298_new_n2339_; 
wire _abc_40298_new_n2340_; 
wire _abc_40298_new_n2342_; 
wire _abc_40298_new_n2343_; 
wire _abc_40298_new_n2344_; 
wire _abc_40298_new_n2345_; 
wire _abc_40298_new_n2346_; 
wire _abc_40298_new_n2347_; 
wire _abc_40298_new_n2349_; 
wire _abc_40298_new_n2350_; 
wire _abc_40298_new_n2351_; 
wire _abc_40298_new_n2352_; 
wire _abc_40298_new_n2353_; 
wire _abc_40298_new_n2354_; 
wire _abc_40298_new_n2355_; 
wire _abc_40298_new_n2356_; 
wire _abc_40298_new_n2358_; 
wire _abc_40298_new_n2359_; 
wire _abc_40298_new_n2360_; 
wire _abc_40298_new_n2361_; 
wire _abc_40298_new_n2362_; 
wire _abc_40298_new_n2364_; 
wire _abc_40298_new_n2365_; 
wire _abc_40298_new_n2366_; 
wire _abc_40298_new_n2367_; 
wire _abc_40298_new_n2369_; 
wire _abc_40298_new_n2370_; 
wire _abc_40298_new_n2371_; 
wire _abc_40298_new_n2373_; 
wire _abc_40298_new_n2374_; 
wire _abc_40298_new_n2375_; 
wire _abc_40298_new_n2377_; 
wire _abc_40298_new_n2378_; 
wire _abc_40298_new_n2379_; 
wire _abc_40298_new_n2381_; 
wire _abc_40298_new_n2382_; 
wire _abc_40298_new_n2383_; 
wire _abc_40298_new_n2385_; 
wire _abc_40298_new_n2386_; 
wire _abc_40298_new_n2387_; 
wire _abc_40298_new_n2388_; 
wire _abc_40298_new_n2389_; 
wire _abc_40298_new_n2390_; 
wire _abc_40298_new_n2392_; 
wire _abc_40298_new_n2393_; 
wire _abc_40298_new_n2394_; 
wire _abc_40298_new_n2395_; 
wire _abc_40298_new_n2396_; 
wire _abc_40298_new_n2397_; 
wire _abc_40298_new_n2399_; 
wire _abc_40298_new_n2400_; 
wire _abc_40298_new_n2401_; 
wire _abc_40298_new_n2402_; 
wire _abc_40298_new_n2403_; 
wire _abc_40298_new_n2404_; 
wire _abc_40298_new_n2406_; 
wire _abc_40298_new_n2407_; 
wire _abc_40298_new_n2408_; 
wire _abc_40298_new_n2409_; 
wire _abc_40298_new_n2410_; 
wire _abc_40298_new_n2411_; 
wire _abc_40298_new_n2413_; 
wire _abc_40298_new_n2414_; 
wire _abc_40298_new_n2415_; 
wire _abc_40298_new_n2416_; 
wire _abc_40298_new_n2417_; 
wire _abc_40298_new_n2418_; 
wire _abc_40298_new_n2420_; 
wire _abc_40298_new_n2421_; 
wire _abc_40298_new_n2422_; 
wire _abc_40298_new_n2423_; 
wire _abc_40298_new_n2424_; 
wire _abc_40298_new_n2425_; 
wire _abc_40298_new_n2427_; 
wire _abc_40298_new_n2428_; 
wire _abc_40298_new_n2429_; 
wire _abc_40298_new_n2430_; 
wire _abc_40298_new_n2431_; 
wire _abc_40298_new_n2432_; 
wire _abc_40298_new_n2434_; 
wire _abc_40298_new_n2435_; 
wire _abc_40298_new_n2436_; 
wire _abc_40298_new_n2437_; 
wire _abc_40298_new_n2438_; 
wire _abc_40298_new_n2439_; 
wire _abc_40298_new_n2441_; 
wire _abc_40298_new_n2442_; 
wire _abc_40298_new_n2443_; 
wire _abc_40298_new_n2444_; 
wire _abc_40298_new_n2445_; 
wire _abc_40298_new_n2446_; 
wire _abc_40298_new_n2448_; 
wire _abc_40298_new_n2449_; 
wire _abc_40298_new_n2450_; 
wire _abc_40298_new_n2451_; 
wire _abc_40298_new_n2452_; 
wire _abc_40298_new_n2453_; 
wire _abc_40298_new_n2455_; 
wire _abc_40298_new_n2456_; 
wire _abc_40298_new_n2457_; 
wire _abc_40298_new_n2458_; 
wire _abc_40298_new_n2459_; 
wire _abc_40298_new_n2460_; 
wire _abc_40298_new_n2461_; 
wire _abc_40298_new_n2463_; 
wire _abc_40298_new_n2464_; 
wire _abc_40298_new_n2465_; 
wire _abc_40298_new_n2466_; 
wire _abc_40298_new_n2467_; 
wire _abc_40298_new_n2468_; 
wire _abc_40298_new_n2470_; 
wire _abc_40298_new_n2471_; 
wire _abc_40298_new_n2472_; 
wire _abc_40298_new_n2473_; 
wire _abc_40298_new_n2474_; 
wire _abc_40298_new_n2475_; 
wire _abc_40298_new_n2476_; 
wire _abc_40298_new_n2478_; 
wire _abc_40298_new_n2479_; 
wire _abc_40298_new_n2480_; 
wire _abc_40298_new_n2481_; 
wire _abc_40298_new_n2482_; 
wire _abc_40298_new_n2483_; 
wire _abc_40298_new_n2484_; 
wire _abc_40298_new_n2486_; 
wire _abc_40298_new_n2487_; 
wire _abc_40298_new_n2488_; 
wire _abc_40298_new_n2489_; 
wire _abc_40298_new_n2490_; 
wire _abc_40298_new_n2491_; 
wire _abc_40298_new_n2493_; 
wire _abc_40298_new_n2494_; 
wire _abc_40298_new_n2495_; 
wire _abc_40298_new_n2496_; 
wire _abc_40298_new_n2497_; 
wire _abc_40298_new_n2498_; 
wire _abc_40298_new_n2500_; 
wire _abc_40298_new_n2501_; 
wire _abc_40298_new_n2502_; 
wire _abc_40298_new_n2503_; 
wire _abc_40298_new_n2505_; 
wire _abc_40298_new_n2506_; 
wire _abc_40298_new_n2507_; 
wire _abc_40298_new_n2510_; 
wire _abc_40298_new_n2511_; 
wire _abc_40298_new_n2513_; 
wire _abc_40298_new_n2514_; 
wire _abc_40298_new_n2515_; 
wire _abc_40298_new_n2516_; 
wire _abc_40298_new_n2518_; 
wire _abc_40298_new_n2519_; 
wire _abc_40298_new_n2520_; 
wire _abc_40298_new_n2521_; 
wire _abc_40298_new_n2522_; 
wire _abc_40298_new_n2524_; 
wire _abc_40298_new_n2530_; 
wire _abc_40298_new_n2532_; 
wire _abc_40298_new_n2535_; 
wire _abc_40298_new_n2537_; 
wire _abc_40298_new_n2542_; 
wire _abc_40298_new_n2544_; 
wire _abc_40298_new_n2547_; 
wire _abc_40298_new_n2559_; 
wire _abc_40298_new_n2562_; 
wire _abc_40298_new_n2567_; 
wire _abc_40298_new_n2568_; 
wire _abc_40298_new_n2569_; 
wire _abc_40298_new_n2570_; 
wire _abc_40298_new_n2571_; 
wire _abc_40298_new_n2572_; 
wire _abc_40298_new_n2573_; 
wire _abc_40298_new_n2574_; 
wire _abc_40298_new_n2575_; 
wire _abc_40298_new_n2576_; 
wire _abc_40298_new_n2577_; 
wire _abc_40298_new_n2578_; 
wire _abc_40298_new_n2579_; 
wire _abc_40298_new_n2580_; 
wire _abc_40298_new_n2581_; 
wire _abc_40298_new_n2582_; 
wire _abc_40298_new_n2584_; 
wire _abc_40298_new_n2585_; 
wire _abc_40298_new_n2586_; 
wire _abc_40298_new_n2587_; 
wire _abc_40298_new_n2588_; 
wire _abc_40298_new_n2589_; 
wire _abc_40298_new_n2590_; 
wire _abc_40298_new_n2592_; 
wire _abc_40298_new_n2593_; 
wire _abc_40298_new_n2594_; 
wire _abc_40298_new_n2595_; 
wire _abc_40298_new_n2596_; 
wire _abc_40298_new_n2597_; 
wire _abc_40298_new_n2598_; 
wire _abc_40298_new_n2600_; 
wire _abc_40298_new_n2601_; 
wire _abc_40298_new_n2602_; 
wire _abc_40298_new_n2603_; 
wire _abc_40298_new_n2604_; 
wire _abc_40298_new_n2605_; 
wire _abc_40298_new_n2607_; 
wire _abc_40298_new_n2608_; 
wire _abc_40298_new_n2609_; 
wire _abc_40298_new_n2610_; 
wire _abc_40298_new_n2611_; 
wire _abc_40298_new_n2612_; 
wire _abc_40298_new_n2613_; 
wire _abc_40298_new_n2614_; 
wire _abc_40298_new_n2615_; 
wire _abc_40298_new_n2616_; 
wire _abc_40298_new_n2618_; 
wire _abc_40298_new_n2619_; 
wire _abc_40298_new_n2620_; 
wire _abc_40298_new_n2621_; 
wire _abc_40298_new_n2622_; 
wire _abc_40298_new_n2623_; 
wire _abc_40298_new_n2624_; 
wire _abc_40298_new_n2626_; 
wire _abc_40298_new_n2627_; 
wire _abc_40298_new_n2628_; 
wire _abc_40298_new_n2629_; 
wire _abc_40298_new_n2630_; 
wire _abc_40298_new_n2631_; 
wire _abc_40298_new_n2632_; 
wire _abc_40298_new_n2634_; 
wire _abc_40298_new_n2635_; 
wire _abc_40298_new_n2636_; 
wire _abc_40298_new_n2637_; 
wire _abc_40298_new_n2638_; 
wire _abc_40298_new_n2639_; 
wire _abc_40298_new_n2640_; 
wire _abc_40298_new_n2642_; 
wire _abc_40298_new_n2643_; 
wire _abc_40298_new_n2644_; 
wire _abc_40298_new_n2645_; 
wire _abc_40298_new_n2646_; 
wire _abc_40298_new_n2647_; 
wire _abc_40298_new_n2648_; 
wire _abc_40298_new_n2650_; 
wire _abc_40298_new_n2651_; 
wire _abc_40298_new_n2652_; 
wire _abc_40298_new_n2653_; 
wire _abc_40298_new_n2654_; 
wire _abc_40298_new_n2655_; 
wire _abc_40298_new_n2656_; 
wire _abc_40298_new_n2658_; 
wire _abc_40298_new_n2659_; 
wire _abc_40298_new_n2660_; 
wire _abc_40298_new_n2661_; 
wire _abc_40298_new_n2662_; 
wire _abc_40298_new_n2663_; 
wire _abc_40298_new_n2664_; 
wire _abc_40298_new_n2666_; 
wire _abc_40298_new_n2667_; 
wire _abc_40298_new_n2668_; 
wire _abc_40298_new_n2669_; 
wire _abc_40298_new_n2670_; 
wire _abc_40298_new_n2671_; 
wire _abc_40298_new_n2672_; 
wire _abc_40298_new_n2674_; 
wire _abc_40298_new_n2675_; 
wire _abc_40298_new_n2676_; 
wire _abc_40298_new_n2677_; 
wire _abc_40298_new_n2678_; 
wire _abc_40298_new_n2679_; 
wire _abc_40298_new_n2680_; 
wire _abc_40298_new_n2681_; 
wire _abc_40298_new_n2683_; 
wire _abc_40298_new_n2684_; 
wire _abc_40298_new_n2685_; 
wire _abc_40298_new_n2686_; 
wire _abc_40298_new_n2687_; 
wire _abc_40298_new_n2688_; 
wire _abc_40298_new_n2689_; 
wire _abc_40298_new_n2690_; 
wire _abc_40298_new_n2692_; 
wire _abc_40298_new_n2693_; 
wire _abc_40298_new_n2694_; 
wire _abc_40298_new_n2695_; 
wire _abc_40298_new_n2696_; 
wire _abc_40298_new_n2697_; 
wire _abc_40298_new_n2698_; 
wire _abc_40298_new_n2699_; 
wire _abc_40298_new_n2701_; 
wire _abc_40298_new_n2702_; 
wire _abc_40298_new_n2703_; 
wire _abc_40298_new_n2704_; 
wire _abc_40298_new_n2705_; 
wire _abc_40298_new_n2706_; 
wire _abc_40298_new_n2707_; 
wire _abc_40298_new_n2708_; 
wire _abc_40298_new_n2710_; 
wire _abc_40298_new_n2711_; 
wire _abc_40298_new_n2712_; 
wire _abc_40298_new_n2713_; 
wire _abc_40298_new_n2714_; 
wire _abc_40298_new_n2715_; 
wire _abc_40298_new_n2716_; 
wire _abc_40298_new_n2717_; 
wire _abc_40298_new_n2719_; 
wire _abc_40298_new_n2720_; 
wire _abc_40298_new_n2721_; 
wire _abc_40298_new_n2722_; 
wire _abc_40298_new_n2723_; 
wire _abc_40298_new_n2724_; 
wire _abc_40298_new_n2725_; 
wire _abc_40298_new_n2726_; 
wire _abc_40298_new_n2728_; 
wire _abc_40298_new_n2729_; 
wire _abc_40298_new_n2730_; 
wire _abc_40298_new_n2731_; 
wire _abc_40298_new_n2732_; 
wire _abc_40298_new_n2733_; 
wire _abc_40298_new_n2734_; 
wire _abc_40298_new_n2735_; 
wire _abc_40298_new_n2737_; 
wire _abc_40298_new_n2738_; 
wire _abc_40298_new_n2739_; 
wire _abc_40298_new_n2740_; 
wire _abc_40298_new_n2741_; 
wire _abc_40298_new_n2742_; 
wire _abc_40298_new_n2743_; 
wire _abc_40298_new_n2744_; 
wire _abc_40298_new_n2746_; 
wire _abc_40298_new_n2747_; 
wire _abc_40298_new_n2748_; 
wire _abc_40298_new_n2749_; 
wire _abc_40298_new_n2750_; 
wire _abc_40298_new_n2751_; 
wire _abc_40298_new_n2752_; 
wire _abc_40298_new_n2754_; 
wire _abc_40298_new_n2755_; 
wire _abc_40298_new_n2756_; 
wire _abc_40298_new_n2757_; 
wire _abc_40298_new_n2758_; 
wire _abc_40298_new_n2759_; 
wire _abc_40298_new_n2760_; 
wire _abc_40298_new_n2762_; 
wire _abc_40298_new_n2763_; 
wire _abc_40298_new_n2764_; 
wire _abc_40298_new_n2765_; 
wire _abc_40298_new_n2766_; 
wire _abc_40298_new_n2767_; 
wire _abc_40298_new_n2768_; 
wire _abc_40298_new_n2770_; 
wire _abc_40298_new_n2771_; 
wire _abc_40298_new_n2772_; 
wire _abc_40298_new_n2773_; 
wire _abc_40298_new_n2774_; 
wire _abc_40298_new_n2775_; 
wire _abc_40298_new_n2776_; 
wire _abc_40298_new_n2778_; 
wire _abc_40298_new_n2779_; 
wire _abc_40298_new_n2780_; 
wire _abc_40298_new_n2781_; 
wire _abc_40298_new_n2782_; 
wire _abc_40298_new_n2783_; 
wire _abc_40298_new_n2784_; 
wire _abc_40298_new_n2786_; 
wire _abc_40298_new_n2787_; 
wire _abc_40298_new_n2788_; 
wire _abc_40298_new_n2789_; 
wire _abc_40298_new_n2790_; 
wire _abc_40298_new_n2791_; 
wire _abc_40298_new_n2792_; 
wire _abc_40298_new_n2794_; 
wire _abc_40298_new_n2795_; 
wire _abc_40298_new_n2796_; 
wire _abc_40298_new_n2797_; 
wire _abc_40298_new_n2798_; 
wire _abc_40298_new_n2799_; 
wire _abc_40298_new_n2800_; 
wire _abc_40298_new_n2802_; 
wire _abc_40298_new_n2803_; 
wire _abc_40298_new_n2804_; 
wire _abc_40298_new_n2805_; 
wire _abc_40298_new_n2806_; 
wire _abc_40298_new_n2807_; 
wire _abc_40298_new_n2808_; 
wire _abc_40298_new_n2810_; 
wire _abc_40298_new_n2811_; 
wire _abc_40298_new_n2812_; 
wire _abc_40298_new_n2813_; 
wire _abc_40298_new_n2814_; 
wire _abc_40298_new_n2815_; 
wire _abc_40298_new_n2816_; 
wire _abc_40298_new_n2817_; 
wire _abc_40298_new_n2819_; 
wire _abc_40298_new_n2820_; 
wire _abc_40298_new_n2821_; 
wire _abc_40298_new_n2822_; 
wire _abc_40298_new_n2823_; 
wire _abc_40298_new_n2824_; 
wire _abc_40298_new_n2825_; 
wire _abc_40298_new_n2826_; 
wire _abc_40298_new_n2828_; 
wire _abc_40298_new_n2829_; 
wire _abc_40298_new_n2830_; 
wire _abc_40298_new_n2831_; 
wire _abc_40298_new_n2832_; 
wire _abc_40298_new_n2833_; 
wire _abc_40298_new_n2834_; 
wire _abc_40298_new_n2835_; 
wire _abc_40298_new_n2837_; 
wire _abc_40298_new_n2838_; 
wire _abc_40298_new_n2839_; 
wire _abc_40298_new_n2840_; 
wire _abc_40298_new_n2841_; 
wire _abc_40298_new_n2842_; 
wire _abc_40298_new_n2843_; 
wire _abc_40298_new_n2844_; 
wire _abc_40298_new_n2846_; 
wire _abc_40298_new_n2847_; 
wire _abc_40298_new_n2848_; 
wire _abc_40298_new_n2849_; 
wire _abc_40298_new_n2850_; 
wire _abc_40298_new_n2851_; 
wire _abc_40298_new_n2852_; 
wire _abc_40298_new_n2853_; 
wire _abc_40298_new_n2855_; 
wire _abc_40298_new_n2856_; 
wire _abc_40298_new_n2857_; 
wire _abc_40298_new_n2858_; 
wire _abc_40298_new_n2859_; 
wire _abc_40298_new_n2860_; 
wire _abc_40298_new_n2861_; 
wire _abc_40298_new_n2862_; 
wire _abc_40298_new_n2864_; 
wire _abc_40298_new_n2865_; 
wire _abc_40298_new_n2866_; 
wire _abc_40298_new_n2867_; 
wire _abc_40298_new_n2868_; 
wire _abc_40298_new_n2869_; 
wire _abc_40298_new_n2870_; 
wire _abc_40298_new_n2871_; 
wire _abc_40298_new_n2873_; 
wire _abc_40298_new_n2874_; 
wire _abc_40298_new_n2875_; 
wire _abc_40298_new_n2876_; 
wire _abc_40298_new_n2877_; 
wire _abc_40298_new_n2878_; 
wire _abc_40298_new_n2879_; 
wire _abc_40298_new_n2880_; 
wire _abc_40298_new_n2882_; 
wire _abc_40298_new_n2883_; 
wire _abc_40298_new_n2884_; 
wire _abc_40298_new_n2885_; 
wire _abc_40298_new_n2886_; 
wire _abc_40298_new_n2888_; 
wire _abc_40298_new_n2889_; 
wire _abc_40298_new_n2891_; 
wire _abc_40298_new_n2892_; 
wire _abc_40298_new_n2893_; 
wire _abc_40298_new_n2895_; 
wire _abc_40298_new_n2896_; 
wire _abc_40298_new_n2898_; 
wire _abc_40298_new_n2900_; 
wire _abc_40298_new_n2901_; 
wire _abc_40298_new_n2902_; 
wire _abc_40298_new_n2903_; 
wire _abc_40298_new_n2904_; 
wire _abc_40298_new_n2905_; 
wire _abc_40298_new_n2906_; 
wire _abc_40298_new_n2907_; 
wire _abc_40298_new_n2908_; 
wire _abc_40298_new_n2909_; 
wire _abc_40298_new_n2911_; 
wire _abc_40298_new_n2912_; 
wire _abc_40298_new_n2913_; 
wire _abc_40298_new_n2914_; 
wire _abc_40298_new_n2915_; 
wire _abc_40298_new_n2916_; 
wire _abc_40298_new_n2917_; 
wire _abc_40298_new_n2918_; 
wire _abc_40298_new_n2920_; 
wire _abc_40298_new_n2921_; 
wire _abc_40298_new_n2922_; 
wire _abc_40298_new_n2923_; 
wire _abc_40298_new_n2924_; 
wire _abc_40298_new_n2925_; 
wire _abc_40298_new_n2927_; 
wire _abc_40298_new_n2928_; 
wire _abc_40298_new_n2929_; 
wire _abc_40298_new_n2930_; 
wire _abc_40298_new_n2931_; 
wire _abc_40298_new_n2932_; 
wire _abc_40298_new_n2933_; 
wire _abc_40298_new_n2934_; 
wire _abc_40298_new_n2935_; 
wire _abc_40298_new_n2936_; 
wire _abc_40298_new_n2937_; 
wire _abc_40298_new_n2938_; 
wire _abc_40298_new_n2940_; 
wire _abc_40298_new_n2941_; 
wire _abc_40298_new_n2942_; 
wire _abc_40298_new_n2943_; 
wire _abc_40298_new_n2944_; 
wire _abc_40298_new_n2945_; 
wire _abc_40298_new_n2946_; 
wire _abc_40298_new_n2948_; 
wire _abc_40298_new_n2949_; 
wire _abc_40298_new_n2950_; 
wire _abc_40298_new_n2951_; 
wire _abc_40298_new_n2952_; 
wire _abc_40298_new_n2953_; 
wire _abc_40298_new_n2954_; 
wire _abc_40298_new_n2955_; 
wire _abc_40298_new_n2956_; 
wire _abc_40298_new_n2958_; 
wire _abc_40298_new_n2959_; 
wire _abc_40298_new_n2960_; 
wire _abc_40298_new_n2961_; 
wire _abc_40298_new_n2962_; 
wire _abc_40298_new_n2963_; 
wire _abc_40298_new_n2964_; 
wire _abc_40298_new_n2965_; 
wire _abc_40298_new_n2966_; 
wire _abc_40298_new_n2968_; 
wire _abc_40298_new_n2969_; 
wire _abc_40298_new_n2970_; 
wire _abc_40298_new_n2971_; 
wire _abc_40298_new_n2972_; 
wire _abc_40298_new_n2973_; 
wire _abc_40298_new_n2974_; 
wire _abc_40298_new_n2976_; 
wire _abc_40298_new_n2977_; 
wire _abc_40298_new_n2978_; 
wire _abc_40298_new_n2979_; 
wire _abc_40298_new_n2980_; 
wire _abc_40298_new_n2981_; 
wire _abc_40298_new_n2982_; 
wire _abc_40298_new_n2983_; 
wire _abc_40298_new_n2984_; 
wire _abc_40298_new_n2986_; 
wire _abc_40298_new_n2987_; 
wire _abc_40298_new_n2988_; 
wire _abc_40298_new_n2989_; 
wire _abc_40298_new_n2990_; 
wire _abc_40298_new_n2991_; 
wire _abc_40298_new_n2992_; 
wire _abc_40298_new_n2994_; 
wire _abc_40298_new_n2995_; 
wire _abc_40298_new_n2996_; 
wire _abc_40298_new_n2997_; 
wire _abc_40298_new_n2998_; 
wire _abc_40298_new_n2999_; 
wire _abc_40298_new_n3000_; 
wire _abc_40298_new_n3001_; 
wire _abc_40298_new_n3002_; 
wire _abc_40298_new_n3003_; 
wire _abc_40298_new_n3004_; 
wire _abc_40298_new_n3005_; 
wire _abc_40298_new_n3006_; 
wire _abc_40298_new_n3007_; 
wire _abc_40298_new_n3008_; 
wire _abc_40298_new_n3010_; 
wire _abc_40298_new_n3011_; 
wire _abc_40298_new_n3012_; 
wire _abc_40298_new_n3013_; 
wire _abc_40298_new_n3014_; 
wire _abc_40298_new_n3015_; 
wire _abc_40298_new_n3016_; 
wire _abc_40298_new_n3017_; 
wire _abc_40298_new_n3018_; 
wire _abc_40298_new_n3019_; 
wire _abc_40298_new_n3020_; 
wire _abc_40298_new_n3021_; 
wire _abc_40298_new_n3023_; 
wire _abc_40298_new_n3024_; 
wire _abc_40298_new_n3025_; 
wire _abc_40298_new_n3026_; 
wire _abc_40298_new_n3027_; 
wire _abc_40298_new_n3028_; 
wire _abc_40298_new_n3029_; 
wire _abc_40298_new_n3030_; 
wire _abc_40298_new_n3032_; 
wire _abc_40298_new_n3033_; 
wire _abc_40298_new_n3034_; 
wire _abc_40298_new_n3035_; 
wire _abc_40298_new_n3036_; 
wire _abc_40298_new_n3037_; 
wire _abc_40298_new_n3038_; 
wire _abc_40298_new_n3039_; 
wire _abc_40298_new_n3040_; 
wire _abc_40298_new_n3041_; 
wire _abc_40298_new_n3042_; 
wire _abc_40298_new_n3043_; 
wire _abc_40298_new_n3045_; 
wire _abc_40298_new_n3046_; 
wire _abc_40298_new_n3047_; 
wire _abc_40298_new_n3048_; 
wire _abc_40298_new_n3049_; 
wire _abc_40298_new_n3050_; 
wire _abc_40298_new_n3051_; 
wire _abc_40298_new_n3052_; 
wire _abc_40298_new_n3053_; 
wire _abc_40298_new_n3054_; 
wire _abc_40298_new_n3055_; 
wire _abc_40298_new_n3056_; 
wire _abc_40298_new_n3057_; 
wire _abc_40298_new_n3058_; 
wire _abc_40298_new_n3059_; 
wire _abc_40298_new_n3061_; 
wire _abc_40298_new_n3062_; 
wire _abc_40298_new_n3063_; 
wire _abc_40298_new_n3064_; 
wire _abc_40298_new_n3066_; 
wire _abc_40298_new_n3067_; 
wire _abc_40298_new_n3068_; 
wire _abc_40298_new_n3069_; 
wire _abc_40298_new_n3070_; 
wire _abc_40298_new_n3071_; 
wire _abc_40298_new_n3072_; 
wire _abc_40298_new_n3073_; 
wire _abc_40298_new_n3075_; 
wire _abc_40298_new_n3076_; 
wire _abc_40298_new_n3077_; 
wire _abc_40298_new_n3078_; 
wire _abc_40298_new_n3079_; 
wire _abc_40298_new_n3080_; 
wire _abc_40298_new_n3082_; 
wire _abc_40298_new_n3083_; 
wire _abc_40298_new_n3084_; 
wire _abc_40298_new_n3085_; 
wire _abc_40298_new_n3086_; 
wire _abc_40298_new_n3087_; 
wire _abc_40298_new_n3088_; 
wire _abc_40298_new_n3089_; 
wire _abc_40298_new_n3090_; 
wire _abc_40298_new_n3091_; 
wire _abc_40298_new_n3092_; 
wire _abc_40298_new_n3093_; 
wire _abc_40298_new_n3094_; 
wire _abc_40298_new_n3095_; 
wire _abc_40298_new_n3097_; 
wire _abc_40298_new_n3098_; 
wire _abc_40298_new_n3099_; 
wire _abc_40298_new_n3100_; 
wire _abc_40298_new_n3101_; 
wire _abc_40298_new_n3102_; 
wire _abc_40298_new_n3104_; 
wire _abc_40298_new_n3105_; 
wire _abc_40298_new_n3106_; 
wire _abc_40298_new_n3107_; 
wire _abc_40298_new_n3108_; 
wire _abc_40298_new_n3109_; 
wire _abc_40298_new_n3110_; 
wire _abc_40298_new_n3111_; 
wire _abc_40298_new_n3112_; 
wire _abc_40298_new_n3114_; 
wire _abc_40298_new_n3115_; 
wire _abc_40298_new_n3116_; 
wire _abc_40298_new_n3117_; 
wire _abc_40298_new_n3118_; 
wire _abc_40298_new_n3119_; 
wire _abc_40298_new_n3120_; 
wire _abc_40298_new_n3122_; 
wire _abc_40298_new_n3123_; 
wire _abc_40298_new_n3124_; 
wire _abc_40298_new_n3125_; 
wire _abc_40298_new_n3126_; 
wire _abc_40298_new_n3127_; 
wire _abc_40298_new_n3128_; 
wire _abc_40298_new_n3129_; 
wire _abc_40298_new_n3130_; 
wire _abc_40298_new_n3131_; 
wire _abc_40298_new_n3132_; 
wire _abc_40298_new_n3133_; 
wire _abc_40298_new_n3135_; 
wire _abc_40298_new_n3136_; 
wire _abc_40298_new_n3137_; 
wire _abc_40298_new_n3138_; 
wire _abc_40298_new_n3139_; 
wire _abc_40298_new_n3140_; 
wire _abc_40298_new_n3141_; 
wire _abc_40298_new_n3142_; 
wire _abc_40298_new_n3143_; 
wire _abc_40298_new_n3145_; 
wire _abc_40298_new_n3146_; 
wire _abc_40298_new_n3147_; 
wire _abc_40298_new_n3148_; 
wire _abc_40298_new_n3149_; 
wire _abc_40298_new_n3150_; 
wire _abc_40298_new_n3151_; 
wire _abc_40298_new_n3152_; 
wire _abc_40298_new_n3153_; 
wire _abc_40298_new_n3155_; 
wire _abc_40298_new_n3156_; 
wire _abc_40298_new_n3157_; 
wire _abc_40298_new_n3158_; 
wire _abc_40298_new_n3159_; 
wire _abc_40298_new_n3161_; 
wire _abc_40298_new_n3162_; 
wire _abc_40298_new_n3163_; 
wire _abc_40298_new_n3164_; 
wire _abc_40298_new_n3165_; 
wire _abc_40298_new_n3166_; 
wire _abc_40298_new_n3167_; 
wire _abc_40298_new_n3168_; 
wire _abc_40298_new_n3169_; 
wire _abc_40298_new_n3170_; 
wire _abc_40298_new_n3172_; 
wire _abc_40298_new_n3173_; 
wire _abc_40298_new_n3174_; 
wire _abc_40298_new_n3175_; 
wire _abc_40298_new_n3177_; 
wire _abc_40298_new_n3178_; 
wire _abc_40298_new_n3179_; 
wire _abc_40298_new_n3180_; 
wire _abc_40298_new_n3181_; 
wire _abc_40298_new_n3182_; 
wire _abc_40298_new_n3183_; 
wire _abc_40298_new_n3184_; 
wire _abc_40298_new_n3185_; 
wire _abc_40298_new_n3186_; 
wire _abc_40298_new_n3187_; 
wire _abc_40298_new_n3188_; 
wire _abc_40298_new_n3190_; 
wire _abc_40298_new_n3191_; 
wire _abc_40298_new_n3192_; 
wire _abc_40298_new_n3193_; 
wire _abc_40298_new_n3194_; 
wire _abc_40298_new_n3195_; 
wire _abc_40298_new_n3198_; 
wire _abc_40298_new_n3200_; 
wire _abc_40298_new_n617_; 
wire _abc_40298_new_n618_; 
wire _abc_40298_new_n619_; 
wire _abc_40298_new_n620_; 
wire _abc_40298_new_n621_; 
wire _abc_40298_new_n622_; 
wire _abc_40298_new_n623_; 
wire _abc_40298_new_n624_; 
wire _abc_40298_new_n625_; 
wire _abc_40298_new_n626_; 
wire _abc_40298_new_n627_; 
wire _abc_40298_new_n628_; 
wire _abc_40298_new_n630_; 
wire _abc_40298_new_n631_; 
wire _abc_40298_new_n632_; 
wire _abc_40298_new_n634_; 
wire _abc_40298_new_n635_; 
wire _abc_40298_new_n636_; 
wire _abc_40298_new_n637_; 
wire _abc_40298_new_n638_; 
wire _abc_40298_new_n639_; 
wire _abc_40298_new_n640_; 
wire _abc_40298_new_n641_; 
wire _abc_40298_new_n642_; 
wire _abc_40298_new_n643_; 
wire _abc_40298_new_n644_; 
wire _abc_40298_new_n645_; 
wire _abc_40298_new_n646_; 
wire _abc_40298_new_n647_; 
wire _abc_40298_new_n648_; 
wire _abc_40298_new_n649_; 
wire _abc_40298_new_n650_; 
wire _abc_40298_new_n651_; 
wire _abc_40298_new_n652_; 
wire _abc_40298_new_n653_; 
wire _abc_40298_new_n654_; 
wire _abc_40298_new_n655_; 
wire _abc_40298_new_n656_; 
wire _abc_40298_new_n657_; 
wire _abc_40298_new_n658_; 
wire _abc_40298_new_n659_; 
wire _abc_40298_new_n660_; 
wire _abc_40298_new_n661_; 
wire _abc_40298_new_n662_; 
wire _abc_40298_new_n663_; 
wire _abc_40298_new_n664_; 
wire _abc_40298_new_n666_; 
wire _abc_40298_new_n667_; 
wire _abc_40298_new_n669_; 
wire _abc_40298_new_n671_; 
wire _abc_40298_new_n672_; 
wire _abc_40298_new_n673_; 
wire _abc_40298_new_n674_; 
wire _abc_40298_new_n675_; 
wire _abc_40298_new_n676_; 
wire _abc_40298_new_n677_; 
wire _abc_40298_new_n678_; 
wire _abc_40298_new_n679_; 
wire _abc_40298_new_n680_; 
wire _abc_40298_new_n681_; 
wire _abc_40298_new_n682_; 
wire _abc_40298_new_n683_; 
wire _abc_40298_new_n684_; 
wire _abc_40298_new_n685_; 
wire _abc_40298_new_n686_; 
wire _abc_40298_new_n687_; 
wire _abc_40298_new_n688_; 
wire _abc_40298_new_n689_; 
wire _abc_40298_new_n690_; 
wire _abc_40298_new_n691_; 
wire _abc_40298_new_n693_; 
wire _abc_40298_new_n694_; 
wire _abc_40298_new_n695_; 
wire _abc_40298_new_n696_; 
wire _abc_40298_new_n697_; 
wire _abc_40298_new_n698_; 
wire _abc_40298_new_n699_; 
wire _abc_40298_new_n700_; 
wire _abc_40298_new_n701_; 
wire _abc_40298_new_n702_; 
wire _abc_40298_new_n703_; 
wire _abc_40298_new_n704_; 
wire _abc_40298_new_n706_; 
wire _abc_40298_new_n707_; 
wire _abc_40298_new_n708_; 
wire _abc_40298_new_n709_; 
wire _abc_40298_new_n710_; 
wire _abc_40298_new_n711_; 
wire _abc_40298_new_n712_; 
wire _abc_40298_new_n713_; 
wire _abc_40298_new_n714_; 
wire _abc_40298_new_n715_; 
wire _abc_40298_new_n717_; 
wire _abc_40298_new_n718_; 
wire _abc_40298_new_n719_; 
wire _abc_40298_new_n720_; 
wire _abc_40298_new_n721_; 
wire _abc_40298_new_n722_; 
wire _abc_40298_new_n723_; 
wire _abc_40298_new_n724_; 
wire _abc_40298_new_n725_; 
wire _abc_40298_new_n726_; 
wire _abc_40298_new_n728_; 
wire _abc_40298_new_n729_; 
wire _abc_40298_new_n730_; 
wire _abc_40298_new_n731_; 
wire _abc_40298_new_n732_; 
wire _abc_40298_new_n733_; 
wire _abc_40298_new_n734_; 
wire _abc_40298_new_n735_; 
wire _abc_40298_new_n737_; 
wire _abc_40298_new_n738_; 
wire _abc_40298_new_n739_; 
wire _abc_40298_new_n740_; 
wire _abc_40298_new_n741_; 
wire _abc_40298_new_n742_; 
wire _abc_40298_new_n743_; 
wire _abc_40298_new_n744_; 
wire _abc_40298_new_n746_; 
wire _abc_40298_new_n747_; 
wire _abc_40298_new_n748_; 
wire _abc_40298_new_n749_; 
wire _abc_40298_new_n750_; 
wire _abc_40298_new_n751_; 
wire _abc_40298_new_n752_; 
wire _abc_40298_new_n753_; 
wire _abc_40298_new_n755_; 
wire _abc_40298_new_n756_; 
wire _abc_40298_new_n757_; 
wire _abc_40298_new_n758_; 
wire _abc_40298_new_n759_; 
wire _abc_40298_new_n760_; 
wire _abc_40298_new_n761_; 
wire _abc_40298_new_n763_; 
wire _abc_40298_new_n764_; 
wire _abc_40298_new_n765_; 
wire _abc_40298_new_n766_; 
wire _abc_40298_new_n767_; 
wire _abc_40298_new_n769_; 
wire _abc_40298_new_n770_; 
wire _abc_40298_new_n771_; 
wire _abc_40298_new_n772_; 
wire _abc_40298_new_n773_; 
wire _abc_40298_new_n775_; 
wire _abc_40298_new_n776_; 
wire _abc_40298_new_n777_; 
wire _abc_40298_new_n778_; 
wire _abc_40298_new_n780_; 
wire _abc_40298_new_n781_; 
wire _abc_40298_new_n782_; 
wire _abc_40298_new_n783_; 
wire _abc_40298_new_n785_; 
wire _abc_40298_new_n786_; 
wire _abc_40298_new_n787_; 
wire _abc_40298_new_n789_; 
wire _abc_40298_new_n790_; 
wire _abc_40298_new_n791_; 
wire _abc_40298_new_n793_; 
wire _abc_40298_new_n794_; 
wire _abc_40298_new_n795_; 
wire _abc_40298_new_n796_; 
wire _abc_40298_new_n797_; 
wire _abc_40298_new_n799_; 
wire _abc_40298_new_n800_; 
wire _abc_40298_new_n801_; 
wire _abc_40298_new_n803_; 
wire _abc_40298_new_n804_; 
wire _abc_40298_new_n805_; 
wire _abc_40298_new_n806_; 
wire _abc_40298_new_n807_; 
wire _abc_40298_new_n809_; 
wire _abc_40298_new_n810_; 
wire _abc_40298_new_n811_; 
wire _abc_40298_new_n812_; 
wire _abc_40298_new_n814_; 
wire _abc_40298_new_n815_; 
wire _abc_40298_new_n816_; 
wire _abc_40298_new_n817_; 
wire _abc_40298_new_n819_; 
wire _abc_40298_new_n820_; 
wire _abc_40298_new_n821_; 
wire _abc_40298_new_n822_; 
wire _abc_40298_new_n824_; 
wire _abc_40298_new_n825_; 
wire _abc_40298_new_n826_; 
wire _abc_40298_new_n827_; 
wire _abc_40298_new_n829_; 
wire _abc_40298_new_n830_; 
wire _abc_40298_new_n831_; 
wire _abc_40298_new_n832_; 
wire _abc_40298_new_n834_; 
wire _abc_40298_new_n835_; 
wire _abc_40298_new_n836_; 
wire _abc_40298_new_n837_; 
wire _abc_40298_new_n839_; 
wire _abc_40298_new_n840_; 
wire _abc_40298_new_n841_; 
wire _abc_40298_new_n842_; 
wire _abc_40298_new_n844_; 
wire _abc_40298_new_n845_; 
wire _abc_40298_new_n846_; 
wire _abc_40298_new_n847_; 
wire _abc_40298_new_n849_; 
wire _abc_40298_new_n850_; 
wire _abc_40298_new_n851_; 
wire _abc_40298_new_n852_; 
wire _abc_40298_new_n854_; 
wire _abc_40298_new_n855_; 
wire _abc_40298_new_n856_; 
wire _abc_40298_new_n857_; 
wire _abc_40298_new_n859_; 
wire _abc_40298_new_n860_; 
wire _abc_40298_new_n861_; 
wire _abc_40298_new_n862_; 
wire _abc_40298_new_n864_; 
wire _abc_40298_new_n865_; 
wire _abc_40298_new_n866_; 
wire _abc_40298_new_n867_; 
wire _abc_40298_new_n869_; 
wire _abc_40298_new_n870_; 
wire _abc_40298_new_n871_; 
wire _abc_40298_new_n872_; 
wire _abc_40298_new_n874_; 
wire _abc_40298_new_n875_; 
wire _abc_40298_new_n876_; 
wire _abc_40298_new_n877_; 
wire _abc_40298_new_n879_; 
wire _abc_40298_new_n880_; 
wire _abc_40298_new_n881_; 
wire _abc_40298_new_n882_; 
wire _abc_40298_new_n885_; 
wire _abc_40298_new_n886_; 
wire _abc_40298_new_n887_; 
wire _abc_40298_new_n888_; 
wire _abc_40298_new_n889_; 
wire _abc_40298_new_n890_; 
wire _abc_40298_new_n891_; 
wire _abc_40298_new_n892_; 
wire _abc_40298_new_n893_; 
wire _abc_40298_new_n894_; 
wire _abc_40298_new_n895_; 
wire _abc_40298_new_n896_; 
wire _abc_40298_new_n897_; 
wire _abc_40298_new_n898_; 
wire _abc_40298_new_n899_; 
wire _abc_40298_new_n900_; 
wire _abc_40298_new_n901_; 
wire _abc_40298_new_n902_; 
wire _abc_40298_new_n903_; 
wire _abc_40298_new_n904_; 
wire _abc_40298_new_n905_; 
wire _abc_40298_new_n906_; 
wire _abc_40298_new_n907_; 
wire _abc_40298_new_n908_; 
wire _abc_40298_new_n909_; 
wire _abc_40298_new_n910_; 
wire _abc_40298_new_n911_; 
wire _abc_40298_new_n912_; 
wire _abc_40298_new_n913_; 
wire _abc_40298_new_n914_; 
wire _abc_40298_new_n915_; 
wire _abc_40298_new_n916_; 
wire _abc_40298_new_n917_; 
wire _abc_40298_new_n918_; 
wire _abc_40298_new_n919_; 
wire _abc_40298_new_n920_; 
wire _abc_40298_new_n921_; 
wire _abc_40298_new_n922_; 
wire _abc_40298_new_n923_; 
wire _abc_40298_new_n924_; 
wire _abc_40298_new_n925_; 
wire _abc_40298_new_n926_; 
wire _abc_40298_new_n927_; 
wire _abc_40298_new_n928_; 
wire _abc_40298_new_n929_; 
wire _abc_40298_new_n930_; 
wire _abc_40298_new_n931_; 
wire _abc_40298_new_n932_; 
wire _abc_40298_new_n933_; 
wire _abc_40298_new_n934_; 
wire _abc_40298_new_n935_; 
wire _abc_40298_new_n936_; 
wire _abc_40298_new_n937_; 
wire _abc_40298_new_n938_; 
wire _abc_40298_new_n939_; 
wire _abc_40298_new_n940_; 
wire _abc_40298_new_n941_; 
wire _abc_40298_new_n942_; 
wire _abc_40298_new_n943_; 
wire _abc_40298_new_n944_; 
wire _abc_40298_new_n945_; 
wire _abc_40298_new_n946_; 
wire _abc_40298_new_n947_; 
wire _abc_40298_new_n948_; 
wire _abc_40298_new_n949_; 
wire _abc_40298_new_n950_; 
wire _abc_40298_new_n951_; 
wire _abc_40298_new_n952_; 
wire _abc_40298_new_n953_; 
wire _abc_40298_new_n954_; 
wire _abc_40298_new_n955_; 
wire _abc_40298_new_n956_; 
wire _abc_40298_new_n957_; 
wire _abc_40298_new_n958_; 
wire _abc_40298_new_n959_; 
wire _abc_40298_new_n960_; 
wire _abc_40298_new_n961_; 
wire _abc_40298_new_n962_; 
wire _abc_40298_new_n963_; 
wire _abc_40298_new_n964_; 
wire _abc_40298_new_n965_; 
wire _abc_40298_new_n966_; 
wire _abc_40298_new_n967_; 
wire _abc_40298_new_n968_; 
wire _abc_40298_new_n969_; 
wire _abc_40298_new_n970_; 
wire _abc_40298_new_n971_; 
wire _abc_40298_new_n972_; 
wire _abc_40298_new_n973_; 
wire _abc_40298_new_n974_; 
wire _abc_40298_new_n975_; 
wire _abc_40298_new_n976_; 
wire _abc_40298_new_n977_; 
wire _abc_40298_new_n978_; 
wire _abc_40298_new_n979_; 
wire _abc_40298_new_n980_; 
wire _abc_40298_new_n981_; 
wire _abc_40298_new_n982_; 
wire _abc_40298_new_n983_; 
wire _abc_40298_new_n984_; 
wire _abc_40298_new_n985_; 
wire _abc_40298_new_n986_; 
wire _abc_40298_new_n987_; 
wire _abc_40298_new_n988_; 
wire _abc_40298_new_n989_; 
wire _abc_40298_new_n990_; 
wire _abc_40298_new_n991_; 
wire _abc_40298_new_n992_; 
wire _abc_40298_new_n993_; 
wire _abc_40298_new_n994_; 
wire _abc_40298_new_n995_; 
wire _abc_40298_new_n996_; 
wire _abc_40298_new_n997_; 
wire _abc_40298_new_n998_; 
wire _abc_40298_new_n999_; 
wire alu__abc_38674_new_n1000_; 
wire alu__abc_38674_new_n1001_; 
wire alu__abc_38674_new_n1002_; 
wire alu__abc_38674_new_n1003_; 
wire alu__abc_38674_new_n1004_; 
wire alu__abc_38674_new_n1005_; 
wire alu__abc_38674_new_n1007_; 
wire alu__abc_38674_new_n1008_; 
wire alu__abc_38674_new_n1009_; 
wire alu__abc_38674_new_n1010_; 
wire alu__abc_38674_new_n1011_; 
wire alu__abc_38674_new_n1012_; 
wire alu__abc_38674_new_n1013_; 
wire alu__abc_38674_new_n1014_; 
wire alu__abc_38674_new_n1015_; 
wire alu__abc_38674_new_n1016_; 
wire alu__abc_38674_new_n1017_; 
wire alu__abc_38674_new_n1018_; 
wire alu__abc_38674_new_n1019_; 
wire alu__abc_38674_new_n1020_; 
wire alu__abc_38674_new_n1021_; 
wire alu__abc_38674_new_n1022_; 
wire alu__abc_38674_new_n1023_; 
wire alu__abc_38674_new_n1024_; 
wire alu__abc_38674_new_n1025_; 
wire alu__abc_38674_new_n1026_; 
wire alu__abc_38674_new_n1027_; 
wire alu__abc_38674_new_n1028_; 
wire alu__abc_38674_new_n1029_; 
wire alu__abc_38674_new_n1030_; 
wire alu__abc_38674_new_n1031_; 
wire alu__abc_38674_new_n1032_; 
wire alu__abc_38674_new_n1033_; 
wire alu__abc_38674_new_n1034_; 
wire alu__abc_38674_new_n1035_; 
wire alu__abc_38674_new_n1036_; 
wire alu__abc_38674_new_n1037_; 
wire alu__abc_38674_new_n1038_; 
wire alu__abc_38674_new_n1039_; 
wire alu__abc_38674_new_n1041_; 
wire alu__abc_38674_new_n1042_; 
wire alu__abc_38674_new_n1043_; 
wire alu__abc_38674_new_n1044_; 
wire alu__abc_38674_new_n1045_; 
wire alu__abc_38674_new_n1046_; 
wire alu__abc_38674_new_n1047_; 
wire alu__abc_38674_new_n1048_; 
wire alu__abc_38674_new_n1049_; 
wire alu__abc_38674_new_n1050_; 
wire alu__abc_38674_new_n1051_; 
wire alu__abc_38674_new_n1052_; 
wire alu__abc_38674_new_n1053_; 
wire alu__abc_38674_new_n1054_; 
wire alu__abc_38674_new_n1055_; 
wire alu__abc_38674_new_n1056_; 
wire alu__abc_38674_new_n1057_; 
wire alu__abc_38674_new_n1058_; 
wire alu__abc_38674_new_n1059_; 
wire alu__abc_38674_new_n1060_; 
wire alu__abc_38674_new_n1061_; 
wire alu__abc_38674_new_n1062_; 
wire alu__abc_38674_new_n1063_; 
wire alu__abc_38674_new_n1064_; 
wire alu__abc_38674_new_n1065_; 
wire alu__abc_38674_new_n1066_; 
wire alu__abc_38674_new_n1067_; 
wire alu__abc_38674_new_n1068_; 
wire alu__abc_38674_new_n1069_; 
wire alu__abc_38674_new_n1070_; 
wire alu__abc_38674_new_n1071_; 
wire alu__abc_38674_new_n1072_; 
wire alu__abc_38674_new_n1073_; 
wire alu__abc_38674_new_n1075_; 
wire alu__abc_38674_new_n1076_; 
wire alu__abc_38674_new_n1077_; 
wire alu__abc_38674_new_n1078_; 
wire alu__abc_38674_new_n1079_; 
wire alu__abc_38674_new_n1080_; 
wire alu__abc_38674_new_n1081_; 
wire alu__abc_38674_new_n1082_; 
wire alu__abc_38674_new_n1083_; 
wire alu__abc_38674_new_n1084_; 
wire alu__abc_38674_new_n1085_; 
wire alu__abc_38674_new_n1086_; 
wire alu__abc_38674_new_n1087_; 
wire alu__abc_38674_new_n1088_; 
wire alu__abc_38674_new_n1089_; 
wire alu__abc_38674_new_n1090_; 
wire alu__abc_38674_new_n1091_; 
wire alu__abc_38674_new_n1092_; 
wire alu__abc_38674_new_n1093_; 
wire alu__abc_38674_new_n1094_; 
wire alu__abc_38674_new_n1095_; 
wire alu__abc_38674_new_n1096_; 
wire alu__abc_38674_new_n1097_; 
wire alu__abc_38674_new_n1098_; 
wire alu__abc_38674_new_n1099_; 
wire alu__abc_38674_new_n1100_; 
wire alu__abc_38674_new_n1101_; 
wire alu__abc_38674_new_n1102_; 
wire alu__abc_38674_new_n1103_; 
wire alu__abc_38674_new_n1104_; 
wire alu__abc_38674_new_n1105_; 
wire alu__abc_38674_new_n1106_; 
wire alu__abc_38674_new_n1107_; 
wire alu__abc_38674_new_n1109_; 
wire alu__abc_38674_new_n110_; 
wire alu__abc_38674_new_n1110_; 
wire alu__abc_38674_new_n1111_; 
wire alu__abc_38674_new_n1112_; 
wire alu__abc_38674_new_n1113_; 
wire alu__abc_38674_new_n1114_; 
wire alu__abc_38674_new_n1115_; 
wire alu__abc_38674_new_n1116_; 
wire alu__abc_38674_new_n1117_; 
wire alu__abc_38674_new_n1118_; 
wire alu__abc_38674_new_n1119_; 
wire alu__abc_38674_new_n111_; 
wire alu__abc_38674_new_n1120_; 
wire alu__abc_38674_new_n1121_; 
wire alu__abc_38674_new_n1122_; 
wire alu__abc_38674_new_n1123_; 
wire alu__abc_38674_new_n1124_; 
wire alu__abc_38674_new_n1125_; 
wire alu__abc_38674_new_n1126_; 
wire alu__abc_38674_new_n1127_; 
wire alu__abc_38674_new_n1128_; 
wire alu__abc_38674_new_n1129_; 
wire alu__abc_38674_new_n112_; 
wire alu__abc_38674_new_n1130_; 
wire alu__abc_38674_new_n1131_; 
wire alu__abc_38674_new_n1132_; 
wire alu__abc_38674_new_n1133_; 
wire alu__abc_38674_new_n1134_; 
wire alu__abc_38674_new_n1135_; 
wire alu__abc_38674_new_n1137_; 
wire alu__abc_38674_new_n1138_; 
wire alu__abc_38674_new_n1139_; 
wire alu__abc_38674_new_n113_; 
wire alu__abc_38674_new_n1140_; 
wire alu__abc_38674_new_n1141_; 
wire alu__abc_38674_new_n1142_; 
wire alu__abc_38674_new_n1143_; 
wire alu__abc_38674_new_n1144_; 
wire alu__abc_38674_new_n1145_; 
wire alu__abc_38674_new_n1146_; 
wire alu__abc_38674_new_n1147_; 
wire alu__abc_38674_new_n1148_; 
wire alu__abc_38674_new_n1149_; 
wire alu__abc_38674_new_n114_; 
wire alu__abc_38674_new_n1150_; 
wire alu__abc_38674_new_n1151_; 
wire alu__abc_38674_new_n1152_; 
wire alu__abc_38674_new_n1153_; 
wire alu__abc_38674_new_n1154_; 
wire alu__abc_38674_new_n1155_; 
wire alu__abc_38674_new_n1156_; 
wire alu__abc_38674_new_n1157_; 
wire alu__abc_38674_new_n1158_; 
wire alu__abc_38674_new_n1159_; 
wire alu__abc_38674_new_n115_; 
wire alu__abc_38674_new_n1160_; 
wire alu__abc_38674_new_n1161_; 
wire alu__abc_38674_new_n1162_; 
wire alu__abc_38674_new_n1163_; 
wire alu__abc_38674_new_n1164_; 
wire alu__abc_38674_new_n1165_; 
wire alu__abc_38674_new_n1166_; 
wire alu__abc_38674_new_n1167_; 
wire alu__abc_38674_new_n1168_; 
wire alu__abc_38674_new_n1169_; 
wire alu__abc_38674_new_n116_; 
wire alu__abc_38674_new_n1171_; 
wire alu__abc_38674_new_n1172_; 
wire alu__abc_38674_new_n1173_; 
wire alu__abc_38674_new_n1174_; 
wire alu__abc_38674_new_n1175_; 
wire alu__abc_38674_new_n1176_; 
wire alu__abc_38674_new_n1177_; 
wire alu__abc_38674_new_n1178_; 
wire alu__abc_38674_new_n1179_; 
wire alu__abc_38674_new_n117_; 
wire alu__abc_38674_new_n1180_; 
wire alu__abc_38674_new_n1181_; 
wire alu__abc_38674_new_n1182_; 
wire alu__abc_38674_new_n1183_; 
wire alu__abc_38674_new_n1184_; 
wire alu__abc_38674_new_n1185_; 
wire alu__abc_38674_new_n1186_; 
wire alu__abc_38674_new_n1187_; 
wire alu__abc_38674_new_n1188_; 
wire alu__abc_38674_new_n1189_; 
wire alu__abc_38674_new_n118_; 
wire alu__abc_38674_new_n1190_; 
wire alu__abc_38674_new_n1191_; 
wire alu__abc_38674_new_n1192_; 
wire alu__abc_38674_new_n1193_; 
wire alu__abc_38674_new_n1194_; 
wire alu__abc_38674_new_n1195_; 
wire alu__abc_38674_new_n1196_; 
wire alu__abc_38674_new_n1197_; 
wire alu__abc_38674_new_n1198_; 
wire alu__abc_38674_new_n119_; 
wire alu__abc_38674_new_n1200_; 
wire alu__abc_38674_new_n1201_; 
wire alu__abc_38674_new_n1202_; 
wire alu__abc_38674_new_n1203_; 
wire alu__abc_38674_new_n1204_; 
wire alu__abc_38674_new_n1205_; 
wire alu__abc_38674_new_n1206_; 
wire alu__abc_38674_new_n1207_; 
wire alu__abc_38674_new_n1208_; 
wire alu__abc_38674_new_n1209_; 
wire alu__abc_38674_new_n120_; 
wire alu__abc_38674_new_n1210_; 
wire alu__abc_38674_new_n1211_; 
wire alu__abc_38674_new_n1212_; 
wire alu__abc_38674_new_n1213_; 
wire alu__abc_38674_new_n1214_; 
wire alu__abc_38674_new_n1215_; 
wire alu__abc_38674_new_n1216_; 
wire alu__abc_38674_new_n1217_; 
wire alu__abc_38674_new_n1218_; 
wire alu__abc_38674_new_n1219_; 
wire alu__abc_38674_new_n121_; 
wire alu__abc_38674_new_n1220_; 
wire alu__abc_38674_new_n1221_; 
wire alu__abc_38674_new_n1222_; 
wire alu__abc_38674_new_n1223_; 
wire alu__abc_38674_new_n1224_; 
wire alu__abc_38674_new_n1225_; 
wire alu__abc_38674_new_n1226_; 
wire alu__abc_38674_new_n1227_; 
wire alu__abc_38674_new_n1228_; 
wire alu__abc_38674_new_n1229_; 
wire alu__abc_38674_new_n122_; 
wire alu__abc_38674_new_n1230_; 
wire alu__abc_38674_new_n1231_; 
wire alu__abc_38674_new_n1232_; 
wire alu__abc_38674_new_n1234_; 
wire alu__abc_38674_new_n1235_; 
wire alu__abc_38674_new_n1236_; 
wire alu__abc_38674_new_n1237_; 
wire alu__abc_38674_new_n1238_; 
wire alu__abc_38674_new_n1239_; 
wire alu__abc_38674_new_n123_; 
wire alu__abc_38674_new_n1240_; 
wire alu__abc_38674_new_n1241_; 
wire alu__abc_38674_new_n1242_; 
wire alu__abc_38674_new_n1243_; 
wire alu__abc_38674_new_n1244_; 
wire alu__abc_38674_new_n1245_; 
wire alu__abc_38674_new_n1246_; 
wire alu__abc_38674_new_n1247_; 
wire alu__abc_38674_new_n1248_; 
wire alu__abc_38674_new_n1249_; 
wire alu__abc_38674_new_n124_; 
wire alu__abc_38674_new_n1250_; 
wire alu__abc_38674_new_n1251_; 
wire alu__abc_38674_new_n1252_; 
wire alu__abc_38674_new_n1253_; 
wire alu__abc_38674_new_n1254_; 
wire alu__abc_38674_new_n1255_; 
wire alu__abc_38674_new_n1256_; 
wire alu__abc_38674_new_n1257_; 
wire alu__abc_38674_new_n1258_; 
wire alu__abc_38674_new_n1259_; 
wire alu__abc_38674_new_n125_; 
wire alu__abc_38674_new_n1260_; 
wire alu__abc_38674_new_n1261_; 
wire alu__abc_38674_new_n1263_; 
wire alu__abc_38674_new_n1264_; 
wire alu__abc_38674_new_n1265_; 
wire alu__abc_38674_new_n1266_; 
wire alu__abc_38674_new_n1267_; 
wire alu__abc_38674_new_n1268_; 
wire alu__abc_38674_new_n1269_; 
wire alu__abc_38674_new_n126_; 
wire alu__abc_38674_new_n1270_; 
wire alu__abc_38674_new_n1271_; 
wire alu__abc_38674_new_n1272_; 
wire alu__abc_38674_new_n1273_; 
wire alu__abc_38674_new_n1274_; 
wire alu__abc_38674_new_n1275_; 
wire alu__abc_38674_new_n1276_; 
wire alu__abc_38674_new_n1277_; 
wire alu__abc_38674_new_n1278_; 
wire alu__abc_38674_new_n1279_; 
wire alu__abc_38674_new_n127_; 
wire alu__abc_38674_new_n1280_; 
wire alu__abc_38674_new_n1281_; 
wire alu__abc_38674_new_n1282_; 
wire alu__abc_38674_new_n1283_; 
wire alu__abc_38674_new_n1284_; 
wire alu__abc_38674_new_n1285_; 
wire alu__abc_38674_new_n1286_; 
wire alu__abc_38674_new_n1287_; 
wire alu__abc_38674_new_n1288_; 
wire alu__abc_38674_new_n1289_; 
wire alu__abc_38674_new_n128_; 
wire alu__abc_38674_new_n1290_; 
wire alu__abc_38674_new_n1291_; 
wire alu__abc_38674_new_n1292_; 
wire alu__abc_38674_new_n1294_; 
wire alu__abc_38674_new_n1295_; 
wire alu__abc_38674_new_n1296_; 
wire alu__abc_38674_new_n1297_; 
wire alu__abc_38674_new_n1298_; 
wire alu__abc_38674_new_n1299_; 
wire alu__abc_38674_new_n129_; 
wire alu__abc_38674_new_n1300_; 
wire alu__abc_38674_new_n1301_; 
wire alu__abc_38674_new_n1302_; 
wire alu__abc_38674_new_n1303_; 
wire alu__abc_38674_new_n1304_; 
wire alu__abc_38674_new_n1305_; 
wire alu__abc_38674_new_n1306_; 
wire alu__abc_38674_new_n1307_; 
wire alu__abc_38674_new_n1308_; 
wire alu__abc_38674_new_n1309_; 
wire alu__abc_38674_new_n130_; 
wire alu__abc_38674_new_n1310_; 
wire alu__abc_38674_new_n1311_; 
wire alu__abc_38674_new_n1312_; 
wire alu__abc_38674_new_n1313_; 
wire alu__abc_38674_new_n1314_; 
wire alu__abc_38674_new_n1315_; 
wire alu__abc_38674_new_n1316_; 
wire alu__abc_38674_new_n1317_; 
wire alu__abc_38674_new_n1318_; 
wire alu__abc_38674_new_n1319_; 
wire alu__abc_38674_new_n131_; 
wire alu__abc_38674_new_n1320_; 
wire alu__abc_38674_new_n1321_; 
wire alu__abc_38674_new_n1322_; 
wire alu__abc_38674_new_n1323_; 
wire alu__abc_38674_new_n1324_; 
wire alu__abc_38674_new_n1325_; 
wire alu__abc_38674_new_n1327_; 
wire alu__abc_38674_new_n1328_; 
wire alu__abc_38674_new_n1329_; 
wire alu__abc_38674_new_n132_; 
wire alu__abc_38674_new_n1330_; 
wire alu__abc_38674_new_n1331_; 
wire alu__abc_38674_new_n1332_; 
wire alu__abc_38674_new_n1333_; 
wire alu__abc_38674_new_n1334_; 
wire alu__abc_38674_new_n1335_; 
wire alu__abc_38674_new_n1336_; 
wire alu__abc_38674_new_n1337_; 
wire alu__abc_38674_new_n1338_; 
wire alu__abc_38674_new_n1339_; 
wire alu__abc_38674_new_n133_; 
wire alu__abc_38674_new_n1340_; 
wire alu__abc_38674_new_n1341_; 
wire alu__abc_38674_new_n1342_; 
wire alu__abc_38674_new_n1343_; 
wire alu__abc_38674_new_n1344_; 
wire alu__abc_38674_new_n1345_; 
wire alu__abc_38674_new_n1346_; 
wire alu__abc_38674_new_n1347_; 
wire alu__abc_38674_new_n1348_; 
wire alu__abc_38674_new_n1349_; 
wire alu__abc_38674_new_n134_; 
wire alu__abc_38674_new_n1350_; 
wire alu__abc_38674_new_n1351_; 
wire alu__abc_38674_new_n1352_; 
wire alu__abc_38674_new_n1353_; 
wire alu__abc_38674_new_n1354_; 
wire alu__abc_38674_new_n1355_; 
wire alu__abc_38674_new_n1356_; 
wire alu__abc_38674_new_n1358_; 
wire alu__abc_38674_new_n1359_; 
wire alu__abc_38674_new_n135_; 
wire alu__abc_38674_new_n1360_; 
wire alu__abc_38674_new_n1361_; 
wire alu__abc_38674_new_n1362_; 
wire alu__abc_38674_new_n1363_; 
wire alu__abc_38674_new_n1364_; 
wire alu__abc_38674_new_n1365_; 
wire alu__abc_38674_new_n1366_; 
wire alu__abc_38674_new_n1367_; 
wire alu__abc_38674_new_n1368_; 
wire alu__abc_38674_new_n1369_; 
wire alu__abc_38674_new_n136_; 
wire alu__abc_38674_new_n1370_; 
wire alu__abc_38674_new_n1371_; 
wire alu__abc_38674_new_n1372_; 
wire alu__abc_38674_new_n1373_; 
wire alu__abc_38674_new_n1374_; 
wire alu__abc_38674_new_n1375_; 
wire alu__abc_38674_new_n1376_; 
wire alu__abc_38674_new_n1377_; 
wire alu__abc_38674_new_n1378_; 
wire alu__abc_38674_new_n1379_; 
wire alu__abc_38674_new_n137_; 
wire alu__abc_38674_new_n1380_; 
wire alu__abc_38674_new_n1381_; 
wire alu__abc_38674_new_n1382_; 
wire alu__abc_38674_new_n1384_; 
wire alu__abc_38674_new_n1385_; 
wire alu__abc_38674_new_n1386_; 
wire alu__abc_38674_new_n1387_; 
wire alu__abc_38674_new_n1388_; 
wire alu__abc_38674_new_n1389_; 
wire alu__abc_38674_new_n138_; 
wire alu__abc_38674_new_n1390_; 
wire alu__abc_38674_new_n1391_; 
wire alu__abc_38674_new_n1392_; 
wire alu__abc_38674_new_n1393_; 
wire alu__abc_38674_new_n1394_; 
wire alu__abc_38674_new_n1395_; 
wire alu__abc_38674_new_n1396_; 
wire alu__abc_38674_new_n1397_; 
wire alu__abc_38674_new_n1398_; 
wire alu__abc_38674_new_n1399_; 
wire alu__abc_38674_new_n139_; 
wire alu__abc_38674_new_n1400_; 
wire alu__abc_38674_new_n1401_; 
wire alu__abc_38674_new_n1402_; 
wire alu__abc_38674_new_n1403_; 
wire alu__abc_38674_new_n1404_; 
wire alu__abc_38674_new_n1405_; 
wire alu__abc_38674_new_n1406_; 
wire alu__abc_38674_new_n1407_; 
wire alu__abc_38674_new_n1408_; 
wire alu__abc_38674_new_n1409_; 
wire alu__abc_38674_new_n140_; 
wire alu__abc_38674_new_n1411_; 
wire alu__abc_38674_new_n1412_; 
wire alu__abc_38674_new_n1413_; 
wire alu__abc_38674_new_n1414_; 
wire alu__abc_38674_new_n1415_; 
wire alu__abc_38674_new_n1416_; 
wire alu__abc_38674_new_n1417_; 
wire alu__abc_38674_new_n1418_; 
wire alu__abc_38674_new_n1419_; 
wire alu__abc_38674_new_n141_; 
wire alu__abc_38674_new_n1420_; 
wire alu__abc_38674_new_n1421_; 
wire alu__abc_38674_new_n1422_; 
wire alu__abc_38674_new_n1423_; 
wire alu__abc_38674_new_n1424_; 
wire alu__abc_38674_new_n1425_; 
wire alu__abc_38674_new_n1426_; 
wire alu__abc_38674_new_n1427_; 
wire alu__abc_38674_new_n1428_; 
wire alu__abc_38674_new_n1429_; 
wire alu__abc_38674_new_n142_; 
wire alu__abc_38674_new_n1430_; 
wire alu__abc_38674_new_n1431_; 
wire alu__abc_38674_new_n1432_; 
wire alu__abc_38674_new_n1433_; 
wire alu__abc_38674_new_n1434_; 
wire alu__abc_38674_new_n1435_; 
wire alu__abc_38674_new_n1436_; 
wire alu__abc_38674_new_n1437_; 
wire alu__abc_38674_new_n1438_; 
wire alu__abc_38674_new_n1439_; 
wire alu__abc_38674_new_n143_; 
wire alu__abc_38674_new_n1440_; 
wire alu__abc_38674_new_n1442_; 
wire alu__abc_38674_new_n1443_; 
wire alu__abc_38674_new_n1444_; 
wire alu__abc_38674_new_n1445_; 
wire alu__abc_38674_new_n1446_; 
wire alu__abc_38674_new_n1447_; 
wire alu__abc_38674_new_n1448_; 
wire alu__abc_38674_new_n1449_; 
wire alu__abc_38674_new_n144_; 
wire alu__abc_38674_new_n1450_; 
wire alu__abc_38674_new_n1451_; 
wire alu__abc_38674_new_n1452_; 
wire alu__abc_38674_new_n1453_; 
wire alu__abc_38674_new_n1454_; 
wire alu__abc_38674_new_n1455_; 
wire alu__abc_38674_new_n1456_; 
wire alu__abc_38674_new_n1457_; 
wire alu__abc_38674_new_n1458_; 
wire alu__abc_38674_new_n1459_; 
wire alu__abc_38674_new_n145_; 
wire alu__abc_38674_new_n1460_; 
wire alu__abc_38674_new_n1461_; 
wire alu__abc_38674_new_n1462_; 
wire alu__abc_38674_new_n1463_; 
wire alu__abc_38674_new_n1464_; 
wire alu__abc_38674_new_n1465_; 
wire alu__abc_38674_new_n1466_; 
wire alu__abc_38674_new_n1467_; 
wire alu__abc_38674_new_n1468_; 
wire alu__abc_38674_new_n146_; 
wire alu__abc_38674_new_n1470_; 
wire alu__abc_38674_new_n1471_; 
wire alu__abc_38674_new_n1472_; 
wire alu__abc_38674_new_n1473_; 
wire alu__abc_38674_new_n1474_; 
wire alu__abc_38674_new_n1475_; 
wire alu__abc_38674_new_n1476_; 
wire alu__abc_38674_new_n1477_; 
wire alu__abc_38674_new_n1478_; 
wire alu__abc_38674_new_n1479_; 
wire alu__abc_38674_new_n147_; 
wire alu__abc_38674_new_n1480_; 
wire alu__abc_38674_new_n1481_; 
wire alu__abc_38674_new_n1482_; 
wire alu__abc_38674_new_n1483_; 
wire alu__abc_38674_new_n1484_; 
wire alu__abc_38674_new_n1485_; 
wire alu__abc_38674_new_n1486_; 
wire alu__abc_38674_new_n1487_; 
wire alu__abc_38674_new_n1488_; 
wire alu__abc_38674_new_n1489_; 
wire alu__abc_38674_new_n148_; 
wire alu__abc_38674_new_n1490_; 
wire alu__abc_38674_new_n1491_; 
wire alu__abc_38674_new_n1492_; 
wire alu__abc_38674_new_n1493_; 
wire alu__abc_38674_new_n1494_; 
wire alu__abc_38674_new_n1495_; 
wire alu__abc_38674_new_n1497_; 
wire alu__abc_38674_new_n1498_; 
wire alu__abc_38674_new_n1499_; 
wire alu__abc_38674_new_n149_; 
wire alu__abc_38674_new_n1500_; 
wire alu__abc_38674_new_n1501_; 
wire alu__abc_38674_new_n1502_; 
wire alu__abc_38674_new_n1503_; 
wire alu__abc_38674_new_n1504_; 
wire alu__abc_38674_new_n1505_; 
wire alu__abc_38674_new_n1506_; 
wire alu__abc_38674_new_n1507_; 
wire alu__abc_38674_new_n1508_; 
wire alu__abc_38674_new_n1509_; 
wire alu__abc_38674_new_n150_; 
wire alu__abc_38674_new_n1510_; 
wire alu__abc_38674_new_n1511_; 
wire alu__abc_38674_new_n1512_; 
wire alu__abc_38674_new_n1513_; 
wire alu__abc_38674_new_n1514_; 
wire alu__abc_38674_new_n1515_; 
wire alu__abc_38674_new_n1516_; 
wire alu__abc_38674_new_n1517_; 
wire alu__abc_38674_new_n1518_; 
wire alu__abc_38674_new_n1519_; 
wire alu__abc_38674_new_n151_; 
wire alu__abc_38674_new_n1520_; 
wire alu__abc_38674_new_n1521_; 
wire alu__abc_38674_new_n1522_; 
wire alu__abc_38674_new_n1524_; 
wire alu__abc_38674_new_n1525_; 
wire alu__abc_38674_new_n1526_; 
wire alu__abc_38674_new_n1527_; 
wire alu__abc_38674_new_n1528_; 
wire alu__abc_38674_new_n1529_; 
wire alu__abc_38674_new_n152_; 
wire alu__abc_38674_new_n1530_; 
wire alu__abc_38674_new_n1531_; 
wire alu__abc_38674_new_n1532_; 
wire alu__abc_38674_new_n1533_; 
wire alu__abc_38674_new_n1534_; 
wire alu__abc_38674_new_n1535_; 
wire alu__abc_38674_new_n1536_; 
wire alu__abc_38674_new_n1537_; 
wire alu__abc_38674_new_n1538_; 
wire alu__abc_38674_new_n1539_; 
wire alu__abc_38674_new_n153_; 
wire alu__abc_38674_new_n1540_; 
wire alu__abc_38674_new_n1541_; 
wire alu__abc_38674_new_n1542_; 
wire alu__abc_38674_new_n1543_; 
wire alu__abc_38674_new_n1544_; 
wire alu__abc_38674_new_n1545_; 
wire alu__abc_38674_new_n1547_; 
wire alu__abc_38674_new_n1548_; 
wire alu__abc_38674_new_n1549_; 
wire alu__abc_38674_new_n154_; 
wire alu__abc_38674_new_n1550_; 
wire alu__abc_38674_new_n1551_; 
wire alu__abc_38674_new_n1552_; 
wire alu__abc_38674_new_n1553_; 
wire alu__abc_38674_new_n1554_; 
wire alu__abc_38674_new_n1555_; 
wire alu__abc_38674_new_n1556_; 
wire alu__abc_38674_new_n1557_; 
wire alu__abc_38674_new_n1558_; 
wire alu__abc_38674_new_n1559_; 
wire alu__abc_38674_new_n155_; 
wire alu__abc_38674_new_n1560_; 
wire alu__abc_38674_new_n1561_; 
wire alu__abc_38674_new_n1562_; 
wire alu__abc_38674_new_n1563_; 
wire alu__abc_38674_new_n1564_; 
wire alu__abc_38674_new_n1565_; 
wire alu__abc_38674_new_n1566_; 
wire alu__abc_38674_new_n1567_; 
wire alu__abc_38674_new_n1568_; 
wire alu__abc_38674_new_n1569_; 
wire alu__abc_38674_new_n156_; 
wire alu__abc_38674_new_n1570_; 
wire alu__abc_38674_new_n1572_; 
wire alu__abc_38674_new_n1573_; 
wire alu__abc_38674_new_n1574_; 
wire alu__abc_38674_new_n1575_; 
wire alu__abc_38674_new_n1576_; 
wire alu__abc_38674_new_n1577_; 
wire alu__abc_38674_new_n1578_; 
wire alu__abc_38674_new_n1579_; 
wire alu__abc_38674_new_n157_; 
wire alu__abc_38674_new_n1580_; 
wire alu__abc_38674_new_n1581_; 
wire alu__abc_38674_new_n1582_; 
wire alu__abc_38674_new_n1583_; 
wire alu__abc_38674_new_n1584_; 
wire alu__abc_38674_new_n1585_; 
wire alu__abc_38674_new_n1586_; 
wire alu__abc_38674_new_n1587_; 
wire alu__abc_38674_new_n1588_; 
wire alu__abc_38674_new_n1589_; 
wire alu__abc_38674_new_n158_; 
wire alu__abc_38674_new_n1590_; 
wire alu__abc_38674_new_n1591_; 
wire alu__abc_38674_new_n1592_; 
wire alu__abc_38674_new_n1593_; 
wire alu__abc_38674_new_n1594_; 
wire alu__abc_38674_new_n1595_; 
wire alu__abc_38674_new_n1596_; 
wire alu__abc_38674_new_n1597_; 
wire alu__abc_38674_new_n1598_; 
wire alu__abc_38674_new_n1599_; 
wire alu__abc_38674_new_n159_; 
wire alu__abc_38674_new_n1601_; 
wire alu__abc_38674_new_n1602_; 
wire alu__abc_38674_new_n1603_; 
wire alu__abc_38674_new_n1604_; 
wire alu__abc_38674_new_n1605_; 
wire alu__abc_38674_new_n1606_; 
wire alu__abc_38674_new_n1607_; 
wire alu__abc_38674_new_n1608_; 
wire alu__abc_38674_new_n1609_; 
wire alu__abc_38674_new_n160_; 
wire alu__abc_38674_new_n1610_; 
wire alu__abc_38674_new_n1611_; 
wire alu__abc_38674_new_n1612_; 
wire alu__abc_38674_new_n1613_; 
wire alu__abc_38674_new_n1614_; 
wire alu__abc_38674_new_n1615_; 
wire alu__abc_38674_new_n1616_; 
wire alu__abc_38674_new_n1617_; 
wire alu__abc_38674_new_n1618_; 
wire alu__abc_38674_new_n1619_; 
wire alu__abc_38674_new_n161_; 
wire alu__abc_38674_new_n1620_; 
wire alu__abc_38674_new_n1621_; 
wire alu__abc_38674_new_n1622_; 
wire alu__abc_38674_new_n1624_; 
wire alu__abc_38674_new_n1625_; 
wire alu__abc_38674_new_n1626_; 
wire alu__abc_38674_new_n1627_; 
wire alu__abc_38674_new_n1628_; 
wire alu__abc_38674_new_n1629_; 
wire alu__abc_38674_new_n162_; 
wire alu__abc_38674_new_n1630_; 
wire alu__abc_38674_new_n1631_; 
wire alu__abc_38674_new_n1632_; 
wire alu__abc_38674_new_n1633_; 
wire alu__abc_38674_new_n1634_; 
wire alu__abc_38674_new_n1635_; 
wire alu__abc_38674_new_n1636_; 
wire alu__abc_38674_new_n1637_; 
wire alu__abc_38674_new_n1638_; 
wire alu__abc_38674_new_n1639_; 
wire alu__abc_38674_new_n163_; 
wire alu__abc_38674_new_n1640_; 
wire alu__abc_38674_new_n1641_; 
wire alu__abc_38674_new_n1642_; 
wire alu__abc_38674_new_n1643_; 
wire alu__abc_38674_new_n1644_; 
wire alu__abc_38674_new_n1645_; 
wire alu__abc_38674_new_n1646_; 
wire alu__abc_38674_new_n1647_; 
wire alu__abc_38674_new_n1649_; 
wire alu__abc_38674_new_n164_; 
wire alu__abc_38674_new_n1650_; 
wire alu__abc_38674_new_n1651_; 
wire alu__abc_38674_new_n1652_; 
wire alu__abc_38674_new_n1653_; 
wire alu__abc_38674_new_n1654_; 
wire alu__abc_38674_new_n1655_; 
wire alu__abc_38674_new_n1656_; 
wire alu__abc_38674_new_n1657_; 
wire alu__abc_38674_new_n1658_; 
wire alu__abc_38674_new_n1659_; 
wire alu__abc_38674_new_n165_; 
wire alu__abc_38674_new_n1660_; 
wire alu__abc_38674_new_n1661_; 
wire alu__abc_38674_new_n1662_; 
wire alu__abc_38674_new_n1663_; 
wire alu__abc_38674_new_n1664_; 
wire alu__abc_38674_new_n1665_; 
wire alu__abc_38674_new_n1666_; 
wire alu__abc_38674_new_n1667_; 
wire alu__abc_38674_new_n1668_; 
wire alu__abc_38674_new_n1669_; 
wire alu__abc_38674_new_n166_; 
wire alu__abc_38674_new_n1671_; 
wire alu__abc_38674_new_n1672_; 
wire alu__abc_38674_new_n1673_; 
wire alu__abc_38674_new_n1674_; 
wire alu__abc_38674_new_n1675_; 
wire alu__abc_38674_new_n1676_; 
wire alu__abc_38674_new_n1677_; 
wire alu__abc_38674_new_n1678_; 
wire alu__abc_38674_new_n1679_; 
wire alu__abc_38674_new_n167_; 
wire alu__abc_38674_new_n1680_; 
wire alu__abc_38674_new_n1681_; 
wire alu__abc_38674_new_n1682_; 
wire alu__abc_38674_new_n1683_; 
wire alu__abc_38674_new_n1684_; 
wire alu__abc_38674_new_n1685_; 
wire alu__abc_38674_new_n1686_; 
wire alu__abc_38674_new_n1687_; 
wire alu__abc_38674_new_n1688_; 
wire alu__abc_38674_new_n1689_; 
wire alu__abc_38674_new_n168_; 
wire alu__abc_38674_new_n1690_; 
wire alu__abc_38674_new_n1691_; 
wire alu__abc_38674_new_n1692_; 
wire alu__abc_38674_new_n1693_; 
wire alu__abc_38674_new_n1695_; 
wire alu__abc_38674_new_n1696_; 
wire alu__abc_38674_new_n1697_; 
wire alu__abc_38674_new_n1698_; 
wire alu__abc_38674_new_n1699_; 
wire alu__abc_38674_new_n169_; 
wire alu__abc_38674_new_n1700_; 
wire alu__abc_38674_new_n1701_; 
wire alu__abc_38674_new_n1702_; 
wire alu__abc_38674_new_n1703_; 
wire alu__abc_38674_new_n1704_; 
wire alu__abc_38674_new_n1705_; 
wire alu__abc_38674_new_n1706_; 
wire alu__abc_38674_new_n1707_; 
wire alu__abc_38674_new_n1708_; 
wire alu__abc_38674_new_n1709_; 
wire alu__abc_38674_new_n170_; 
wire alu__abc_38674_new_n1710_; 
wire alu__abc_38674_new_n1711_; 
wire alu__abc_38674_new_n1712_; 
wire alu__abc_38674_new_n1713_; 
wire alu__abc_38674_new_n1714_; 
wire alu__abc_38674_new_n1715_; 
wire alu__abc_38674_new_n1716_; 
wire alu__abc_38674_new_n1717_; 
wire alu__abc_38674_new_n1718_; 
wire alu__abc_38674_new_n1719_; 
wire alu__abc_38674_new_n171_; 
wire alu__abc_38674_new_n1720_; 
wire alu__abc_38674_new_n1723_; 
wire alu__abc_38674_new_n1724_; 
wire alu__abc_38674_new_n1725_; 
wire alu__abc_38674_new_n1726_; 
wire alu__abc_38674_new_n1727_; 
wire alu__abc_38674_new_n1728_; 
wire alu__abc_38674_new_n1729_; 
wire alu__abc_38674_new_n172_; 
wire alu__abc_38674_new_n1730_; 
wire alu__abc_38674_new_n173_; 
wire alu__abc_38674_new_n174_; 
wire alu__abc_38674_new_n175_; 
wire alu__abc_38674_new_n176_; 
wire alu__abc_38674_new_n177_; 
wire alu__abc_38674_new_n178_; 
wire alu__abc_38674_new_n179_; 
wire alu__abc_38674_new_n180_; 
wire alu__abc_38674_new_n181_; 
wire alu__abc_38674_new_n182_; 
wire alu__abc_38674_new_n183_; 
wire alu__abc_38674_new_n184_; 
wire alu__abc_38674_new_n185_; 
wire alu__abc_38674_new_n186_; 
wire alu__abc_38674_new_n187_; 
wire alu__abc_38674_new_n188_; 
wire alu__abc_38674_new_n189_; 
wire alu__abc_38674_new_n190_; 
wire alu__abc_38674_new_n191_; 
wire alu__abc_38674_new_n192_; 
wire alu__abc_38674_new_n193_; 
wire alu__abc_38674_new_n194_; 
wire alu__abc_38674_new_n195_; 
wire alu__abc_38674_new_n196_; 
wire alu__abc_38674_new_n197_; 
wire alu__abc_38674_new_n198_; 
wire alu__abc_38674_new_n199_; 
wire alu__abc_38674_new_n200_; 
wire alu__abc_38674_new_n201_; 
wire alu__abc_38674_new_n202_; 
wire alu__abc_38674_new_n203_; 
wire alu__abc_38674_new_n204_; 
wire alu__abc_38674_new_n205_; 
wire alu__abc_38674_new_n206_; 
wire alu__abc_38674_new_n207_; 
wire alu__abc_38674_new_n208_; 
wire alu__abc_38674_new_n209_; 
wire alu__abc_38674_new_n210_; 
wire alu__abc_38674_new_n211_; 
wire alu__abc_38674_new_n212_; 
wire alu__abc_38674_new_n213_; 
wire alu__abc_38674_new_n214_; 
wire alu__abc_38674_new_n215_; 
wire alu__abc_38674_new_n216_; 
wire alu__abc_38674_new_n217_; 
wire alu__abc_38674_new_n218_; 
wire alu__abc_38674_new_n219_; 
wire alu__abc_38674_new_n220_; 
wire alu__abc_38674_new_n221_; 
wire alu__abc_38674_new_n222_; 
wire alu__abc_38674_new_n223_; 
wire alu__abc_38674_new_n224_; 
wire alu__abc_38674_new_n225_; 
wire alu__abc_38674_new_n226_; 
wire alu__abc_38674_new_n227_; 
wire alu__abc_38674_new_n228_; 
wire alu__abc_38674_new_n229_; 
wire alu__abc_38674_new_n230_; 
wire alu__abc_38674_new_n231_; 
wire alu__abc_38674_new_n232_; 
wire alu__abc_38674_new_n233_; 
wire alu__abc_38674_new_n234_; 
wire alu__abc_38674_new_n235_; 
wire alu__abc_38674_new_n236_; 
wire alu__abc_38674_new_n237_; 
wire alu__abc_38674_new_n238_; 
wire alu__abc_38674_new_n239_; 
wire alu__abc_38674_new_n240_; 
wire alu__abc_38674_new_n241_; 
wire alu__abc_38674_new_n242_; 
wire alu__abc_38674_new_n243_; 
wire alu__abc_38674_new_n244_; 
wire alu__abc_38674_new_n245_; 
wire alu__abc_38674_new_n246_; 
wire alu__abc_38674_new_n247_; 
wire alu__abc_38674_new_n248_; 
wire alu__abc_38674_new_n249_; 
wire alu__abc_38674_new_n250_; 
wire alu__abc_38674_new_n251_; 
wire alu__abc_38674_new_n252_; 
wire alu__abc_38674_new_n253_; 
wire alu__abc_38674_new_n254_; 
wire alu__abc_38674_new_n255_; 
wire alu__abc_38674_new_n256_; 
wire alu__abc_38674_new_n257_; 
wire alu__abc_38674_new_n258_; 
wire alu__abc_38674_new_n259_; 
wire alu__abc_38674_new_n260_; 
wire alu__abc_38674_new_n261_; 
wire alu__abc_38674_new_n262_; 
wire alu__abc_38674_new_n263_; 
wire alu__abc_38674_new_n264_; 
wire alu__abc_38674_new_n265_; 
wire alu__abc_38674_new_n266_; 
wire alu__abc_38674_new_n267_; 
wire alu__abc_38674_new_n268_; 
wire alu__abc_38674_new_n269_; 
wire alu__abc_38674_new_n270_; 
wire alu__abc_38674_new_n271_; 
wire alu__abc_38674_new_n272_; 
wire alu__abc_38674_new_n273_; 
wire alu__abc_38674_new_n274_; 
wire alu__abc_38674_new_n275_; 
wire alu__abc_38674_new_n277_; 
wire alu__abc_38674_new_n278_; 
wire alu__abc_38674_new_n279_; 
wire alu__abc_38674_new_n280_; 
wire alu__abc_38674_new_n281_; 
wire alu__abc_38674_new_n282_; 
wire alu__abc_38674_new_n283_; 
wire alu__abc_38674_new_n284_; 
wire alu__abc_38674_new_n285_; 
wire alu__abc_38674_new_n286_; 
wire alu__abc_38674_new_n288_; 
wire alu__abc_38674_new_n289_; 
wire alu__abc_38674_new_n290_; 
wire alu__abc_38674_new_n291_; 
wire alu__abc_38674_new_n292_; 
wire alu__abc_38674_new_n294_; 
wire alu__abc_38674_new_n295_; 
wire alu__abc_38674_new_n296_; 
wire alu__abc_38674_new_n297_; 
wire alu__abc_38674_new_n298_; 
wire alu__abc_38674_new_n299_; 
wire alu__abc_38674_new_n300_; 
wire alu__abc_38674_new_n301_; 
wire alu__abc_38674_new_n302_; 
wire alu__abc_38674_new_n303_; 
wire alu__abc_38674_new_n304_; 
wire alu__abc_38674_new_n305_; 
wire alu__abc_38674_new_n306_; 
wire alu__abc_38674_new_n307_; 
wire alu__abc_38674_new_n308_; 
wire alu__abc_38674_new_n309_; 
wire alu__abc_38674_new_n310_; 
wire alu__abc_38674_new_n311_; 
wire alu__abc_38674_new_n312_; 
wire alu__abc_38674_new_n313_; 
wire alu__abc_38674_new_n314_; 
wire alu__abc_38674_new_n315_; 
wire alu__abc_38674_new_n316_; 
wire alu__abc_38674_new_n317_; 
wire alu__abc_38674_new_n318_; 
wire alu__abc_38674_new_n319_; 
wire alu__abc_38674_new_n320_; 
wire alu__abc_38674_new_n321_; 
wire alu__abc_38674_new_n322_; 
wire alu__abc_38674_new_n323_; 
wire alu__abc_38674_new_n324_; 
wire alu__abc_38674_new_n325_; 
wire alu__abc_38674_new_n326_; 
wire alu__abc_38674_new_n327_; 
wire alu__abc_38674_new_n328_; 
wire alu__abc_38674_new_n329_; 
wire alu__abc_38674_new_n330_; 
wire alu__abc_38674_new_n331_; 
wire alu__abc_38674_new_n332_; 
wire alu__abc_38674_new_n333_; 
wire alu__abc_38674_new_n334_; 
wire alu__abc_38674_new_n335_; 
wire alu__abc_38674_new_n336_; 
wire alu__abc_38674_new_n337_; 
wire alu__abc_38674_new_n338_; 
wire alu__abc_38674_new_n339_; 
wire alu__abc_38674_new_n340_; 
wire alu__abc_38674_new_n341_; 
wire alu__abc_38674_new_n342_; 
wire alu__abc_38674_new_n343_; 
wire alu__abc_38674_new_n344_; 
wire alu__abc_38674_new_n345_; 
wire alu__abc_38674_new_n346_; 
wire alu__abc_38674_new_n347_; 
wire alu__abc_38674_new_n348_; 
wire alu__abc_38674_new_n349_; 
wire alu__abc_38674_new_n350_; 
wire alu__abc_38674_new_n351_; 
wire alu__abc_38674_new_n352_; 
wire alu__abc_38674_new_n353_; 
wire alu__abc_38674_new_n354_; 
wire alu__abc_38674_new_n355_; 
wire alu__abc_38674_new_n356_; 
wire alu__abc_38674_new_n357_; 
wire alu__abc_38674_new_n358_; 
wire alu__abc_38674_new_n359_; 
wire alu__abc_38674_new_n360_; 
wire alu__abc_38674_new_n361_; 
wire alu__abc_38674_new_n362_; 
wire alu__abc_38674_new_n363_; 
wire alu__abc_38674_new_n364_; 
wire alu__abc_38674_new_n365_; 
wire alu__abc_38674_new_n366_; 
wire alu__abc_38674_new_n367_; 
wire alu__abc_38674_new_n368_; 
wire alu__abc_38674_new_n369_; 
wire alu__abc_38674_new_n370_; 
wire alu__abc_38674_new_n371_; 
wire alu__abc_38674_new_n372_; 
wire alu__abc_38674_new_n373_; 
wire alu__abc_38674_new_n374_; 
wire alu__abc_38674_new_n375_; 
wire alu__abc_38674_new_n376_; 
wire alu__abc_38674_new_n377_; 
wire alu__abc_38674_new_n378_; 
wire alu__abc_38674_new_n379_; 
wire alu__abc_38674_new_n381_; 
wire alu__abc_38674_new_n382_; 
wire alu__abc_38674_new_n383_; 
wire alu__abc_38674_new_n384_; 
wire alu__abc_38674_new_n385_; 
wire alu__abc_38674_new_n386_; 
wire alu__abc_38674_new_n387_; 
wire alu__abc_38674_new_n388_; 
wire alu__abc_38674_new_n389_; 
wire alu__abc_38674_new_n390_; 
wire alu__abc_38674_new_n391_; 
wire alu__abc_38674_new_n392_; 
wire alu__abc_38674_new_n393_; 
wire alu__abc_38674_new_n394_; 
wire alu__abc_38674_new_n395_; 
wire alu__abc_38674_new_n396_; 
wire alu__abc_38674_new_n397_; 
wire alu__abc_38674_new_n398_; 
wire alu__abc_38674_new_n399_; 
wire alu__abc_38674_new_n400_; 
wire alu__abc_38674_new_n401_; 
wire alu__abc_38674_new_n402_; 
wire alu__abc_38674_new_n403_; 
wire alu__abc_38674_new_n404_; 
wire alu__abc_38674_new_n405_; 
wire alu__abc_38674_new_n406_; 
wire alu__abc_38674_new_n407_; 
wire alu__abc_38674_new_n408_; 
wire alu__abc_38674_new_n409_; 
wire alu__abc_38674_new_n410_; 
wire alu__abc_38674_new_n411_; 
wire alu__abc_38674_new_n412_; 
wire alu__abc_38674_new_n413_; 
wire alu__abc_38674_new_n414_; 
wire alu__abc_38674_new_n415_; 
wire alu__abc_38674_new_n416_; 
wire alu__abc_38674_new_n417_; 
wire alu__abc_38674_new_n418_; 
wire alu__abc_38674_new_n419_; 
wire alu__abc_38674_new_n420_; 
wire alu__abc_38674_new_n421_; 
wire alu__abc_38674_new_n422_; 
wire alu__abc_38674_new_n423_; 
wire alu__abc_38674_new_n424_; 
wire alu__abc_38674_new_n425_; 
wire alu__abc_38674_new_n426_; 
wire alu__abc_38674_new_n427_; 
wire alu__abc_38674_new_n428_; 
wire alu__abc_38674_new_n429_; 
wire alu__abc_38674_new_n430_; 
wire alu__abc_38674_new_n431_; 
wire alu__abc_38674_new_n432_; 
wire alu__abc_38674_new_n433_; 
wire alu__abc_38674_new_n434_; 
wire alu__abc_38674_new_n435_; 
wire alu__abc_38674_new_n436_; 
wire alu__abc_38674_new_n437_; 
wire alu__abc_38674_new_n438_; 
wire alu__abc_38674_new_n439_; 
wire alu__abc_38674_new_n440_; 
wire alu__abc_38674_new_n441_; 
wire alu__abc_38674_new_n442_; 
wire alu__abc_38674_new_n443_; 
wire alu__abc_38674_new_n444_; 
wire alu__abc_38674_new_n445_; 
wire alu__abc_38674_new_n446_; 
wire alu__abc_38674_new_n447_; 
wire alu__abc_38674_new_n448_; 
wire alu__abc_38674_new_n449_; 
wire alu__abc_38674_new_n450_; 
wire alu__abc_38674_new_n451_; 
wire alu__abc_38674_new_n452_; 
wire alu__abc_38674_new_n453_; 
wire alu__abc_38674_new_n454_; 
wire alu__abc_38674_new_n455_; 
wire alu__abc_38674_new_n456_; 
wire alu__abc_38674_new_n457_; 
wire alu__abc_38674_new_n458_; 
wire alu__abc_38674_new_n459_; 
wire alu__abc_38674_new_n460_; 
wire alu__abc_38674_new_n461_; 
wire alu__abc_38674_new_n462_; 
wire alu__abc_38674_new_n463_; 
wire alu__abc_38674_new_n464_; 
wire alu__abc_38674_new_n465_; 
wire alu__abc_38674_new_n466_; 
wire alu__abc_38674_new_n467_; 
wire alu__abc_38674_new_n468_; 
wire alu__abc_38674_new_n469_; 
wire alu__abc_38674_new_n470_; 
wire alu__abc_38674_new_n471_; 
wire alu__abc_38674_new_n472_; 
wire alu__abc_38674_new_n473_; 
wire alu__abc_38674_new_n474_; 
wire alu__abc_38674_new_n475_; 
wire alu__abc_38674_new_n476_; 
wire alu__abc_38674_new_n477_; 
wire alu__abc_38674_new_n478_; 
wire alu__abc_38674_new_n479_; 
wire alu__abc_38674_new_n480_; 
wire alu__abc_38674_new_n481_; 
wire alu__abc_38674_new_n482_; 
wire alu__abc_38674_new_n483_; 
wire alu__abc_38674_new_n484_; 
wire alu__abc_38674_new_n485_; 
wire alu__abc_38674_new_n486_; 
wire alu__abc_38674_new_n487_; 
wire alu__abc_38674_new_n488_; 
wire alu__abc_38674_new_n489_; 
wire alu__abc_38674_new_n490_; 
wire alu__abc_38674_new_n491_; 
wire alu__abc_38674_new_n492_; 
wire alu__abc_38674_new_n493_; 
wire alu__abc_38674_new_n494_; 
wire alu__abc_38674_new_n495_; 
wire alu__abc_38674_new_n496_; 
wire alu__abc_38674_new_n497_; 
wire alu__abc_38674_new_n498_; 
wire alu__abc_38674_new_n499_; 
wire alu__abc_38674_new_n500_; 
wire alu__abc_38674_new_n501_; 
wire alu__abc_38674_new_n502_; 
wire alu__abc_38674_new_n503_; 
wire alu__abc_38674_new_n504_; 
wire alu__abc_38674_new_n505_; 
wire alu__abc_38674_new_n506_; 
wire alu__abc_38674_new_n507_; 
wire alu__abc_38674_new_n508_; 
wire alu__abc_38674_new_n509_; 
wire alu__abc_38674_new_n510_; 
wire alu__abc_38674_new_n511_; 
wire alu__abc_38674_new_n512_; 
wire alu__abc_38674_new_n513_; 
wire alu__abc_38674_new_n514_; 
wire alu__abc_38674_new_n515_; 
wire alu__abc_38674_new_n516_; 
wire alu__abc_38674_new_n517_; 
wire alu__abc_38674_new_n518_; 
wire alu__abc_38674_new_n519_; 
wire alu__abc_38674_new_n520_; 
wire alu__abc_38674_new_n521_; 
wire alu__abc_38674_new_n522_; 
wire alu__abc_38674_new_n523_; 
wire alu__abc_38674_new_n524_; 
wire alu__abc_38674_new_n525_; 
wire alu__abc_38674_new_n526_; 
wire alu__abc_38674_new_n527_; 
wire alu__abc_38674_new_n528_; 
wire alu__abc_38674_new_n529_; 
wire alu__abc_38674_new_n530_; 
wire alu__abc_38674_new_n531_; 
wire alu__abc_38674_new_n532_; 
wire alu__abc_38674_new_n533_; 
wire alu__abc_38674_new_n534_; 
wire alu__abc_38674_new_n535_; 
wire alu__abc_38674_new_n536_; 
wire alu__abc_38674_new_n537_; 
wire alu__abc_38674_new_n538_; 
wire alu__abc_38674_new_n539_; 
wire alu__abc_38674_new_n540_; 
wire alu__abc_38674_new_n541_; 
wire alu__abc_38674_new_n542_; 
wire alu__abc_38674_new_n543_; 
wire alu__abc_38674_new_n544_; 
wire alu__abc_38674_new_n545_; 
wire alu__abc_38674_new_n546_; 
wire alu__abc_38674_new_n547_; 
wire alu__abc_38674_new_n548_; 
wire alu__abc_38674_new_n549_; 
wire alu__abc_38674_new_n550_; 
wire alu__abc_38674_new_n551_; 
wire alu__abc_38674_new_n552_; 
wire alu__abc_38674_new_n553_; 
wire alu__abc_38674_new_n554_; 
wire alu__abc_38674_new_n555_; 
wire alu__abc_38674_new_n556_; 
wire alu__abc_38674_new_n557_; 
wire alu__abc_38674_new_n558_; 
wire alu__abc_38674_new_n559_; 
wire alu__abc_38674_new_n560_; 
wire alu__abc_38674_new_n561_; 
wire alu__abc_38674_new_n562_; 
wire alu__abc_38674_new_n563_; 
wire alu__abc_38674_new_n564_; 
wire alu__abc_38674_new_n565_; 
wire alu__abc_38674_new_n566_; 
wire alu__abc_38674_new_n567_; 
wire alu__abc_38674_new_n568_; 
wire alu__abc_38674_new_n569_; 
wire alu__abc_38674_new_n570_; 
wire alu__abc_38674_new_n571_; 
wire alu__abc_38674_new_n572_; 
wire alu__abc_38674_new_n573_; 
wire alu__abc_38674_new_n574_; 
wire alu__abc_38674_new_n575_; 
wire alu__abc_38674_new_n576_; 
wire alu__abc_38674_new_n577_; 
wire alu__abc_38674_new_n578_; 
wire alu__abc_38674_new_n579_; 
wire alu__abc_38674_new_n580_; 
wire alu__abc_38674_new_n581_; 
wire alu__abc_38674_new_n582_; 
wire alu__abc_38674_new_n583_; 
wire alu__abc_38674_new_n584_; 
wire alu__abc_38674_new_n585_; 
wire alu__abc_38674_new_n586_; 
wire alu__abc_38674_new_n587_; 
wire alu__abc_38674_new_n588_; 
wire alu__abc_38674_new_n589_; 
wire alu__abc_38674_new_n590_; 
wire alu__abc_38674_new_n591_; 
wire alu__abc_38674_new_n592_; 
wire alu__abc_38674_new_n593_; 
wire alu__abc_38674_new_n594_; 
wire alu__abc_38674_new_n595_; 
wire alu__abc_38674_new_n596_; 
wire alu__abc_38674_new_n597_; 
wire alu__abc_38674_new_n598_; 
wire alu__abc_38674_new_n599_; 
wire alu__abc_38674_new_n600_; 
wire alu__abc_38674_new_n601_; 
wire alu__abc_38674_new_n602_; 
wire alu__abc_38674_new_n603_; 
wire alu__abc_38674_new_n604_; 
wire alu__abc_38674_new_n605_; 
wire alu__abc_38674_new_n606_; 
wire alu__abc_38674_new_n607_; 
wire alu__abc_38674_new_n608_; 
wire alu__abc_38674_new_n609_; 
wire alu__abc_38674_new_n610_; 
wire alu__abc_38674_new_n611_; 
wire alu__abc_38674_new_n612_; 
wire alu__abc_38674_new_n613_; 
wire alu__abc_38674_new_n614_; 
wire alu__abc_38674_new_n615_; 
wire alu__abc_38674_new_n616_; 
wire alu__abc_38674_new_n617_; 
wire alu__abc_38674_new_n618_; 
wire alu__abc_38674_new_n619_; 
wire alu__abc_38674_new_n620_; 
wire alu__abc_38674_new_n621_; 
wire alu__abc_38674_new_n622_; 
wire alu__abc_38674_new_n623_; 
wire alu__abc_38674_new_n624_; 
wire alu__abc_38674_new_n625_; 
wire alu__abc_38674_new_n626_; 
wire alu__abc_38674_new_n627_; 
wire alu__abc_38674_new_n629_; 
wire alu__abc_38674_new_n630_; 
wire alu__abc_38674_new_n631_; 
wire alu__abc_38674_new_n632_; 
wire alu__abc_38674_new_n633_; 
wire alu__abc_38674_new_n634_; 
wire alu__abc_38674_new_n635_; 
wire alu__abc_38674_new_n636_; 
wire alu__abc_38674_new_n637_; 
wire alu__abc_38674_new_n638_; 
wire alu__abc_38674_new_n639_; 
wire alu__abc_38674_new_n640_; 
wire alu__abc_38674_new_n641_; 
wire alu__abc_38674_new_n642_; 
wire alu__abc_38674_new_n643_; 
wire alu__abc_38674_new_n644_; 
wire alu__abc_38674_new_n645_; 
wire alu__abc_38674_new_n646_; 
wire alu__abc_38674_new_n647_; 
wire alu__abc_38674_new_n648_; 
wire alu__abc_38674_new_n649_; 
wire alu__abc_38674_new_n650_; 
wire alu__abc_38674_new_n651_; 
wire alu__abc_38674_new_n652_; 
wire alu__abc_38674_new_n653_; 
wire alu__abc_38674_new_n654_; 
wire alu__abc_38674_new_n655_; 
wire alu__abc_38674_new_n656_; 
wire alu__abc_38674_new_n657_; 
wire alu__abc_38674_new_n658_; 
wire alu__abc_38674_new_n659_; 
wire alu__abc_38674_new_n660_; 
wire alu__abc_38674_new_n661_; 
wire alu__abc_38674_new_n662_; 
wire alu__abc_38674_new_n663_; 
wire alu__abc_38674_new_n664_; 
wire alu__abc_38674_new_n665_; 
wire alu__abc_38674_new_n666_; 
wire alu__abc_38674_new_n667_; 
wire alu__abc_38674_new_n668_; 
wire alu__abc_38674_new_n669_; 
wire alu__abc_38674_new_n670_; 
wire alu__abc_38674_new_n671_; 
wire alu__abc_38674_new_n672_; 
wire alu__abc_38674_new_n673_; 
wire alu__abc_38674_new_n674_; 
wire alu__abc_38674_new_n675_; 
wire alu__abc_38674_new_n676_; 
wire alu__abc_38674_new_n677_; 
wire alu__abc_38674_new_n678_; 
wire alu__abc_38674_new_n679_; 
wire alu__abc_38674_new_n680_; 
wire alu__abc_38674_new_n681_; 
wire alu__abc_38674_new_n682_; 
wire alu__abc_38674_new_n683_; 
wire alu__abc_38674_new_n684_; 
wire alu__abc_38674_new_n685_; 
wire alu__abc_38674_new_n686_; 
wire alu__abc_38674_new_n687_; 
wire alu__abc_38674_new_n688_; 
wire alu__abc_38674_new_n689_; 
wire alu__abc_38674_new_n690_; 
wire alu__abc_38674_new_n691_; 
wire alu__abc_38674_new_n692_; 
wire alu__abc_38674_new_n693_; 
wire alu__abc_38674_new_n694_; 
wire alu__abc_38674_new_n695_; 
wire alu__abc_38674_new_n696_; 
wire alu__abc_38674_new_n697_; 
wire alu__abc_38674_new_n698_; 
wire alu__abc_38674_new_n699_; 
wire alu__abc_38674_new_n700_; 
wire alu__abc_38674_new_n701_; 
wire alu__abc_38674_new_n702_; 
wire alu__abc_38674_new_n703_; 
wire alu__abc_38674_new_n704_; 
wire alu__abc_38674_new_n705_; 
wire alu__abc_38674_new_n706_; 
wire alu__abc_38674_new_n707_; 
wire alu__abc_38674_new_n708_; 
wire alu__abc_38674_new_n709_; 
wire alu__abc_38674_new_n710_; 
wire alu__abc_38674_new_n711_; 
wire alu__abc_38674_new_n712_; 
wire alu__abc_38674_new_n713_; 
wire alu__abc_38674_new_n714_; 
wire alu__abc_38674_new_n715_; 
wire alu__abc_38674_new_n717_; 
wire alu__abc_38674_new_n718_; 
wire alu__abc_38674_new_n719_; 
wire alu__abc_38674_new_n720_; 
wire alu__abc_38674_new_n721_; 
wire alu__abc_38674_new_n722_; 
wire alu__abc_38674_new_n723_; 
wire alu__abc_38674_new_n724_; 
wire alu__abc_38674_new_n725_; 
wire alu__abc_38674_new_n726_; 
wire alu__abc_38674_new_n727_; 
wire alu__abc_38674_new_n728_; 
wire alu__abc_38674_new_n729_; 
wire alu__abc_38674_new_n730_; 
wire alu__abc_38674_new_n731_; 
wire alu__abc_38674_new_n732_; 
wire alu__abc_38674_new_n733_; 
wire alu__abc_38674_new_n734_; 
wire alu__abc_38674_new_n735_; 
wire alu__abc_38674_new_n736_; 
wire alu__abc_38674_new_n737_; 
wire alu__abc_38674_new_n738_; 
wire alu__abc_38674_new_n739_; 
wire alu__abc_38674_new_n740_; 
wire alu__abc_38674_new_n741_; 
wire alu__abc_38674_new_n742_; 
wire alu__abc_38674_new_n743_; 
wire alu__abc_38674_new_n744_; 
wire alu__abc_38674_new_n745_; 
wire alu__abc_38674_new_n746_; 
wire alu__abc_38674_new_n747_; 
wire alu__abc_38674_new_n748_; 
wire alu__abc_38674_new_n749_; 
wire alu__abc_38674_new_n750_; 
wire alu__abc_38674_new_n751_; 
wire alu__abc_38674_new_n752_; 
wire alu__abc_38674_new_n753_; 
wire alu__abc_38674_new_n754_; 
wire alu__abc_38674_new_n755_; 
wire alu__abc_38674_new_n756_; 
wire alu__abc_38674_new_n757_; 
wire alu__abc_38674_new_n758_; 
wire alu__abc_38674_new_n759_; 
wire alu__abc_38674_new_n760_; 
wire alu__abc_38674_new_n761_; 
wire alu__abc_38674_new_n762_; 
wire alu__abc_38674_new_n763_; 
wire alu__abc_38674_new_n764_; 
wire alu__abc_38674_new_n765_; 
wire alu__abc_38674_new_n766_; 
wire alu__abc_38674_new_n767_; 
wire alu__abc_38674_new_n768_; 
wire alu__abc_38674_new_n769_; 
wire alu__abc_38674_new_n770_; 
wire alu__abc_38674_new_n771_; 
wire alu__abc_38674_new_n772_; 
wire alu__abc_38674_new_n773_; 
wire alu__abc_38674_new_n774_; 
wire alu__abc_38674_new_n775_; 
wire alu__abc_38674_new_n776_; 
wire alu__abc_38674_new_n777_; 
wire alu__abc_38674_new_n778_; 
wire alu__abc_38674_new_n779_; 
wire alu__abc_38674_new_n780_; 
wire alu__abc_38674_new_n781_; 
wire alu__abc_38674_new_n782_; 
wire alu__abc_38674_new_n783_; 
wire alu__abc_38674_new_n784_; 
wire alu__abc_38674_new_n785_; 
wire alu__abc_38674_new_n786_; 
wire alu__abc_38674_new_n787_; 
wire alu__abc_38674_new_n788_; 
wire alu__abc_38674_new_n789_; 
wire alu__abc_38674_new_n790_; 
wire alu__abc_38674_new_n791_; 
wire alu__abc_38674_new_n792_; 
wire alu__abc_38674_new_n793_; 
wire alu__abc_38674_new_n794_; 
wire alu__abc_38674_new_n795_; 
wire alu__abc_38674_new_n796_; 
wire alu__abc_38674_new_n798_; 
wire alu__abc_38674_new_n799_; 
wire alu__abc_38674_new_n800_; 
wire alu__abc_38674_new_n801_; 
wire alu__abc_38674_new_n802_; 
wire alu__abc_38674_new_n803_; 
wire alu__abc_38674_new_n804_; 
wire alu__abc_38674_new_n805_; 
wire alu__abc_38674_new_n806_; 
wire alu__abc_38674_new_n807_; 
wire alu__abc_38674_new_n808_; 
wire alu__abc_38674_new_n809_; 
wire alu__abc_38674_new_n810_; 
wire alu__abc_38674_new_n811_; 
wire alu__abc_38674_new_n812_; 
wire alu__abc_38674_new_n813_; 
wire alu__abc_38674_new_n814_; 
wire alu__abc_38674_new_n815_; 
wire alu__abc_38674_new_n816_; 
wire alu__abc_38674_new_n817_; 
wire alu__abc_38674_new_n818_; 
wire alu__abc_38674_new_n819_; 
wire alu__abc_38674_new_n820_; 
wire alu__abc_38674_new_n821_; 
wire alu__abc_38674_new_n822_; 
wire alu__abc_38674_new_n823_; 
wire alu__abc_38674_new_n824_; 
wire alu__abc_38674_new_n825_; 
wire alu__abc_38674_new_n826_; 
wire alu__abc_38674_new_n827_; 
wire alu__abc_38674_new_n828_; 
wire alu__abc_38674_new_n829_; 
wire alu__abc_38674_new_n830_; 
wire alu__abc_38674_new_n831_; 
wire alu__abc_38674_new_n832_; 
wire alu__abc_38674_new_n833_; 
wire alu__abc_38674_new_n834_; 
wire alu__abc_38674_new_n835_; 
wire alu__abc_38674_new_n836_; 
wire alu__abc_38674_new_n837_; 
wire alu__abc_38674_new_n838_; 
wire alu__abc_38674_new_n839_; 
wire alu__abc_38674_new_n840_; 
wire alu__abc_38674_new_n841_; 
wire alu__abc_38674_new_n842_; 
wire alu__abc_38674_new_n843_; 
wire alu__abc_38674_new_n844_; 
wire alu__abc_38674_new_n845_; 
wire alu__abc_38674_new_n846_; 
wire alu__abc_38674_new_n847_; 
wire alu__abc_38674_new_n848_; 
wire alu__abc_38674_new_n849_; 
wire alu__abc_38674_new_n851_; 
wire alu__abc_38674_new_n852_; 
wire alu__abc_38674_new_n853_; 
wire alu__abc_38674_new_n854_; 
wire alu__abc_38674_new_n855_; 
wire alu__abc_38674_new_n856_; 
wire alu__abc_38674_new_n857_; 
wire alu__abc_38674_new_n858_; 
wire alu__abc_38674_new_n859_; 
wire alu__abc_38674_new_n860_; 
wire alu__abc_38674_new_n861_; 
wire alu__abc_38674_new_n862_; 
wire alu__abc_38674_new_n863_; 
wire alu__abc_38674_new_n864_; 
wire alu__abc_38674_new_n865_; 
wire alu__abc_38674_new_n866_; 
wire alu__abc_38674_new_n867_; 
wire alu__abc_38674_new_n868_; 
wire alu__abc_38674_new_n869_; 
wire alu__abc_38674_new_n870_; 
wire alu__abc_38674_new_n871_; 
wire alu__abc_38674_new_n872_; 
wire alu__abc_38674_new_n873_; 
wire alu__abc_38674_new_n874_; 
wire alu__abc_38674_new_n875_; 
wire alu__abc_38674_new_n876_; 
wire alu__abc_38674_new_n877_; 
wire alu__abc_38674_new_n878_; 
wire alu__abc_38674_new_n879_; 
wire alu__abc_38674_new_n880_; 
wire alu__abc_38674_new_n881_; 
wire alu__abc_38674_new_n882_; 
wire alu__abc_38674_new_n883_; 
wire alu__abc_38674_new_n884_; 
wire alu__abc_38674_new_n885_; 
wire alu__abc_38674_new_n886_; 
wire alu__abc_38674_new_n887_; 
wire alu__abc_38674_new_n888_; 
wire alu__abc_38674_new_n889_; 
wire alu__abc_38674_new_n890_; 
wire alu__abc_38674_new_n891_; 
wire alu__abc_38674_new_n892_; 
wire alu__abc_38674_new_n893_; 
wire alu__abc_38674_new_n894_; 
wire alu__abc_38674_new_n895_; 
wire alu__abc_38674_new_n896_; 
wire alu__abc_38674_new_n897_; 
wire alu__abc_38674_new_n898_; 
wire alu__abc_38674_new_n899_; 
wire alu__abc_38674_new_n900_; 
wire alu__abc_38674_new_n902_; 
wire alu__abc_38674_new_n903_; 
wire alu__abc_38674_new_n904_; 
wire alu__abc_38674_new_n905_; 
wire alu__abc_38674_new_n906_; 
wire alu__abc_38674_new_n907_; 
wire alu__abc_38674_new_n908_; 
wire alu__abc_38674_new_n909_; 
wire alu__abc_38674_new_n910_; 
wire alu__abc_38674_new_n911_; 
wire alu__abc_38674_new_n912_; 
wire alu__abc_38674_new_n913_; 
wire alu__abc_38674_new_n914_; 
wire alu__abc_38674_new_n915_; 
wire alu__abc_38674_new_n916_; 
wire alu__abc_38674_new_n917_; 
wire alu__abc_38674_new_n918_; 
wire alu__abc_38674_new_n919_; 
wire alu__abc_38674_new_n920_; 
wire alu__abc_38674_new_n921_; 
wire alu__abc_38674_new_n922_; 
wire alu__abc_38674_new_n923_; 
wire alu__abc_38674_new_n924_; 
wire alu__abc_38674_new_n925_; 
wire alu__abc_38674_new_n926_; 
wire alu__abc_38674_new_n927_; 
wire alu__abc_38674_new_n928_; 
wire alu__abc_38674_new_n929_; 
wire alu__abc_38674_new_n930_; 
wire alu__abc_38674_new_n931_; 
wire alu__abc_38674_new_n932_; 
wire alu__abc_38674_new_n933_; 
wire alu__abc_38674_new_n934_; 
wire alu__abc_38674_new_n935_; 
wire alu__abc_38674_new_n936_; 
wire alu__abc_38674_new_n937_; 
wire alu__abc_38674_new_n938_; 
wire alu__abc_38674_new_n939_; 
wire alu__abc_38674_new_n941_; 
wire alu__abc_38674_new_n942_; 
wire alu__abc_38674_new_n943_; 
wire alu__abc_38674_new_n944_; 
wire alu__abc_38674_new_n945_; 
wire alu__abc_38674_new_n946_; 
wire alu__abc_38674_new_n947_; 
wire alu__abc_38674_new_n948_; 
wire alu__abc_38674_new_n949_; 
wire alu__abc_38674_new_n950_; 
wire alu__abc_38674_new_n951_; 
wire alu__abc_38674_new_n952_; 
wire alu__abc_38674_new_n953_; 
wire alu__abc_38674_new_n954_; 
wire alu__abc_38674_new_n955_; 
wire alu__abc_38674_new_n956_; 
wire alu__abc_38674_new_n957_; 
wire alu__abc_38674_new_n958_; 
wire alu__abc_38674_new_n959_; 
wire alu__abc_38674_new_n960_; 
wire alu__abc_38674_new_n961_; 
wire alu__abc_38674_new_n962_; 
wire alu__abc_38674_new_n963_; 
wire alu__abc_38674_new_n964_; 
wire alu__abc_38674_new_n965_; 
wire alu__abc_38674_new_n966_; 
wire alu__abc_38674_new_n967_; 
wire alu__abc_38674_new_n968_; 
wire alu__abc_38674_new_n969_; 
wire alu__abc_38674_new_n970_; 
wire alu__abc_38674_new_n971_; 
wire alu__abc_38674_new_n972_; 
wire alu__abc_38674_new_n973_; 
wire alu__abc_38674_new_n974_; 
wire alu__abc_38674_new_n976_; 
wire alu__abc_38674_new_n977_; 
wire alu__abc_38674_new_n978_; 
wire alu__abc_38674_new_n979_; 
wire alu__abc_38674_new_n980_; 
wire alu__abc_38674_new_n981_; 
wire alu__abc_38674_new_n982_; 
wire alu__abc_38674_new_n983_; 
wire alu__abc_38674_new_n984_; 
wire alu__abc_38674_new_n985_; 
wire alu__abc_38674_new_n986_; 
wire alu__abc_38674_new_n987_; 
wire alu__abc_38674_new_n988_; 
wire alu__abc_38674_new_n989_; 
wire alu__abc_38674_new_n990_; 
wire alu__abc_38674_new_n991_; 
wire alu__abc_38674_new_n992_; 
wire alu__abc_38674_new_n993_; 
wire alu__abc_38674_new_n994_; 
wire alu__abc_38674_new_n995_; 
wire alu__abc_38674_new_n996_; 
wire alu__abc_38674_new_n997_; 
wire alu__abc_38674_new_n998_; 
wire alu__abc_38674_new_n999_; 
wire alu_a_i_0_; 
wire alu_a_i_10_; 
wire alu_a_i_11_; 
wire alu_a_i_12_; 
wire alu_a_i_13_; 
wire alu_a_i_14_; 
wire alu_a_i_15_; 
wire alu_a_i_16_; 
wire alu_a_i_17_; 
wire alu_a_i_18_; 
wire alu_a_i_19_; 
wire alu_a_i_1_; 
wire alu_a_i_20_; 
wire alu_a_i_21_; 
wire alu_a_i_22_; 
wire alu_a_i_23_; 
wire alu_a_i_24_; 
wire alu_a_i_25_; 
wire alu_a_i_26_; 
wire alu_a_i_27_; 
wire alu_a_i_28_; 
wire alu_a_i_29_; 
wire alu_a_i_2_; 
wire alu_a_i_30_; 
wire alu_a_i_31_; 
wire alu_a_i_3_; 
wire alu_a_i_4_; 
wire alu_a_i_5_; 
wire alu_a_i_6_; 
wire alu_a_i_7_; 
wire alu_a_i_8_; 
wire alu_a_i_9_; 
wire alu_b_i_0_; 
wire alu_b_i_10_; 
wire alu_b_i_11_; 
wire alu_b_i_12_; 
wire alu_b_i_13_; 
wire alu_b_i_14_; 
wire alu_b_i_15_; 
wire alu_b_i_16_; 
wire alu_b_i_17_; 
wire alu_b_i_18_; 
wire alu_b_i_19_; 
wire alu_b_i_1_; 
wire alu_b_i_20_; 
wire alu_b_i_21_; 
wire alu_b_i_22_; 
wire alu_b_i_23_; 
wire alu_b_i_24_; 
wire alu_b_i_25_; 
wire alu_b_i_26_; 
wire alu_b_i_27_; 
wire alu_b_i_28_; 
wire alu_b_i_29_; 
wire alu_b_i_2_; 
wire alu_b_i_30_; 
wire alu_b_i_31_; 
wire alu_b_i_3_; 
wire alu_b_i_4_; 
wire alu_b_i_5_; 
wire alu_b_i_6_; 
wire alu_b_i_7_; 
wire alu_b_i_8_; 
wire alu_b_i_9_; 
wire alu_c_i; 
wire alu_c_o; 
wire alu_c_update_o; 
wire alu_equal_o; 
wire alu_flag_update_o; 
wire alu_func_r_0_; 
wire alu_func_r_1_; 
wire alu_func_r_2_; 
wire alu_func_r_3_; 
wire alu_greater_than_o; 
wire alu_greater_than_signed_o; 
wire alu_input_a_r_0_; 
wire alu_input_a_r_10_; 
wire alu_input_a_r_11_; 
wire alu_input_a_r_12_; 
wire alu_input_a_r_13_; 
wire alu_input_a_r_14_; 
wire alu_input_a_r_15_; 
wire alu_input_a_r_16_; 
wire alu_input_a_r_17_; 
wire alu_input_a_r_18_; 
wire alu_input_a_r_19_; 
wire alu_input_a_r_1_; 
wire alu_input_a_r_20_; 
wire alu_input_a_r_21_; 
wire alu_input_a_r_22_; 
wire alu_input_a_r_23_; 
wire alu_input_a_r_24_; 
wire alu_input_a_r_25_; 
wire alu_input_a_r_26_; 
wire alu_input_a_r_27_; 
wire alu_input_a_r_28_; 
wire alu_input_a_r_29_; 
wire alu_input_a_r_2_; 
wire alu_input_a_r_30_; 
wire alu_input_a_r_31_; 
wire alu_input_a_r_3_; 
wire alu_input_a_r_4_; 
wire alu_input_a_r_5_; 
wire alu_input_a_r_6_; 
wire alu_input_a_r_7_; 
wire alu_input_a_r_8_; 
wire alu_input_a_r_9_; 
wire alu_input_b_r_0_; 
wire alu_input_b_r_10_; 
wire alu_input_b_r_11_; 
wire alu_input_b_r_12_; 
wire alu_input_b_r_13_; 
wire alu_input_b_r_14_; 
wire alu_input_b_r_15_; 
wire alu_input_b_r_16_; 
wire alu_input_b_r_17_; 
wire alu_input_b_r_18_; 
wire alu_input_b_r_19_; 
wire alu_input_b_r_1_; 
wire alu_input_b_r_20_; 
wire alu_input_b_r_21_; 
wire alu_input_b_r_22_; 
wire alu_input_b_r_23_; 
wire alu_input_b_r_24_; 
wire alu_input_b_r_25_; 
wire alu_input_b_r_26_; 
wire alu_input_b_r_27_; 
wire alu_input_b_r_28_; 
wire alu_input_b_r_29_; 
wire alu_input_b_r_2_; 
wire alu_input_b_r_30_; 
wire alu_input_b_r_31_; 
wire alu_input_b_r_3_; 
wire alu_input_b_r_4_; 
wire alu_input_b_r_5_; 
wire alu_input_b_r_6_; 
wire alu_input_b_r_7_; 
wire alu_input_b_r_8_; 
wire alu_input_b_r_9_; 
wire alu_less_than_o; 
wire alu_less_than_signed_o; 
wire alu_op_i_0_; 
wire alu_op_i_1_; 
wire alu_op_i_2_; 
wire alu_op_i_3_; 
wire alu_op_r_0_; 
wire alu_op_r_1_; 
wire alu_op_r_2_; 
wire alu_op_r_3_; 
wire alu_op_r_4_; 
wire alu_op_r_5_; 
wire alu_op_r_6_; 
wire alu_op_r_7_; 
wire alu_p_o_0_; 
wire alu_p_o_10_; 
wire alu_p_o_11_; 
wire alu_p_o_12_; 
wire alu_p_o_13_; 
wire alu_p_o_14_; 
wire alu_p_o_15_; 
wire alu_p_o_16_; 
wire alu_p_o_17_; 
wire alu_p_o_18_; 
wire alu_p_o_19_; 
wire alu_p_o_1_; 
wire alu_p_o_20_; 
wire alu_p_o_21_; 
wire alu_p_o_22_; 
wire alu_p_o_23_; 
wire alu_p_o_24_; 
wire alu_p_o_25_; 
wire alu_p_o_26_; 
wire alu_p_o_27_; 
wire alu_p_o_28_; 
wire alu_p_o_29_; 
wire alu_p_o_2_; 
wire alu_p_o_30_; 
wire alu_p_o_31_; 
wire alu_p_o_3_; 
wire alu_p_o_4_; 
wire alu_p_o_5_; 
wire alu_p_o_6_; 
wire alu_p_o_7_; 
wire alu_p_o_8_; 
wire alu_p_o_9_; 
output break_o;
input clk_i;
input enable_i;
wire epc_q_0_; 
wire epc_q_10_; 
wire epc_q_11_; 
wire epc_q_12_; 
wire epc_q_13_; 
wire epc_q_14_; 
wire epc_q_15_; 
wire epc_q_16_; 
wire epc_q_17_; 
wire epc_q_18_; 
wire epc_q_19_; 
wire epc_q_1_; 
wire epc_q_20_; 
wire epc_q_21_; 
wire epc_q_22_; 
wire epc_q_23_; 
wire epc_q_24_; 
wire epc_q_25_; 
wire epc_q_26_; 
wire epc_q_27_; 
wire epc_q_28_; 
wire epc_q_29_; 
wire epc_q_2_; 
wire epc_q_30_; 
wire epc_q_31_; 
wire epc_q_3_; 
wire epc_q_4_; 
wire epc_q_5_; 
wire epc_q_6_; 
wire epc_q_7_; 
wire epc_q_8_; 
wire epc_q_9_; 
wire esr_q_10_; 
wire esr_q_2_; 
wire esr_q_9_; 
output fault_o;
wire inst_r_0_; 
wire inst_r_1_; 
wire inst_r_2_; 
wire inst_r_3_; 
wire inst_r_4_; 
wire inst_r_5_; 
wire inst_trap_w; 
wire int32_r_10_; 
wire int32_r_4_; 
wire int32_r_5_; 
input intr_i;
input mem_ack_i;
output \mem_addr_o[0] ;
output \mem_addr_o[10] ;
output \mem_addr_o[11] ;
output \mem_addr_o[12] ;
output \mem_addr_o[13] ;
output \mem_addr_o[14] ;
output \mem_addr_o[15] ;
output \mem_addr_o[16] ;
output \mem_addr_o[17] ;
output \mem_addr_o[18] ;
output \mem_addr_o[19] ;
output \mem_addr_o[1] ;
output \mem_addr_o[20] ;
output \mem_addr_o[21] ;
output \mem_addr_o[22] ;
output \mem_addr_o[23] ;
output \mem_addr_o[24] ;
output \mem_addr_o[25] ;
output \mem_addr_o[26] ;
output \mem_addr_o[27] ;
output \mem_addr_o[28] ;
output \mem_addr_o[29] ;
output \mem_addr_o[2] ;
output \mem_addr_o[30] ;
output \mem_addr_o[31] ;
output \mem_addr_o[3] ;
output \mem_addr_o[4] ;
output \mem_addr_o[5] ;
output \mem_addr_o[6] ;
output \mem_addr_o[7] ;
output \mem_addr_o[8] ;
output \mem_addr_o[9] ;
output \mem_cti_o[0] ;
output \mem_cti_o[1] ;
output \mem_cti_o[2] ;
output mem_cyc_o;
input \mem_dat_i[0] ;
input \mem_dat_i[10] ;
input \mem_dat_i[11] ;
input \mem_dat_i[12] ;
input \mem_dat_i[13] ;
input \mem_dat_i[14] ;
input \mem_dat_i[15] ;
input \mem_dat_i[16] ;
input \mem_dat_i[17] ;
input \mem_dat_i[18] ;
input \mem_dat_i[19] ;
input \mem_dat_i[1] ;
input \mem_dat_i[20] ;
input \mem_dat_i[21] ;
input \mem_dat_i[22] ;
input \mem_dat_i[23] ;
input \mem_dat_i[24] ;
input \mem_dat_i[25] ;
input \mem_dat_i[26] ;
input \mem_dat_i[27] ;
input \mem_dat_i[28] ;
input \mem_dat_i[29] ;
input \mem_dat_i[2] ;
input \mem_dat_i[30] ;
input \mem_dat_i[31] ;
input \mem_dat_i[3] ;
input \mem_dat_i[4] ;
input \mem_dat_i[5] ;
input \mem_dat_i[6] ;
input \mem_dat_i[7] ;
input \mem_dat_i[8] ;
input \mem_dat_i[9] ;
output \mem_dat_o[0] ;
output \mem_dat_o[10] ;
output \mem_dat_o[11] ;
output \mem_dat_o[12] ;
output \mem_dat_o[13] ;
output \mem_dat_o[14] ;
output \mem_dat_o[15] ;
output \mem_dat_o[16] ;
output \mem_dat_o[17] ;
output \mem_dat_o[18] ;
output \mem_dat_o[19] ;
output \mem_dat_o[1] ;
output \mem_dat_o[20] ;
output \mem_dat_o[21] ;
output \mem_dat_o[22] ;
output \mem_dat_o[23] ;
output \mem_dat_o[24] ;
output \mem_dat_o[25] ;
output \mem_dat_o[26] ;
output \mem_dat_o[27] ;
output \mem_dat_o[28] ;
output \mem_dat_o[29] ;
output \mem_dat_o[2] ;
output \mem_dat_o[30] ;
output \mem_dat_o[31] ;
output \mem_dat_o[3] ;
output \mem_dat_o[4] ;
output \mem_dat_o[5] ;
output \mem_dat_o[6] ;
output \mem_dat_o[7] ;
output \mem_dat_o[8] ;
output \mem_dat_o[9] ;
wire mem_offset_q_0_; 
wire mem_offset_q_1_; 
output \mem_sel_o[0] ;
output \mem_sel_o[1] ;
output \mem_sel_o[2] ;
output \mem_sel_o[3] ;
input mem_stall_i;
output mem_stb_o;
output mem_we_o;
wire next_pc_r_0_; 
wire next_pc_r_1_; 
input nmi_i;
wire nmi_q; 
wire opcode_q_21_; 
wire opcode_q_22_; 
wire opcode_q_23_; 
wire opcode_q_24_; 
wire opcode_q_25_; 
wire pc_q_10_; 
wire pc_q_11_; 
wire pc_q_12_; 
wire pc_q_13_; 
wire pc_q_14_; 
wire pc_q_15_; 
wire pc_q_16_; 
wire pc_q_17_; 
wire pc_q_18_; 
wire pc_q_19_; 
wire pc_q_20_; 
wire pc_q_21_; 
wire pc_q_22_; 
wire pc_q_23_; 
wire pc_q_24_; 
wire pc_q_25_; 
wire pc_q_26_; 
wire pc_q_27_; 
wire pc_q_28_; 
wire pc_q_29_; 
wire pc_q_2_; 
wire pc_q_30_; 
wire pc_q_31_; 
wire pc_q_3_; 
wire pc_q_4_; 
wire pc_q_5_; 
wire pc_q_6_; 
wire pc_q_7_; 
wire pc_q_8_; 
wire pc_q_9_; 
input rst_i;
wire sr_q_2_; 
wire sr_q_9_; 
wire state_q_0_; 
wire state_q_1_; 
wire state_q_2_; 
wire state_q_3_; 
wire state_q_4_; 
wire state_q_5_; 
AND2X2 AND2X2_1 ( .A(_abc_40298_new_n686_), .B(_abc_40298_new_n674_), .Y(_abc_40298_new_n688_));
AND2X2 AND2X2_10 ( .A(_abc_40298_new_n1096_), .B(_abc_40298_new_n942_), .Y(_abc_40298_new_n1097_));
AND2X2 AND2X2_100 ( .A(alu__abc_38674_new_n376_), .B(alu__abc_38674_new_n383_), .Y(alu__abc_38674_new_n1675_));
AND2X2 AND2X2_101 ( .A(alu__abc_38674_new_n1690_), .B(alu__abc_38674_new_n1679_), .Y(alu__abc_38674_new_n1691_));
AND2X2 AND2X2_11 ( .A(_abc_40298_new_n1061_), .B(_abc_40298_new_n1145_), .Y(_abc_40298_new_n1149_));
AND2X2 AND2X2_12 ( .A(_abc_40298_new_n1151_), .B(_abc_40298_new_n1148_), .Y(_abc_40298_new_n1152_));
AND2X2 AND2X2_13 ( .A(pc_q_2_), .B(pc_q_3_), .Y(_abc_40298_new_n1242_));
AND2X2 AND2X2_14 ( .A(_abc_40298_new_n1261_), .B(_abc_40298_new_n1264_), .Y(_abc_40298_new_n1265_));
AND2X2 AND2X2_15 ( .A(_abc_40298_new_n1305_), .B(_abc_40298_new_n1303_), .Y(_abc_40298_new_n1306_));
AND2X2 AND2X2_16 ( .A(_abc_40298_new_n1264_), .B(_abc_40298_new_n1281_), .Y(_abc_40298_new_n1310_));
AND2X2 AND2X2_17 ( .A(_abc_40298_new_n1373_), .B(_abc_40298_new_n1376_), .Y(_abc_40298_new_n1377_));
AND2X2 AND2X2_18 ( .A(_abc_40298_new_n1406_), .B(_abc_40298_new_n1175_), .Y(_abc_40298_new_n1407_));
AND2X2 AND2X2_19 ( .A(_abc_40298_new_n1433_), .B(_abc_40298_new_n1434_), .Y(_abc_40298_new_n1435_));
AND2X2 AND2X2_2 ( .A(_abc_40298_new_n904_), .B(_abc_40298_new_n893_), .Y(_abc_40298_new_n905_));
AND2X2 AND2X2_20 ( .A(_abc_40298_new_n1464_), .B(_abc_40298_new_n1175_), .Y(_abc_40298_new_n1465_));
AND2X2 AND2X2_21 ( .A(_abc_40298_new_n1474_), .B(_abc_40298_new_n1475_), .Y(_abc_40298_new_n1476_));
AND2X2 AND2X2_22 ( .A(_abc_40298_new_n1515_), .B(_abc_40298_new_n1493_), .Y(_abc_40298_new_n1516_));
AND2X2 AND2X2_23 ( .A(_abc_40298_new_n1565_), .B(_abc_40298_new_n1563_), .Y(_abc_40298_new_n1566_));
AND2X2 AND2X2_24 ( .A(_abc_40298_new_n1588_), .B(_abc_40298_new_n1589_), .Y(_abc_40298_new_n1590_));
AND2X2 AND2X2_25 ( .A(_abc_40298_new_n1546_), .B(_abc_40298_new_n1573_), .Y(_abc_40298_new_n1593_));
AND2X2 AND2X2_26 ( .A(_abc_40298_new_n1516_), .B(_abc_40298_new_n1593_), .Y(_abc_40298_new_n1594_));
AND2X2 AND2X2_27 ( .A(_abc_40298_new_n1484_), .B(_abc_40298_new_n1594_), .Y(_abc_40298_new_n1595_));
AND2X2 AND2X2_28 ( .A(_abc_40298_new_n1621_), .B(_abc_40298_new_n1622_), .Y(_abc_40298_new_n1623_));
AND2X2 AND2X2_29 ( .A(_abc_40298_new_n1681_), .B(_abc_40298_new_n1685_), .Y(_abc_40298_new_n1686_));
AND2X2 AND2X2_3 ( .A(_abc_40298_new_n927_), .B(_abc_40298_new_n922_), .Y(_abc_40298_new_n928_));
AND2X2 AND2X2_30 ( .A(_abc_40298_new_n1710_), .B(_abc_40298_new_n1714_), .Y(_abc_40298_new_n1715_));
AND2X2 AND2X2_31 ( .A(_abc_40298_new_n1728_), .B(_abc_40298_new_n1727_), .Y(_abc_40298_new_n1729_));
AND2X2 AND2X2_32 ( .A(_abc_40298_new_n1789_), .B(_abc_40298_new_n1793_), .Y(_abc_40298_new_n1794_));
AND2X2 AND2X2_33 ( .A(_abc_40298_new_n1820_), .B(_abc_40298_new_n1817_), .Y(_abc_40298_new_n1826_));
AND2X2 AND2X2_34 ( .A(_abc_40298_new_n1065_), .B(epc_q_25_), .Y(_abc_40298_new_n1850_));
AND2X2 AND2X2_35 ( .A(_abc_40298_new_n1865_), .B(_abc_40298_new_n1863_), .Y(_abc_40298_new_n1866_));
AND2X2 AND2X2_36 ( .A(_abc_40298_new_n1065_), .B(epc_q_26_), .Y(_abc_40298_new_n1881_));
AND2X2 AND2X2_37 ( .A(_abc_40298_new_n1912_), .B(_abc_40298_new_n1913_), .Y(_abc_40298_new_n1914_));
AND2X2 AND2X2_38 ( .A(_abc_40298_new_n1870_), .B(_abc_40298_new_n1918_), .Y(_abc_40298_new_n1919_));
AND2X2 AND2X2_39 ( .A(_abc_40298_new_n1925_), .B(_abc_40298_new_n1928_), .Y(_abc_40298_new_n1930_));
AND2X2 AND2X2_4 ( .A(_abc_40298_new_n941_), .B(_abc_40298_new_n950_), .Y(_abc_40298_new_n951_));
AND2X2 AND2X2_40 ( .A(_abc_40298_new_n1943_), .B(_abc_40298_new_n1945_), .Y(_abc_40298_new_n1946_));
AND2X2 AND2X2_41 ( .A(_abc_40298_new_n1964_), .B(_abc_40298_new_n1962_), .Y(_abc_40298_new_n1965_));
AND2X2 AND2X2_42 ( .A(_abc_40298_new_n1928_), .B(_abc_40298_new_n1944_), .Y(_abc_40298_new_n1968_));
AND2X2 AND2X2_43 ( .A(_abc_40298_new_n1065_), .B(epc_q_30_), .Y(_abc_40298_new_n1978_));
AND2X2 AND2X2_44 ( .A(_abc_40298_new_n1991_), .B(pc_q_31_), .Y(_abc_40298_new_n1992_));
AND2X2 AND2X2_45 ( .A(_abc_40298_new_n2003_), .B(_abc_40298_new_n2004_), .Y(_abc_40298_new_n2010_));
AND2X2 AND2X2_46 ( .A(_abc_40298_new_n2040_), .B(enable_i), .Y(_abc_40298_new_n2041_));
AND2X2 AND2X2_47 ( .A(_abc_40298_new_n2129_), .B(_abc_40298_new_n2120_), .Y(_abc_40298_new_n2130_));
AND2X2 AND2X2_48 ( .A(_abc_40298_new_n2150_), .B(_abc_40298_new_n2147_), .Y(_abc_40298_new_n2151_));
AND2X2 AND2X2_49 ( .A(_abc_40298_new_n2166_), .B(_abc_40298_new_n892_), .Y(_abc_40298_new_n2167_));
AND2X2 AND2X2_5 ( .A(_abc_40298_new_n937_), .B(_abc_40298_new_n967_), .Y(_abc_40298_new_n968_));
AND2X2 AND2X2_50 ( .A(_abc_40298_new_n2168_), .B(_abc_40298_new_n2170_), .Y(_abc_40298_new_n2171_));
AND2X2 AND2X2_51 ( .A(_abc_40298_new_n2148_), .B(_abc_40298_new_n2173_), .Y(_abc_40298_new_n2505_));
AND2X2 AND2X2_52 ( .A(_abc_40298_new_n932_), .B(_abc_40298_new_n2170_), .Y(_abc_40298_new_n2506_));
AND2X2 AND2X2_53 ( .A(_abc_40298_new_n2905_), .B(_abc_40298_new_n2903_), .Y(_abc_40298_new_n2907_));
AND2X2 AND2X2_54 ( .A(_abc_40298_new_n2952_), .B(_abc_40298_new_n2902_), .Y(_abc_40298_new_n2953_));
AND2X2 AND2X2_55 ( .A(_abc_40298_new_n2986_), .B(_abc_40298_new_n2989_), .Y(_abc_40298_new_n2990_));
AND2X2 AND2X2_56 ( .A(_abc_40298_new_n3085_), .B(_abc_40298_new_n3086_), .Y(_abc_40298_new_n3087_));
AND2X2 AND2X2_57 ( .A(_abc_40298_new_n3089_), .B(_abc_40298_new_n3092_), .Y(_abc_40298_new_n3093_));
AND2X2 AND2X2_58 ( .A(_abc_40298_new_n3128_), .B(_abc_40298_new_n3130_), .Y(_abc_40298_new_n3131_));
AND2X2 AND2X2_59 ( .A(_abc_40298_new_n3136_), .B(_abc_40298_new_n3138_), .Y(_abc_40298_new_n3139_));
AND2X2 AND2X2_6 ( .A(_abc_40298_new_n998_), .B(_abc_40298_new_n999_), .Y(_abc_40298_new_n1000_));
AND2X2 AND2X2_60 ( .A(_abc_40298_new_n1166_), .B(state_q_0_), .Y(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2382));
AND2X2 AND2X2_61 ( .A(alu_b_i_17_), .B(alu_a_i_17_), .Y(alu__abc_38674_new_n138_));
AND2X2 AND2X2_62 ( .A(alu_b_i_19_), .B(alu_a_i_19_), .Y(alu__abc_38674_new_n147_));
AND2X2 AND2X2_63 ( .A(alu_b_i_31_), .B(alu_a_i_31_), .Y(alu__abc_38674_new_n160_));
AND2X2 AND2X2_64 ( .A(alu_b_i_25_), .B(alu_a_i_25_), .Y(alu__abc_38674_new_n181_));
AND2X2 AND2X2_65 ( .A(alu_b_i_15_), .B(alu_a_i_15_), .Y(alu__abc_38674_new_n205_));
AND2X2 AND2X2_66 ( .A(alu_b_i_7_), .B(alu_a_i_7_), .Y(alu__abc_38674_new_n248_));
AND2X2 AND2X2_67 ( .A(alu_b_i_4_), .B(alu_a_i_4_), .Y(alu__abc_38674_new_n254_));
AND2X2 AND2X2_68 ( .A(alu_a_i_2_), .B(alu_b_i_2_), .Y(alu__abc_38674_new_n266_));
AND2X2 AND2X2_69 ( .A(alu_a_i_3_), .B(alu_b_i_3_), .Y(alu__abc_38674_new_n269_));
AND2X2 AND2X2_7 ( .A(_abc_40298_new_n1031_), .B(_abc_40298_new_n1032_), .Y(_abc_40298_new_n1033_));
AND2X2 AND2X2_70 ( .A(alu__abc_38674_new_n277_), .B(alu_op_i_3_), .Y(alu__abc_38674_new_n291_));
AND2X2 AND2X2_71 ( .A(alu__abc_38674_new_n241_), .B(alu__abc_38674_new_n354_), .Y(alu__abc_38674_new_n355_));
AND2X2 AND2X2_72 ( .A(alu_b_i_6_), .B(alu_a_i_6_), .Y(alu__abc_38674_new_n426_));
AND2X2 AND2X2_73 ( .A(alu_b_i_5_), .B(alu_a_i_5_), .Y(alu__abc_38674_new_n431_));
AND2X2 AND2X2_74 ( .A(alu__abc_38674_new_n447_), .B(alu__abc_38674_new_n237_), .Y(alu__abc_38674_new_n448_));
AND2X2 AND2X2_75 ( .A(alu__abc_38674_new_n514_), .B(alu__abc_38674_new_n448_), .Y(alu__abc_38674_new_n515_));
AND2X2 AND2X2_76 ( .A(alu__abc_38674_new_n534_), .B(alu__abc_38674_new_n528_), .Y(alu__abc_38674_new_n535_));
AND2X2 AND2X2_77 ( .A(alu__abc_38674_new_n421_), .B(alu__abc_38674_new_n268_), .Y(alu__abc_38674_new_n556_));
AND2X2 AND2X2_78 ( .A(alu__abc_38674_new_n587_), .B(alu__abc_38674_new_n593_), .Y(alu__abc_38674_new_n594_));
AND2X2 AND2X2_79 ( .A(alu__abc_38674_new_n613_), .B(alu__abc_38674_new_n614_), .Y(alu__abc_38674_new_n615_));
AND2X2 AND2X2_8 ( .A(_abc_40298_new_n1049_), .B(_abc_40298_new_n1050_), .Y(_abc_40298_new_n1051_));
AND2X2 AND2X2_80 ( .A(alu__abc_38674_new_n563_), .B(alu__abc_38674_new_n420_), .Y(alu__abc_38674_new_n692_));
AND2X2 AND2X2_81 ( .A(alu__abc_38674_new_n381_), .B(alu__abc_38674_new_n564_), .Y(alu__abc_38674_new_n693_));
AND2X2 AND2X2_82 ( .A(alu__abc_38674_new_n707_), .B(alu__abc_38674_new_n704_), .Y(alu__abc_38674_new_n708_));
AND2X2 AND2X2_83 ( .A(alu__abc_38674_new_n840_), .B(alu__abc_38674_new_n340_), .Y(alu__abc_38674_new_n841_));
AND2X2 AND2X2_84 ( .A(alu__abc_38674_new_n846_), .B(alu__abc_38674_new_n843_), .Y(alu__abc_38674_new_n847_));
AND2X2 AND2X2_85 ( .A(alu__abc_38674_new_n767_), .B(alu__abc_38674_new_n798_), .Y(alu__abc_38674_new_n851_));
AND2X2 AND2X2_86 ( .A(alu__abc_38674_new_n546_), .B(alu__abc_38674_new_n542_), .Y(alu__abc_38674_new_n979_));
AND2X2 AND2X2_87 ( .A(alu__abc_38674_new_n998_), .B(alu__abc_38674_new_n340_), .Y(alu__abc_38674_new_n999_));
AND2X2 AND2X2_88 ( .A(alu__abc_38674_new_n1100_), .B(alu__abc_38674_new_n230_), .Y(alu__abc_38674_new_n1101_));
AND2X2 AND2X2_89 ( .A(alu__abc_38674_new_n1106_), .B(alu__abc_38674_new_n1095_), .Y(alu__abc_38674_new_n1107_));
AND2X2 AND2X2_9 ( .A(_abc_40298_new_n1078_), .B(_abc_40298_new_n1076_), .Y(_abc_40298_new_n1079_));
AND2X2 AND2X2_90 ( .A(alu__abc_38674_new_n1121_), .B(alu__abc_38674_new_n1132_), .Y(alu__abc_38674_new_n1133_));
AND2X2 AND2X2_91 ( .A(alu__abc_38674_new_n949_), .B(alu__abc_38674_new_n340_), .Y(alu__abc_38674_new_n1212_));
AND2X2 AND2X2_92 ( .A(alu__abc_38674_new_n944_), .B(alu_b_i_3_), .Y(alu__abc_38674_new_n1213_));
AND2X2 AND2X2_93 ( .A(alu__abc_38674_new_n844_), .B(alu__abc_38674_new_n218_), .Y(alu__abc_38674_new_n1226_));
AND2X2 AND2X2_94 ( .A(alu__abc_38674_new_n1446_), .B(alu__abc_38674_new_n496_), .Y(alu__abc_38674_new_n1470_));
AND2X2 AND2X2_95 ( .A(alu__abc_38674_new_n1487_), .B(alu__abc_38674_new_n115_), .Y(alu__abc_38674_new_n1488_));
AND2X2 AND2X2_96 ( .A(alu__abc_38674_new_n1503_), .B(alu__abc_38674_new_n321_), .Y(alu__abc_38674_new_n1504_));
AND2X2 AND2X2_97 ( .A(alu__abc_38674_new_n1579_), .B(alu__abc_38674_new_n191_), .Y(alu__abc_38674_new_n1580_));
AND2X2 AND2X2_98 ( .A(alu__abc_38674_new_n1604_), .B(alu__abc_38674_new_n395_), .Y(alu__abc_38674_new_n1605_));
AND2X2 AND2X2_99 ( .A(alu__abc_38674_new_n1644_), .B(alu__abc_38674_new_n1632_), .Y(alu__abc_38674_new_n1645_));
AOI21X1 AOI21X1_1 ( .A(_abc_40298_new_n689_), .B(_abc_40298_new_n655_), .C(_abc_40298_new_n631_), .Y(_abc_40298_new_n690_));
AOI21X1 AOI21X1_10 ( .A(_abc_40298_new_n750_), .B(_abc_40298_new_n751_), .C(_abc_40298_new_n655_), .Y(_abc_40298_new_n752_));
AOI21X1 AOI21X1_100 ( .A(_abc_40298_new_n1706_), .B(_abc_40298_new_n1813_), .C(_abc_40298_new_n1816_), .Y(_abc_40298_new_n1817_));
AOI21X1 AOI21X1_101 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1836_), .C(_abc_40298_new_n1071_), .Y(_abc_40298_new_n1837_));
AOI21X1 AOI21X1_102 ( .A(_abc_40298_new_n1838_), .B(_abc_40298_new_n1810_), .C(_abc_40298_new_n1839_), .Y(_0epc_q_31_0__24_));
AOI21X1 AOI21X1_103 ( .A(_abc_40298_new_n1853_), .B(_abc_40298_new_n1176_), .C(_abc_40298_new_n1232_), .Y(_abc_40298_new_n1854_));
AOI21X1 AOI21X1_104 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1857_), .C(_abc_40298_new_n1071_), .Y(_abc_40298_new_n1858_));
AOI21X1 AOI21X1_105 ( .A(_abc_40298_new_n1859_), .B(_abc_40298_new_n1842_), .C(_abc_40298_new_n1860_), .Y(_0epc_q_31_0__25_));
AOI21X1 AOI21X1_106 ( .A(_abc_40298_new_n1821_), .B(_abc_40298_new_n1870_), .C(_abc_40298_new_n1873_), .Y(_abc_40298_new_n1874_));
AOI21X1 AOI21X1_107 ( .A(_abc_40298_new_n1874_), .B(_abc_40298_new_n1878_), .C(_abc_40298_new_n1879_), .Y(_abc_40298_new_n1880_));
AOI21X1 AOI21X1_108 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1886_), .C(_abc_40298_new_n1071_), .Y(_abc_40298_new_n1887_));
AOI21X1 AOI21X1_109 ( .A(_abc_40298_new_n1888_), .B(_abc_40298_new_n1867_), .C(_abc_40298_new_n1889_), .Y(_0epc_q_31_0__26_));
AOI21X1 AOI21X1_11 ( .A(_abc_40298_new_n749_), .B(_abc_40298_new_n655_), .C(_abc_40298_new_n752_), .Y(_abc_40298_new_n753_));
AOI21X1 AOI21X1_110 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1906_), .C(_abc_40298_new_n1071_), .Y(_abc_40298_new_n1907_));
AOI21X1 AOI21X1_111 ( .A(_abc_40298_new_n1908_), .B(_abc_40298_new_n1893_), .C(_abc_40298_new_n1909_), .Y(_0epc_q_31_0__27_));
AOI21X1 AOI21X1_112 ( .A(_abc_40298_new_n1820_), .B(_abc_40298_new_n1817_), .C(_abc_40298_new_n1920_), .Y(_abc_40298_new_n1921_));
AOI21X1 AOI21X1_113 ( .A(_abc_40298_new_n1897_), .B(_abc_40298_new_n1876_), .C(_abc_40298_new_n1896_), .Y(_abc_40298_new_n1923_));
AOI21X1 AOI21X1_114 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1936_), .C(_abc_40298_new_n1071_), .Y(_abc_40298_new_n1937_));
AOI21X1 AOI21X1_115 ( .A(_abc_40298_new_n1938_), .B(_abc_40298_new_n1915_), .C(_abc_40298_new_n1939_), .Y(_0epc_q_31_0__28_));
AOI21X1 AOI21X1_116 ( .A(_abc_40298_new_n1065_), .B(epc_q_29_), .C(_abc_40298_new_n1176_), .Y(_abc_40298_new_n1948_));
AOI21X1 AOI21X1_117 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1955_), .C(_abc_40298_new_n1071_), .Y(_abc_40298_new_n1956_));
AOI21X1 AOI21X1_118 ( .A(_abc_40298_new_n1957_), .B(_abc_40298_new_n1942_), .C(_abc_40298_new_n1958_), .Y(_0epc_q_31_0__29_));
AOI21X1 AOI21X1_119 ( .A(_abc_40298_new_n1971_), .B(_abc_40298_new_n1975_), .C(_abc_40298_new_n1976_), .Y(_abc_40298_new_n1977_));
AOI21X1 AOI21X1_12 ( .A(_abc_40298_new_n686_), .B(_abc_40298_new_n675_), .C(_abc_40298_new_n654_), .Y(_abc_40298_new_n764_));
AOI21X1 AOI21X1_120 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1984_), .C(_abc_40298_new_n1071_), .Y(_abc_40298_new_n1985_));
AOI21X1 AOI21X1_121 ( .A(_abc_40298_new_n1986_), .B(_abc_40298_new_n1966_), .C(_abc_40298_new_n1987_), .Y(_0epc_q_31_0__30_));
AOI21X1 AOI21X1_122 ( .A(_abc_40298_new_n1065_), .B(epc_q_31_), .C(_abc_40298_new_n1176_), .Y(_abc_40298_new_n1994_));
AOI21X1 AOI21X1_123 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n2007_), .C(_abc_40298_new_n1071_), .Y(_abc_40298_new_n2008_));
AOI21X1 AOI21X1_124 ( .A(_abc_40298_new_n2010_), .B(_abc_40298_new_n1071_), .C(_abc_40298_new_n1138_), .Y(_abc_40298_new_n2011_));
AOI21X1 AOI21X1_125 ( .A(_abc_40298_new_n2009_), .B(_abc_40298_new_n2011_), .C(_abc_40298_new_n2012_), .Y(_0epc_q_31_0__31_));
AOI21X1 AOI21X1_126 ( .A(_abc_40298_new_n2015_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n2016_), .Y(_0pc_q_31_0__0_));
AOI21X1 AOI21X1_127 ( .A(_abc_40298_new_n2018_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n2019_), .Y(_0pc_q_31_0__1_));
AOI21X1 AOI21X1_128 ( .A(_abc_40298_new_n2021_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n2022_), .Y(_0pc_q_31_0__2_));
AOI21X1 AOI21X1_129 ( .A(_abc_40298_new_n2028_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n2029_), .Y(_0pc_q_31_0__4_));
AOI21X1 AOI21X1_13 ( .A(_abc_40298_new_n766_), .B(_abc_40298_new_n757_), .C(_abc_40298_new_n631_), .Y(_abc_40298_new_n767_));
AOI21X1 AOI21X1_130 ( .A(_abc_40298_new_n2034_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n2035_), .Y(_0pc_q_31_0__6_));
AOI21X1 AOI21X1_131 ( .A(_abc_40298_new_n1409_), .B(_abc_40298_new_n1168_), .C(_abc_40298_new_n888_), .Y(_abc_40298_new_n2044_));
AOI21X1 AOI21X1_132 ( .A(_abc_40298_new_n1024_), .B(_abc_40298_new_n954_), .C(_abc_40298_new_n1138_), .Y(_abc_40298_new_n2046_));
AOI21X1 AOI21X1_133 ( .A(_abc_40298_new_n2045_), .B(_abc_40298_new_n2046_), .C(_abc_40298_new_n2047_), .Y(_0pc_q_31_0__9_));
AOI21X1 AOI21X1_134 ( .A(_abc_40298_new_n2055_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n2056_), .Y(_0pc_q_31_0__11_));
AOI21X1 AOI21X1_135 ( .A(_abc_40298_new_n2061_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n2062_), .Y(_0pc_q_31_0__13_));
AOI21X1 AOI21X1_136 ( .A(_abc_40298_new_n2064_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n2065_), .Y(_0pc_q_31_0__14_));
AOI21X1 AOI21X1_137 ( .A(_abc_40298_new_n2067_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n2068_), .Y(_0pc_q_31_0__15_));
AOI21X1 AOI21X1_138 ( .A(_abc_40298_new_n2073_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n2074_), .Y(_0pc_q_31_0__17_));
AOI21X1 AOI21X1_139 ( .A(_abc_40298_new_n2076_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n2077_), .Y(_0pc_q_31_0__18_));
AOI21X1 AOI21X1_14 ( .A(_abc_40298_new_n686_), .B(_abc_40298_new_n729_), .C(_abc_40298_new_n654_), .Y(_abc_40298_new_n786_));
AOI21X1 AOI21X1_140 ( .A(_abc_40298_new_n2079_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n2080_), .Y(_0pc_q_31_0__19_));
AOI21X1 AOI21X1_141 ( .A(_abc_40298_new_n2082_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n2083_), .Y(_0pc_q_31_0__20_));
AOI21X1 AOI21X1_142 ( .A(_abc_40298_new_n2085_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n2086_), .Y(_0pc_q_31_0__21_));
AOI21X1 AOI21X1_143 ( .A(_abc_40298_new_n2088_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n2089_), .Y(_0pc_q_31_0__22_));
AOI21X1 AOI21X1_144 ( .A(_abc_40298_new_n2091_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n2092_), .Y(_0pc_q_31_0__23_));
AOI21X1 AOI21X1_145 ( .A(_abc_40298_new_n2103_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n2104_), .Y(_0pc_q_31_0__27_));
AOI21X1 AOI21X1_146 ( .A(_abc_40298_new_n2106_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n2107_), .Y(_0pc_q_31_0__28_));
AOI21X1 AOI21X1_147 ( .A(_abc_40298_new_n2109_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n2110_), .Y(_0pc_q_31_0__29_));
AOI21X1 AOI21X1_148 ( .A(_abc_40298_new_n2112_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n2113_), .Y(_0pc_q_31_0__30_));
AOI21X1 AOI21X1_149 ( .A(_abc_40298_new_n2116_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n2117_), .Y(_0pc_q_31_0__31_));
AOI21X1 AOI21X1_15 ( .A(_abc_40298_new_n686_), .B(_abc_40298_new_n738_), .C(_abc_40298_new_n654_), .Y(_abc_40298_new_n790_));
AOI21X1 AOI21X1_150 ( .A(_abc_40298_new_n1001_), .B(_abc_40298_new_n2121_), .C(_abc_40298_new_n2128_), .Y(_abc_40298_new_n2129_));
AOI21X1 AOI21X1_151 ( .A(_abc_40298_new_n2142_), .B(_abc_40298_new_n973_), .C(_abc_40298_new_n1015_), .Y(_abc_40298_new_n2143_));
AOI21X1 AOI21X1_152 ( .A(_abc_40298_new_n959_), .B(REGFILE_SIM_reg_bank_rb_i_4_), .C(_abc_40298_new_n931_), .Y(_abc_40298_new_n2197_));
AOI21X1 AOI21X1_153 ( .A(_abc_40298_new_n2196_), .B(_abc_40298_new_n931_), .C(_abc_40298_new_n2197_), .Y(_abc_40298_new_n2198_));
AOI21X1 AOI21X1_154 ( .A(_abc_40298_new_n2159_), .B(_abc_40298_new_n1628_), .C(_abc_40298_new_n2175_), .Y(_abc_40298_new_n2199_));
AOI21X1 AOI21X1_155 ( .A(_abc_40298_new_n2207_), .B(_abc_40298_new_n2204_), .C(_abc_40298_new_n2203_), .Y(_abc_40298_new_n2208_));
AOI21X1 AOI21X1_156 ( .A(_abc_40298_new_n2212_), .B(_abc_40298_new_n2204_), .C(_abc_40298_new_n2203_), .Y(_abc_40298_new_n2213_));
AOI21X1 AOI21X1_157 ( .A(_abc_40298_new_n2217_), .B(_abc_40298_new_n2204_), .C(_abc_40298_new_n2203_), .Y(_abc_40298_new_n2218_));
AOI21X1 AOI21X1_158 ( .A(_abc_40298_new_n2222_), .B(_abc_40298_new_n2204_), .C(_abc_40298_new_n2203_), .Y(_abc_40298_new_n2223_));
AOI21X1 AOI21X1_159 ( .A(_abc_40298_new_n2227_), .B(_abc_40298_new_n2204_), .C(_abc_40298_new_n2203_), .Y(_abc_40298_new_n2228_));
AOI21X1 AOI21X1_16 ( .A(_abc_40298_new_n686_), .B(_abc_40298_new_n755_), .C(_abc_40298_new_n654_), .Y(_abc_40298_new_n800_));
AOI21X1 AOI21X1_160 ( .A(_abc_40298_new_n2232_), .B(_abc_40298_new_n2204_), .C(_abc_40298_new_n2203_), .Y(_abc_40298_new_n2233_));
AOI21X1 AOI21X1_161 ( .A(_abc_40298_new_n2237_), .B(_abc_40298_new_n2204_), .C(_abc_40298_new_n2203_), .Y(_abc_40298_new_n2238_));
AOI21X1 AOI21X1_162 ( .A(_abc_40298_new_n2242_), .B(_abc_40298_new_n2204_), .C(_abc_40298_new_n2203_), .Y(_abc_40298_new_n2243_));
AOI21X1 AOI21X1_163 ( .A(_abc_40298_new_n2247_), .B(_abc_40298_new_n2204_), .C(_abc_40298_new_n2203_), .Y(_abc_40298_new_n2248_));
AOI21X1 AOI21X1_164 ( .A(_abc_40298_new_n2251_), .B(_abc_40298_new_n2204_), .C(_abc_40298_new_n2203_), .Y(_abc_40298_new_n2252_));
AOI21X1 AOI21X1_165 ( .A(_abc_40298_new_n2255_), .B(_abc_40298_new_n2204_), .C(_abc_40298_new_n2203_), .Y(_abc_40298_new_n2256_));
AOI21X1 AOI21X1_166 ( .A(_abc_40298_new_n2259_), .B(_abc_40298_new_n2204_), .C(_abc_40298_new_n2203_), .Y(_abc_40298_new_n2260_));
AOI21X1 AOI21X1_167 ( .A(_abc_40298_new_n2264_), .B(_abc_40298_new_n2204_), .C(_abc_40298_new_n2203_), .Y(_abc_40298_new_n2265_));
AOI21X1 AOI21X1_168 ( .A(_abc_40298_new_n2269_), .B(_abc_40298_new_n2204_), .C(_abc_40298_new_n2203_), .Y(_abc_40298_new_n2270_));
AOI21X1 AOI21X1_169 ( .A(_abc_40298_new_n2273_), .B(_abc_40298_new_n2204_), .C(_abc_40298_new_n2203_), .Y(_abc_40298_new_n2274_));
AOI21X1 AOI21X1_17 ( .A(_abc_40298_new_n918_), .B(_abc_40298_new_n955_), .C(_abc_40298_new_n961_), .Y(_abc_40298_new_n962_));
AOI21X1 AOI21X1_170 ( .A(_abc_40298_new_n2277_), .B(_abc_40298_new_n2204_), .C(_abc_40298_new_n2203_), .Y(_abc_40298_new_n2278_));
AOI21X1 AOI21X1_171 ( .A(_abc_40298_new_n2301_), .B(_abc_40298_new_n1001_), .C(_abc_40298_new_n2303_), .Y(_abc_40298_new_n2304_));
AOI21X1 AOI21X1_172 ( .A(_abc_40298_new_n2286_), .B(REGFILE_SIM_reg_bank_reg_ra_o_5_), .C(_abc_40298_new_n1001_), .Y(_abc_40298_new_n2322_));
AOI21X1 AOI21X1_173 ( .A(_abc_40298_new_n1186_), .B(epc_q_5_), .C(_abc_40298_new_n1002_), .Y(_abc_40298_new_n2323_));
AOI21X1 AOI21X1_174 ( .A(_abc_40298_new_n1081_), .B(esr_q_9_), .C(_abc_40298_new_n1002_), .Y(_abc_40298_new_n2349_));
AOI21X1 AOI21X1_175 ( .A(_abc_40298_new_n1132_), .B(_abc_40298_new_n1124_), .C(_abc_40298_new_n1061_), .Y(_abc_40298_new_n2351_));
AOI21X1 AOI21X1_176 ( .A(_abc_40298_new_n1152_), .B(_abc_40298_new_n1060_), .C(_abc_40298_new_n2359_), .Y(_abc_40298_new_n2360_));
AOI21X1 AOI21X1_177 ( .A(_abc_40298_new_n1012_), .B(_abc_40298_new_n1419_), .C(_abc_40298_new_n2361_), .Y(_abc_40298_new_n2362_));
AOI21X1 AOI21X1_178 ( .A(_abc_40298_new_n1186_), .B(epc_q_11_), .C(_abc_40298_new_n1002_), .Y(_abc_40298_new_n2364_));
AOI21X1 AOI21X1_179 ( .A(_abc_40298_new_n2286_), .B(REGFILE_SIM_reg_bank_reg_ra_o_11_), .C(_abc_40298_new_n1001_), .Y(_abc_40298_new_n2365_));
AOI21X1 AOI21X1_18 ( .A(_abc_40298_new_n933_), .B(_abc_40298_new_n1008_), .C(_abc_40298_new_n1017_), .Y(_abc_40298_new_n1018_));
AOI21X1 AOI21X1_180 ( .A(_abc_40298_new_n1012_), .B(_abc_40298_new_n1509_), .C(_abc_40298_new_n2374_), .Y(_abc_40298_new_n2375_));
AOI21X1 AOI21X1_181 ( .A(_abc_40298_new_n1537_), .B(_abc_40298_new_n1012_), .C(_abc_40298_new_n2378_), .Y(_abc_40298_new_n2379_));
AOI21X1 AOI21X1_182 ( .A(_abc_40298_new_n897_), .B(_abc_40298_new_n976_), .C(_abc_40298_new_n2500_), .Y(_abc_40298_new_n2501_));
AOI21X1 AOI21X1_183 ( .A(_abc_40298_new_n905_), .B(_abc_40298_new_n907_), .C(_abc_40298_new_n961_), .Y(_abc_40298_new_n2503_));
AOI21X1 AOI21X1_184 ( .A(_abc_40298_new_n907_), .B(_abc_40298_new_n926_), .C(_abc_40298_new_n1015_), .Y(_abc_40298_new_n2511_));
AOI21X1 AOI21X1_185 ( .A(_abc_40298_new_n855_), .B(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2420), .C(_abc_40298_new_n2559_), .Y(_0opcode_q_31_0__26_));
AOI21X1 AOI21X1_186 ( .A(_abc_40298_new_n865_), .B(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2420), .C(_abc_40298_new_n2562_), .Y(_0opcode_q_31_0__28_));
AOI21X1 AOI21X1_187 ( .A(_abc_40298_new_n2571_), .B(_abc_40298_new_n2516_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2589_));
AOI21X1 AOI21X1_188 ( .A(\mem_dat_o[0] ), .B(_abc_40298_new_n2515_), .C(_abc_40298_new_n2608_), .Y(_abc_40298_new_n2609_));
AOI21X1 AOI21X1_189 ( .A(_abc_40298_new_n2614_), .B(_abc_40298_new_n2608_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2615_));
AOI21X1 AOI21X1_19 ( .A(_abc_40298_new_n1066_), .B(sr_q_2_), .C(_abc_40298_new_n993_), .Y(_abc_40298_new_n1067_));
AOI21X1 AOI21X1_190 ( .A(\mem_dat_o[1] ), .B(_abc_40298_new_n2515_), .C(_abc_40298_new_n2608_), .Y(_abc_40298_new_n2619_));
AOI21X1 AOI21X1_191 ( .A(_abc_40298_new_n2622_), .B(_abc_40298_new_n2608_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2623_));
AOI21X1 AOI21X1_192 ( .A(\mem_dat_o[2] ), .B(_abc_40298_new_n2515_), .C(_abc_40298_new_n2608_), .Y(_abc_40298_new_n2627_));
AOI21X1 AOI21X1_193 ( .A(_abc_40298_new_n2630_), .B(_abc_40298_new_n2608_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2631_));
AOI21X1 AOI21X1_194 ( .A(\mem_dat_o[3] ), .B(_abc_40298_new_n2515_), .C(_abc_40298_new_n2608_), .Y(_abc_40298_new_n2635_));
AOI21X1 AOI21X1_195 ( .A(_abc_40298_new_n2638_), .B(_abc_40298_new_n2608_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2639_));
AOI21X1 AOI21X1_196 ( .A(\mem_dat_o[4] ), .B(_abc_40298_new_n2515_), .C(_abc_40298_new_n2608_), .Y(_abc_40298_new_n2643_));
AOI21X1 AOI21X1_197 ( .A(_abc_40298_new_n2646_), .B(_abc_40298_new_n2608_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2647_));
AOI21X1 AOI21X1_198 ( .A(\mem_dat_o[5] ), .B(_abc_40298_new_n2515_), .C(_abc_40298_new_n2608_), .Y(_abc_40298_new_n2651_));
AOI21X1 AOI21X1_199 ( .A(_abc_40298_new_n2654_), .B(_abc_40298_new_n2608_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2655_));
AOI21X1 AOI21X1_2 ( .A(_abc_40298_new_n698_), .B(_abc_40298_new_n702_), .C(_abc_40298_new_n655_), .Y(_abc_40298_new_n703_));
AOI21X1 AOI21X1_20 ( .A(_abc_40298_new_n1086_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n1087_), .Y(_0esr_q_31_0__2_));
AOI21X1 AOI21X1_200 ( .A(\mem_dat_o[6] ), .B(_abc_40298_new_n2515_), .C(_abc_40298_new_n2608_), .Y(_abc_40298_new_n2659_));
AOI21X1 AOI21X1_201 ( .A(_abc_40298_new_n2662_), .B(_abc_40298_new_n2608_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2663_));
AOI21X1 AOI21X1_202 ( .A(\mem_dat_o[7] ), .B(_abc_40298_new_n2515_), .C(_abc_40298_new_n2608_), .Y(_abc_40298_new_n2667_));
AOI21X1 AOI21X1_203 ( .A(_abc_40298_new_n2670_), .B(_abc_40298_new_n2608_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2671_));
AOI21X1 AOI21X1_204 ( .A(\mem_dat_o[8] ), .B(_abc_40298_new_n2515_), .C(_abc_40298_new_n2608_), .Y(_abc_40298_new_n2677_));
AOI21X1 AOI21X1_205 ( .A(_abc_40298_new_n2678_), .B(_abc_40298_new_n2676_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2679_));
AOI21X1 AOI21X1_206 ( .A(\mem_dat_o[9] ), .B(_abc_40298_new_n2515_), .C(_abc_40298_new_n2608_), .Y(_abc_40298_new_n2686_));
AOI21X1 AOI21X1_207 ( .A(_abc_40298_new_n2687_), .B(_abc_40298_new_n2685_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2688_));
AOI21X1 AOI21X1_208 ( .A(\mem_dat_o[10] ), .B(_abc_40298_new_n2515_), .C(_abc_40298_new_n2608_), .Y(_abc_40298_new_n2695_));
AOI21X1 AOI21X1_209 ( .A(_abc_40298_new_n2696_), .B(_abc_40298_new_n2694_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2697_));
AOI21X1 AOI21X1_21 ( .A(_abc_40298_new_n1094_), .B(_abc_40298_new_n1097_), .C(_abc_40298_new_n1099_), .Y(_abc_40298_new_n1100_));
AOI21X1 AOI21X1_210 ( .A(\mem_dat_o[11] ), .B(_abc_40298_new_n2515_), .C(_abc_40298_new_n2608_), .Y(_abc_40298_new_n2704_));
AOI21X1 AOI21X1_211 ( .A(_abc_40298_new_n2705_), .B(_abc_40298_new_n2703_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2706_));
AOI21X1 AOI21X1_212 ( .A(\mem_dat_o[12] ), .B(_abc_40298_new_n2515_), .C(_abc_40298_new_n2608_), .Y(_abc_40298_new_n2713_));
AOI21X1 AOI21X1_213 ( .A(_abc_40298_new_n2714_), .B(_abc_40298_new_n2712_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2715_));
AOI21X1 AOI21X1_214 ( .A(\mem_dat_o[13] ), .B(_abc_40298_new_n2515_), .C(_abc_40298_new_n2608_), .Y(_abc_40298_new_n2722_));
AOI21X1 AOI21X1_215 ( .A(_abc_40298_new_n2723_), .B(_abc_40298_new_n2721_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2724_));
AOI21X1 AOI21X1_216 ( .A(\mem_dat_o[14] ), .B(_abc_40298_new_n2515_), .C(_abc_40298_new_n2608_), .Y(_abc_40298_new_n2731_));
AOI21X1 AOI21X1_217 ( .A(_abc_40298_new_n2732_), .B(_abc_40298_new_n2730_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2733_));
AOI21X1 AOI21X1_218 ( .A(\mem_dat_o[15] ), .B(_abc_40298_new_n2515_), .C(_abc_40298_new_n2608_), .Y(_abc_40298_new_n2740_));
AOI21X1 AOI21X1_219 ( .A(_abc_40298_new_n2741_), .B(_abc_40298_new_n2739_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2742_));
AOI21X1 AOI21X1_22 ( .A(_abc_40298_new_n1110_), .B(_abc_40298_new_n1111_), .C(_abc_40298_new_n1116_), .Y(_abc_40298_new_n1117_));
AOI21X1 AOI21X1_220 ( .A(\mem_dat_o[16] ), .B(_abc_40298_new_n2515_), .C(_abc_40298_new_n2608_), .Y(_abc_40298_new_n2747_));
AOI21X1 AOI21X1_221 ( .A(_abc_40298_new_n2750_), .B(_abc_40298_new_n2608_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2751_));
AOI21X1 AOI21X1_222 ( .A(\mem_dat_o[17] ), .B(_abc_40298_new_n2515_), .C(_abc_40298_new_n2608_), .Y(_abc_40298_new_n2755_));
AOI21X1 AOI21X1_223 ( .A(_abc_40298_new_n2758_), .B(_abc_40298_new_n2608_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2759_));
AOI21X1 AOI21X1_224 ( .A(\mem_dat_o[18] ), .B(_abc_40298_new_n2515_), .C(_abc_40298_new_n2608_), .Y(_abc_40298_new_n2763_));
AOI21X1 AOI21X1_225 ( .A(_abc_40298_new_n2766_), .B(_abc_40298_new_n2608_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2767_));
AOI21X1 AOI21X1_226 ( .A(\mem_dat_o[19] ), .B(_abc_40298_new_n2515_), .C(_abc_40298_new_n2608_), .Y(_abc_40298_new_n2771_));
AOI21X1 AOI21X1_227 ( .A(_abc_40298_new_n2774_), .B(_abc_40298_new_n2608_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2775_));
AOI21X1 AOI21X1_228 ( .A(\mem_dat_o[20] ), .B(_abc_40298_new_n2515_), .C(_abc_40298_new_n2608_), .Y(_abc_40298_new_n2779_));
AOI21X1 AOI21X1_229 ( .A(_abc_40298_new_n2782_), .B(_abc_40298_new_n2608_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2783_));
AOI21X1 AOI21X1_23 ( .A(_abc_40298_new_n1092_), .B(_abc_40298_new_n1118_), .C(_abc_40298_new_n1112_), .Y(_abc_40298_new_n1119_));
AOI21X1 AOI21X1_230 ( .A(\mem_dat_o[21] ), .B(_abc_40298_new_n2515_), .C(_abc_40298_new_n2608_), .Y(_abc_40298_new_n2787_));
AOI21X1 AOI21X1_231 ( .A(_abc_40298_new_n2790_), .B(_abc_40298_new_n2608_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2791_));
AOI21X1 AOI21X1_232 ( .A(\mem_dat_o[22] ), .B(_abc_40298_new_n2515_), .C(_abc_40298_new_n2608_), .Y(_abc_40298_new_n2795_));
AOI21X1 AOI21X1_233 ( .A(_abc_40298_new_n2798_), .B(_abc_40298_new_n2608_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2799_));
AOI21X1 AOI21X1_234 ( .A(\mem_dat_o[23] ), .B(_abc_40298_new_n2515_), .C(_abc_40298_new_n2608_), .Y(_abc_40298_new_n2803_));
AOI21X1 AOI21X1_235 ( .A(_abc_40298_new_n2806_), .B(_abc_40298_new_n2608_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2807_));
AOI21X1 AOI21X1_236 ( .A(\mem_dat_o[24] ), .B(_abc_40298_new_n2515_), .C(_abc_40298_new_n2608_), .Y(_abc_40298_new_n2813_));
AOI21X1 AOI21X1_237 ( .A(_abc_40298_new_n2814_), .B(_abc_40298_new_n2812_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2815_));
AOI21X1 AOI21X1_238 ( .A(\mem_dat_o[25] ), .B(_abc_40298_new_n2515_), .C(_abc_40298_new_n2608_), .Y(_abc_40298_new_n2822_));
AOI21X1 AOI21X1_239 ( .A(_abc_40298_new_n2823_), .B(_abc_40298_new_n2821_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2824_));
AOI21X1 AOI21X1_24 ( .A(_abc_40298_new_n1120_), .B(_abc_40298_new_n1126_), .C(_abc_40298_new_n933_), .Y(_abc_40298_new_n1127_));
AOI21X1 AOI21X1_240 ( .A(\mem_dat_o[26] ), .B(_abc_40298_new_n2515_), .C(_abc_40298_new_n2608_), .Y(_abc_40298_new_n2831_));
AOI21X1 AOI21X1_241 ( .A(_abc_40298_new_n2832_), .B(_abc_40298_new_n2830_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2833_));
AOI21X1 AOI21X1_242 ( .A(\mem_dat_o[27] ), .B(_abc_40298_new_n2515_), .C(_abc_40298_new_n2608_), .Y(_abc_40298_new_n2840_));
AOI21X1 AOI21X1_243 ( .A(_abc_40298_new_n2841_), .B(_abc_40298_new_n2839_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2842_));
AOI21X1 AOI21X1_244 ( .A(\mem_dat_o[28] ), .B(_abc_40298_new_n2515_), .C(_abc_40298_new_n2608_), .Y(_abc_40298_new_n2849_));
AOI21X1 AOI21X1_245 ( .A(_abc_40298_new_n2850_), .B(_abc_40298_new_n2848_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2851_));
AOI21X1 AOI21X1_246 ( .A(\mem_dat_o[29] ), .B(_abc_40298_new_n2515_), .C(_abc_40298_new_n2608_), .Y(_abc_40298_new_n2858_));
AOI21X1 AOI21X1_247 ( .A(_abc_40298_new_n2859_), .B(_abc_40298_new_n2857_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2860_));
AOI21X1 AOI21X1_248 ( .A(\mem_dat_o[30] ), .B(_abc_40298_new_n2515_), .C(_abc_40298_new_n2608_), .Y(_abc_40298_new_n2867_));
AOI21X1 AOI21X1_249 ( .A(_abc_40298_new_n2868_), .B(_abc_40298_new_n2866_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2869_));
AOI21X1 AOI21X1_25 ( .A(_abc_40298_new_n1135_), .B(_abc_40298_new_n1141_), .C(_abc_40298_new_n1138_), .Y(_abc_40298_new_n1142_));
AOI21X1 AOI21X1_250 ( .A(\mem_dat_o[31] ), .B(_abc_40298_new_n2515_), .C(_abc_40298_new_n2608_), .Y(_abc_40298_new_n2876_));
AOI21X1 AOI21X1_251 ( .A(_abc_40298_new_n2877_), .B(_abc_40298_new_n2875_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2878_));
AOI21X1 AOI21X1_252 ( .A(mem_stb_o), .B(mem_stall_i), .C(state_q_3_), .Y(_abc_40298_new_n2889_));
AOI21X1 AOI21X1_253 ( .A(_abc_40298_new_n2892_), .B(mem_cyc_o), .C(state_q_3_), .Y(_abc_40298_new_n2893_));
AOI21X1 AOI21X1_254 ( .A(_abc_40298_new_n2913_), .B(_abc_40298_new_n2915_), .C(_abc_40298_new_n663_), .Y(_abc_40298_new_n2916_));
AOI21X1 AOI21X1_255 ( .A(_abc_40298_new_n2927_), .B(_abc_40298_new_n2932_), .C(_abc_40298_new_n2933_), .Y(_abc_40298_new_n2934_));
AOI21X1 AOI21X1_256 ( .A(_abc_40298_new_n2949_), .B(_abc_40298_new_n2941_), .C(_abc_40298_new_n2948_), .Y(_abc_40298_new_n2959_));
AOI21X1 AOI21X1_257 ( .A(_abc_40298_new_n2981_), .B(_abc_40298_new_n2980_), .C(_abc_40298_new_n663_), .Y(_abc_40298_new_n2982_));
AOI21X1 AOI21X1_258 ( .A(_abc_40298_new_n2970_), .B(_abc_40298_new_n2961_), .C(_abc_40298_new_n2969_), .Y(_abc_40298_new_n2997_));
AOI21X1 AOI21X1_259 ( .A(_abc_40298_new_n2989_), .B(_abc_40298_new_n2976_), .C(_abc_40298_new_n2998_), .Y(_abc_40298_new_n2999_));
AOI21X1 AOI21X1_26 ( .A(_abc_40298_new_n1137_), .B(_abc_40298_new_n1142_), .C(_abc_40298_new_n1143_), .Y(_0esr_q_31_0__9_));
AOI21X1 AOI21X1_260 ( .A(_abc_40298_new_n2960_), .B(_abc_40298_new_n2996_), .C(_abc_40298_new_n3000_), .Y(_abc_40298_new_n3001_));
AOI21X1 AOI21X1_261 ( .A(_abc_40298_new_n3045_), .B(_abc_40298_new_n3046_), .C(_abc_40298_new_n3047_), .Y(_abc_40298_new_n3048_));
AOI21X1 AOI21X1_262 ( .A(_abc_40298_new_n3051_), .B(_abc_40298_new_n3068_), .C(_abc_40298_new_n3067_), .Y(_abc_40298_new_n3069_));
AOI21X1 AOI21X1_263 ( .A(_abc_40298_new_n3075_), .B(_abc_40298_new_n3076_), .C(_abc_40298_new_n3077_), .Y(_abc_40298_new_n3078_));
AOI21X1 AOI21X1_264 ( .A(_abc_40298_new_n3097_), .B(_abc_40298_new_n3098_), .C(_abc_40298_new_n3099_), .Y(_abc_40298_new_n3100_));
AOI21X1 AOI21X1_265 ( .A(_abc_40298_new_n3110_), .B(_abc_40298_new_n3114_), .C(_abc_40298_new_n3116_), .Y(_abc_40298_new_n3117_));
AOI21X1 AOI21X1_266 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_23_), .B(_abc_40298_new_n3036_), .C(_abc_40298_new_n3123_), .Y(_abc_40298_new_n3124_));
AOI21X1 AOI21X1_267 ( .A(_abc_40298_new_n3051_), .B(_abc_40298_new_n3127_), .C(_abc_40298_new_n3126_), .Y(_abc_40298_new_n3128_));
AOI21X1 AOI21X1_268 ( .A(_abc_40298_new_n3148_), .B(_abc_40298_new_n3149_), .C(_abc_40298_new_n669_), .Y(_abc_40298_new_n3150_));
AOI21X1 AOI21X1_269 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_27_), .B(_abc_40298_new_n3036_), .C(_abc_40298_new_n3163_), .Y(_abc_40298_new_n3164_));
AOI21X1 AOI21X1_27 ( .A(_abc_40298_new_n1156_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n1157_), .Y(_0esr_q_31_0__10_));
AOI21X1 AOI21X1_270 ( .A(_abc_40298_new_n3184_), .B(_abc_40298_new_n3185_), .C(_abc_40298_new_n663_), .Y(_abc_40298_new_n3186_));
AOI21X1 AOI21X1_271 ( .A(_abc_40298_new_n3190_), .B(_abc_40298_new_n3191_), .C(_abc_40298_new_n3192_), .Y(_abc_40298_new_n3193_));
AOI21X1 AOI21X1_272 ( .A(_abc_40298_new_n1027_), .B(REGFILE_SIM_reg_bank_wr_i), .C(fault_o), .Y(_abc_40298_new_n3200_));
AOI21X1 AOI21X1_273 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2100_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2604_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__0_));
AOI21X1 AOI21X1_274 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2109_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2606_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__1_));
AOI21X1 AOI21X1_275 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2112_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2608_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__2_));
AOI21X1 AOI21X1_276 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2115_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2610_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__3_));
AOI21X1 AOI21X1_277 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2118_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2612_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__4_));
AOI21X1 AOI21X1_278 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2121_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2614_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__5_));
AOI21X1 AOI21X1_279 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2124_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2616_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__6_));
AOI21X1 AOI21X1_28 ( .A(_abc_40298_new_n1160_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n1161_), .Y(_0sr_q_31_0__2_));
AOI21X1 AOI21X1_280 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2127_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2618_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__7_));
AOI21X1 AOI21X1_281 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2130_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2620_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__8_));
AOI21X1 AOI21X1_282 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2133_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2622_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__9_));
AOI21X1 AOI21X1_283 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2136_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2624_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__10_));
AOI21X1 AOI21X1_284 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2139_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2626_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__11_));
AOI21X1 AOI21X1_285 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2142_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2628_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__12_));
AOI21X1 AOI21X1_286 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2145_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2630_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__13_));
AOI21X1 AOI21X1_287 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2148_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2632_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__14_));
AOI21X1 AOI21X1_288 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2151_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2634_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__15_));
AOI21X1 AOI21X1_289 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2154_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2636_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__16_));
AOI21X1 AOI21X1_29 ( .A(_abc_40298_new_n1163_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n1164_), .Y(_0sr_q_31_0__9_));
AOI21X1 AOI21X1_290 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2157_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2638_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__17_));
AOI21X1 AOI21X1_291 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2160_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2640_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__18_));
AOI21X1 AOI21X1_292 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2163_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2642_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__19_));
AOI21X1 AOI21X1_293 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2166_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2644_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__20_));
AOI21X1 AOI21X1_294 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2169_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2646_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__21_));
AOI21X1 AOI21X1_295 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2172_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2648_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__22_));
AOI21X1 AOI21X1_296 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2175_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2650_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__23_));
AOI21X1 AOI21X1_297 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2178_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2652_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__24_));
AOI21X1 AOI21X1_298 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2181_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2654_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__25_));
AOI21X1 AOI21X1_299 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2184_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2656_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__26_));
AOI21X1 AOI21X1_3 ( .A(_abc_40298_new_n697_), .B(_abc_40298_new_n655_), .C(_abc_40298_new_n703_), .Y(_abc_40298_new_n704_));
AOI21X1 AOI21X1_30 ( .A(_abc_40298_new_n1171_), .B(_abc_40298_new_n1167_), .C(_abc_40298_new_n1166_), .Y(_0sr_q_31_0__10_));
AOI21X1 AOI21X1_300 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2187_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2658_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__27_));
AOI21X1 AOI21X1_301 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2190_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2660_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__28_));
AOI21X1 AOI21X1_302 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2193_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2662_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__29_));
AOI21X1 AOI21X1_303 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2196_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2664_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__30_));
AOI21X1 AOI21X1_304 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2199_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2666_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__31_));
AOI21X1 AOI21X1_305 ( .A(REGFILE_SIM_reg_bank_reg_r22_0_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4233_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4236_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4237_));
AOI21X1 AOI21X1_306 ( .A(REGFILE_SIM_reg_bank_reg_r22_1_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4233_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4276_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4277_));
AOI21X1 AOI21X1_307 ( .A(REGFILE_SIM_reg_bank_reg_r22_2_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4233_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4308_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4309_));
AOI21X1 AOI21X1_308 ( .A(REGFILE_SIM_reg_bank_reg_r22_3_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4233_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4340_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4341_));
AOI21X1 AOI21X1_309 ( .A(REGFILE_SIM_reg_bank_reg_r22_4_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4233_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4372_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4373_));
AOI21X1 AOI21X1_31 ( .A(_abc_40298_new_n1192_), .B(_abc_40298_new_n1193_), .C(_abc_40298_new_n1194_), .Y(_0epc_q_31_0__0_));
AOI21X1 AOI21X1_310 ( .A(REGFILE_SIM_reg_bank_reg_r22_5_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4233_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4404_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4405_));
AOI21X1 AOI21X1_311 ( .A(REGFILE_SIM_reg_bank_reg_r22_6_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4233_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4436_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4437_));
AOI21X1 AOI21X1_312 ( .A(REGFILE_SIM_reg_bank_reg_r22_7_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4233_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4468_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4469_));
AOI21X1 AOI21X1_313 ( .A(REGFILE_SIM_reg_bank_reg_r22_8_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4233_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4500_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4501_));
AOI21X1 AOI21X1_314 ( .A(REGFILE_SIM_reg_bank_reg_r22_9_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4233_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4532_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4533_));
AOI21X1 AOI21X1_315 ( .A(REGFILE_SIM_reg_bank_reg_r22_10_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4233_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4564_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4565_));
AOI21X1 AOI21X1_316 ( .A(REGFILE_SIM_reg_bank_reg_r22_11_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4233_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4596_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4597_));
AOI21X1 AOI21X1_317 ( .A(REGFILE_SIM_reg_bank_reg_r22_12_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4233_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4628_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4629_));
AOI21X1 AOI21X1_318 ( .A(REGFILE_SIM_reg_bank_reg_r22_13_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4233_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4660_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4661_));
AOI21X1 AOI21X1_319 ( .A(REGFILE_SIM_reg_bank_reg_r22_14_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4233_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4692_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4693_));
AOI21X1 AOI21X1_32 ( .A(_abc_40298_new_n1204_), .B(_abc_40298_new_n1205_), .C(_abc_40298_new_n1206_), .Y(_0epc_q_31_0__1_));
AOI21X1 AOI21X1_320 ( .A(REGFILE_SIM_reg_bank_reg_r22_15_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4233_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4724_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4725_));
AOI21X1 AOI21X1_321 ( .A(REGFILE_SIM_reg_bank_reg_r22_16_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4233_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4756_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4757_));
AOI21X1 AOI21X1_322 ( .A(REGFILE_SIM_reg_bank_reg_r22_17_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4233_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4788_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4789_));
AOI21X1 AOI21X1_323 ( .A(REGFILE_SIM_reg_bank_reg_r22_18_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4233_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4820_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4821_));
AOI21X1 AOI21X1_324 ( .A(REGFILE_SIM_reg_bank_reg_r22_19_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4233_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4852_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4853_));
AOI21X1 AOI21X1_325 ( .A(REGFILE_SIM_reg_bank_reg_r22_20_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4233_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4884_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4885_));
AOI21X1 AOI21X1_326 ( .A(REGFILE_SIM_reg_bank_reg_r22_21_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4233_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4916_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4917_));
AOI21X1 AOI21X1_327 ( .A(REGFILE_SIM_reg_bank_reg_r22_22_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4233_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4948_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4949_));
AOI21X1 AOI21X1_328 ( .A(REGFILE_SIM_reg_bank_reg_r22_23_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4233_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4980_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4981_));
AOI21X1 AOI21X1_329 ( .A(REGFILE_SIM_reg_bank_reg_r22_24_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4233_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5012_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5013_));
AOI21X1 AOI21X1_33 ( .A(_abc_40298_new_n1065_), .B(epc_q_2_), .C(_abc_40298_new_n1176_), .Y(_abc_40298_new_n1219_));
AOI21X1 AOI21X1_330 ( .A(REGFILE_SIM_reg_bank_reg_r22_25_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4233_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5044_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5045_));
AOI21X1 AOI21X1_331 ( .A(REGFILE_SIM_reg_bank_reg_r22_26_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4233_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5076_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5077_));
AOI21X1 AOI21X1_332 ( .A(REGFILE_SIM_reg_bank_reg_r22_27_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4233_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5108_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5109_));
AOI21X1 AOI21X1_333 ( .A(REGFILE_SIM_reg_bank_reg_r22_28_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4233_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5140_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5141_));
AOI21X1 AOI21X1_334 ( .A(REGFILE_SIM_reg_bank_reg_r22_29_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4233_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5172_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5173_));
AOI21X1 AOI21X1_335 ( .A(REGFILE_SIM_reg_bank_reg_r22_30_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4233_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5204_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5205_));
AOI21X1 AOI21X1_336 ( .A(REGFILE_SIM_reg_bank_reg_r22_31_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4233_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5236_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5237_));
AOI21X1 AOI21X1_337 ( .A(REGFILE_SIM_reg_bank_reg_r22_0_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5305_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5308_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5309_));
AOI21X1 AOI21X1_338 ( .A(REGFILE_SIM_reg_bank_reg_r22_1_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5305_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5348_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5349_));
AOI21X1 AOI21X1_339 ( .A(REGFILE_SIM_reg_bank_reg_r22_2_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5305_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5380_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5381_));
AOI21X1 AOI21X1_34 ( .A(_abc_40298_new_n1226_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n1227_), .Y(_0epc_q_31_0__2_));
AOI21X1 AOI21X1_340 ( .A(REGFILE_SIM_reg_bank_reg_r22_3_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5305_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5412_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5413_));
AOI21X1 AOI21X1_341 ( .A(REGFILE_SIM_reg_bank_reg_r22_4_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5305_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5444_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5445_));
AOI21X1 AOI21X1_342 ( .A(REGFILE_SIM_reg_bank_reg_r22_5_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5305_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5476_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5477_));
AOI21X1 AOI21X1_343 ( .A(REGFILE_SIM_reg_bank_reg_r22_6_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5305_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5508_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5509_));
AOI21X1 AOI21X1_344 ( .A(REGFILE_SIM_reg_bank_reg_r22_7_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5305_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5540_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5541_));
AOI21X1 AOI21X1_345 ( .A(REGFILE_SIM_reg_bank_reg_r22_8_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5305_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5572_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5573_));
AOI21X1 AOI21X1_346 ( .A(REGFILE_SIM_reg_bank_reg_r22_9_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5305_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5604_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5605_));
AOI21X1 AOI21X1_347 ( .A(REGFILE_SIM_reg_bank_reg_r22_10_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5305_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5636_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5637_));
AOI21X1 AOI21X1_348 ( .A(REGFILE_SIM_reg_bank_reg_r22_11_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5305_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5668_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5669_));
AOI21X1 AOI21X1_349 ( .A(REGFILE_SIM_reg_bank_reg_r22_12_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5305_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5700_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5701_));
AOI21X1 AOI21X1_35 ( .A(_abc_40298_new_n1249_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n1250_), .Y(_0epc_q_31_0__3_));
AOI21X1 AOI21X1_350 ( .A(REGFILE_SIM_reg_bank_reg_r22_13_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5305_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5732_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5733_));
AOI21X1 AOI21X1_351 ( .A(REGFILE_SIM_reg_bank_reg_r22_14_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5305_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5764_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5765_));
AOI21X1 AOI21X1_352 ( .A(REGFILE_SIM_reg_bank_reg_r22_15_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5305_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5796_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5797_));
AOI21X1 AOI21X1_353 ( .A(REGFILE_SIM_reg_bank_reg_r22_16_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5305_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5828_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5829_));
AOI21X1 AOI21X1_354 ( .A(REGFILE_SIM_reg_bank_reg_r22_17_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5305_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5860_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5861_));
AOI21X1 AOI21X1_355 ( .A(REGFILE_SIM_reg_bank_reg_r22_18_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5305_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5892_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5893_));
AOI21X1 AOI21X1_356 ( .A(REGFILE_SIM_reg_bank_reg_r22_19_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5305_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5924_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5925_));
AOI21X1 AOI21X1_357 ( .A(REGFILE_SIM_reg_bank_reg_r22_20_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5305_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5956_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5957_));
AOI21X1 AOI21X1_358 ( .A(REGFILE_SIM_reg_bank_reg_r22_21_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5305_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5988_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5989_));
AOI21X1 AOI21X1_359 ( .A(REGFILE_SIM_reg_bank_reg_r22_22_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5305_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n6020_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6021_));
AOI21X1 AOI21X1_36 ( .A(_abc_40298_new_n1065_), .B(epc_q_4_), .C(_abc_40298_new_n1176_), .Y(_abc_40298_new_n1268_));
AOI21X1 AOI21X1_360 ( .A(REGFILE_SIM_reg_bank_reg_r22_23_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5305_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n6052_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6053_));
AOI21X1 AOI21X1_361 ( .A(REGFILE_SIM_reg_bank_reg_r22_24_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5305_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n6084_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6085_));
AOI21X1 AOI21X1_362 ( .A(REGFILE_SIM_reg_bank_reg_r22_25_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5305_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n6116_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6117_));
AOI21X1 AOI21X1_363 ( .A(REGFILE_SIM_reg_bank_reg_r22_26_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5305_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n6148_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6149_));
AOI21X1 AOI21X1_364 ( .A(REGFILE_SIM_reg_bank_reg_r22_27_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5305_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n6180_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6181_));
AOI21X1 AOI21X1_365 ( .A(REGFILE_SIM_reg_bank_reg_r22_28_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5305_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n6212_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6213_));
AOI21X1 AOI21X1_366 ( .A(REGFILE_SIM_reg_bank_reg_r22_29_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5305_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n6244_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6245_));
AOI21X1 AOI21X1_367 ( .A(REGFILE_SIM_reg_bank_reg_r22_30_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5305_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n6276_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6277_));
AOI21X1 AOI21X1_368 ( .A(REGFILE_SIM_reg_bank_reg_r22_31_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5305_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n6308_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6309_));
AOI21X1 AOI21X1_369 ( .A(alu__abc_38674_new_n150_), .B(alu__abc_38674_new_n314_), .C(alu__abc_38674_new_n313_), .Y(alu__abc_38674_new_n315_));
AOI21X1 AOI21X1_37 ( .A(_abc_40298_new_n1275_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n1276_), .Y(_0epc_q_31_0__4_));
AOI21X1 AOI21X1_370 ( .A(alu__abc_38674_new_n311_), .B(alu__abc_38674_new_n315_), .C(alu__abc_38674_new_n133_), .Y(alu__abc_38674_new_n316_));
AOI21X1 AOI21X1_371 ( .A(alu__abc_38674_new_n322_), .B(alu__abc_38674_new_n324_), .C(alu__abc_38674_new_n323_), .Y(alu__abc_38674_new_n325_));
AOI21X1 AOI21X1_372 ( .A(alu__abc_38674_new_n337_), .B(alu__abc_38674_new_n272_), .C(alu__abc_38674_new_n342_), .Y(alu__abc_38674_new_n343_));
AOI21X1 AOI21X1_373 ( .A(alu__abc_38674_new_n348_), .B(alu__abc_38674_new_n328_), .C(alu__abc_38674_new_n333_), .Y(alu__abc_38674_new_n349_));
AOI21X1 AOI21X1_374 ( .A(alu__abc_38674_new_n360_), .B(alu__abc_38674_new_n363_), .C(alu__abc_38674_new_n367_), .Y(alu__abc_38674_new_n368_));
AOI21X1 AOI21X1_375 ( .A(alu__abc_38674_new_n370_), .B(alu__abc_38674_new_n327_), .C(alu__abc_38674_new_n198_), .Y(alu__abc_38674_new_n371_));
AOI21X1 AOI21X1_376 ( .A(alu__abc_38674_new_n169_), .B(alu__abc_38674_new_n374_), .C(alu__abc_38674_new_n373_), .Y(alu__abc_38674_new_n375_));
AOI21X1 AOI21X1_377 ( .A(alu__abc_38674_new_n183_), .B(alu__abc_38674_new_n179_), .C(alu__abc_38674_new_n181_), .Y(alu__abc_38674_new_n399_));
AOI21X1 AOI21X1_378 ( .A(alu__abc_38674_new_n398_), .B(alu__abc_38674_new_n400_), .C(alu__abc_38674_new_n397_), .Y(alu__abc_38674_new_n401_));
AOI21X1 AOI21X1_379 ( .A(alu__abc_38674_new_n162_), .B(alu__abc_38674_new_n157_), .C(alu__abc_38674_new_n160_), .Y(alu__abc_38674_new_n402_));
AOI21X1 AOI21X1_38 ( .A(_abc_40298_new_n1299_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n1300_), .Y(_0epc_q_31_0__5_));
AOI21X1 AOI21X1_380 ( .A(alu__abc_38674_new_n385_), .B(alu__abc_38674_new_n388_), .C(alu__abc_38674_new_n403_), .Y(alu__abc_38674_new_n404_));
AOI21X1 AOI21X1_381 ( .A(alu__abc_38674_new_n140_), .B(alu__abc_38674_new_n136_), .C(alu__abc_38674_new_n138_), .Y(alu__abc_38674_new_n414_));
AOI21X1 AOI21X1_382 ( .A(alu__abc_38674_new_n145_), .B(alu__abc_38674_new_n415_), .C(alu__abc_38674_new_n147_), .Y(alu__abc_38674_new_n416_));
AOI21X1 AOI21X1_383 ( .A(alu__abc_38674_new_n321_), .B(alu__abc_38674_new_n112_), .C(alu__abc_38674_new_n118_), .Y(alu__abc_38674_new_n419_));
AOI21X1 AOI21X1_384 ( .A(alu__abc_38674_new_n423_), .B(alu__abc_38674_new_n266_), .C(alu__abc_38674_new_n269_), .Y(alu__abc_38674_new_n424_));
AOI21X1 AOI21X1_385 ( .A(alu__abc_38674_new_n439_), .B(alu__abc_38674_new_n426_), .C(alu__abc_38674_new_n248_), .Y(alu__abc_38674_new_n440_));
AOI21X1 AOI21X1_386 ( .A(alu__abc_38674_new_n435_), .B(alu__abc_38674_new_n425_), .C(alu__abc_38674_new_n441_), .Y(alu__abc_38674_new_n442_));
AOI21X1 AOI21X1_387 ( .A(alu__abc_38674_new_n207_), .B(alu__abc_38674_new_n203_), .C(alu__abc_38674_new_n205_), .Y(alu__abc_38674_new_n450_));
AOI21X1 AOI21X1_388 ( .A(alu__abc_38674_new_n451_), .B(alu__abc_38674_new_n212_), .C(alu__abc_38674_new_n218_), .Y(alu__abc_38674_new_n452_));
AOI21X1 AOI21X1_389 ( .A(alu__abc_38674_new_n449_), .B(alu__abc_38674_new_n457_), .C(alu__abc_38674_new_n455_), .Y(alu__abc_38674_new_n458_));
AOI21X1 AOI21X1_39 ( .A(_abc_40298_new_n1281_), .B(_abc_40298_new_n1263_), .C(_abc_40298_new_n1280_), .Y(_abc_40298_new_n1312_));
AOI21X1 AOI21X1_390 ( .A(alu__abc_38674_new_n406_), .B(alu__abc_38674_new_n409_), .C(alu__abc_38674_new_n469_), .Y(alu__abc_38674_new_n470_));
AOI21X1 AOI21X1_391 ( .A(alu__abc_38674_new_n464_), .B(alu__abc_38674_new_n487_), .C(alu__abc_38674_new_n486_), .Y(alu__abc_38674_new_n488_));
AOI21X1 AOI21X1_392 ( .A(alu__abc_38674_new_n464_), .B(alu__abc_38674_new_n467_), .C(alu__abc_38674_new_n417_), .Y(alu__abc_38674_new_n491_));
AOI21X1 AOI21X1_393 ( .A(alu__abc_38674_new_n422_), .B(alu__abc_38674_new_n424_), .C(alu__abc_38674_new_n523_), .Y(alu__abc_38674_new_n524_));
AOI21X1 AOI21X1_394 ( .A(alu__abc_38674_new_n525_), .B(alu__abc_38674_new_n515_), .C(alu__abc_38674_new_n456_), .Y(alu__abc_38674_new_n526_));
AOI21X1 AOI21X1_395 ( .A(alu__abc_38674_new_n531_), .B(alu__abc_38674_new_n530_), .C(alu__abc_38674_new_n513_), .Y(alu__abc_38674_new_n532_));
AOI21X1 AOI21X1_396 ( .A(alu__abc_38674_new_n422_), .B(alu__abc_38674_new_n424_), .C(alu__abc_38674_new_n434_), .Y(alu__abc_38674_new_n541_));
AOI21X1 AOI21X1_397 ( .A(alu__abc_38674_new_n422_), .B(alu__abc_38674_new_n424_), .C(alu__abc_38674_new_n521_), .Y(alu__abc_38674_new_n550_));
AOI21X1 AOI21X1_398 ( .A(alu__abc_38674_new_n421_), .B(alu__abc_38674_new_n268_), .C(alu__abc_38674_new_n266_), .Y(alu__abc_38674_new_n553_));
AOI21X1 AOI21X1_399 ( .A(alu__abc_38674_new_n525_), .B(alu__abc_38674_new_n515_), .C(alu__abc_38674_new_n215_), .Y(alu__abc_38674_new_n582_));
AOI21X1 AOI21X1_4 ( .A(_abc_40298_new_n710_), .B(_abc_40298_new_n713_), .C(_abc_40298_new_n655_), .Y(_abc_40298_new_n714_));
AOI21X1 AOI21X1_40 ( .A(_abc_40298_new_n1313_), .B(_abc_40298_new_n1318_), .C(_abc_40298_new_n984_), .Y(_abc_40298_new_n1319_));
AOI21X1 AOI21X1_400 ( .A(alu__abc_38674_new_n589_), .B(alu__abc_38674_new_n445_), .C(alu__abc_38674_new_n235_), .Y(alu__abc_38674_new_n590_));
AOI21X1 AOI21X1_401 ( .A(alu__abc_38674_new_n480_), .B(alu__abc_38674_new_n391_), .C(alu__abc_38674_new_n388_), .Y(alu__abc_38674_new_n611_));
AOI21X1 AOI21X1_402 ( .A(alu__abc_38674_new_n652_), .B(alu_b_i_2_), .C(alu_b_i_3_), .Y(alu__abc_38674_new_n653_));
AOI21X1 AOI21X1_403 ( .A(alu__abc_38674_new_n294_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n659_), .Y(alu__abc_38674_new_n660_));
AOI21X1 AOI21X1_404 ( .A(alu__abc_38674_new_n689_), .B(alu_b_i_4_), .C(alu__abc_38674_new_n658_), .Y(alu__abc_38674_new_n690_));
AOI21X1 AOI21X1_405 ( .A(alu__abc_38674_new_n786_), .B(alu__abc_38674_new_n564_), .C(alu__abc_38674_new_n382_), .Y(alu__abc_38674_new_n793_));
AOI21X1 AOI21X1_406 ( .A(alu_a_i_1_), .B(alu__abc_38674_new_n712_), .C(alu__abc_38674_new_n795_), .Y(alu__abc_38674_new_n796_));
AOI21X1 AOI21X1_407 ( .A(alu__abc_38674_new_n828_), .B(alu_b_i_3_), .C(alu_b_i_4_), .Y(alu__abc_38674_new_n829_));
AOI21X1 AOI21X1_408 ( .A(alu__abc_38674_new_n337_), .B(alu__abc_38674_new_n834_), .C(alu__abc_38674_new_n782_), .Y(alu__abc_38674_new_n835_));
AOI21X1 AOI21X1_409 ( .A(alu__abc_38674_new_n266_), .B(alu__abc_38674_new_n844_), .C(alu__abc_38674_new_n845_), .Y(alu__abc_38674_new_n846_));
AOI21X1 AOI21X1_41 ( .A(_abc_40298_new_n1321_), .B(_abc_40298_new_n1175_), .C(_abc_40298_new_n1323_), .Y(_abc_40298_new_n1324_));
AOI21X1 AOI21X1_410 ( .A(alu__abc_38674_new_n832_), .B(alu__abc_38674_new_n833_), .C(alu__abc_38674_new_n848_), .Y(alu__abc_38674_new_n849_));
AOI21X1 AOI21X1_411 ( .A(alu__abc_38674_new_n878_), .B(alu__abc_38674_new_n519_), .C(alu__abc_38674_new_n658_), .Y(alu__abc_38674_new_n879_));
AOI21X1 AOI21X1_412 ( .A(alu__abc_38674_new_n570_), .B(alu__abc_38674_new_n558_), .C(alu__abc_38674_new_n382_), .Y(alu__abc_38674_new_n881_));
AOI21X1 AOI21X1_413 ( .A(alu__abc_38674_new_n641_), .B(alu__abc_38674_new_n562_), .C(alu__abc_38674_new_n718_), .Y(alu__abc_38674_new_n885_));
AOI21X1 AOI21X1_414 ( .A(alu__abc_38674_new_n889_), .B(alu__abc_38674_new_n701_), .C(alu__abc_38674_new_n891_), .Y(alu__abc_38674_new_n892_));
AOI21X1 AOI21X1_415 ( .A(alu__abc_38674_new_n555_), .B(alu__abc_38674_new_n896_), .C(alu__abc_38674_new_n897_), .Y(alu__abc_38674_new_n898_));
AOI21X1 AOI21X1_416 ( .A(alu__abc_38674_new_n343_), .B(alu__abc_38674_new_n335_), .C(alu__abc_38674_new_n782_), .Y(alu__abc_38674_new_n906_));
AOI21X1 AOI21X1_417 ( .A(alu__abc_38674_new_n932_), .B(alu__abc_38674_new_n701_), .C(alu__abc_38674_new_n936_), .Y(alu__abc_38674_new_n937_));
AOI21X1 AOI21X1_418 ( .A(alu__abc_38674_new_n908_), .B(alu__abc_38674_new_n924_), .C(alu__abc_38674_new_n938_), .Y(alu__abc_38674_new_n939_));
AOI21X1 AOI21X1_419 ( .A(alu__abc_38674_new_n771_), .B(alu__abc_38674_new_n338_), .C(alu__abc_38674_new_n941_), .Y(alu__abc_38674_new_n942_));
AOI21X1 AOI21X1_42 ( .A(_abc_40298_new_n1232_), .B(_abc_40298_new_n1308_), .C(_abc_40298_new_n1324_), .Y(_abc_40298_new_n1325_));
AOI21X1 AOI21X1_420 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n947_), .C(alu__abc_38674_new_n950_), .Y(alu__abc_38674_new_n951_));
AOI21X1 AOI21X1_421 ( .A(alu__abc_38674_new_n946_), .B(alu_b_i_4_), .C(alu__abc_38674_new_n951_), .Y(alu__abc_38674_new_n952_));
AOI21X1 AOI21X1_422 ( .A(alu__abc_38674_new_n960_), .B(alu__abc_38674_new_n701_), .C(alu__abc_38674_new_n963_), .Y(alu__abc_38674_new_n964_));
AOI21X1 AOI21X1_423 ( .A(alu__abc_38674_new_n952_), .B(alu__abc_38674_new_n908_), .C(alu__abc_38674_new_n965_), .Y(alu__abc_38674_new_n966_));
AOI21X1 AOI21X1_424 ( .A(alu__abc_38674_new_n976_), .B(alu__abc_38674_new_n428_), .C(alu__abc_38674_new_n782_), .Y(alu__abc_38674_new_n977_));
AOI21X1 AOI21X1_425 ( .A(alu__abc_38674_new_n246_), .B(alu__abc_38674_new_n703_), .C(alu__abc_38674_new_n1000_), .Y(alu__abc_38674_new_n1001_));
AOI21X1 AOI21X1_426 ( .A(alu__abc_38674_new_n999_), .B(alu__abc_38674_new_n701_), .C(alu__abc_38674_new_n1002_), .Y(alu__abc_38674_new_n1003_));
AOI21X1 AOI21X1_427 ( .A(alu__abc_38674_new_n908_), .B(alu__abc_38674_new_n992_), .C(alu__abc_38674_new_n1004_), .Y(alu__abc_38674_new_n1005_));
AOI21X1 AOI21X1_428 ( .A(alu__abc_38674_new_n1008_), .B(alu__abc_38674_new_n517_), .C(alu__abc_38674_new_n782_), .Y(alu__abc_38674_new_n1009_));
AOI21X1 AOI21X1_429 ( .A(alu__abc_38674_new_n573_), .B(alu__abc_38674_new_n544_), .C(alu__abc_38674_new_n382_), .Y(alu__abc_38674_new_n1011_));
AOI21X1 AOI21X1_43 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1326_), .C(_abc_40298_new_n1071_), .Y(_abc_40298_new_n1327_));
AOI21X1 AOI21X1_430 ( .A(alu_a_i_7_), .B(alu__abc_38674_new_n712_), .C(alu__abc_38674_new_n1034_), .Y(alu__abc_38674_new_n1035_));
AOI21X1 AOI21X1_431 ( .A(alu__abc_38674_new_n248_), .B(alu__abc_38674_new_n844_), .C(alu__abc_38674_new_n1036_), .Y(alu__abc_38674_new_n1037_));
AOI21X1 AOI21X1_432 ( .A(alu__abc_38674_new_n282_), .B(alu__abc_38674_new_n544_), .C(alu__abc_38674_new_n1038_), .Y(alu__abc_38674_new_n1039_));
AOI21X1 AOI21X1_433 ( .A(alu__abc_38674_new_n349_), .B(alu__abc_38674_new_n539_), .C(alu__abc_38674_new_n782_), .Y(alu__abc_38674_new_n1041_));
AOI21X1 AOI21X1_434 ( .A(alu__abc_38674_new_n1054_), .B(alu_b_i_4_), .C(alu__abc_38674_new_n658_), .Y(alu__abc_38674_new_n1055_));
AOI21X1 AOI21X1_435 ( .A(alu_a_i_8_), .B(alu__abc_38674_new_n712_), .C(alu__abc_38674_new_n1070_), .Y(alu__abc_38674_new_n1071_));
AOI21X1 AOI21X1_436 ( .A(alu__abc_38674_new_n282_), .B(alu__abc_38674_new_n540_), .C(alu__abc_38674_new_n1072_), .Y(alu__abc_38674_new_n1073_));
AOI21X1 AOI21X1_437 ( .A(alu__abc_38674_new_n773_), .B(alu__abc_38674_new_n340_), .C(alu__abc_38674_new_n1079_), .Y(alu__abc_38674_new_n1080_));
AOI21X1 AOI21X1_438 ( .A(alu__abc_38674_new_n1109_), .B(alu__abc_38674_new_n236_), .C(alu__abc_38674_new_n782_), .Y(alu__abc_38674_new_n1110_));
AOI21X1 AOI21X1_439 ( .A(alu__abc_38674_new_n1119_), .B(alu_b_i_4_), .C(alu__abc_38674_new_n658_), .Y(alu__abc_38674_new_n1120_));
AOI21X1 AOI21X1_44 ( .A(_abc_40298_new_n1328_), .B(_abc_40298_new_n1307_), .C(_abc_40298_new_n1329_), .Y(_0epc_q_31_0__6_));
AOI21X1 AOI21X1_440 ( .A(alu__abc_38674_new_n1129_), .B(alu__abc_38674_new_n701_), .C(alu__abc_38674_new_n1131_), .Y(alu__abc_38674_new_n1132_));
AOI21X1 AOI21X1_441 ( .A(alu__abc_38674_new_n234_), .B(alu__abc_38674_new_n703_), .C(alu__abc_38674_new_n1134_), .Y(alu__abc_38674_new_n1135_));
AOI21X1 AOI21X1_442 ( .A(alu__abc_38674_new_n1138_), .B(alu__abc_38674_new_n239_), .C(alu__abc_38674_new_n782_), .Y(alu__abc_38674_new_n1139_));
AOI21X1 AOI21X1_443 ( .A(alu__abc_38674_new_n1112_), .B(alu__abc_38674_new_n592_), .C(alu__abc_38674_new_n382_), .Y(alu__abc_38674_new_n1141_));
AOI21X1 AOI21X1_444 ( .A(alu__abc_38674_new_n240_), .B(alu__abc_38674_new_n705_), .C(alu__abc_38674_new_n1164_), .Y(alu__abc_38674_new_n1165_));
AOI21X1 AOI21X1_445 ( .A(alu__abc_38674_new_n1162_), .B(alu__abc_38674_new_n701_), .C(alu__abc_38674_new_n1166_), .Y(alu__abc_38674_new_n1167_));
AOI21X1 AOI21X1_446 ( .A(alu__abc_38674_new_n282_), .B(alu__abc_38674_new_n1145_), .C(alu__abc_38674_new_n1168_), .Y(alu__abc_38674_new_n1169_));
AOI21X1 AOI21X1_447 ( .A(alu__abc_38674_new_n1171_), .B(alu__abc_38674_new_n215_), .C(alu__abc_38674_new_n782_), .Y(alu__abc_38674_new_n1172_));
AOI21X1 AOI21X1_448 ( .A(alu_a_i_12_), .B(alu__abc_38674_new_n712_), .C(alu__abc_38674_new_n1188_), .Y(alu__abc_38674_new_n1189_));
AOI21X1 AOI21X1_449 ( .A(alu__abc_38674_new_n282_), .B(alu__abc_38674_new_n595_), .C(alu__abc_38674_new_n1197_), .Y(alu__abc_38674_new_n1198_));
AOI21X1 AOI21X1_45 ( .A(_abc_40298_new_n1316_), .B(_abc_40298_new_n1343_), .C(_abc_40298_new_n984_), .Y(_abc_40298_new_n1351_));
AOI21X1 AOI21X1_450 ( .A(alu__abc_38674_new_n1215_), .B(alu_b_i_4_), .C(alu__abc_38674_new_n658_), .Y(alu__abc_38674_new_n1216_));
AOI21X1 AOI21X1_451 ( .A(alu__abc_38674_new_n451_), .B(alu__abc_38674_new_n705_), .C(alu__abc_38674_new_n1226_), .Y(alu__abc_38674_new_n1227_));
AOI21X1 AOI21X1_452 ( .A(alu_a_i_13_), .B(alu__abc_38674_new_n712_), .C(alu__abc_38674_new_n1228_), .Y(alu__abc_38674_new_n1229_));
AOI21X1 AOI21X1_453 ( .A(alu__abc_38674_new_n1214_), .B(alu__abc_38674_new_n1216_), .C(alu__abc_38674_new_n1230_), .Y(alu__abc_38674_new_n1231_));
AOI21X1 AOI21X1_454 ( .A(alu__abc_38674_new_n1204_), .B(alu__abc_38674_new_n576_), .C(alu__abc_38674_new_n382_), .Y(alu__abc_38674_new_n1238_));
AOI21X1 AOI21X1_455 ( .A(alu__abc_38674_new_n989_), .B(alu__abc_38674_new_n340_), .C(alu__abc_38674_new_n1079_), .Y(alu__abc_38674_new_n1241_));
AOI21X1 AOI21X1_456 ( .A(alu__abc_38674_new_n453_), .B(alu__abc_38674_new_n705_), .C(alu__abc_38674_new_n1256_), .Y(alu__abc_38674_new_n1257_));
AOI21X1 AOI21X1_457 ( .A(alu__abc_38674_new_n1255_), .B(alu__abc_38674_new_n701_), .C(alu__abc_38674_new_n1258_), .Y(alu__abc_38674_new_n1259_));
AOI21X1 AOI21X1_458 ( .A(alu__abc_38674_new_n282_), .B(alu__abc_38674_new_n1240_), .C(alu__abc_38674_new_n1260_), .Y(alu__abc_38674_new_n1261_));
AOI21X1 AOI21X1_459 ( .A(alu__abc_38674_new_n1263_), .B(alu__abc_38674_new_n208_), .C(alu__abc_38674_new_n782_), .Y(alu__abc_38674_new_n1264_));
AOI21X1 AOI21X1_46 ( .A(_abc_40298_new_n1335_), .B(_abc_40298_new_n1359_), .C(_abc_40298_new_n1360_), .Y(_0epc_q_31_0__7_));
AOI21X1 AOI21X1_460 ( .A(alu_a_i_15_), .B(alu__abc_38674_new_n712_), .C(alu__abc_38674_new_n1289_), .Y(alu__abc_38674_new_n1290_));
AOI21X1 AOI21X1_461 ( .A(alu__abc_38674_new_n1278_), .B(alu__abc_38674_new_n908_), .C(alu__abc_38674_new_n1291_), .Y(alu__abc_38674_new_n1292_));
AOI21X1 AOI21X1_462 ( .A(alu__abc_38674_new_n1301_), .B(alu__abc_38674_new_n465_), .C(alu__abc_38674_new_n782_), .Y(alu__abc_38674_new_n1302_));
AOI21X1 AOI21X1_463 ( .A(alu__abc_38674_new_n465_), .B(alu__abc_38674_new_n705_), .C(alu__abc_38674_new_n1320_), .Y(alu__abc_38674_new_n1321_));
AOI21X1 AOI21X1_464 ( .A(alu_a_i_16_), .B(alu__abc_38674_new_n712_), .C(alu__abc_38674_new_n1322_), .Y(alu__abc_38674_new_n1323_));
AOI21X1 AOI21X1_465 ( .A(alu__abc_38674_new_n1306_), .B(alu__abc_38674_new_n1307_), .C(alu__abc_38674_new_n1324_), .Y(alu__abc_38674_new_n1325_));
AOI21X1 AOI21X1_466 ( .A(alu_a_i_17_), .B(alu__abc_38674_new_n712_), .C(alu__abc_38674_new_n1353_), .Y(alu__abc_38674_new_n1354_));
AOI21X1 AOI21X1_467 ( .A(alu__abc_38674_new_n1306_), .B(alu__abc_38674_new_n1341_), .C(alu__abc_38674_new_n1355_), .Y(alu__abc_38674_new_n1356_));
AOI21X1 AOI21X1_468 ( .A(alu__abc_38674_new_n1363_), .B(alu__abc_38674_new_n306_), .C(alu__abc_38674_new_n782_), .Y(alu__abc_38674_new_n1364_));
AOI21X1 AOI21X1_469 ( .A(alu__abc_38674_new_n814_), .B(alu__abc_38674_new_n519_), .C(alu__abc_38674_new_n1305_), .Y(alu__abc_38674_new_n1366_));
AOI21X1 AOI21X1_47 ( .A(_abc_40298_new_n1313_), .B(_abc_40298_new_n1349_), .C(_abc_40298_new_n1371_), .Y(_abc_40298_new_n1372_));
AOI21X1 AOI21X1_470 ( .A(alu__abc_38674_new_n1375_), .B(alu_b_i_3_), .C(alu_b_i_4_), .Y(alu__abc_38674_new_n1376_));
AOI21X1 AOI21X1_471 ( .A(alu_a_i_18_), .B(alu__abc_38674_new_n712_), .C(alu__abc_38674_new_n1379_), .Y(alu__abc_38674_new_n1380_));
AOI21X1 AOI21X1_472 ( .A(alu__abc_38674_new_n1403_), .B(alu__abc_38674_new_n150_), .C(alu__abc_38674_new_n782_), .Y(alu__abc_38674_new_n1404_));
AOI21X1 AOI21X1_473 ( .A(alu__abc_38674_new_n1413_), .B(alu__abc_38674_new_n1414_), .C(alu__abc_38674_new_n1296_), .Y(alu__abc_38674_new_n1415_));
AOI21X1 AOI21X1_474 ( .A(alu__abc_38674_new_n1422_), .B(alu__abc_38674_new_n125_), .C(alu__abc_38674_new_n782_), .Y(alu__abc_38674_new_n1423_));
AOI21X1 AOI21X1_475 ( .A(alu__abc_38674_new_n1185_), .B(alu_b_i_3_), .C(alu_b_i_4_), .Y(alu__abc_38674_new_n1431_));
AOI21X1 AOI21X1_476 ( .A(alu_a_i_20_), .B(alu__abc_38674_new_n712_), .C(alu__abc_38674_new_n1434_), .Y(alu__abc_38674_new_n1435_));
AOI21X1 AOI21X1_477 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n1457_), .C(alu__abc_38674_new_n1458_), .Y(alu__abc_38674_new_n1459_));
AOI21X1 AOI21X1_478 ( .A(alu_a_i_21_), .B(alu__abc_38674_new_n712_), .C(alu__abc_38674_new_n1462_), .Y(alu__abc_38674_new_n1463_));
AOI21X1 AOI21X1_479 ( .A(alu__abc_38674_new_n1306_), .B(alu__abc_38674_new_n1452_), .C(alu__abc_38674_new_n1464_), .Y(alu__abc_38674_new_n1465_));
AOI21X1 AOI21X1_48 ( .A(_abc_40298_new_n1387_), .B(_abc_40298_new_n1028_), .C(_abc_40298_new_n1366_), .Y(_abc_40298_new_n1388_));
AOI21X1 AOI21X1_480 ( .A(alu__abc_38674_new_n1450_), .B(alu__abc_38674_new_n706_), .C(alu__abc_38674_new_n1467_), .Y(alu__abc_38674_new_n1468_));
AOI21X1 AOI21X1_481 ( .A(alu__abc_38674_new_n1472_), .B(alu__abc_38674_new_n381_), .C(alu__abc_38674_new_n1471_), .Y(alu__abc_38674_new_n1473_));
AOI21X1 AOI21X1_482 ( .A(alu__abc_38674_new_n1512_), .B(alu_b_i_3_), .C(alu_b_i_4_), .Y(alu__abc_38674_new_n1513_));
AOI21X1 AOI21X1_483 ( .A(alu__abc_38674_new_n1033_), .B(alu_b_i_4_), .C(alu__abc_38674_new_n700_), .Y(alu__abc_38674_new_n1515_));
AOI21X1 AOI21X1_484 ( .A(alu__abc_38674_new_n1023_), .B(alu__abc_38674_new_n519_), .C(alu__abc_38674_new_n1305_), .Y(alu__abc_38674_new_n1516_));
AOI21X1 AOI21X1_485 ( .A(alu__abc_38674_new_n118_), .B(alu__abc_38674_new_n844_), .C(alu__abc_38674_new_n1517_), .Y(alu__abc_38674_new_n1518_));
AOI21X1 AOI21X1_486 ( .A(alu__abc_38674_new_n1514_), .B(alu__abc_38674_new_n1515_), .C(alu__abc_38674_new_n1520_), .Y(alu__abc_38674_new_n1521_));
AOI21X1 AOI21X1_487 ( .A(alu__abc_38674_new_n1529_), .B(alu__abc_38674_new_n471_), .C(alu__abc_38674_new_n782_), .Y(alu__abc_38674_new_n1530_));
AOI21X1 AOI21X1_488 ( .A(alu__abc_38674_new_n471_), .B(alu__abc_38674_new_n705_), .C(alu__abc_38674_new_n1540_), .Y(alu__abc_38674_new_n1541_));
AOI21X1 AOI21X1_489 ( .A(alu__abc_38674_new_n1539_), .B(alu__abc_38674_new_n701_), .C(alu__abc_38674_new_n1542_), .Y(alu__abc_38674_new_n1543_));
AOI21X1 AOI21X1_49 ( .A(_abc_40298_new_n1402_), .B(_abc_40298_new_n1404_), .C(inst_trap_w), .Y(_abc_40298_new_n1405_));
AOI21X1 AOI21X1_490 ( .A(alu__abc_38674_new_n1306_), .B(alu__abc_38674_new_n1532_), .C(alu__abc_38674_new_n1544_), .Y(alu__abc_38674_new_n1545_));
AOI21X1 AOI21X1_491 ( .A(alu__abc_38674_new_n1554_), .B(alu__abc_38674_new_n338_), .C(alu_b_i_3_), .Y(alu__abc_38674_new_n1555_));
AOI21X1 AOI21X1_492 ( .A(alu_a_i_25_), .B(alu__abc_38674_new_n712_), .C(alu__abc_38674_new_n1565_), .Y(alu__abc_38674_new_n1566_));
AOI21X1 AOI21X1_493 ( .A(alu__abc_38674_new_n1563_), .B(alu__abc_38674_new_n1306_), .C(alu__abc_38674_new_n1567_), .Y(alu__abc_38674_new_n1568_));
AOI21X1 AOI21X1_494 ( .A(alu__abc_38674_new_n282_), .B(alu__abc_38674_new_n503_), .C(alu__abc_38674_new_n1569_), .Y(alu__abc_38674_new_n1570_));
AOI21X1 AOI21X1_495 ( .A(alu_a_i_26_), .B(alu__abc_38674_new_n712_), .C(alu__abc_38674_new_n1596_), .Y(alu__abc_38674_new_n1597_));
AOI21X1 AOI21X1_496 ( .A(alu__abc_38674_new_n1583_), .B(alu__abc_38674_new_n1306_), .C(alu__abc_38674_new_n1598_), .Y(alu__abc_38674_new_n1599_));
AOI21X1 AOI21X1_497 ( .A(alu_a_i_27_), .B(alu__abc_38674_new_n712_), .C(alu__abc_38674_new_n1615_), .Y(alu__abc_38674_new_n1616_));
AOI21X1 AOI21X1_498 ( .A(alu__abc_38674_new_n1162_), .B(alu__abc_38674_new_n1317_), .C(alu__abc_38674_new_n1617_), .Y(alu__abc_38674_new_n1618_));
AOI21X1 AOI21X1_499 ( .A(alu__abc_38674_new_n701_), .B(alu__abc_38674_new_n1613_), .C(alu__abc_38674_new_n1619_), .Y(alu__abc_38674_new_n1620_));
AOI21X1 AOI21X1_5 ( .A(_abc_40298_new_n709_), .B(_abc_40298_new_n655_), .C(_abc_40298_new_n714_), .Y(_abc_40298_new_n715_));
AOI21X1 AOI21X1_50 ( .A(_abc_40298_new_n1411_), .B(_abc_40298_new_n1392_), .C(_abc_40298_new_n1412_), .Y(_0epc_q_31_0__9_));
AOI21X1 AOI21X1_500 ( .A(alu__abc_38674_new_n282_), .B(alu__abc_38674_new_n619_), .C(alu__abc_38674_new_n1621_), .Y(alu__abc_38674_new_n1622_));
AOI21X1 AOI21X1_501 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n1637_), .C(alu__abc_38674_new_n702_), .Y(alu__abc_38674_new_n1638_));
AOI21X1 AOI21X1_502 ( .A(alu_a_i_28_), .B(alu__abc_38674_new_n712_), .C(alu__abc_38674_new_n1641_), .Y(alu__abc_38674_new_n1642_));
AOI21X1 AOI21X1_503 ( .A(alu__abc_38674_new_n1633_), .B(alu__abc_38674_new_n1638_), .C(alu__abc_38674_new_n1643_), .Y(alu__abc_38674_new_n1644_));
AOI21X1 AOI21X1_504 ( .A(alu__abc_38674_new_n1652_), .B(alu__abc_38674_new_n169_), .C(alu__abc_38674_new_n782_), .Y(alu__abc_38674_new_n1653_));
AOI21X1 AOI21X1_505 ( .A(alu__abc_38674_new_n1660_), .B(alu__abc_38674_new_n519_), .C(alu__abc_38674_new_n700_), .Y(alu__abc_38674_new_n1661_));
AOI21X1 AOI21X1_506 ( .A(alu__abc_38674_new_n168_), .B(alu__abc_38674_new_n705_), .C(alu__abc_38674_new_n1664_), .Y(alu__abc_38674_new_n1665_));
AOI21X1 AOI21X1_507 ( .A(alu__abc_38674_new_n1663_), .B(alu__abc_38674_new_n1306_), .C(alu__abc_38674_new_n1666_), .Y(alu__abc_38674_new_n1667_));
AOI21X1 AOI21X1_508 ( .A(alu__abc_38674_new_n282_), .B(alu__abc_38674_new_n483_), .C(alu__abc_38674_new_n1668_), .Y(alu__abc_38674_new_n1669_));
AOI21X1 AOI21X1_509 ( .A(alu__abc_38674_new_n165_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n659_), .Y(alu__abc_38674_new_n1680_));
AOI21X1 AOI21X1_51 ( .A(_abc_40298_new_n1065_), .B(_abc_40298_new_n1437_), .C(_abc_40298_new_n1176_), .Y(_abc_40298_new_n1438_));
AOI21X1 AOI21X1_510 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n1683_), .C(alu__abc_38674_new_n1684_), .Y(alu__abc_38674_new_n1685_));
AOI21X1 AOI21X1_511 ( .A(alu_b_i_4_), .B(alu__abc_38674_new_n1254_), .C(alu__abc_38674_new_n1685_), .Y(alu__abc_38674_new_n1686_));
AOI21X1 AOI21X1_512 ( .A(alu_a_i_30_), .B(alu__abc_38674_new_n712_), .C(alu__abc_38674_new_n1687_), .Y(alu__abc_38674_new_n1688_));
AOI21X1 AOI21X1_513 ( .A(alu__abc_38674_new_n1686_), .B(alu__abc_38674_new_n699_), .C(alu__abc_38674_new_n1689_), .Y(alu__abc_38674_new_n1690_));
AOI21X1 AOI21X1_514 ( .A(alu__abc_38674_new_n162_), .B(alu__abc_38674_new_n705_), .C(alu__abc_38674_new_n1713_), .Y(alu__abc_38674_new_n1714_));
AOI21X1 AOI21X1_515 ( .A(alu__abc_38674_new_n1286_), .B(alu__abc_38674_new_n1317_), .C(alu__abc_38674_new_n1715_), .Y(alu__abc_38674_new_n1716_));
AOI21X1 AOI21X1_516 ( .A(alu__abc_38674_new_n1704_), .B(alu__abc_38674_new_n1306_), .C(alu__abc_38674_new_n1717_), .Y(alu__abc_38674_new_n1718_));
AOI21X1 AOI21X1_517 ( .A(alu__abc_38674_new_n282_), .B(alu__abc_38674_new_n615_), .C(alu__abc_38674_new_n1719_), .Y(alu__abc_38674_new_n1720_));
AOI21X1 AOI21X1_518 ( .A(alu__abc_38674_new_n1726_), .B(alu__abc_38674_new_n163_), .C(alu__abc_38674_new_n1728_), .Y(alu__abc_38674_new_n1729_));
AOI21X1 AOI21X1_52 ( .A(_abc_40298_new_n1443_), .B(_abc_40298_new_n1420_), .C(_abc_40298_new_n1444_), .Y(_0epc_q_31_0__10_));
AOI21X1 AOI21X1_53 ( .A(_abc_40298_new_n1456_), .B(_abc_40298_new_n1461_), .C(_abc_40298_new_n984_), .Y(_abc_40298_new_n1462_));
AOI21X1 AOI21X1_54 ( .A(_abc_40298_new_n1470_), .B(_abc_40298_new_n1451_), .C(_abc_40298_new_n1471_), .Y(_0epc_q_31_0__11_));
AOI21X1 AOI21X1_55 ( .A(_abc_40298_new_n1429_), .B(_abc_40298_new_n1458_), .C(_abc_40298_new_n1482_), .Y(_abc_40298_new_n1483_));
AOI21X1 AOI21X1_56 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1504_), .C(_abc_40298_new_n1071_), .Y(_abc_40298_new_n1505_));
AOI21X1 AOI21X1_57 ( .A(_abc_40298_new_n1506_), .B(_abc_40298_new_n1477_), .C(_abc_40298_new_n1507_), .Y(_0epc_q_31_0__12_));
AOI21X1 AOI21X1_58 ( .A(_abc_40298_new_n1494_), .B(_abc_40298_new_n1518_), .C(_abc_40298_new_n1520_), .Y(_abc_40298_new_n1521_));
AOI21X1 AOI21X1_59 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_13_), .B(_abc_40298_new_n1176_), .C(_abc_40298_new_n1523_), .Y(_abc_40298_new_n1524_));
AOI21X1 AOI21X1_6 ( .A(_abc_40298_new_n721_), .B(_abc_40298_new_n724_), .C(_abc_40298_new_n655_), .Y(_abc_40298_new_n725_));
AOI21X1 AOI21X1_60 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1527_), .C(_abc_40298_new_n1071_), .Y(_abc_40298_new_n1528_));
AOI21X1 AOI21X1_61 ( .A(_abc_40298_new_n1529_), .B(_abc_40298_new_n1510_), .C(_abc_40298_new_n1530_), .Y(_0epc_q_31_0__13_));
AOI21X1 AOI21X1_62 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_14_), .B(_abc_40298_new_n1176_), .C(_abc_40298_new_n1232_), .Y(_abc_40298_new_n1554_));
AOI21X1 AOI21X1_63 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1556_), .C(_abc_40298_new_n1071_), .Y(_abc_40298_new_n1557_));
AOI21X1 AOI21X1_64 ( .A(_abc_40298_new_n1558_), .B(_abc_40298_new_n1538_), .C(_abc_40298_new_n1559_), .Y(_0epc_q_31_0__14_));
AOI21X1 AOI21X1_65 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_15_), .B(_abc_40298_new_n1176_), .C(_abc_40298_new_n1232_), .Y(_abc_40298_new_n1580_));
AOI21X1 AOI21X1_66 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1582_), .C(_abc_40298_new_n1071_), .Y(_abc_40298_new_n1583_));
AOI21X1 AOI21X1_67 ( .A(_abc_40298_new_n1584_), .B(_abc_40298_new_n1567_), .C(_abc_40298_new_n1585_), .Y(_0epc_q_31_0__15_));
AOI21X1 AOI21X1_68 ( .A(_abc_40298_new_n1573_), .B(_abc_40298_new_n1545_), .C(_abc_40298_new_n1572_), .Y(_abc_40298_new_n1597_));
AOI21X1 AOI21X1_69 ( .A(_abc_40298_new_n1602_), .B(_abc_40298_new_n1607_), .C(_abc_40298_new_n1608_), .Y(_abc_40298_new_n1609_));
AOI21X1 AOI21X1_7 ( .A(_abc_40298_new_n720_), .B(_abc_40298_new_n655_), .C(_abc_40298_new_n725_), .Y(_abc_40298_new_n726_));
AOI21X1 AOI21X1_70 ( .A(epc_q_16_), .B(_abc_40298_new_n1065_), .C(_abc_40298_new_n1609_), .Y(_abc_40298_new_n1610_));
AOI21X1 AOI21X1_71 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1615_), .C(_abc_40298_new_n1071_), .Y(_abc_40298_new_n1616_));
AOI21X1 AOI21X1_72 ( .A(_abc_40298_new_n1617_), .B(_abc_40298_new_n1591_), .C(_abc_40298_new_n1618_), .Y(_0epc_q_31_0__16_));
AOI21X1 AOI21X1_73 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_17_), .B(_abc_40298_new_n1176_), .C(_abc_40298_new_n1232_), .Y(_abc_40298_new_n1637_));
AOI21X1 AOI21X1_74 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1639_), .C(_abc_40298_new_n1071_), .Y(_abc_40298_new_n1640_));
AOI21X1 AOI21X1_75 ( .A(_abc_40298_new_n1641_), .B(_abc_40298_new_n1624_), .C(_abc_40298_new_n1642_), .Y(_0epc_q_31_0__17_));
AOI21X1 AOI21X1_76 ( .A(_abc_40298_new_n1630_), .B(_abc_40298_new_n1605_), .C(_abc_40298_new_n1629_), .Y(_abc_40298_new_n1654_));
AOI21X1 AOI21X1_77 ( .A(_abc_40298_new_n1652_), .B(_abc_40298_new_n1653_), .C(_abc_40298_new_n1655_), .Y(_abc_40298_new_n1656_));
AOI21X1 AOI21X1_78 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_18_), .B(_abc_40298_new_n1176_), .C(_abc_40298_new_n1232_), .Y(_abc_40298_new_n1667_));
AOI21X1 AOI21X1_79 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1669_), .C(_abc_40298_new_n1071_), .Y(_abc_40298_new_n1670_));
AOI21X1 AOI21X1_8 ( .A(_abc_40298_new_n733_), .B(_abc_40298_new_n655_), .C(_abc_40298_new_n631_), .Y(_abc_40298_new_n734_));
AOI21X1 AOI21X1_80 ( .A(_abc_40298_new_n1671_), .B(_abc_40298_new_n1650_), .C(_abc_40298_new_n1672_), .Y(_0epc_q_31_0__18_));
AOI21X1 AOI21X1_81 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_19_), .B(_abc_40298_new_n1176_), .C(_abc_40298_new_n1232_), .Y(_abc_40298_new_n1690_));
AOI21X1 AOI21X1_82 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1692_), .C(_abc_40298_new_n1071_), .Y(_abc_40298_new_n1693_));
AOI21X1 AOI21X1_83 ( .A(_abc_40298_new_n1694_), .B(_abc_40298_new_n1678_), .C(_abc_40298_new_n1695_), .Y(_0epc_q_31_0__19_));
AOI21X1 AOI21X1_84 ( .A(_abc_40298_new_n1685_), .B(_abc_40298_new_n1659_), .C(_abc_40298_new_n1684_), .Y(_abc_40298_new_n1705_));
AOI21X1 AOI21X1_85 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_20_), .B(_abc_40298_new_n1176_), .C(_abc_40298_new_n1232_), .Y(_abc_40298_new_n1719_));
AOI21X1 AOI21X1_86 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1721_), .C(_abc_40298_new_n1071_), .Y(_abc_40298_new_n1722_));
AOI21X1 AOI21X1_87 ( .A(_abc_40298_new_n1723_), .B(_abc_40298_new_n1702_), .C(_abc_40298_new_n1724_), .Y(_0epc_q_31_0__20_));
AOI21X1 AOI21X1_88 ( .A(_abc_40298_new_n1713_), .B(_abc_40298_new_n1740_), .C(_abc_40298_new_n984_), .Y(_abc_40298_new_n1742_));
AOI21X1 AOI21X1_89 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_21_), .B(_abc_40298_new_n1176_), .C(_abc_40298_new_n1232_), .Y(_abc_40298_new_n1746_));
AOI21X1 AOI21X1_9 ( .A(_abc_40298_new_n742_), .B(_abc_40298_new_n655_), .C(_abc_40298_new_n631_), .Y(_abc_40298_new_n743_));
AOI21X1 AOI21X1_90 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1748_), .C(_abc_40298_new_n1071_), .Y(_abc_40298_new_n1749_));
AOI21X1 AOI21X1_91 ( .A(_abc_40298_new_n1750_), .B(_abc_40298_new_n1730_), .C(_abc_40298_new_n1751_), .Y(_0epc_q_31_0__21_));
AOI21X1 AOI21X1_92 ( .A(_abc_40298_new_n1710_), .B(_abc_40298_new_n1761_), .C(_abc_40298_new_n1763_), .Y(_abc_40298_new_n1764_));
AOI21X1 AOI21X1_93 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_22_), .B(_abc_40298_new_n1176_), .C(_abc_40298_new_n1232_), .Y(_abc_40298_new_n1775_));
AOI21X1 AOI21X1_94 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1777_), .C(_abc_40298_new_n1071_), .Y(_abc_40298_new_n1778_));
AOI21X1 AOI21X1_95 ( .A(_abc_40298_new_n1779_), .B(_abc_40298_new_n1759_), .C(_abc_40298_new_n1780_), .Y(_0epc_q_31_0__22_));
AOI21X1 AOI21X1_96 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_23_), .B(_abc_40298_new_n1176_), .C(_abc_40298_new_n1232_), .Y(_abc_40298_new_n1798_));
AOI21X1 AOI21X1_97 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1800_), .C(_abc_40298_new_n1071_), .Y(_abc_40298_new_n1801_));
AOI21X1 AOI21X1_98 ( .A(_abc_40298_new_n1802_), .B(_abc_40298_new_n1786_), .C(_abc_40298_new_n1803_), .Y(_0epc_q_31_0__23_));
AOI21X1 AOI21X1_99 ( .A(_abc_40298_new_n1792_), .B(_abc_40298_new_n1767_), .C(_abc_40298_new_n1791_), .Y(_abc_40298_new_n1815_));
AOI22X1 AOI22X1_1 ( .A(\mem_dat_i[24] ), .B(_abc_40298_new_n674_), .C(\mem_dat_i[8] ), .D(_abc_40298_new_n673_), .Y(_abc_40298_new_n675_));
AOI22X1 AOI22X1_10 ( .A(_abc_40298_new_n673_), .B(\mem_dat_i[14] ), .C(\mem_dat_i[22] ), .D(_abc_40298_new_n677_), .Y(_abc_40298_new_n750_));
AOI22X1 AOI22X1_100 ( .A(state_q_3_), .B(pc_q_14_), .C(\mem_addr_o[14] ), .D(_abc_40298_new_n2883_), .Y(_abc_40298_new_n3030_));
AOI22X1 AOI22X1_101 ( .A(state_q_3_), .B(pc_q_15_), .C(\mem_addr_o[15] ), .D(_abc_40298_new_n2895_), .Y(_abc_40298_new_n3043_));
AOI22X1 AOI22X1_102 ( .A(state_q_3_), .B(pc_q_16_), .C(\mem_addr_o[16] ), .D(_abc_40298_new_n2895_), .Y(_abc_40298_new_n3059_));
AOI22X1 AOI22X1_103 ( .A(state_q_3_), .B(pc_q_17_), .C(\mem_addr_o[17] ), .D(_abc_40298_new_n2895_), .Y(_abc_40298_new_n3064_));
AOI22X1 AOI22X1_104 ( .A(state_q_3_), .B(pc_q_18_), .C(\mem_addr_o[18] ), .D(_abc_40298_new_n2895_), .Y(_abc_40298_new_n3073_));
AOI22X1 AOI22X1_105 ( .A(state_q_3_), .B(pc_q_19_), .C(\mem_addr_o[19] ), .D(_abc_40298_new_n2883_), .Y(_abc_40298_new_n3080_));
AOI22X1 AOI22X1_106 ( .A(state_q_3_), .B(pc_q_20_), .C(\mem_addr_o[20] ), .D(_abc_40298_new_n2895_), .Y(_abc_40298_new_n3095_));
AOI22X1 AOI22X1_107 ( .A(state_q_3_), .B(pc_q_21_), .C(\mem_addr_o[21] ), .D(_abc_40298_new_n2883_), .Y(_abc_40298_new_n3102_));
AOI22X1 AOI22X1_108 ( .A(state_q_3_), .B(pc_q_22_), .C(\mem_addr_o[22] ), .D(_abc_40298_new_n2895_), .Y(_abc_40298_new_n3112_));
AOI22X1 AOI22X1_109 ( .A(state_q_3_), .B(pc_q_23_), .C(\mem_addr_o[23] ), .D(_abc_40298_new_n2895_), .Y(_abc_40298_new_n3120_));
AOI22X1 AOI22X1_11 ( .A(\mem_dat_i[30] ), .B(_abc_40298_new_n674_), .C(\mem_dat_i[6] ), .D(_abc_40298_new_n679_), .Y(_abc_40298_new_n751_));
AOI22X1 AOI22X1_110 ( .A(state_q_3_), .B(pc_q_24_), .C(\mem_addr_o[24] ), .D(_abc_40298_new_n2895_), .Y(_abc_40298_new_n3133_));
AOI22X1 AOI22X1_111 ( .A(state_q_3_), .B(pc_q_25_), .C(\mem_addr_o[25] ), .D(_abc_40298_new_n2883_), .Y(_abc_40298_new_n3143_));
AOI22X1 AOI22X1_112 ( .A(state_q_3_), .B(pc_q_27_), .C(\mem_addr_o[27] ), .D(_abc_40298_new_n2895_), .Y(_abc_40298_new_n3159_));
AOI22X1 AOI22X1_113 ( .A(state_q_3_), .B(pc_q_28_), .C(\mem_addr_o[28] ), .D(_abc_40298_new_n2895_), .Y(_abc_40298_new_n3170_));
AOI22X1 AOI22X1_114 ( .A(state_q_3_), .B(pc_q_29_), .C(\mem_addr_o[29] ), .D(_abc_40298_new_n2895_), .Y(_abc_40298_new_n3175_));
AOI22X1 AOI22X1_115 ( .A(_abc_40298_new_n3036_), .B(_abc_40298_new_n3180_), .C(_abc_40298_new_n3182_), .D(_abc_40298_new_n3165_), .Y(_abc_40298_new_n3183_));
AOI22X1 AOI22X1_116 ( .A(state_q_3_), .B(pc_q_30_), .C(\mem_addr_o[30] ), .D(_abc_40298_new_n2883_), .Y(_abc_40298_new_n3188_));
AOI22X1 AOI22X1_117 ( .A(state_q_3_), .B(pc_q_31_), .C(\mem_addr_o[31] ), .D(_abc_40298_new_n2883_), .Y(_abc_40298_new_n3195_));
AOI22X1 AOI22X1_118 ( .A(alu__abc_38674_new_n282_), .B(alu__abc_38674_new_n692_), .C(alu__abc_38674_new_n563_), .D(alu__abc_38674_new_n703_), .Y(alu__abc_38674_new_n704_));
AOI22X1 AOI22X1_119 ( .A(alu__abc_38674_new_n269_), .B(alu__abc_38674_new_n844_), .C(alu__abc_38674_new_n271_), .D(alu__abc_38674_new_n705_), .Y(alu__abc_38674_new_n890_));
AOI22X1 AOI22X1_12 ( .A(\mem_dat_i[31] ), .B(_abc_40298_new_n674_), .C(\mem_dat_i[15] ), .D(_abc_40298_new_n673_), .Y(_abc_40298_new_n755_));
AOI22X1 AOI22X1_120 ( .A(alu__abc_38674_new_n703_), .B(alu__abc_38674_new_n520_), .C(alu__abc_38674_new_n335_), .D(alu__abc_38674_new_n705_), .Y(alu__abc_38674_new_n934_));
AOI22X1 AOI22X1_121 ( .A(alu__abc_38674_new_n431_), .B(alu__abc_38674_new_n844_), .C(alu__abc_38674_new_n252_), .D(alu__abc_38674_new_n961_), .Y(alu__abc_38674_new_n962_));
AOI22X1 AOI22X1_122 ( .A(alu__abc_38674_new_n703_), .B(alu__abc_38674_new_n224_), .C(alu__abc_38674_new_n539_), .D(alu__abc_38674_new_n705_), .Y(alu__abc_38674_new_n1069_));
AOI22X1 AOI22X1_123 ( .A(alu__abc_38674_new_n446_), .B(alu__abc_38674_new_n844_), .C(alu__abc_38674_new_n236_), .D(alu__abc_38674_new_n705_), .Y(alu__abc_38674_new_n1130_));
AOI22X1 AOI22X1_124 ( .A(alu__abc_38674_new_n703_), .B(alu__abc_38674_new_n1351_), .C(alu__abc_38674_new_n140_), .D(alu__abc_38674_new_n705_), .Y(alu__abc_38674_new_n1352_));
AOI22X1 AOI22X1_125 ( .A(alu__abc_38674_new_n699_), .B(alu__abc_38674_new_n1398_), .C(alu__abc_38674_new_n1306_), .D(alu__abc_38674_new_n1399_), .Y(alu__abc_38674_new_n1400_));
AOI22X1 AOI22X1_126 ( .A(alu__abc_38674_new_n703_), .B(alu__abc_38674_new_n415_), .C(alu__abc_38674_new_n149_), .D(alu__abc_38674_new_n705_), .Y(alu__abc_38674_new_n1406_));
AOI22X1 AOI22X1_127 ( .A(alu__abc_38674_new_n1306_), .B(alu__abc_38674_new_n1484_), .C(alu__abc_38674_new_n699_), .D(alu__abc_38674_new_n1483_), .Y(alu__abc_38674_new_n1485_));
AOI22X1 AOI22X1_128 ( .A(alu__abc_38674_new_n703_), .B(alu__abc_38674_new_n1492_), .C(alu__abc_38674_new_n114_), .D(alu__abc_38674_new_n705_), .Y(alu__abc_38674_new_n1493_));
AOI22X1 AOI22X1_129 ( .A(alu__abc_38674_new_n1550_), .B(alu__abc_38674_new_n1555_), .C(alu_b_i_3_), .D(alu__abc_38674_new_n1345_), .Y(alu__abc_38674_new_n1556_));
AOI22X1 AOI22X1_13 ( .A(_abc_40298_new_n677_), .B(\mem_dat_i[23] ), .C(\mem_dat_i[7] ), .D(_abc_40298_new_n679_), .Y(_abc_40298_new_n756_));
AOI22X1 AOI22X1_130 ( .A(alu__abc_38674_new_n181_), .B(alu__abc_38674_new_n844_), .C(alu__abc_38674_new_n183_), .D(alu__abc_38674_new_n705_), .Y(alu__abc_38674_new_n1564_));
AOI22X1 AOI22X1_131 ( .A(alu__abc_38674_new_n282_), .B(alu__abc_38674_new_n499_), .C(alu__abc_38674_new_n381_), .D(alu__abc_38674_new_n1577_), .Y(alu__abc_38674_new_n1578_));
AOI22X1 AOI22X1_132 ( .A(alu__abc_38674_new_n188_), .B(alu__abc_38674_new_n844_), .C(alu__abc_38674_new_n190_), .D(alu__abc_38674_new_n705_), .Y(alu__abc_38674_new_n1595_));
AOI22X1 AOI22X1_133 ( .A(alu__abc_38674_new_n844_), .B(alu__abc_38674_new_n172_), .C(alu__abc_38674_new_n1639_), .D(alu__abc_38674_new_n703_), .Y(alu__abc_38674_new_n1640_));
AOI22X1 AOI22X1_134 ( .A(alu__abc_38674_new_n613_), .B(alu__abc_38674_new_n614_), .C(alu__abc_38674_new_n616_), .D(alu__abc_38674_new_n1696_), .Y(alu__abc_38674_new_n1697_));
AOI22X1 AOI22X1_14 ( .A(\mem_dat_i[7] ), .B(_abc_40298_new_n687_), .C(\mem_dat_i[23] ), .D(_abc_40298_new_n688_), .Y(_abc_40298_new_n758_));
AOI22X1 AOI22X1_15 ( .A(_abc_40298_new_n631_), .B(_abc_40298_new_n763_), .C(_abc_40298_new_n767_), .D(_abc_40298_new_n765_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_8_));
AOI22X1 AOI22X1_16 ( .A(_abc_40298_new_n631_), .B(_abc_40298_new_n769_), .C(_abc_40298_new_n767_), .D(_abc_40298_new_n773_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_9_));
AOI22X1 AOI22X1_17 ( .A(_abc_40298_new_n631_), .B(_abc_40298_new_n775_), .C(_abc_40298_new_n767_), .D(_abc_40298_new_n778_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_10_));
AOI22X1 AOI22X1_18 ( .A(_abc_40298_new_n631_), .B(_abc_40298_new_n780_), .C(_abc_40298_new_n767_), .D(_abc_40298_new_n783_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_11_));
AOI22X1 AOI22X1_19 ( .A(_abc_40298_new_n631_), .B(_abc_40298_new_n785_), .C(_abc_40298_new_n767_), .D(_abc_40298_new_n787_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_12_));
AOI22X1 AOI22X1_2 ( .A(\mem_dat_i[0] ), .B(_abc_40298_new_n687_), .C(\mem_dat_i[16] ), .D(_abc_40298_new_n688_), .Y(_abc_40298_new_n689_));
AOI22X1 AOI22X1_20 ( .A(_abc_40298_new_n631_), .B(_abc_40298_new_n789_), .C(_abc_40298_new_n767_), .D(_abc_40298_new_n791_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_13_));
AOI22X1 AOI22X1_21 ( .A(_abc_40298_new_n631_), .B(_abc_40298_new_n793_), .C(_abc_40298_new_n767_), .D(_abc_40298_new_n797_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_14_));
AOI22X1 AOI22X1_22 ( .A(_abc_40298_new_n631_), .B(_abc_40298_new_n799_), .C(_abc_40298_new_n767_), .D(_abc_40298_new_n801_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_15_));
AOI22X1 AOI22X1_23 ( .A(_abc_40298_new_n631_), .B(_abc_40298_new_n803_), .C(_abc_40298_new_n767_), .D(_abc_40298_new_n807_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_16_));
AOI22X1 AOI22X1_24 ( .A(_abc_40298_new_n631_), .B(_abc_40298_new_n809_), .C(_abc_40298_new_n767_), .D(_abc_40298_new_n812_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_17_));
AOI22X1 AOI22X1_25 ( .A(_abc_40298_new_n631_), .B(_abc_40298_new_n814_), .C(_abc_40298_new_n767_), .D(_abc_40298_new_n817_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_18_));
AOI22X1 AOI22X1_26 ( .A(_abc_40298_new_n631_), .B(_abc_40298_new_n819_), .C(_abc_40298_new_n767_), .D(_abc_40298_new_n822_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_19_));
AOI22X1 AOI22X1_27 ( .A(_abc_40298_new_n631_), .B(_abc_40298_new_n824_), .C(_abc_40298_new_n767_), .D(_abc_40298_new_n827_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_20_));
AOI22X1 AOI22X1_28 ( .A(_abc_40298_new_n631_), .B(_abc_40298_new_n829_), .C(_abc_40298_new_n767_), .D(_abc_40298_new_n832_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_21_));
AOI22X1 AOI22X1_29 ( .A(_abc_40298_new_n631_), .B(_abc_40298_new_n834_), .C(_abc_40298_new_n767_), .D(_abc_40298_new_n837_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_22_));
AOI22X1 AOI22X1_3 ( .A(_abc_40298_new_n673_), .B(\mem_dat_i[9] ), .C(\mem_dat_i[17] ), .D(_abc_40298_new_n677_), .Y(_abc_40298_new_n700_));
AOI22X1 AOI22X1_30 ( .A(_abc_40298_new_n631_), .B(_abc_40298_new_n839_), .C(_abc_40298_new_n767_), .D(_abc_40298_new_n842_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_23_));
AOI22X1 AOI22X1_31 ( .A(_abc_40298_new_n631_), .B(_abc_40298_new_n844_), .C(_abc_40298_new_n767_), .D(_abc_40298_new_n847_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_24_));
AOI22X1 AOI22X1_32 ( .A(_abc_40298_new_n631_), .B(_abc_40298_new_n849_), .C(_abc_40298_new_n767_), .D(_abc_40298_new_n852_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_25_));
AOI22X1 AOI22X1_33 ( .A(_abc_40298_new_n631_), .B(_abc_40298_new_n854_), .C(_abc_40298_new_n767_), .D(_abc_40298_new_n857_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_26_));
AOI22X1 AOI22X1_34 ( .A(_abc_40298_new_n631_), .B(_abc_40298_new_n859_), .C(_abc_40298_new_n767_), .D(_abc_40298_new_n862_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_27_));
AOI22X1 AOI22X1_35 ( .A(_abc_40298_new_n631_), .B(_abc_40298_new_n864_), .C(_abc_40298_new_n767_), .D(_abc_40298_new_n867_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_28_));
AOI22X1 AOI22X1_36 ( .A(_abc_40298_new_n631_), .B(_abc_40298_new_n869_), .C(_abc_40298_new_n767_), .D(_abc_40298_new_n872_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_29_));
AOI22X1 AOI22X1_37 ( .A(_abc_40298_new_n631_), .B(_abc_40298_new_n874_), .C(_abc_40298_new_n767_), .D(_abc_40298_new_n877_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_30_));
AOI22X1 AOI22X1_38 ( .A(_abc_40298_new_n631_), .B(_abc_40298_new_n879_), .C(_abc_40298_new_n767_), .D(_abc_40298_new_n882_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_31_));
AOI22X1 AOI22X1_39 ( .A(_abc_40298_new_n964_), .B(_abc_40298_new_n1006_), .C(alu_greater_than_signed_o), .D(_abc_40298_new_n1107_), .Y(_abc_40298_new_n1111_));
AOI22X1 AOI22X1_4 ( .A(_abc_40298_new_n673_), .B(\mem_dat_i[10] ), .C(\mem_dat_i[18] ), .D(_abc_40298_new_n677_), .Y(_abc_40298_new_n711_));
AOI22X1 AOI22X1_40 ( .A(epc_q_0_), .B(_abc_40298_new_n1065_), .C(next_pc_r_0_), .D(_abc_40298_new_n985_), .Y(_abc_40298_new_n1174_));
AOI22X1 AOI22X1_41 ( .A(epc_q_1_), .B(_abc_40298_new_n1065_), .C(next_pc_r_1_), .D(_abc_40298_new_n985_), .Y(_abc_40298_new_n1196_));
AOI22X1 AOI22X1_42 ( .A(_abc_40298_new_n1030_), .B(_abc_40298_new_n1176_), .C(_abc_40298_new_n1219_), .D(_abc_40298_new_n1218_), .Y(_abc_40298_new_n1220_));
AOI22X1 AOI22X1_43 ( .A(_abc_40298_new_n1260_), .B(_abc_40298_new_n1176_), .C(_abc_40298_new_n1268_), .D(_abc_40298_new_n1267_), .Y(_abc_40298_new_n1269_));
AOI22X1 AOI22X1_44 ( .A(epc_q_5_), .B(_abc_40298_new_n1065_), .C(_abc_40298_new_n985_), .D(_abc_40298_new_n1283_), .Y(_abc_40298_new_n1284_));
AOI22X1 AOI22X1_45 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_10_), .B(_abc_40298_new_n1176_), .C(_abc_40298_new_n1438_), .D(_abc_40298_new_n1436_), .Y(_abc_40298_new_n1439_));
AOI22X1 AOI22X1_46 ( .A(epc_q_13_), .B(_abc_40298_new_n1065_), .C(_abc_40298_new_n1517_), .D(_abc_40298_new_n1521_), .Y(_abc_40298_new_n1522_));
AOI22X1 AOI22X1_47 ( .A(_abc_40298_new_n1232_), .B(_abc_40298_new_n1536_), .C(_abc_40298_new_n1554_), .D(_abc_40298_new_n1553_), .Y(_abc_40298_new_n1555_));
AOI22X1 AOI22X1_48 ( .A(_abc_40298_new_n1232_), .B(_abc_40298_new_n1568_), .C(_abc_40298_new_n1580_), .D(_abc_40298_new_n1579_), .Y(_abc_40298_new_n1581_));
AOI22X1 AOI22X1_49 ( .A(_abc_40298_new_n1232_), .B(_abc_40298_new_n1625_), .C(_abc_40298_new_n1637_), .D(_abc_40298_new_n1636_), .Y(_abc_40298_new_n1638_));
AOI22X1 AOI22X1_5 ( .A(_abc_40298_new_n673_), .B(\mem_dat_i[11] ), .C(\mem_dat_i[19] ), .D(_abc_40298_new_n677_), .Y(_abc_40298_new_n722_));
AOI22X1 AOI22X1_50 ( .A(_abc_40298_new_n1232_), .B(_abc_40298_new_n1648_), .C(_abc_40298_new_n1667_), .D(_abc_40298_new_n1666_), .Y(_abc_40298_new_n1668_));
AOI22X1 AOI22X1_51 ( .A(_abc_40298_new_n1232_), .B(_abc_40298_new_n1679_), .C(_abc_40298_new_n1690_), .D(_abc_40298_new_n1689_), .Y(_abc_40298_new_n1691_));
AOI22X1 AOI22X1_52 ( .A(_abc_40298_new_n1232_), .B(_abc_40298_new_n1700_), .C(_abc_40298_new_n1719_), .D(_abc_40298_new_n1718_), .Y(_abc_40298_new_n1720_));
AOI22X1 AOI22X1_53 ( .A(_abc_40298_new_n1232_), .B(_abc_40298_new_n1731_), .C(_abc_40298_new_n1746_), .D(_abc_40298_new_n1745_), .Y(_abc_40298_new_n1747_));
AOI22X1 AOI22X1_54 ( .A(_abc_40298_new_n1232_), .B(_abc_40298_new_n1757_), .C(_abc_40298_new_n1775_), .D(_abc_40298_new_n1774_), .Y(_abc_40298_new_n1776_));
AOI22X1 AOI22X1_55 ( .A(_abc_40298_new_n1232_), .B(_abc_40298_new_n1787_), .C(_abc_40298_new_n1798_), .D(_abc_40298_new_n1797_), .Y(_abc_40298_new_n1799_));
AOI22X1 AOI22X1_56 ( .A(_abc_40298_new_n1232_), .B(_abc_40298_new_n1841_), .C(_abc_40298_new_n1854_), .D(_abc_40298_new_n1852_), .Y(_abc_40298_new_n1855_));
AOI22X1 AOI22X1_57 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_6_), .B(_abc_40298_new_n931_), .C(alu_op_r_4_), .D(_abc_40298_new_n2160_), .Y(_abc_40298_new_n2161_));
AOI22X1 AOI22X1_58 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_7_), .B(_abc_40298_new_n931_), .C(alu_op_r_5_), .D(_abc_40298_new_n2160_), .Y(_abc_40298_new_n2178_));
AOI22X1 AOI22X1_59 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_8_), .B(_abc_40298_new_n931_), .C(alu_op_r_6_), .D(_abc_40298_new_n2160_), .Y(_abc_40298_new_n2180_));
AOI22X1 AOI22X1_6 ( .A(\mem_dat_i[28] ), .B(_abc_40298_new_n674_), .C(\mem_dat_i[12] ), .D(_abc_40298_new_n673_), .Y(_abc_40298_new_n729_));
AOI22X1 AOI22X1_60 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_9_), .B(_abc_40298_new_n931_), .C(alu_op_r_7_), .D(_abc_40298_new_n2160_), .Y(_abc_40298_new_n2182_));
AOI22X1 AOI22X1_61 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_10_), .B(_abc_40298_new_n931_), .C(int32_r_10_), .D(_abc_40298_new_n2160_), .Y(_abc_40298_new_n2184_));
AOI22X1 AOI22X1_62 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_11_), .B(_abc_40298_new_n931_), .C(REGFILE_SIM_reg_bank_rb_i_0_), .D(_abc_40298_new_n2160_), .Y(_abc_40298_new_n2186_));
AOI22X1 AOI22X1_63 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_12_), .B(_abc_40298_new_n931_), .C(REGFILE_SIM_reg_bank_rb_i_1_), .D(_abc_40298_new_n2160_), .Y(_abc_40298_new_n2188_));
AOI22X1 AOI22X1_64 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_13_), .B(_abc_40298_new_n931_), .C(REGFILE_SIM_reg_bank_rb_i_2_), .D(_abc_40298_new_n2160_), .Y(_abc_40298_new_n2191_));
AOI22X1 AOI22X1_65 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_14_), .B(_abc_40298_new_n931_), .C(REGFILE_SIM_reg_bank_rb_i_3_), .D(_abc_40298_new_n2160_), .Y(_abc_40298_new_n2194_));
AOI22X1 AOI22X1_66 ( .A(_abc_40298_new_n1186_), .B(_abc_40298_new_n2287_), .C(REGFILE_SIM_reg_bank_reg_ra_o_0_), .D(_abc_40298_new_n2286_), .Y(_abc_40298_new_n2288_));
AOI22X1 AOI22X1_67 ( .A(_abc_40298_new_n1186_), .B(_abc_40298_new_n2294_), .C(REGFILE_SIM_reg_bank_reg_ra_o_1_), .D(_abc_40298_new_n2286_), .Y(_abc_40298_new_n2295_));
AOI22X1 AOI22X1_68 ( .A(_abc_40298_new_n1081_), .B(esr_q_2_), .C(epc_q_2_), .D(_abc_40298_new_n1186_), .Y(_abc_40298_new_n2300_));
AOI22X1 AOI22X1_69 ( .A(_abc_40298_new_n1012_), .B(_abc_40298_new_n1476_), .C(_abc_40298_new_n2370_), .D(_abc_40298_new_n2369_), .Y(_abc_40298_new_n2371_));
AOI22X1 AOI22X1_7 ( .A(\mem_dat_i[4] ), .B(_abc_40298_new_n687_), .C(\mem_dat_i[20] ), .D(_abc_40298_new_n688_), .Y(_abc_40298_new_n733_));
AOI22X1 AOI22X1_70 ( .A(_abc_40298_new_n2381_), .B(_abc_40298_new_n2382_), .C(_abc_40298_new_n1012_), .D(_abc_40298_new_n1566_), .Y(_abc_40298_new_n2383_));
AOI22X1 AOI22X1_71 ( .A(_abc_40298_new_n635_), .B(_abc_40298_new_n2567_), .C(_abc_40298_new_n2582_), .D(_abc_40298_new_n2575_), .Y(_0mem_sel_o_3_0__0_));
AOI22X1 AOI22X1_72 ( .A(_abc_40298_new_n635_), .B(_abc_40298_new_n2584_), .C(_abc_40298_new_n2576_), .D(_abc_40298_new_n2590_), .Y(_0mem_sel_o_3_0__1_));
AOI22X1 AOI22X1_73 ( .A(_abc_40298_new_n635_), .B(_abc_40298_new_n2592_), .C(_abc_40298_new_n2596_), .D(_abc_40298_new_n2598_), .Y(_0mem_sel_o_3_0__2_));
AOI22X1 AOI22X1_74 ( .A(_abc_40298_new_n635_), .B(_abc_40298_new_n2600_), .C(_abc_40298_new_n2576_), .D(_abc_40298_new_n2605_), .Y(_0mem_sel_o_3_0__3_));
AOI22X1 AOI22X1_75 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_0_), .B(_abc_40298_new_n2581_), .C(_abc_40298_new_n2615_), .D(_abc_40298_new_n2610_), .Y(_abc_40298_new_n2616_));
AOI22X1 AOI22X1_76 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_1_), .B(_abc_40298_new_n2581_), .C(_abc_40298_new_n2623_), .D(_abc_40298_new_n2620_), .Y(_abc_40298_new_n2624_));
AOI22X1 AOI22X1_77 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_2_), .B(_abc_40298_new_n2581_), .C(_abc_40298_new_n2631_), .D(_abc_40298_new_n2628_), .Y(_abc_40298_new_n2632_));
AOI22X1 AOI22X1_78 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_3_), .B(_abc_40298_new_n2581_), .C(_abc_40298_new_n2639_), .D(_abc_40298_new_n2636_), .Y(_abc_40298_new_n2640_));
AOI22X1 AOI22X1_79 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_4_), .B(_abc_40298_new_n2581_), .C(_abc_40298_new_n2647_), .D(_abc_40298_new_n2644_), .Y(_abc_40298_new_n2648_));
AOI22X1 AOI22X1_8 ( .A(\mem_dat_i[29] ), .B(_abc_40298_new_n674_), .C(\mem_dat_i[13] ), .D(_abc_40298_new_n673_), .Y(_abc_40298_new_n738_));
AOI22X1 AOI22X1_80 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_5_), .B(_abc_40298_new_n2581_), .C(_abc_40298_new_n2655_), .D(_abc_40298_new_n2652_), .Y(_abc_40298_new_n2656_));
AOI22X1 AOI22X1_81 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_6_), .B(_abc_40298_new_n2581_), .C(_abc_40298_new_n2663_), .D(_abc_40298_new_n2660_), .Y(_abc_40298_new_n2664_));
AOI22X1 AOI22X1_82 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_7_), .B(_abc_40298_new_n2581_), .C(_abc_40298_new_n2671_), .D(_abc_40298_new_n2668_), .Y(_abc_40298_new_n2672_));
AOI22X1 AOI22X1_83 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_0_), .B(_abc_40298_new_n2597_), .C(_abc_40298_new_n2751_), .D(_abc_40298_new_n2748_), .Y(_abc_40298_new_n2752_));
AOI22X1 AOI22X1_84 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_1_), .B(_abc_40298_new_n2597_), .C(_abc_40298_new_n2759_), .D(_abc_40298_new_n2756_), .Y(_abc_40298_new_n2760_));
AOI22X1 AOI22X1_85 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_2_), .B(_abc_40298_new_n2597_), .C(_abc_40298_new_n2767_), .D(_abc_40298_new_n2764_), .Y(_abc_40298_new_n2768_));
AOI22X1 AOI22X1_86 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_3_), .B(_abc_40298_new_n2597_), .C(_abc_40298_new_n2775_), .D(_abc_40298_new_n2772_), .Y(_abc_40298_new_n2776_));
AOI22X1 AOI22X1_87 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_4_), .B(_abc_40298_new_n2597_), .C(_abc_40298_new_n2783_), .D(_abc_40298_new_n2780_), .Y(_abc_40298_new_n2784_));
AOI22X1 AOI22X1_88 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_5_), .B(_abc_40298_new_n2597_), .C(_abc_40298_new_n2791_), .D(_abc_40298_new_n2788_), .Y(_abc_40298_new_n2792_));
AOI22X1 AOI22X1_89 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_6_), .B(_abc_40298_new_n2597_), .C(_abc_40298_new_n2799_), .D(_abc_40298_new_n2796_), .Y(_abc_40298_new_n2800_));
AOI22X1 AOI22X1_9 ( .A(\mem_dat_i[5] ), .B(_abc_40298_new_n687_), .C(\mem_dat_i[21] ), .D(_abc_40298_new_n688_), .Y(_abc_40298_new_n742_));
AOI22X1 AOI22X1_90 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_7_), .B(_abc_40298_new_n2597_), .C(_abc_40298_new_n2807_), .D(_abc_40298_new_n2804_), .Y(_abc_40298_new_n2808_));
AOI22X1 AOI22X1_91 ( .A(state_q_3_), .B(pc_q_3_), .C(\mem_addr_o[3] ), .D(_abc_40298_new_n2883_), .Y(_abc_40298_new_n2918_));
AOI22X1 AOI22X1_92 ( .A(state_q_3_), .B(pc_q_4_), .C(\mem_addr_o[4] ), .D(_abc_40298_new_n2895_), .Y(_abc_40298_new_n2925_));
AOI22X1 AOI22X1_93 ( .A(state_q_3_), .B(pc_q_5_), .C(\mem_addr_o[5] ), .D(_abc_40298_new_n2883_), .Y(_abc_40298_new_n2938_));
AOI22X1 AOI22X1_94 ( .A(state_q_3_), .B(pc_q_6_), .C(\mem_addr_o[6] ), .D(_abc_40298_new_n2895_), .Y(_abc_40298_new_n2946_));
AOI22X1 AOI22X1_95 ( .A(state_q_3_), .B(pc_q_8_), .C(\mem_addr_o[8] ), .D(_abc_40298_new_n2895_), .Y(_abc_40298_new_n2966_));
AOI22X1 AOI22X1_96 ( .A(state_q_3_), .B(pc_q_9_), .C(\mem_addr_o[9] ), .D(_abc_40298_new_n2883_), .Y(_abc_40298_new_n2974_));
AOI22X1 AOI22X1_97 ( .A(state_q_3_), .B(pc_q_10_), .C(\mem_addr_o[10] ), .D(_abc_40298_new_n2883_), .Y(_abc_40298_new_n2984_));
AOI22X1 AOI22X1_98 ( .A(state_q_3_), .B(pc_q_11_), .C(\mem_addr_o[11] ), .D(_abc_40298_new_n2895_), .Y(_abc_40298_new_n2992_));
AOI22X1 AOI22X1_99 ( .A(state_q_3_), .B(pc_q_12_), .C(\mem_addr_o[12] ), .D(_abc_40298_new_n2895_), .Y(_abc_40298_new_n3008_));
DFFSR DFFSR_1 ( .CLK(clk_i), .D(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2382), .Q(state_q_0_), .R(1'h1), .S(_abc_40298_auto_rtlil_cc_1942_NotGate_33938));
DFFSR DFFSR_10 ( .CLK(clk_i), .D(_0pc_q_31_0__1_), .Q(next_pc_r_1_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_100 ( .CLK(clk_i), .D(alu_input_a_r_15_), .Q(alu_a_i_15_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_1000 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r24_6_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1001 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r24_7_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1002 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r24_8_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1003 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r24_9_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1004 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r24_10_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1005 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r24_11_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1006 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r24_12_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1007 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r24_13_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1008 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r24_14_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1009 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r24_15_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_101 ( .CLK(clk_i), .D(alu_input_a_r_16_), .Q(alu_a_i_16_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_1010 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r24_16_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1011 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r24_17_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1012 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r24_18_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1013 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r24_19_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1014 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r24_20_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1015 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r24_21_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1016 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r24_22_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1017 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r24_23_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1018 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r24_24_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1019 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r24_25_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_102 ( .CLK(clk_i), .D(alu_input_a_r_17_), .Q(alu_a_i_17_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_1020 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r24_26_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1021 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r24_27_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1022 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r24_28_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1023 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r24_29_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1024 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r24_30_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1025 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r24_31_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1026 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r25_0_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1027 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r25_1_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1028 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r25_2_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1029 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r25_3_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_103 ( .CLK(clk_i), .D(alu_input_a_r_18_), .Q(alu_a_i_18_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_1030 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r25_4_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1031 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r25_5_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1032 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r25_6_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1033 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r25_7_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1034 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r25_8_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1035 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r25_9_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1036 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r25_10_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1037 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r25_11_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1038 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r25_12_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1039 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r25_13_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_104 ( .CLK(clk_i), .D(alu_input_a_r_19_), .Q(alu_a_i_19_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_1040 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r25_14_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1041 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r25_15_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1042 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r25_16_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1043 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r25_17_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1044 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r25_18_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1045 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r25_19_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1046 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r25_20_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1047 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r25_21_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1048 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r25_22_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1049 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r25_23_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_105 ( .CLK(clk_i), .D(alu_input_a_r_20_), .Q(alu_a_i_20_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_1050 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r25_24_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1051 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r25_25_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1052 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r25_26_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1053 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r25_27_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1054 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r25_28_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1055 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r25_29_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1056 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r25_30_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1057 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r25_31_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1058 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r26_0_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1059 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r26_1_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_106 ( .CLK(clk_i), .D(alu_input_a_r_21_), .Q(alu_a_i_21_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_1060 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r26_2_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1061 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r26_3_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1062 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r26_4_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1063 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r26_5_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1064 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r26_6_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1065 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r26_7_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1066 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r26_8_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1067 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r26_9_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1068 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r26_10_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1069 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r26_11_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_107 ( .CLK(clk_i), .D(alu_input_a_r_22_), .Q(alu_a_i_22_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_1070 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r26_12_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1071 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r26_13_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1072 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r26_14_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1073 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r26_15_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1074 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r26_16_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1075 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r26_17_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1076 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r26_18_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1077 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r26_19_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1078 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r26_20_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1079 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r26_21_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_108 ( .CLK(clk_i), .D(alu_input_a_r_23_), .Q(alu_a_i_23_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_1080 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r26_22_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1081 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r26_23_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1082 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r26_24_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1083 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r26_25_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1084 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r26_26_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1085 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r26_27_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1086 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r26_28_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1087 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r26_29_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1088 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r26_30_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1089 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r26_31_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_109 ( .CLK(clk_i), .D(alu_input_a_r_24_), .Q(alu_a_i_24_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_1090 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r27_0_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1091 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r27_1_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1092 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r27_2_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1093 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r27_3_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1094 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r27_4_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1095 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r27_5_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1096 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r27_6_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1097 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r27_7_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1098 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r27_8_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1099 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r27_9_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_11 ( .CLK(clk_i), .D(_0pc_q_31_0__2_), .Q(pc_q_2_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_110 ( .CLK(clk_i), .D(alu_input_a_r_25_), .Q(alu_a_i_25_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_1100 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r27_10_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1101 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r27_11_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1102 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r27_12_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1103 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r27_13_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1104 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r27_14_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1105 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r27_15_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1106 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r27_16_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1107 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r27_17_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1108 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r27_18_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1109 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r27_19_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_111 ( .CLK(clk_i), .D(alu_input_a_r_26_), .Q(alu_a_i_26_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_1110 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r27_20_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1111 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r27_21_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1112 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r27_22_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1113 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r27_23_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1114 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r27_24_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1115 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r27_25_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1116 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r27_26_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1117 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r27_27_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1118 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r27_28_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1119 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r27_29_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_112 ( .CLK(clk_i), .D(alu_input_a_r_27_), .Q(alu_a_i_27_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_1120 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r27_30_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1121 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r27_31_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1122 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r28_0_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1123 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r28_1_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1124 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r28_2_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1125 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r28_3_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1126 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r28_4_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1127 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r28_5_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1128 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r28_6_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1129 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r28_7_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_113 ( .CLK(clk_i), .D(alu_input_a_r_28_), .Q(alu_a_i_28_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_1130 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r28_8_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1131 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r28_9_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1132 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r28_10_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1133 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r28_11_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1134 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r28_12_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1135 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r28_13_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1136 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r28_14_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1137 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r28_15_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1138 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r28_16_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1139 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r28_17_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_114 ( .CLK(clk_i), .D(alu_input_a_r_29_), .Q(alu_a_i_29_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_1140 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r28_18_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1141 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r28_19_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1142 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r28_20_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1143 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r28_21_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1144 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r28_22_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1145 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r28_23_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1146 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r28_24_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1147 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r28_25_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1148 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r28_26_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1149 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r28_27_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_115 ( .CLK(clk_i), .D(alu_input_a_r_30_), .Q(alu_a_i_30_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_1150 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r28_28_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1151 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r28_29_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1152 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r28_30_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1153 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r28_31_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1154 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r29_0_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1155 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r29_1_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1156 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r29_2_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1157 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r29_3_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1158 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r29_4_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1159 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r29_5_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_116 ( .CLK(clk_i), .D(alu_input_a_r_31_), .Q(alu_a_i_31_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_1160 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r29_6_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1161 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r29_7_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1162 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r29_8_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1163 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r29_9_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1164 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r29_10_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1165 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r29_11_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1166 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r29_12_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1167 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r29_13_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1168 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r29_14_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1169 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r29_15_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_117 ( .CLK(clk_i), .D(alu_input_b_r_0_), .Q(alu_b_i_0_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_1170 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r29_16_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1171 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r29_17_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1172 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r29_18_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1173 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r29_19_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1174 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r29_20_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1175 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r29_21_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1176 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r29_22_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1177 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r29_23_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1178 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r29_24_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1179 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r29_25_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_118 ( .CLK(clk_i), .D(alu_input_b_r_1_), .Q(alu_b_i_1_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_1180 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r29_26_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1181 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r29_27_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1182 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r29_28_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1183 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r29_29_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1184 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r29_30_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1185 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r29_31_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1186 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r30_0_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1187 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r30_1_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1188 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r30_2_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1189 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r30_3_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_119 ( .CLK(clk_i), .D(alu_input_b_r_2_), .Q(alu_b_i_2_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_1190 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r30_4_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1191 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r30_5_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1192 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r30_6_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1193 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r30_7_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1194 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r30_8_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1195 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r30_9_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1196 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r30_10_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1197 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r30_11_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1198 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r30_12_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1199 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r30_13_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_12 ( .CLK(clk_i), .D(_0pc_q_31_0__3_), .Q(pc_q_3_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_120 ( .CLK(clk_i), .D(alu_input_b_r_3_), .Q(alu_b_i_3_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_1200 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r30_14_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1201 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r30_15_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1202 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r30_16_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1203 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r30_17_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1204 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r30_18_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1205 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r30_19_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1206 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r30_20_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1207 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r30_21_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1208 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r30_22_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1209 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r30_23_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_121 ( .CLK(clk_i), .D(alu_input_b_r_4_), .Q(alu_b_i_4_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_1210 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r30_24_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1211 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r30_25_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1212 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r30_26_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1213 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r30_27_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1214 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r30_28_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1215 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r30_29_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1216 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r30_30_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1217 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r30_31_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1218 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r31_0_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1219 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r31_1_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_122 ( .CLK(clk_i), .D(alu_input_b_r_5_), .Q(alu_b_i_5_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_1220 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r31_2_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1221 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r31_3_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1222 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r31_4_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1223 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r31_5_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1224 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r31_6_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1225 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r31_7_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1226 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r31_8_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1227 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r31_9_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1228 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r31_10_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1229 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r31_11_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_123 ( .CLK(clk_i), .D(alu_input_b_r_6_), .Q(alu_b_i_6_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_1230 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r31_12_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1231 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r31_13_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1232 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r31_14_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1233 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r31_15_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1234 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r31_16_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1235 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r31_17_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1236 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r31_18_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1237 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r31_19_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1238 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r31_20_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1239 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r31_21_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_124 ( .CLK(clk_i), .D(alu_input_b_r_7_), .Q(alu_b_i_7_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_1240 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r31_22_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1241 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r31_23_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1242 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r31_24_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1243 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r31_25_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1244 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r31_26_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1245 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r31_27_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1246 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r31_28_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1247 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r31_29_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1248 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r31_30_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_1249 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r31_31_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_125 ( .CLK(clk_i), .D(alu_input_b_r_8_), .Q(alu_b_i_8_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_126 ( .CLK(clk_i), .D(alu_input_b_r_9_), .Q(alu_b_i_9_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_127 ( .CLK(clk_i), .D(alu_input_b_r_10_), .Q(alu_b_i_10_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_128 ( .CLK(clk_i), .D(alu_input_b_r_11_), .Q(alu_b_i_11_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_129 ( .CLK(clk_i), .D(alu_input_b_r_12_), .Q(alu_b_i_12_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_13 ( .CLK(clk_i), .D(_0pc_q_31_0__4_), .Q(pc_q_4_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_130 ( .CLK(clk_i), .D(alu_input_b_r_13_), .Q(alu_b_i_13_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_131 ( .CLK(clk_i), .D(alu_input_b_r_14_), .Q(alu_b_i_14_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_132 ( .CLK(clk_i), .D(alu_input_b_r_15_), .Q(alu_b_i_15_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_133 ( .CLK(clk_i), .D(alu_input_b_r_16_), .Q(alu_b_i_16_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_134 ( .CLK(clk_i), .D(alu_input_b_r_17_), .Q(alu_b_i_17_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_135 ( .CLK(clk_i), .D(alu_input_b_r_18_), .Q(alu_b_i_18_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_136 ( .CLK(clk_i), .D(alu_input_b_r_19_), .Q(alu_b_i_19_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_137 ( .CLK(clk_i), .D(alu_input_b_r_20_), .Q(alu_b_i_20_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_138 ( .CLK(clk_i), .D(alu_input_b_r_21_), .Q(alu_b_i_21_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_139 ( .CLK(clk_i), .D(alu_input_b_r_22_), .Q(alu_b_i_22_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_14 ( .CLK(clk_i), .D(_0pc_q_31_0__5_), .Q(pc_q_5_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_140 ( .CLK(clk_i), .D(alu_input_b_r_23_), .Q(alu_b_i_23_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_141 ( .CLK(clk_i), .D(alu_input_b_r_24_), .Q(alu_b_i_24_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_142 ( .CLK(clk_i), .D(alu_input_b_r_25_), .Q(alu_b_i_25_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_143 ( .CLK(clk_i), .D(alu_input_b_r_26_), .Q(alu_b_i_26_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_144 ( .CLK(clk_i), .D(alu_input_b_r_27_), .Q(alu_b_i_27_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_145 ( .CLK(clk_i), .D(alu_input_b_r_28_), .Q(alu_b_i_28_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_146 ( .CLK(clk_i), .D(alu_input_b_r_29_), .Q(alu_b_i_29_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_147 ( .CLK(clk_i), .D(alu_input_b_r_30_), .Q(alu_b_i_30_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_148 ( .CLK(clk_i), .D(alu_input_b_r_31_), .Q(alu_b_i_31_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_149 ( .CLK(clk_i), .D(alu_func_r_0_), .Q(alu_op_i_0_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_15 ( .CLK(clk_i), .D(_0pc_q_31_0__6_), .Q(pc_q_6_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_150 ( .CLK(clk_i), .D(alu_func_r_1_), .Q(alu_op_i_1_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_151 ( .CLK(clk_i), .D(alu_func_r_2_), .Q(alu_op_i_2_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_152 ( .CLK(clk_i), .D(alu_func_r_3_), .Q(alu_op_i_3_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_153 ( .CLK(clk_i), .D(_0mem_addr_o_31_0__0_), .Q(\mem_addr_o[0] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_154 ( .CLK(clk_i), .D(_0mem_addr_o_31_0__1_), .Q(\mem_addr_o[1] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_155 ( .CLK(clk_i), .D(_0mem_addr_o_31_0__2_), .Q(\mem_addr_o[2] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_156 ( .CLK(clk_i), .D(_0mem_addr_o_31_0__3_), .Q(\mem_addr_o[3] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_157 ( .CLK(clk_i), .D(_0mem_addr_o_31_0__4_), .Q(\mem_addr_o[4] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_158 ( .CLK(clk_i), .D(_0mem_addr_o_31_0__5_), .Q(\mem_addr_o[5] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_159 ( .CLK(clk_i), .D(_0mem_addr_o_31_0__6_), .Q(\mem_addr_o[6] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_16 ( .CLK(clk_i), .D(_0pc_q_31_0__7_), .Q(pc_q_7_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_160 ( .CLK(clk_i), .D(_0mem_addr_o_31_0__7_), .Q(\mem_addr_o[7] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_161 ( .CLK(clk_i), .D(_0mem_addr_o_31_0__8_), .Q(\mem_addr_o[8] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_162 ( .CLK(clk_i), .D(_0mem_addr_o_31_0__9_), .Q(\mem_addr_o[9] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_163 ( .CLK(clk_i), .D(_0mem_addr_o_31_0__10_), .Q(\mem_addr_o[10] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_164 ( .CLK(clk_i), .D(_0mem_addr_o_31_0__11_), .Q(\mem_addr_o[11] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_165 ( .CLK(clk_i), .D(_0mem_addr_o_31_0__12_), .Q(\mem_addr_o[12] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_166 ( .CLK(clk_i), .D(_0mem_addr_o_31_0__13_), .Q(\mem_addr_o[13] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_167 ( .CLK(clk_i), .D(_0mem_addr_o_31_0__14_), .Q(\mem_addr_o[14] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_168 ( .CLK(clk_i), .D(_0mem_addr_o_31_0__15_), .Q(\mem_addr_o[15] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_169 ( .CLK(clk_i), .D(_0mem_addr_o_31_0__16_), .Q(\mem_addr_o[16] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_17 ( .CLK(clk_i), .D(_0pc_q_31_0__8_), .Q(pc_q_8_), .R(1'h1), .S(_abc_40298_auto_rtlil_cc_1942_NotGate_33938));
DFFSR DFFSR_170 ( .CLK(clk_i), .D(_0mem_addr_o_31_0__17_), .Q(\mem_addr_o[17] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_171 ( .CLK(clk_i), .D(_0mem_addr_o_31_0__18_), .Q(\mem_addr_o[18] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_172 ( .CLK(clk_i), .D(_0mem_addr_o_31_0__19_), .Q(\mem_addr_o[19] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_173 ( .CLK(clk_i), .D(_0mem_addr_o_31_0__20_), .Q(\mem_addr_o[20] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_174 ( .CLK(clk_i), .D(_0mem_addr_o_31_0__21_), .Q(\mem_addr_o[21] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_175 ( .CLK(clk_i), .D(_0mem_addr_o_31_0__22_), .Q(\mem_addr_o[22] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_176 ( .CLK(clk_i), .D(_0mem_addr_o_31_0__23_), .Q(\mem_addr_o[23] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_177 ( .CLK(clk_i), .D(_0mem_addr_o_31_0__24_), .Q(\mem_addr_o[24] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_178 ( .CLK(clk_i), .D(_0mem_addr_o_31_0__25_), .Q(\mem_addr_o[25] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_179 ( .CLK(clk_i), .D(_0mem_addr_o_31_0__26_), .Q(\mem_addr_o[26] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_18 ( .CLK(clk_i), .D(_0pc_q_31_0__9_), .Q(pc_q_9_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_180 ( .CLK(clk_i), .D(_0mem_addr_o_31_0__27_), .Q(\mem_addr_o[27] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_181 ( .CLK(clk_i), .D(_0mem_addr_o_31_0__28_), .Q(\mem_addr_o[28] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_182 ( .CLK(clk_i), .D(_0mem_addr_o_31_0__29_), .Q(\mem_addr_o[29] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_183 ( .CLK(clk_i), .D(_0mem_addr_o_31_0__30_), .Q(\mem_addr_o[30] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_184 ( .CLK(clk_i), .D(_0mem_addr_o_31_0__31_), .Q(\mem_addr_o[31] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_185 ( .CLK(clk_i), .D(_0mem_dat_o_31_0__0_), .Q(\mem_dat_o[0] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_186 ( .CLK(clk_i), .D(_0mem_dat_o_31_0__1_), .Q(\mem_dat_o[1] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_187 ( .CLK(clk_i), .D(_0mem_dat_o_31_0__2_), .Q(\mem_dat_o[2] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_188 ( .CLK(clk_i), .D(_0mem_dat_o_31_0__3_), .Q(\mem_dat_o[3] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_189 ( .CLK(clk_i), .D(_0mem_dat_o_31_0__4_), .Q(\mem_dat_o[4] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_19 ( .CLK(clk_i), .D(_0pc_q_31_0__10_), .Q(pc_q_10_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_190 ( .CLK(clk_i), .D(_0mem_dat_o_31_0__5_), .Q(\mem_dat_o[5] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_191 ( .CLK(clk_i), .D(_0mem_dat_o_31_0__6_), .Q(\mem_dat_o[6] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_192 ( .CLK(clk_i), .D(_0mem_dat_o_31_0__7_), .Q(\mem_dat_o[7] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_193 ( .CLK(clk_i), .D(_0mem_dat_o_31_0__8_), .Q(\mem_dat_o[8] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_194 ( .CLK(clk_i), .D(_0mem_dat_o_31_0__9_), .Q(\mem_dat_o[9] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_195 ( .CLK(clk_i), .D(_0mem_dat_o_31_0__10_), .Q(\mem_dat_o[10] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_196 ( .CLK(clk_i), .D(_0mem_dat_o_31_0__11_), .Q(\mem_dat_o[11] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_197 ( .CLK(clk_i), .D(_0mem_dat_o_31_0__12_), .Q(\mem_dat_o[12] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_198 ( .CLK(clk_i), .D(_0mem_dat_o_31_0__13_), .Q(\mem_dat_o[13] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_199 ( .CLK(clk_i), .D(_0mem_dat_o_31_0__14_), .Q(\mem_dat_o[14] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_2 ( .CLK(clk_i), .D(_abc_27663_auto_fsm_map_cc_170_map_fsm_2376_1_), .Q(state_q_1_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_20 ( .CLK(clk_i), .D(_0pc_q_31_0__11_), .Q(pc_q_11_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_200 ( .CLK(clk_i), .D(_0mem_dat_o_31_0__15_), .Q(\mem_dat_o[15] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_201 ( .CLK(clk_i), .D(_0mem_dat_o_31_0__16_), .Q(\mem_dat_o[16] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_202 ( .CLK(clk_i), .D(_0mem_dat_o_31_0__17_), .Q(\mem_dat_o[17] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_203 ( .CLK(clk_i), .D(_0mem_dat_o_31_0__18_), .Q(\mem_dat_o[18] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_204 ( .CLK(clk_i), .D(_0mem_dat_o_31_0__19_), .Q(\mem_dat_o[19] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_205 ( .CLK(clk_i), .D(_0mem_dat_o_31_0__20_), .Q(\mem_dat_o[20] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_206 ( .CLK(clk_i), .D(_0mem_dat_o_31_0__21_), .Q(\mem_dat_o[21] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_207 ( .CLK(clk_i), .D(_0mem_dat_o_31_0__22_), .Q(\mem_dat_o[22] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_208 ( .CLK(clk_i), .D(_0mem_dat_o_31_0__23_), .Q(\mem_dat_o[23] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_209 ( .CLK(clk_i), .D(_0mem_dat_o_31_0__24_), .Q(\mem_dat_o[24] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_21 ( .CLK(clk_i), .D(_0pc_q_31_0__12_), .Q(pc_q_12_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_210 ( .CLK(clk_i), .D(_0mem_dat_o_31_0__25_), .Q(\mem_dat_o[25] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_211 ( .CLK(clk_i), .D(_0mem_dat_o_31_0__26_), .Q(\mem_dat_o[26] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_212 ( .CLK(clk_i), .D(_0mem_dat_o_31_0__27_), .Q(\mem_dat_o[27] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_213 ( .CLK(clk_i), .D(_0mem_dat_o_31_0__28_), .Q(\mem_dat_o[28] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_214 ( .CLK(clk_i), .D(_0mem_dat_o_31_0__29_), .Q(\mem_dat_o[29] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_215 ( .CLK(clk_i), .D(_0mem_dat_o_31_0__30_), .Q(\mem_dat_o[30] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_216 ( .CLK(clk_i), .D(_0mem_dat_o_31_0__31_), .Q(\mem_dat_o[31] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_217 ( .CLK(clk_i), .D(_0mem_cyc_o_0_0_), .Q(mem_cyc_o), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_218 ( .CLK(clk_i), .D(_0mem_stb_o_0_0_), .Q(mem_stb_o), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_219 ( .CLK(clk_i), .D(_0mem_we_o_0_0_), .Q(mem_we_o), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_22 ( .CLK(clk_i), .D(_0pc_q_31_0__13_), .Q(pc_q_13_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_220 ( .CLK(clk_i), .D(_0mem_sel_o_3_0__0_), .Q(\mem_sel_o[0] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_221 ( .CLK(clk_i), .D(_0mem_sel_o_3_0__1_), .Q(\mem_sel_o[1] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_222 ( .CLK(clk_i), .D(_0mem_sel_o_3_0__2_), .Q(\mem_sel_o[2] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_223 ( .CLK(clk_i), .D(_0mem_sel_o_3_0__3_), .Q(\mem_sel_o[3] ), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_224 ( .CLK(clk_i), .D(_0opcode_q_31_0__0_), .Q(alu_op_r_0_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_225 ( .CLK(clk_i), .D(_0opcode_q_31_0__1_), .Q(alu_op_r_1_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_226 ( .CLK(clk_i), .D(_0opcode_q_31_0__2_), .Q(alu_op_r_2_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_227 ( .CLK(clk_i), .D(_0opcode_q_31_0__3_), .Q(alu_op_r_3_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_228 ( .CLK(clk_i), .D(_0opcode_q_31_0__4_), .Q(int32_r_4_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_229 ( .CLK(clk_i), .D(_0opcode_q_31_0__5_), .Q(int32_r_5_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_23 ( .CLK(clk_i), .D(_0pc_q_31_0__14_), .Q(pc_q_14_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_230 ( .CLK(clk_i), .D(_0opcode_q_31_0__6_), .Q(alu_op_r_4_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_231 ( .CLK(clk_i), .D(_0opcode_q_31_0__7_), .Q(alu_op_r_5_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_232 ( .CLK(clk_i), .D(_0opcode_q_31_0__8_), .Q(alu_op_r_6_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_233 ( .CLK(clk_i), .D(_0opcode_q_31_0__9_), .Q(alu_op_r_7_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_234 ( .CLK(clk_i), .D(_0opcode_q_31_0__10_), .Q(int32_r_10_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_235 ( .CLK(clk_i), .D(_0opcode_q_31_0__11_), .Q(REGFILE_SIM_reg_bank_rb_i_0_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_236 ( .CLK(clk_i), .D(_0opcode_q_31_0__12_), .Q(REGFILE_SIM_reg_bank_rb_i_1_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_237 ( .CLK(clk_i), .D(_0opcode_q_31_0__13_), .Q(REGFILE_SIM_reg_bank_rb_i_2_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_238 ( .CLK(clk_i), .D(_0opcode_q_31_0__14_), .Q(REGFILE_SIM_reg_bank_rb_i_3_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_239 ( .CLK(clk_i), .D(_0opcode_q_31_0__15_), .Q(REGFILE_SIM_reg_bank_rb_i_4_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_24 ( .CLK(clk_i), .D(_0pc_q_31_0__15_), .Q(pc_q_15_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_240 ( .CLK(clk_i), .D(_0opcode_q_31_0__16_), .Q(REGFILE_SIM_reg_bank_ra_i_0_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_241 ( .CLK(clk_i), .D(_0opcode_q_31_0__17_), .Q(REGFILE_SIM_reg_bank_ra_i_1_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_242 ( .CLK(clk_i), .D(_0opcode_q_31_0__18_), .Q(REGFILE_SIM_reg_bank_ra_i_2_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_243 ( .CLK(clk_i), .D(_0opcode_q_31_0__19_), .Q(REGFILE_SIM_reg_bank_ra_i_3_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_244 ( .CLK(clk_i), .D(_0opcode_q_31_0__20_), .Q(REGFILE_SIM_reg_bank_ra_i_4_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_245 ( .CLK(clk_i), .D(_0opcode_q_31_0__21_), .Q(opcode_q_21_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_246 ( .CLK(clk_i), .D(_0opcode_q_31_0__22_), .Q(opcode_q_22_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_247 ( .CLK(clk_i), .D(_0opcode_q_31_0__23_), .Q(opcode_q_23_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_248 ( .CLK(clk_i), .D(_0opcode_q_31_0__24_), .Q(opcode_q_24_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_249 ( .CLK(clk_i), .D(_0opcode_q_31_0__25_), .Q(opcode_q_25_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_25 ( .CLK(clk_i), .D(_0pc_q_31_0__16_), .Q(pc_q_16_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_250 ( .CLK(clk_i), .D(_0opcode_q_31_0__26_), .Q(inst_r_0_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_251 ( .CLK(clk_i), .D(_0opcode_q_31_0__27_), .Q(inst_r_1_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_252 ( .CLK(clk_i), .D(_0opcode_q_31_0__28_), .Q(inst_r_2_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_253 ( .CLK(clk_i), .D(_0opcode_q_31_0__29_), .Q(inst_r_3_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_254 ( .CLK(clk_i), .D(_0opcode_q_31_0__30_), .Q(inst_r_4_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_255 ( .CLK(clk_i), .D(_0opcode_q_31_0__31_), .Q(inst_r_5_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_256 ( .CLK(clk_i), .D(_0mem_offset_q_1_0__0_), .Q(mem_offset_q_0_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_257 ( .CLK(clk_i), .D(_0mem_offset_q_1_0__1_), .Q(mem_offset_q_1_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_258 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_0_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_259 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_1_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_26 ( .CLK(clk_i), .D(_0pc_q_31_0__17_), .Q(pc_q_17_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_260 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_2_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_261 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_3_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_262 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_4_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_263 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_5_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_264 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_6_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_265 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_7_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_266 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_8_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_267 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_9_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_268 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_10_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_269 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_11_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_27 ( .CLK(clk_i), .D(_0pc_q_31_0__18_), .Q(pc_q_18_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_270 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_12_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_271 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_13_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_272 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_14_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_273 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_15_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_274 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_16_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_275 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_17_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_276 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_18_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_277 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_19_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_278 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_20_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_279 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_21_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_28 ( .CLK(clk_i), .D(_0pc_q_31_0__19_), .Q(pc_q_19_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_280 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_22_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_281 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_23_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_282 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_24_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_283 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_25_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_284 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_26_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_285 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_27_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_286 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_28_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_287 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_29_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_288 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_30_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_289 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_31_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_29 ( .CLK(clk_i), .D(_0pc_q_31_0__20_), .Q(pc_q_20_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_290 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r3_0_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_291 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r3_1_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_292 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r3_2_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_293 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r3_3_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_294 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r3_4_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_295 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r3_5_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_296 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r3_6_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_297 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r3_7_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_298 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r3_8_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_299 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r3_9_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_3 ( .CLK(clk_i), .D(_abc_27663_auto_fsm_map_cc_170_map_fsm_2376_2_), .Q(state_q_2_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_30 ( .CLK(clk_i), .D(_0pc_q_31_0__21_), .Q(pc_q_21_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_300 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r3_10_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_301 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r3_11_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_302 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r3_12_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_303 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r3_13_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_304 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r3_14_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_305 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r3_15_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_306 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r3_16_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_307 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r3_17_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_308 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r3_18_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_309 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r3_19_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_31 ( .CLK(clk_i), .D(_0pc_q_31_0__22_), .Q(pc_q_22_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_310 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r3_20_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_311 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r3_21_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_312 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r3_22_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_313 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r3_23_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_314 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r3_24_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_315 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r3_25_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_316 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r3_26_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_317 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r3_27_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_318 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r3_28_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_319 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r3_29_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_32 ( .CLK(clk_i), .D(_0pc_q_31_0__23_), .Q(pc_q_23_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_320 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r3_30_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_321 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r3_31_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_322 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r4_0_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_323 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r4_1_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_324 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r4_2_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_325 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r4_3_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_326 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r4_4_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_327 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r4_5_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_328 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r4_6_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_329 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r4_7_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_33 ( .CLK(clk_i), .D(_0pc_q_31_0__24_), .Q(pc_q_24_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_330 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r4_8_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_331 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r4_9_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_332 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r4_10_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_333 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r4_11_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_334 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r4_12_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_335 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r4_13_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_336 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r4_14_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_337 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r4_15_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_338 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r4_16_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_339 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r4_17_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_34 ( .CLK(clk_i), .D(_0pc_q_31_0__25_), .Q(pc_q_25_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_340 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r4_18_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_341 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r4_19_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_342 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r4_20_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_343 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r4_21_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_344 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r4_22_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_345 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r4_23_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_346 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r4_24_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_347 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r4_25_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_348 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r4_26_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_349 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r4_27_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_35 ( .CLK(clk_i), .D(_0pc_q_31_0__26_), .Q(pc_q_26_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_350 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r4_28_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_351 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r4_29_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_352 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r4_30_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_353 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r4_31_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_354 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r5_0_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_355 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r5_1_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_356 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r5_2_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_357 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r5_3_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_358 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r5_4_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_359 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r5_5_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_36 ( .CLK(clk_i), .D(_0pc_q_31_0__27_), .Q(pc_q_27_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_360 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r5_6_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_361 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r5_7_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_362 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r5_8_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_363 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r5_9_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_364 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r5_10_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_365 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r5_11_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_366 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r5_12_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_367 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r5_13_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_368 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r5_14_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_369 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r5_15_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_37 ( .CLK(clk_i), .D(_0pc_q_31_0__28_), .Q(pc_q_28_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_370 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r5_16_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_371 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r5_17_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_372 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r5_18_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_373 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r5_19_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_374 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r5_20_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_375 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r5_21_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_376 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r5_22_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_377 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r5_23_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_378 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r5_24_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_379 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r5_25_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_38 ( .CLK(clk_i), .D(_0pc_q_31_0__29_), .Q(pc_q_29_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_380 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r5_26_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_381 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r5_27_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_382 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r5_28_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_383 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r5_29_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_384 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r5_30_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_385 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r5_31_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_386 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r6_0_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_387 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r6_1_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_388 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r6_2_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_389 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r6_3_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_39 ( .CLK(clk_i), .D(_0pc_q_31_0__30_), .Q(pc_q_30_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_390 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r6_4_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_391 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r6_5_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_392 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r6_6_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_393 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r6_7_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_394 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r6_8_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_395 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r6_9_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_396 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r6_10_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_397 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r6_11_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_398 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r6_12_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_399 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r6_13_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_4 ( .CLK(clk_i), .D(_abc_27663_auto_fsm_map_cc_170_map_fsm_2376_3_), .Q(state_q_3_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_40 ( .CLK(clk_i), .D(_0pc_q_31_0__31_), .Q(pc_q_31_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_400 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r6_14_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_401 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r6_15_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_402 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r6_16_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_403 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r6_17_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_404 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r6_18_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_405 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r6_19_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_406 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r6_20_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_407 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r6_21_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_408 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r6_22_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_409 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r6_23_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_41 ( .CLK(clk_i), .D(_0epc_q_31_0__0_), .Q(epc_q_0_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_410 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r6_24_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_411 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r6_25_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_412 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r6_26_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_413 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r6_27_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_414 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r6_28_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_415 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r6_29_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_416 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r6_30_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_417 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r6_31_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_418 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r7_0_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_419 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r7_1_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_42 ( .CLK(clk_i), .D(_0epc_q_31_0__1_), .Q(epc_q_1_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_420 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r7_2_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_421 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r7_3_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_422 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r7_4_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_423 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r7_5_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_424 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r7_6_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_425 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r7_7_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_426 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r7_8_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_427 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r7_9_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_428 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r7_10_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_429 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r7_11_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_43 ( .CLK(clk_i), .D(_0epc_q_31_0__2_), .Q(epc_q_2_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_430 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r7_12_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_431 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r7_13_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_432 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r7_14_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_433 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r7_15_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_434 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r7_16_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_435 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r7_17_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_436 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r7_18_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_437 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r7_19_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_438 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r7_20_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_439 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r7_21_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_44 ( .CLK(clk_i), .D(_0epc_q_31_0__3_), .Q(epc_q_3_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_440 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r7_22_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_441 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r7_23_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_442 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r7_24_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_443 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r7_25_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_444 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r7_26_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_445 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r7_27_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_446 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r7_28_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_447 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r7_29_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_448 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r7_30_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_449 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r7_31_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_45 ( .CLK(clk_i), .D(_0epc_q_31_0__4_), .Q(epc_q_4_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_450 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r8_0_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_451 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r8_1_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_452 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r8_2_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_453 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r8_3_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_454 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r8_4_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_455 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r8_5_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_456 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r8_6_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_457 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r8_7_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_458 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r8_8_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_459 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r8_9_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_46 ( .CLK(clk_i), .D(_0epc_q_31_0__5_), .Q(epc_q_5_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_460 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r8_10_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_461 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r8_11_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_462 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r8_12_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_463 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r8_13_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_464 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r8_14_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_465 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r8_15_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_466 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r8_16_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_467 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r8_17_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_468 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r8_18_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_469 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r8_19_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_47 ( .CLK(clk_i), .D(_0epc_q_31_0__6_), .Q(epc_q_6_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_470 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r8_20_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_471 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r8_21_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_472 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r8_22_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_473 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r8_23_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_474 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r8_24_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_475 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r8_25_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_476 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r8_26_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_477 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r8_27_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_478 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r8_28_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_479 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r8_29_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_48 ( .CLK(clk_i), .D(_0epc_q_31_0__7_), .Q(epc_q_7_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_480 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r8_30_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_481 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r8_31_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_482 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_0_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_483 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_1_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_484 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_2_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_485 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_3_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_486 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_4_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_487 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_5_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_488 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_6_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_489 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_7_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_49 ( .CLK(clk_i), .D(_0epc_q_31_0__8_), .Q(epc_q_8_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_490 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_8_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_491 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_9_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_492 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_10_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_493 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_11_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_494 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_12_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_495 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_13_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_496 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_14_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_497 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_15_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_498 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_16_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_499 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_17_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_5 ( .CLK(clk_i), .D(_abc_27663_auto_fsm_map_cc_170_map_fsm_2376_4_), .Q(state_q_4_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_50 ( .CLK(clk_i), .D(_0epc_q_31_0__9_), .Q(epc_q_9_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_500 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_18_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_501 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_19_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_502 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_20_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_503 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_21_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_504 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_22_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_505 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_23_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_506 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_24_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_507 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_25_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_508 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_26_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_509 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_27_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_51 ( .CLK(clk_i), .D(_0epc_q_31_0__10_), .Q(epc_q_10_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_510 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_28_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_511 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_29_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_512 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_30_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_513 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_31_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_514 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_0_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_515 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_1_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_516 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_2_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_517 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_3_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_518 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_4_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_519 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_5_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_52 ( .CLK(clk_i), .D(_0epc_q_31_0__11_), .Q(epc_q_11_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_520 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_6_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_521 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_7_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_522 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_8_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_523 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_9_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_524 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_10_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_525 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_11_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_526 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_12_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_527 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_13_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_528 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_14_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_529 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_15_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_53 ( .CLK(clk_i), .D(_0epc_q_31_0__12_), .Q(epc_q_12_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_530 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_16_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_531 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_17_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_532 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_18_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_533 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_19_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_534 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_20_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_535 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_21_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_536 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_22_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_537 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_23_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_538 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_24_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_539 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_25_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_54 ( .CLK(clk_i), .D(_0epc_q_31_0__13_), .Q(epc_q_13_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_540 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_26_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_541 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_27_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_542 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_28_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_543 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_29_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_544 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_30_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_545 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_31_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_546 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r10_0_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_547 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r10_1_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_548 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r10_2_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_549 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r10_3_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_55 ( .CLK(clk_i), .D(_0epc_q_31_0__14_), .Q(epc_q_14_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_550 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r10_4_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_551 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r10_5_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_552 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r10_6_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_553 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r10_7_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_554 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r10_8_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_555 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r10_9_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_556 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r10_10_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_557 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r10_11_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_558 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r10_12_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_559 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r10_13_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_56 ( .CLK(clk_i), .D(_0epc_q_31_0__15_), .Q(epc_q_15_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_560 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r10_14_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_561 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r10_15_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_562 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r10_16_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_563 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r10_17_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_564 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r10_18_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_565 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r10_19_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_566 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r10_20_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_567 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r10_21_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_568 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r10_22_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_569 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r10_23_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_57 ( .CLK(clk_i), .D(_0epc_q_31_0__16_), .Q(epc_q_16_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_570 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r10_24_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_571 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r10_25_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_572 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r10_26_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_573 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r10_27_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_574 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r10_28_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_575 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r10_29_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_576 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r10_30_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_577 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r10_31_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_578 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r11_0_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_579 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r11_1_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_58 ( .CLK(clk_i), .D(_0epc_q_31_0__17_), .Q(epc_q_17_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_580 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r11_2_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_581 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r11_3_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_582 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r11_4_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_583 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r11_5_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_584 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r11_6_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_585 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r11_7_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_586 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r11_8_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_587 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r11_9_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_588 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r11_10_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_589 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r11_11_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_59 ( .CLK(clk_i), .D(_0epc_q_31_0__18_), .Q(epc_q_18_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_590 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r11_12_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_591 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r11_13_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_592 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r11_14_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_593 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r11_15_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_594 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r11_16_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_595 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r11_17_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_596 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r11_18_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_597 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r11_19_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_598 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r11_20_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_599 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r11_21_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_6 ( .CLK(clk_i), .D(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2420), .Q(state_q_5_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_60 ( .CLK(clk_i), .D(_0epc_q_31_0__19_), .Q(epc_q_19_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_600 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r11_22_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_601 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r11_23_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_602 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r11_24_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_603 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r11_25_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_604 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r11_26_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_605 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r11_27_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_606 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r11_28_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_607 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r11_29_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_608 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r11_30_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_609 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r11_31_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_61 ( .CLK(clk_i), .D(_0epc_q_31_0__20_), .Q(epc_q_20_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_610 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r12_0_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_611 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r12_1_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_612 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r12_2_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_613 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r12_3_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_614 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r12_4_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_615 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r12_5_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_616 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r12_6_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_617 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r12_7_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_618 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r12_8_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_619 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r12_9_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_62 ( .CLK(clk_i), .D(_0epc_q_31_0__21_), .Q(epc_q_21_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_620 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r12_10_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_621 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r12_11_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_622 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r12_12_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_623 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r12_13_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_624 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r12_14_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_625 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r12_15_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_626 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r12_16_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_627 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r12_17_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_628 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r12_18_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_629 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r12_19_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_63 ( .CLK(clk_i), .D(_0epc_q_31_0__22_), .Q(epc_q_22_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_630 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r12_20_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_631 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r12_21_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_632 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r12_22_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_633 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r12_23_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_634 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r12_24_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_635 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r12_25_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_636 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r12_26_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_637 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r12_27_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_638 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r12_28_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_639 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r12_29_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_64 ( .CLK(clk_i), .D(_0epc_q_31_0__23_), .Q(epc_q_23_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_640 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r12_30_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_641 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r12_31_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_642 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r13_0_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_643 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r13_1_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_644 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r13_2_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_645 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r13_3_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_646 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r13_4_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_647 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r13_5_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_648 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r13_6_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_649 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r13_7_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_65 ( .CLK(clk_i), .D(_0epc_q_31_0__24_), .Q(epc_q_24_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_650 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r13_8_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_651 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r13_9_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_652 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r13_10_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_653 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r13_11_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_654 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r13_12_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_655 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r13_13_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_656 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r13_14_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_657 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r13_15_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_658 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r13_16_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_659 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r13_17_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_66 ( .CLK(clk_i), .D(_0epc_q_31_0__25_), .Q(epc_q_25_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_660 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r13_18_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_661 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r13_19_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_662 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r13_20_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_663 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r13_21_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_664 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r13_22_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_665 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r13_23_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_666 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r13_24_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_667 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r13_25_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_668 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r13_26_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_669 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r13_27_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_67 ( .CLK(clk_i), .D(_0epc_q_31_0__26_), .Q(epc_q_26_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_670 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r13_28_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_671 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r13_29_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_672 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r13_30_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_673 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r13_31_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_674 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r14_0_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_675 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r14_1_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_676 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r14_2_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_677 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r14_3_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_678 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r14_4_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_679 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r14_5_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_68 ( .CLK(clk_i), .D(_0epc_q_31_0__27_), .Q(epc_q_27_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_680 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r14_6_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_681 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r14_7_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_682 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r14_8_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_683 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r14_9_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_684 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r14_10_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_685 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r14_11_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_686 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r14_12_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_687 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r14_13_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_688 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r14_14_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_689 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r14_15_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_69 ( .CLK(clk_i), .D(_0epc_q_31_0__28_), .Q(epc_q_28_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_690 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r14_16_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_691 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r14_17_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_692 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r14_18_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_693 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r14_19_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_694 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r14_20_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_695 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r14_21_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_696 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r14_22_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_697 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r14_23_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_698 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r14_24_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_699 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r14_25_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_7 ( .CLK(clk_i), .D(inst_trap_w), .Q(break_o), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_70 ( .CLK(clk_i), .D(_0epc_q_31_0__29_), .Q(epc_q_29_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_700 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r14_26_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_701 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r14_27_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_702 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r14_28_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_703 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r14_29_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_704 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r14_30_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_705 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r14_31_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_706 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r15_0_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_707 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r15_1_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_708 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r15_2_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_709 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r15_3_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_71 ( .CLK(clk_i), .D(_0epc_q_31_0__30_), .Q(epc_q_30_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_710 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r15_4_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_711 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r15_5_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_712 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r15_6_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_713 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r15_7_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_714 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r15_8_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_715 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r15_9_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_716 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r15_10_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_717 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r15_11_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_718 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r15_12_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_719 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r15_13_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_72 ( .CLK(clk_i), .D(_0epc_q_31_0__31_), .Q(epc_q_31_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_720 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r15_14_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_721 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r15_15_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_722 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r15_16_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_723 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r15_17_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_724 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r15_18_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_725 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r15_19_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_726 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r15_20_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_727 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r15_21_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_728 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r15_22_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_729 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r15_23_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_73 ( .CLK(clk_i), .D(_0sr_q_31_0__2_), .Q(sr_q_2_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_730 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r15_24_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_731 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r15_25_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_732 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r15_26_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_733 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r15_27_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_734 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r15_28_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_735 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r15_29_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_736 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r15_30_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_737 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r15_31_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_738 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r16_0_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_739 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r16_1_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_74 ( .CLK(clk_i), .D(_0sr_q_31_0__9_), .Q(sr_q_9_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_740 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r16_2_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_741 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r16_3_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_742 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r16_4_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_743 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r16_5_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_744 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r16_6_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_745 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r16_7_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_746 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r16_8_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_747 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r16_9_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_748 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r16_10_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_749 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r16_11_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_75 ( .CLK(clk_i), .D(_0sr_q_31_0__10_), .Q(alu_c_i), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_750 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r16_12_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_751 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r16_13_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_752 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r16_14_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_753 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r16_15_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_754 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r16_16_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_755 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r16_17_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_756 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r16_18_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_757 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r16_19_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_758 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r16_20_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_759 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r16_21_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_76 ( .CLK(clk_i), .D(_0esr_q_31_0__2_), .Q(esr_q_2_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_760 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r16_22_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_761 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r16_23_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_762 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r16_24_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_763 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r16_25_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_764 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r16_26_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_765 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r16_27_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_766 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r16_28_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_767 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r16_29_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_768 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r16_30_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_769 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r16_31_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_77 ( .CLK(clk_i), .D(_0esr_q_31_0__9_), .Q(esr_q_9_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_770 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r17_0_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_771 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r17_1_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_772 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r17_2_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_773 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r17_3_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_774 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r17_4_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_775 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r17_5_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_776 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r17_6_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_777 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r17_7_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_778 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r17_8_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_779 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r17_9_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_78 ( .CLK(clk_i), .D(_0esr_q_31_0__10_), .Q(esr_q_10_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_780 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r17_10_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_781 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r17_11_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_782 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r17_12_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_783 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r17_13_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_784 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r17_14_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_785 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r17_15_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_786 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r17_16_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_787 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r17_17_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_788 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r17_18_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_789 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r17_19_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_79 ( .CLK(clk_i), .D(_0nmi_q_0_0_), .Q(nmi_q), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_790 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r17_20_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_791 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r17_21_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_792 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r17_22_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_793 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r17_23_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_794 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r17_24_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_795 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r17_25_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_796 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r17_26_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_797 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r17_27_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_798 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r17_28_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_799 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r17_29_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_8 ( .CLK(clk_i), .D(_0fault_o_0_0_), .Q(fault_o), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_80 ( .CLK(clk_i), .D(_0ex_rd_q_4_0__0_), .Q(REGFILE_SIM_reg_bank_rd_i_0_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_800 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r17_30_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_801 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r17_31_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_802 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r18_0_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_803 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r18_1_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_804 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r18_2_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_805 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r18_3_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_806 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r18_4_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_807 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r18_5_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_808 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r18_6_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_809 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r18_7_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_81 ( .CLK(clk_i), .D(_0ex_rd_q_4_0__1_), .Q(REGFILE_SIM_reg_bank_rd_i_1_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_810 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r18_8_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_811 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r18_9_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_812 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r18_10_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_813 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r18_11_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_814 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r18_12_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_815 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r18_13_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_816 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r18_14_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_817 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r18_15_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_818 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r18_16_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_819 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r18_17_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_82 ( .CLK(clk_i), .D(_0ex_rd_q_4_0__2_), .Q(REGFILE_SIM_reg_bank_rd_i_2_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_820 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r18_18_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_821 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r18_19_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_822 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r18_20_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_823 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r18_21_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_824 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r18_22_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_825 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r18_23_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_826 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r18_24_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_827 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r18_25_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_828 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r18_26_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_829 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r18_27_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_83 ( .CLK(clk_i), .D(_0ex_rd_q_4_0__3_), .Q(REGFILE_SIM_reg_bank_rd_i_3_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_830 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r18_28_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_831 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r18_29_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_832 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r18_30_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_833 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r18_31_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_834 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r19_0_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_835 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r19_1_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_836 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r19_2_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_837 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r19_3_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_838 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r19_4_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_839 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r19_5_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_84 ( .CLK(clk_i), .D(_0ex_rd_q_4_0__4_), .Q(REGFILE_SIM_reg_bank_rd_i_4_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_840 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r19_6_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_841 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r19_7_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_842 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r19_8_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_843 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r19_9_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_844 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r19_10_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_845 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r19_11_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_846 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r19_12_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_847 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r19_13_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_848 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r19_14_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_849 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r19_15_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_85 ( .CLK(clk_i), .D(alu_input_a_r_0_), .Q(alu_a_i_0_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_850 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r19_16_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_851 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r19_17_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_852 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r19_18_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_853 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r19_19_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_854 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r19_20_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_855 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r19_21_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_856 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r19_22_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_857 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r19_23_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_858 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r19_24_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_859 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r19_25_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_86 ( .CLK(clk_i), .D(alu_input_a_r_1_), .Q(alu_a_i_1_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_860 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r19_26_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_861 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r19_27_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_862 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r19_28_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_863 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r19_29_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_864 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r19_30_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_865 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r19_31_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_866 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r20_0_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_867 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r20_1_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_868 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r20_2_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_869 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r20_3_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_87 ( .CLK(clk_i), .D(alu_input_a_r_2_), .Q(alu_a_i_2_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_870 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r20_4_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_871 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r20_5_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_872 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r20_6_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_873 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r20_7_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_874 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r20_8_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_875 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r20_9_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_876 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r20_10_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_877 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r20_11_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_878 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r20_12_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_879 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r20_13_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_88 ( .CLK(clk_i), .D(alu_input_a_r_3_), .Q(alu_a_i_3_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_880 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r20_14_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_881 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r20_15_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_882 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r20_16_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_883 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r20_17_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_884 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r20_18_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_885 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r20_19_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_886 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r20_20_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_887 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r20_21_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_888 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r20_22_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_889 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r20_23_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_89 ( .CLK(clk_i), .D(alu_input_a_r_4_), .Q(alu_a_i_4_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_890 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r20_24_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_891 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r20_25_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_892 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r20_26_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_893 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r20_27_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_894 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r20_28_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_895 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r20_29_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_896 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r20_30_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_897 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r20_31_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_898 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r21_0_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_899 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r21_1_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_9 ( .CLK(clk_i), .D(_0pc_q_31_0__0_), .Q(next_pc_r_0_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_90 ( .CLK(clk_i), .D(alu_input_a_r_5_), .Q(alu_a_i_5_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_900 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r21_2_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_901 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r21_3_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_902 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r21_4_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_903 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r21_5_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_904 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r21_6_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_905 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r21_7_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_906 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r21_8_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_907 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r21_9_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_908 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r21_10_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_909 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r21_11_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_91 ( .CLK(clk_i), .D(alu_input_a_r_6_), .Q(alu_a_i_6_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_910 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r21_12_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_911 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r21_13_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_912 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r21_14_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_913 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r21_15_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_914 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r21_16_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_915 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r21_17_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_916 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r21_18_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_917 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r21_19_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_918 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r21_20_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_919 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r21_21_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_92 ( .CLK(clk_i), .D(alu_input_a_r_7_), .Q(alu_a_i_7_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_920 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r21_22_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_921 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r21_23_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_922 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r21_24_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_923 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r21_25_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_924 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r21_26_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_925 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r21_27_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_926 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r21_28_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_927 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r21_29_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_928 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r21_30_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_929 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r21_31_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_93 ( .CLK(clk_i), .D(alu_input_a_r_8_), .Q(alu_a_i_8_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_930 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r22_0_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_931 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r22_1_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_932 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r22_2_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_933 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r22_3_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_934 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r22_4_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_935 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r22_5_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_936 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r22_6_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_937 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r22_7_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_938 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r22_8_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_939 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r22_9_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_94 ( .CLK(clk_i), .D(alu_input_a_r_9_), .Q(alu_a_i_9_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_940 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r22_10_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_941 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r22_11_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_942 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r22_12_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_943 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r22_13_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_944 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r22_14_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_945 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r22_15_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_946 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r22_16_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_947 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r22_17_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_948 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r22_18_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_949 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r22_19_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_95 ( .CLK(clk_i), .D(alu_input_a_r_10_), .Q(alu_a_i_10_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_950 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r22_20_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_951 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r22_21_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_952 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r22_22_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_953 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r22_23_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_954 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r22_24_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_955 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r22_25_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_956 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r22_26_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_957 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r22_27_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_958 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r22_28_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_959 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r22_29_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_96 ( .CLK(clk_i), .D(alu_input_a_r_11_), .Q(alu_a_i_11_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_960 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r22_30_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_961 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r22_31_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_962 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r23_0_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_963 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r23_1_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_964 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r23_2_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_965 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r23_3_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_966 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r23_4_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_967 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r23_5_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_968 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r23_6_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_969 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r23_7_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_97 ( .CLK(clk_i), .D(alu_input_a_r_12_), .Q(alu_a_i_12_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_970 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r23_8_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_971 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r23_9_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_972 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r23_10_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_973 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r23_11_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_974 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r23_12_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_975 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r23_13_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_976 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r23_14_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_977 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r23_15_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_978 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r23_16_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_979 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r23_17_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_98 ( .CLK(clk_i), .D(alu_input_a_r_13_), .Q(alu_a_i_13_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_980 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r23_18_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_981 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r23_19_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_982 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r23_20_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_983 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r23_21_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_984 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r23_22_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_985 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r23_23_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_986 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r23_24_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_987 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r23_25_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_988 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r23_26_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_989 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r23_27_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_99 ( .CLK(clk_i), .D(alu_input_a_r_14_), .Q(alu_a_i_14_), .R(_abc_40298_auto_rtlil_cc_1942_NotGate_33938), .S(1'h1));
DFFSR DFFSR_990 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r23_28_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_991 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r23_29_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_992 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r23_30_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_993 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r23_31_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_994 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r24_0_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_995 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r24_1_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_996 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r24_2_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_997 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r24_3_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_998 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r24_4_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
DFFSR DFFSR_999 ( .CLK(clk_i), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r24_5_), .R(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954), .S(1'h1));
INVX1 INVX1_1 ( .A(_abc_40298_new_n617_), .Y(_abc_40298_new_n618_));
INVX1 INVX1_10 ( .A(state_q_5_), .Y(_abc_40298_new_n635_));
INVX1 INVX1_100 ( .A(_abc_40298_new_n940_), .Y(_abc_40298_new_n941_));
INVX1 INVX1_1000 ( .A(REGFILE_SIM_reg_bank_reg_r14_8_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3281_));
INVX1 INVX1_1001 ( .A(REGFILE_SIM_reg_bank_reg_r14_9_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3283_));
INVX1 INVX1_1002 ( .A(REGFILE_SIM_reg_bank_reg_r14_10_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3285_));
INVX1 INVX1_1003 ( .A(REGFILE_SIM_reg_bank_reg_r14_11_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3287_));
INVX1 INVX1_1004 ( .A(REGFILE_SIM_reg_bank_reg_r14_12_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3289_));
INVX1 INVX1_1005 ( .A(REGFILE_SIM_reg_bank_reg_r14_13_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3291_));
INVX1 INVX1_1006 ( .A(REGFILE_SIM_reg_bank_reg_r14_14_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3293_));
INVX1 INVX1_1007 ( .A(REGFILE_SIM_reg_bank_reg_r14_15_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3295_));
INVX1 INVX1_1008 ( .A(REGFILE_SIM_reg_bank_reg_r14_16_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3297_));
INVX1 INVX1_1009 ( .A(REGFILE_SIM_reg_bank_reg_r14_17_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3299_));
INVX1 INVX1_101 ( .A(_abc_40298_new_n937_), .Y(_abc_40298_new_n943_));
INVX1 INVX1_1010 ( .A(REGFILE_SIM_reg_bank_reg_r14_18_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3301_));
INVX1 INVX1_1011 ( .A(REGFILE_SIM_reg_bank_reg_r14_19_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3303_));
INVX1 INVX1_1012 ( .A(REGFILE_SIM_reg_bank_reg_r14_20_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3305_));
INVX1 INVX1_1013 ( .A(REGFILE_SIM_reg_bank_reg_r14_21_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3307_));
INVX1 INVX1_1014 ( .A(REGFILE_SIM_reg_bank_reg_r14_22_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3309_));
INVX1 INVX1_1015 ( .A(REGFILE_SIM_reg_bank_reg_r14_23_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3311_));
INVX1 INVX1_1016 ( .A(REGFILE_SIM_reg_bank_reg_r14_24_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3313_));
INVX1 INVX1_1017 ( .A(REGFILE_SIM_reg_bank_reg_r14_25_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3315_));
INVX1 INVX1_1018 ( .A(REGFILE_SIM_reg_bank_reg_r14_26_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3317_));
INVX1 INVX1_1019 ( .A(REGFILE_SIM_reg_bank_reg_r14_27_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3319_));
INVX1 INVX1_102 ( .A(opcode_q_22_), .Y(_abc_40298_new_n944_));
INVX1 INVX1_1020 ( .A(REGFILE_SIM_reg_bank_reg_r14_28_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3321_));
INVX1 INVX1_1021 ( .A(REGFILE_SIM_reg_bank_reg_r14_29_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3323_));
INVX1 INVX1_1022 ( .A(REGFILE_SIM_reg_bank_reg_r14_30_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3325_));
INVX1 INVX1_1023 ( .A(REGFILE_SIM_reg_bank_reg_r14_31_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3327_));
INVX1 INVX1_1024 ( .A(REGFILE_SIM_reg_bank_reg_r13_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3329_));
INVX1 INVX1_1025 ( .A(REGFILE_SIM_reg_bank_reg_r13_1_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3332_));
INVX1 INVX1_1026 ( .A(REGFILE_SIM_reg_bank_reg_r13_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3334_));
INVX1 INVX1_1027 ( .A(REGFILE_SIM_reg_bank_reg_r13_3_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3336_));
INVX1 INVX1_1028 ( .A(REGFILE_SIM_reg_bank_reg_r13_4_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3338_));
INVX1 INVX1_1029 ( .A(REGFILE_SIM_reg_bank_reg_r13_5_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3340_));
INVX1 INVX1_103 ( .A(opcode_q_21_), .Y(_abc_40298_new_n949_));
INVX1 INVX1_1030 ( .A(REGFILE_SIM_reg_bank_reg_r13_6_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3342_));
INVX1 INVX1_1031 ( .A(REGFILE_SIM_reg_bank_reg_r13_7_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3344_));
INVX1 INVX1_1032 ( .A(REGFILE_SIM_reg_bank_reg_r13_8_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3346_));
INVX1 INVX1_1033 ( .A(REGFILE_SIM_reg_bank_reg_r13_9_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3348_));
INVX1 INVX1_1034 ( .A(REGFILE_SIM_reg_bank_reg_r13_10_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3350_));
INVX1 INVX1_1035 ( .A(REGFILE_SIM_reg_bank_reg_r13_11_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3352_));
INVX1 INVX1_1036 ( .A(REGFILE_SIM_reg_bank_reg_r13_12_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3354_));
INVX1 INVX1_1037 ( .A(REGFILE_SIM_reg_bank_reg_r13_13_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3356_));
INVX1 INVX1_1038 ( .A(REGFILE_SIM_reg_bank_reg_r13_14_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3358_));
INVX1 INVX1_1039 ( .A(REGFILE_SIM_reg_bank_reg_r13_15_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3360_));
INVX1 INVX1_104 ( .A(_abc_40298_new_n955_), .Y(_abc_40298_new_n956_));
INVX1 INVX1_1040 ( .A(REGFILE_SIM_reg_bank_reg_r13_16_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3362_));
INVX1 INVX1_1041 ( .A(REGFILE_SIM_reg_bank_reg_r13_17_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3364_));
INVX1 INVX1_1042 ( .A(REGFILE_SIM_reg_bank_reg_r13_18_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3366_));
INVX1 INVX1_1043 ( .A(REGFILE_SIM_reg_bank_reg_r13_19_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3368_));
INVX1 INVX1_1044 ( .A(REGFILE_SIM_reg_bank_reg_r13_20_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3370_));
INVX1 INVX1_1045 ( .A(REGFILE_SIM_reg_bank_reg_r13_21_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3372_));
INVX1 INVX1_1046 ( .A(REGFILE_SIM_reg_bank_reg_r13_22_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3374_));
INVX1 INVX1_1047 ( .A(REGFILE_SIM_reg_bank_reg_r13_23_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3376_));
INVX1 INVX1_1048 ( .A(REGFILE_SIM_reg_bank_reg_r13_24_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3378_));
INVX1 INVX1_1049 ( .A(REGFILE_SIM_reg_bank_reg_r13_25_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3380_));
INVX1 INVX1_105 ( .A(_abc_40298_new_n957_), .Y(_abc_40298_new_n958_));
INVX1 INVX1_1050 ( .A(REGFILE_SIM_reg_bank_reg_r13_26_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3382_));
INVX1 INVX1_1051 ( .A(REGFILE_SIM_reg_bank_reg_r13_27_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3384_));
INVX1 INVX1_1052 ( .A(REGFILE_SIM_reg_bank_reg_r13_28_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3386_));
INVX1 INVX1_1053 ( .A(REGFILE_SIM_reg_bank_reg_r13_29_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3388_));
INVX1 INVX1_1054 ( .A(REGFILE_SIM_reg_bank_reg_r13_30_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3390_));
INVX1 INVX1_1055 ( .A(REGFILE_SIM_reg_bank_reg_r13_31_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3392_));
INVX1 INVX1_1056 ( .A(REGFILE_SIM_reg_bank_reg_r12_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3394_));
INVX1 INVX1_1057 ( .A(REGFILE_SIM_reg_bank_reg_r12_1_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3398_));
INVX1 INVX1_1058 ( .A(REGFILE_SIM_reg_bank_reg_r12_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3400_));
INVX1 INVX1_1059 ( .A(REGFILE_SIM_reg_bank_reg_r12_3_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3402_));
INVX1 INVX1_106 ( .A(_abc_40298_new_n959_), .Y(_abc_40298_new_n960_));
INVX1 INVX1_1060 ( .A(REGFILE_SIM_reg_bank_reg_r12_4_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3404_));
INVX1 INVX1_1061 ( .A(REGFILE_SIM_reg_bank_reg_r12_5_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3406_));
INVX1 INVX1_1062 ( .A(REGFILE_SIM_reg_bank_reg_r12_6_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3408_));
INVX1 INVX1_1063 ( .A(REGFILE_SIM_reg_bank_reg_r12_7_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3410_));
INVX1 INVX1_1064 ( .A(REGFILE_SIM_reg_bank_reg_r12_8_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3412_));
INVX1 INVX1_1065 ( .A(REGFILE_SIM_reg_bank_reg_r12_9_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3414_));
INVX1 INVX1_1066 ( .A(REGFILE_SIM_reg_bank_reg_r12_10_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3416_));
INVX1 INVX1_1067 ( .A(REGFILE_SIM_reg_bank_reg_r12_11_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3418_));
INVX1 INVX1_1068 ( .A(REGFILE_SIM_reg_bank_reg_r12_12_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3420_));
INVX1 INVX1_1069 ( .A(REGFILE_SIM_reg_bank_reg_r12_13_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3422_));
INVX1 INVX1_107 ( .A(_abc_40298_new_n969_), .Y(_abc_40298_new_n970_));
INVX1 INVX1_1070 ( .A(REGFILE_SIM_reg_bank_reg_r12_14_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3424_));
INVX1 INVX1_1071 ( .A(REGFILE_SIM_reg_bank_reg_r12_15_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3426_));
INVX1 INVX1_1072 ( .A(REGFILE_SIM_reg_bank_reg_r12_16_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3428_));
INVX1 INVX1_1073 ( .A(REGFILE_SIM_reg_bank_reg_r12_17_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3430_));
INVX1 INVX1_1074 ( .A(REGFILE_SIM_reg_bank_reg_r12_18_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3432_));
INVX1 INVX1_1075 ( .A(REGFILE_SIM_reg_bank_reg_r12_19_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3434_));
INVX1 INVX1_1076 ( .A(REGFILE_SIM_reg_bank_reg_r12_20_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3436_));
INVX1 INVX1_1077 ( .A(REGFILE_SIM_reg_bank_reg_r12_21_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3438_));
INVX1 INVX1_1078 ( .A(REGFILE_SIM_reg_bank_reg_r12_22_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3440_));
INVX1 INVX1_1079 ( .A(REGFILE_SIM_reg_bank_reg_r12_23_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3442_));
INVX1 INVX1_108 ( .A(alu_op_r_5_), .Y(_abc_40298_new_n973_));
INVX1 INVX1_1080 ( .A(REGFILE_SIM_reg_bank_reg_r12_24_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3444_));
INVX1 INVX1_1081 ( .A(REGFILE_SIM_reg_bank_reg_r12_25_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3446_));
INVX1 INVX1_1082 ( .A(REGFILE_SIM_reg_bank_reg_r12_26_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3448_));
INVX1 INVX1_1083 ( .A(REGFILE_SIM_reg_bank_reg_r12_27_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3450_));
INVX1 INVX1_1084 ( .A(REGFILE_SIM_reg_bank_reg_r12_28_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3452_));
INVX1 INVX1_1085 ( .A(REGFILE_SIM_reg_bank_reg_r12_29_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3454_));
INVX1 INVX1_1086 ( .A(REGFILE_SIM_reg_bank_reg_r12_30_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3456_));
INVX1 INVX1_1087 ( .A(REGFILE_SIM_reg_bank_reg_r12_31_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3458_));
INVX1 INVX1_1088 ( .A(REGFILE_SIM_reg_bank_reg_r11_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3460_));
INVX1 INVX1_1089 ( .A(REGFILE_SIM_reg_bank_reg_r11_1_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3463_));
INVX1 INVX1_109 ( .A(_abc_40298_new_n974_), .Y(_abc_40298_new_n975_));
INVX1 INVX1_1090 ( .A(REGFILE_SIM_reg_bank_reg_r11_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3465_));
INVX1 INVX1_1091 ( .A(REGFILE_SIM_reg_bank_reg_r11_3_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3467_));
INVX1 INVX1_1092 ( .A(REGFILE_SIM_reg_bank_reg_r11_4_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3469_));
INVX1 INVX1_1093 ( .A(REGFILE_SIM_reg_bank_reg_r11_5_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3471_));
INVX1 INVX1_1094 ( .A(REGFILE_SIM_reg_bank_reg_r11_6_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3473_));
INVX1 INVX1_1095 ( .A(REGFILE_SIM_reg_bank_reg_r11_7_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3475_));
INVX1 INVX1_1096 ( .A(REGFILE_SIM_reg_bank_reg_r11_8_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3477_));
INVX1 INVX1_1097 ( .A(REGFILE_SIM_reg_bank_reg_r11_9_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3479_));
INVX1 INVX1_1098 ( .A(REGFILE_SIM_reg_bank_reg_r11_10_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3481_));
INVX1 INVX1_1099 ( .A(REGFILE_SIM_reg_bank_reg_r11_11_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3483_));
INVX1 INVX1_11 ( .A(inst_r_4_), .Y(_abc_40298_new_n637_));
INVX1 INVX1_110 ( .A(_abc_40298_new_n646_), .Y(_abc_40298_new_n978_));
INVX1 INVX1_1100 ( .A(REGFILE_SIM_reg_bank_reg_r11_12_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3485_));
INVX1 INVX1_1101 ( .A(REGFILE_SIM_reg_bank_reg_r11_13_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3487_));
INVX1 INVX1_1102 ( .A(REGFILE_SIM_reg_bank_reg_r11_14_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3489_));
INVX1 INVX1_1103 ( .A(REGFILE_SIM_reg_bank_reg_r11_15_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3491_));
INVX1 INVX1_1104 ( .A(REGFILE_SIM_reg_bank_reg_r11_16_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3493_));
INVX1 INVX1_1105 ( .A(REGFILE_SIM_reg_bank_reg_r11_17_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3495_));
INVX1 INVX1_1106 ( .A(REGFILE_SIM_reg_bank_reg_r11_18_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3497_));
INVX1 INVX1_1107 ( .A(REGFILE_SIM_reg_bank_reg_r11_19_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3499_));
INVX1 INVX1_1108 ( .A(REGFILE_SIM_reg_bank_reg_r11_20_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3501_));
INVX1 INVX1_1109 ( .A(REGFILE_SIM_reg_bank_reg_r11_21_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3503_));
INVX1 INVX1_111 ( .A(_abc_40298_new_n981_), .Y(_abc_40298_new_n982_));
INVX1 INVX1_1110 ( .A(REGFILE_SIM_reg_bank_reg_r11_22_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3505_));
INVX1 INVX1_1111 ( .A(REGFILE_SIM_reg_bank_reg_r11_23_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3507_));
INVX1 INVX1_1112 ( .A(REGFILE_SIM_reg_bank_reg_r11_24_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3509_));
INVX1 INVX1_1113 ( .A(REGFILE_SIM_reg_bank_reg_r11_25_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3511_));
INVX1 INVX1_1114 ( .A(REGFILE_SIM_reg_bank_reg_r11_26_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3513_));
INVX1 INVX1_1115 ( .A(REGFILE_SIM_reg_bank_reg_r11_27_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3515_));
INVX1 INVX1_1116 ( .A(REGFILE_SIM_reg_bank_reg_r11_28_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3517_));
INVX1 INVX1_1117 ( .A(REGFILE_SIM_reg_bank_reg_r11_29_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3519_));
INVX1 INVX1_1118 ( .A(REGFILE_SIM_reg_bank_reg_r11_30_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3521_));
INVX1 INVX1_1119 ( .A(REGFILE_SIM_reg_bank_reg_r11_31_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3523_));
INVX1 INVX1_112 ( .A(_abc_40298_new_n622_), .Y(_abc_40298_new_n983_));
INVX1 INVX1_1120 ( .A(REGFILE_SIM_reg_bank_reg_r10_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3525_));
INVX1 INVX1_1121 ( .A(REGFILE_SIM_reg_bank_reg_r10_1_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3528_));
INVX1 INVX1_1122 ( .A(REGFILE_SIM_reg_bank_reg_r10_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3530_));
INVX1 INVX1_1123 ( .A(REGFILE_SIM_reg_bank_reg_r10_3_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3532_));
INVX1 INVX1_1124 ( .A(REGFILE_SIM_reg_bank_reg_r10_4_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3534_));
INVX1 INVX1_1125 ( .A(REGFILE_SIM_reg_bank_reg_r10_5_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3536_));
INVX1 INVX1_1126 ( .A(REGFILE_SIM_reg_bank_reg_r10_6_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3538_));
INVX1 INVX1_1127 ( .A(REGFILE_SIM_reg_bank_reg_r10_7_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3540_));
INVX1 INVX1_1128 ( .A(REGFILE_SIM_reg_bank_reg_r10_8_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3542_));
INVX1 INVX1_1129 ( .A(REGFILE_SIM_reg_bank_reg_r10_9_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3544_));
INVX1 INVX1_113 ( .A(_abc_40298_new_n984_), .Y(_abc_40298_new_n985_));
INVX1 INVX1_1130 ( .A(REGFILE_SIM_reg_bank_reg_r10_10_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3546_));
INVX1 INVX1_1131 ( .A(REGFILE_SIM_reg_bank_reg_r10_11_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3548_));
INVX1 INVX1_1132 ( .A(REGFILE_SIM_reg_bank_reg_r10_12_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3550_));
INVX1 INVX1_1133 ( .A(REGFILE_SIM_reg_bank_reg_r10_13_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3552_));
INVX1 INVX1_1134 ( .A(REGFILE_SIM_reg_bank_reg_r10_14_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3554_));
INVX1 INVX1_1135 ( .A(REGFILE_SIM_reg_bank_reg_r10_15_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3556_));
INVX1 INVX1_1136 ( .A(REGFILE_SIM_reg_bank_reg_r10_16_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3558_));
INVX1 INVX1_1137 ( .A(REGFILE_SIM_reg_bank_reg_r10_17_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3560_));
INVX1 INVX1_1138 ( .A(REGFILE_SIM_reg_bank_reg_r10_18_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3562_));
INVX1 INVX1_1139 ( .A(REGFILE_SIM_reg_bank_reg_r10_19_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3564_));
INVX1 INVX1_114 ( .A(_abc_40298_new_n934_), .Y(_abc_40298_new_n987_));
INVX1 INVX1_1140 ( .A(REGFILE_SIM_reg_bank_reg_r10_20_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3566_));
INVX1 INVX1_1141 ( .A(REGFILE_SIM_reg_bank_reg_r10_21_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3568_));
INVX1 INVX1_1142 ( .A(REGFILE_SIM_reg_bank_reg_r10_22_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3570_));
INVX1 INVX1_1143 ( .A(REGFILE_SIM_reg_bank_reg_r10_23_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3572_));
INVX1 INVX1_1144 ( .A(REGFILE_SIM_reg_bank_reg_r10_24_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3574_));
INVX1 INVX1_1145 ( .A(REGFILE_SIM_reg_bank_reg_r10_25_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3576_));
INVX1 INVX1_1146 ( .A(REGFILE_SIM_reg_bank_reg_r10_26_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3578_));
INVX1 INVX1_1147 ( .A(REGFILE_SIM_reg_bank_reg_r10_27_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3580_));
INVX1 INVX1_1148 ( .A(REGFILE_SIM_reg_bank_reg_r10_28_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3582_));
INVX1 INVX1_1149 ( .A(REGFILE_SIM_reg_bank_reg_r10_29_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3584_));
INVX1 INVX1_115 ( .A(_abc_40298_new_n992_), .Y(_abc_40298_new_n993_));
INVX1 INVX1_1150 ( .A(REGFILE_SIM_reg_bank_reg_r10_30_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3586_));
INVX1 INVX1_1151 ( .A(REGFILE_SIM_reg_bank_reg_r10_31_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3588_));
INVX1 INVX1_1152 ( .A(REGFILE_SIM_reg_bank_reg_r1_sp_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3590_));
INVX1 INVX1_1153 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3199_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3591_));
INVX1 INVX1_1154 ( .A(REGFILE_SIM_reg_bank_reg_r1_sp_1_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3594_));
INVX1 INVX1_1155 ( .A(REGFILE_SIM_reg_bank_reg_r1_sp_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3596_));
INVX1 INVX1_1156 ( .A(REGFILE_SIM_reg_bank_reg_r1_sp_3_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3598_));
INVX1 INVX1_1157 ( .A(REGFILE_SIM_reg_bank_reg_r1_sp_4_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3600_));
INVX1 INVX1_1158 ( .A(REGFILE_SIM_reg_bank_reg_r1_sp_5_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3602_));
INVX1 INVX1_1159 ( .A(REGFILE_SIM_reg_bank_reg_r1_sp_6_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3604_));
INVX1 INVX1_116 ( .A(_abc_40298_new_n994_), .Y(_abc_40298_new_n995_));
INVX1 INVX1_1160 ( .A(REGFILE_SIM_reg_bank_reg_r1_sp_7_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3606_));
INVX1 INVX1_1161 ( .A(REGFILE_SIM_reg_bank_reg_r1_sp_8_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3608_));
INVX1 INVX1_1162 ( .A(REGFILE_SIM_reg_bank_reg_r1_sp_9_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3610_));
INVX1 INVX1_1163 ( .A(REGFILE_SIM_reg_bank_reg_r1_sp_10_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3612_));
INVX1 INVX1_1164 ( .A(REGFILE_SIM_reg_bank_reg_r1_sp_11_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3614_));
INVX1 INVX1_1165 ( .A(REGFILE_SIM_reg_bank_reg_r1_sp_12_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3616_));
INVX1 INVX1_1166 ( .A(REGFILE_SIM_reg_bank_reg_r1_sp_13_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3618_));
INVX1 INVX1_1167 ( .A(REGFILE_SIM_reg_bank_reg_r1_sp_14_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3620_));
INVX1 INVX1_1168 ( .A(REGFILE_SIM_reg_bank_reg_r1_sp_15_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3622_));
INVX1 INVX1_1169 ( .A(REGFILE_SIM_reg_bank_reg_r1_sp_16_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3624_));
INVX1 INVX1_117 ( .A(_abc_40298_new_n1001_), .Y(_abc_40298_new_n1002_));
INVX1 INVX1_1170 ( .A(REGFILE_SIM_reg_bank_reg_r1_sp_17_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3626_));
INVX1 INVX1_1171 ( .A(REGFILE_SIM_reg_bank_reg_r1_sp_18_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3628_));
INVX1 INVX1_1172 ( .A(REGFILE_SIM_reg_bank_reg_r1_sp_19_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3630_));
INVX1 INVX1_1173 ( .A(REGFILE_SIM_reg_bank_reg_r1_sp_20_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3632_));
INVX1 INVX1_1174 ( .A(REGFILE_SIM_reg_bank_reg_r1_sp_21_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3634_));
INVX1 INVX1_1175 ( .A(REGFILE_SIM_reg_bank_reg_r1_sp_22_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3636_));
INVX1 INVX1_1176 ( .A(REGFILE_SIM_reg_bank_reg_r1_sp_23_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3638_));
INVX1 INVX1_1177 ( .A(REGFILE_SIM_reg_bank_reg_r1_sp_24_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3640_));
INVX1 INVX1_1178 ( .A(REGFILE_SIM_reg_bank_reg_r1_sp_25_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3642_));
INVX1 INVX1_1179 ( .A(REGFILE_SIM_reg_bank_reg_r1_sp_26_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3644_));
INVX1 INVX1_118 ( .A(_abc_40298_new_n998_), .Y(_abc_40298_new_n1009_));
INVX1 INVX1_1180 ( .A(REGFILE_SIM_reg_bank_reg_r1_sp_27_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3646_));
INVX1 INVX1_1181 ( .A(REGFILE_SIM_reg_bank_reg_r1_sp_28_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3648_));
INVX1 INVX1_1182 ( .A(REGFILE_SIM_reg_bank_reg_r1_sp_29_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3650_));
INVX1 INVX1_1183 ( .A(REGFILE_SIM_reg_bank_reg_r1_sp_30_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3652_));
INVX1 INVX1_1184 ( .A(REGFILE_SIM_reg_bank_reg_r1_sp_31_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3654_));
INVX1 INVX1_1185 ( .A(REGFILE_SIM_reg_bank_reg_r9_lr_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3656_));
INVX1 INVX1_1186 ( .A(REGFILE_SIM_reg_bank_reg_r9_lr_1_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3659_));
INVX1 INVX1_1187 ( .A(REGFILE_SIM_reg_bank_reg_r9_lr_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3661_));
INVX1 INVX1_1188 ( .A(REGFILE_SIM_reg_bank_reg_r9_lr_3_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3663_));
INVX1 INVX1_1189 ( .A(REGFILE_SIM_reg_bank_reg_r9_lr_4_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3665_));
INVX1 INVX1_119 ( .A(_abc_40298_new_n1012_), .Y(_abc_40298_new_n1013_));
INVX1 INVX1_1190 ( .A(REGFILE_SIM_reg_bank_reg_r9_lr_5_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3667_));
INVX1 INVX1_1191 ( .A(REGFILE_SIM_reg_bank_reg_r9_lr_6_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3669_));
INVX1 INVX1_1192 ( .A(REGFILE_SIM_reg_bank_reg_r9_lr_7_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3671_));
INVX1 INVX1_1193 ( .A(REGFILE_SIM_reg_bank_reg_r9_lr_8_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3673_));
INVX1 INVX1_1194 ( .A(REGFILE_SIM_reg_bank_reg_r9_lr_9_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3675_));
INVX1 INVX1_1195 ( .A(REGFILE_SIM_reg_bank_reg_r9_lr_10_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3677_));
INVX1 INVX1_1196 ( .A(REGFILE_SIM_reg_bank_reg_r9_lr_11_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3679_));
INVX1 INVX1_1197 ( .A(REGFILE_SIM_reg_bank_reg_r9_lr_12_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3681_));
INVX1 INVX1_1198 ( .A(REGFILE_SIM_reg_bank_reg_r9_lr_13_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3683_));
INVX1 INVX1_1199 ( .A(REGFILE_SIM_reg_bank_reg_r9_lr_14_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3685_));
INVX1 INVX1_12 ( .A(inst_r_5_), .Y(_abc_40298_new_n638_));
INVX1 INVX1_120 ( .A(_abc_40298_new_n1015_), .Y(_abc_40298_new_n1016_));
INVX1 INVX1_1200 ( .A(REGFILE_SIM_reg_bank_reg_r9_lr_15_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3687_));
INVX1 INVX1_1201 ( .A(REGFILE_SIM_reg_bank_reg_r9_lr_16_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3689_));
INVX1 INVX1_1202 ( .A(REGFILE_SIM_reg_bank_reg_r9_lr_17_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3691_));
INVX1 INVX1_1203 ( .A(REGFILE_SIM_reg_bank_reg_r9_lr_18_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3693_));
INVX1 INVX1_1204 ( .A(REGFILE_SIM_reg_bank_reg_r9_lr_19_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3695_));
INVX1 INVX1_1205 ( .A(REGFILE_SIM_reg_bank_reg_r9_lr_20_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3697_));
INVX1 INVX1_1206 ( .A(REGFILE_SIM_reg_bank_reg_r9_lr_21_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3699_));
INVX1 INVX1_1207 ( .A(REGFILE_SIM_reg_bank_reg_r9_lr_22_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3701_));
INVX1 INVX1_1208 ( .A(REGFILE_SIM_reg_bank_reg_r9_lr_23_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3703_));
INVX1 INVX1_1209 ( .A(REGFILE_SIM_reg_bank_reg_r9_lr_24_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3705_));
INVX1 INVX1_121 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_2_), .Y(_abc_40298_new_n1030_));
INVX1 INVX1_1210 ( .A(REGFILE_SIM_reg_bank_reg_r9_lr_25_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3707_));
INVX1 INVX1_1211 ( .A(REGFILE_SIM_reg_bank_reg_r9_lr_26_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3709_));
INVX1 INVX1_1212 ( .A(REGFILE_SIM_reg_bank_reg_r9_lr_27_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3711_));
INVX1 INVX1_1213 ( .A(REGFILE_SIM_reg_bank_reg_r9_lr_28_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3713_));
INVX1 INVX1_1214 ( .A(REGFILE_SIM_reg_bank_reg_r9_lr_29_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3715_));
INVX1 INVX1_1215 ( .A(REGFILE_SIM_reg_bank_reg_r9_lr_30_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3717_));
INVX1 INVX1_1216 ( .A(REGFILE_SIM_reg_bank_reg_r9_lr_31_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3719_));
INVX1 INVX1_1217 ( .A(REGFILE_SIM_reg_bank_reg_r8_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3721_));
INVX1 INVX1_1218 ( .A(REGFILE_SIM_reg_bank_reg_r8_1_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3724_));
INVX1 INVX1_1219 ( .A(REGFILE_SIM_reg_bank_reg_r8_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3726_));
INVX1 INVX1_122 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_12_), .Y(_abc_40298_new_n1034_));
INVX1 INVX1_1220 ( .A(REGFILE_SIM_reg_bank_reg_r8_3_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3728_));
INVX1 INVX1_1221 ( .A(REGFILE_SIM_reg_bank_reg_r8_4_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3730_));
INVX1 INVX1_1222 ( .A(REGFILE_SIM_reg_bank_reg_r8_5_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3732_));
INVX1 INVX1_1223 ( .A(REGFILE_SIM_reg_bank_reg_r8_6_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3734_));
INVX1 INVX1_1224 ( .A(REGFILE_SIM_reg_bank_reg_r8_7_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3736_));
INVX1 INVX1_1225 ( .A(REGFILE_SIM_reg_bank_reg_r8_8_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3738_));
INVX1 INVX1_1226 ( .A(REGFILE_SIM_reg_bank_reg_r8_9_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3740_));
INVX1 INVX1_1227 ( .A(REGFILE_SIM_reg_bank_reg_r8_10_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3742_));
INVX1 INVX1_1228 ( .A(REGFILE_SIM_reg_bank_reg_r8_11_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3744_));
INVX1 INVX1_1229 ( .A(REGFILE_SIM_reg_bank_reg_r8_12_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3746_));
INVX1 INVX1_123 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_15_), .Y(_abc_40298_new_n1035_));
INVX1 INVX1_1230 ( .A(REGFILE_SIM_reg_bank_reg_r8_13_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3748_));
INVX1 INVX1_1231 ( .A(REGFILE_SIM_reg_bank_reg_r8_14_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3750_));
INVX1 INVX1_1232 ( .A(REGFILE_SIM_reg_bank_reg_r8_15_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3752_));
INVX1 INVX1_1233 ( .A(REGFILE_SIM_reg_bank_reg_r8_16_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3754_));
INVX1 INVX1_1234 ( .A(REGFILE_SIM_reg_bank_reg_r8_17_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3756_));
INVX1 INVX1_1235 ( .A(REGFILE_SIM_reg_bank_reg_r8_18_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3758_));
INVX1 INVX1_1236 ( .A(REGFILE_SIM_reg_bank_reg_r8_19_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3760_));
INVX1 INVX1_1237 ( .A(REGFILE_SIM_reg_bank_reg_r8_20_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3762_));
INVX1 INVX1_1238 ( .A(REGFILE_SIM_reg_bank_reg_r8_21_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3764_));
INVX1 INVX1_1239 ( .A(REGFILE_SIM_reg_bank_reg_r8_22_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3766_));
INVX1 INVX1_124 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_14_), .Y(_abc_40298_new_n1036_));
INVX1 INVX1_1240 ( .A(REGFILE_SIM_reg_bank_reg_r8_23_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3768_));
INVX1 INVX1_1241 ( .A(REGFILE_SIM_reg_bank_reg_r8_24_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3770_));
INVX1 INVX1_1242 ( .A(REGFILE_SIM_reg_bank_reg_r8_25_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3772_));
INVX1 INVX1_1243 ( .A(REGFILE_SIM_reg_bank_reg_r8_26_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3774_));
INVX1 INVX1_1244 ( .A(REGFILE_SIM_reg_bank_reg_r8_27_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3776_));
INVX1 INVX1_1245 ( .A(REGFILE_SIM_reg_bank_reg_r8_28_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3778_));
INVX1 INVX1_1246 ( .A(REGFILE_SIM_reg_bank_reg_r8_29_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3780_));
INVX1 INVX1_1247 ( .A(REGFILE_SIM_reg_bank_reg_r8_30_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3782_));
INVX1 INVX1_1248 ( .A(REGFILE_SIM_reg_bank_reg_r8_31_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3784_));
INVX1 INVX1_1249 ( .A(REGFILE_SIM_reg_bank_reg_r7_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3786_));
INVX1 INVX1_125 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_11_), .Y(_abc_40298_new_n1038_));
INVX1 INVX1_1250 ( .A(REGFILE_SIM_reg_bank_reg_r7_1_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3789_));
INVX1 INVX1_1251 ( .A(REGFILE_SIM_reg_bank_reg_r7_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3791_));
INVX1 INVX1_1252 ( .A(REGFILE_SIM_reg_bank_reg_r7_3_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3793_));
INVX1 INVX1_1253 ( .A(REGFILE_SIM_reg_bank_reg_r7_4_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3795_));
INVX1 INVX1_1254 ( .A(REGFILE_SIM_reg_bank_reg_r7_5_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3797_));
INVX1 INVX1_1255 ( .A(REGFILE_SIM_reg_bank_reg_r7_6_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3799_));
INVX1 INVX1_1256 ( .A(REGFILE_SIM_reg_bank_reg_r7_7_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3801_));
INVX1 INVX1_1257 ( .A(REGFILE_SIM_reg_bank_reg_r7_8_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3803_));
INVX1 INVX1_1258 ( .A(REGFILE_SIM_reg_bank_reg_r7_9_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3805_));
INVX1 INVX1_1259 ( .A(REGFILE_SIM_reg_bank_reg_r7_10_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3807_));
INVX1 INVX1_126 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_13_), .Y(_abc_40298_new_n1039_));
INVX1 INVX1_1260 ( .A(REGFILE_SIM_reg_bank_reg_r7_11_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3809_));
INVX1 INVX1_1261 ( .A(REGFILE_SIM_reg_bank_reg_r7_12_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3811_));
INVX1 INVX1_1262 ( .A(REGFILE_SIM_reg_bank_reg_r7_13_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3813_));
INVX1 INVX1_1263 ( .A(REGFILE_SIM_reg_bank_reg_r7_14_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3815_));
INVX1 INVX1_1264 ( .A(REGFILE_SIM_reg_bank_reg_r7_15_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3817_));
INVX1 INVX1_1265 ( .A(REGFILE_SIM_reg_bank_reg_r7_16_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3819_));
INVX1 INVX1_1266 ( .A(REGFILE_SIM_reg_bank_reg_r7_17_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3821_));
INVX1 INVX1_1267 ( .A(REGFILE_SIM_reg_bank_reg_r7_18_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3823_));
INVX1 INVX1_1268 ( .A(REGFILE_SIM_reg_bank_reg_r7_19_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3825_));
INVX1 INVX1_1269 ( .A(REGFILE_SIM_reg_bank_reg_r7_20_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3827_));
INVX1 INVX1_127 ( .A(_abc_40298_new_n1044_), .Y(_abc_40298_new_n1045_));
INVX1 INVX1_1270 ( .A(REGFILE_SIM_reg_bank_reg_r7_21_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3829_));
INVX1 INVX1_1271 ( .A(REGFILE_SIM_reg_bank_reg_r7_22_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3831_));
INVX1 INVX1_1272 ( .A(REGFILE_SIM_reg_bank_reg_r7_23_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3833_));
INVX1 INVX1_1273 ( .A(REGFILE_SIM_reg_bank_reg_r7_24_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3835_));
INVX1 INVX1_1274 ( .A(REGFILE_SIM_reg_bank_reg_r7_25_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3837_));
INVX1 INVX1_1275 ( .A(REGFILE_SIM_reg_bank_reg_r7_26_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3839_));
INVX1 INVX1_1276 ( .A(REGFILE_SIM_reg_bank_reg_r7_27_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3841_));
INVX1 INVX1_1277 ( .A(REGFILE_SIM_reg_bank_reg_r7_28_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3843_));
INVX1 INVX1_1278 ( .A(REGFILE_SIM_reg_bank_reg_r7_29_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3845_));
INVX1 INVX1_1279 ( .A(REGFILE_SIM_reg_bank_reg_r7_30_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3847_));
INVX1 INVX1_128 ( .A(_abc_40298_new_n1048_), .Y(_abc_40298_new_n1049_));
INVX1 INVX1_1280 ( .A(REGFILE_SIM_reg_bank_reg_r7_31_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3849_));
INVX1 INVX1_1281 ( .A(REGFILE_SIM_reg_bank_reg_r6_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3851_));
INVX1 INVX1_1282 ( .A(REGFILE_SIM_reg_bank_reg_r6_1_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3854_));
INVX1 INVX1_1283 ( .A(REGFILE_SIM_reg_bank_reg_r6_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3856_));
INVX1 INVX1_1284 ( .A(REGFILE_SIM_reg_bank_reg_r6_3_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3858_));
INVX1 INVX1_1285 ( .A(REGFILE_SIM_reg_bank_reg_r6_4_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3860_));
INVX1 INVX1_1286 ( .A(REGFILE_SIM_reg_bank_reg_r6_5_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3862_));
INVX1 INVX1_1287 ( .A(REGFILE_SIM_reg_bank_reg_r6_6_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3864_));
INVX1 INVX1_1288 ( .A(REGFILE_SIM_reg_bank_reg_r6_7_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3866_));
INVX1 INVX1_1289 ( .A(REGFILE_SIM_reg_bank_reg_r6_8_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3868_));
INVX1 INVX1_129 ( .A(_abc_40298_new_n1060_), .Y(_abc_40298_new_n1061_));
INVX1 INVX1_1290 ( .A(REGFILE_SIM_reg_bank_reg_r6_9_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3870_));
INVX1 INVX1_1291 ( .A(REGFILE_SIM_reg_bank_reg_r6_10_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3872_));
INVX1 INVX1_1292 ( .A(REGFILE_SIM_reg_bank_reg_r6_11_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3874_));
INVX1 INVX1_1293 ( .A(REGFILE_SIM_reg_bank_reg_r6_12_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3876_));
INVX1 INVX1_1294 ( .A(REGFILE_SIM_reg_bank_reg_r6_13_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3878_));
INVX1 INVX1_1295 ( .A(REGFILE_SIM_reg_bank_reg_r6_14_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3880_));
INVX1 INVX1_1296 ( .A(REGFILE_SIM_reg_bank_reg_r6_15_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3882_));
INVX1 INVX1_1297 ( .A(REGFILE_SIM_reg_bank_reg_r6_16_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3884_));
INVX1 INVX1_1298 ( .A(REGFILE_SIM_reg_bank_reg_r6_17_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3886_));
INVX1 INVX1_1299 ( .A(REGFILE_SIM_reg_bank_reg_r6_18_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3888_));
INVX1 INVX1_13 ( .A(_abc_40298_new_n639_), .Y(_abc_40298_new_n640_));
INVX1 INVX1_130 ( .A(esr_q_2_), .Y(_abc_40298_new_n1064_));
INVX1 INVX1_1300 ( .A(REGFILE_SIM_reg_bank_reg_r6_19_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3890_));
INVX1 INVX1_1301 ( .A(REGFILE_SIM_reg_bank_reg_r6_20_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3892_));
INVX1 INVX1_1302 ( .A(REGFILE_SIM_reg_bank_reg_r6_21_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3894_));
INVX1 INVX1_1303 ( .A(REGFILE_SIM_reg_bank_reg_r6_22_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3896_));
INVX1 INVX1_1304 ( .A(REGFILE_SIM_reg_bank_reg_r6_23_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3898_));
INVX1 INVX1_1305 ( .A(REGFILE_SIM_reg_bank_reg_r6_24_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3900_));
INVX1 INVX1_1306 ( .A(REGFILE_SIM_reg_bank_reg_r6_25_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3902_));
INVX1 INVX1_1307 ( .A(REGFILE_SIM_reg_bank_reg_r6_26_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3904_));
INVX1 INVX1_1308 ( .A(REGFILE_SIM_reg_bank_reg_r6_27_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3906_));
INVX1 INVX1_1309 ( .A(REGFILE_SIM_reg_bank_reg_r6_28_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3908_));
INVX1 INVX1_131 ( .A(_abc_40298_new_n1065_), .Y(_abc_40298_new_n1066_));
INVX1 INVX1_1310 ( .A(REGFILE_SIM_reg_bank_reg_r6_29_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3910_));
INVX1 INVX1_1311 ( .A(REGFILE_SIM_reg_bank_reg_r6_30_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3912_));
INVX1 INVX1_1312 ( .A(REGFILE_SIM_reg_bank_reg_r6_31_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3914_));
INVX1 INVX1_1313 ( .A(REGFILE_SIM_reg_bank_reg_r5_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3916_));
INVX1 INVX1_1314 ( .A(REGFILE_SIM_reg_bank_reg_r5_1_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3919_));
INVX1 INVX1_1315 ( .A(REGFILE_SIM_reg_bank_reg_r5_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3921_));
INVX1 INVX1_1316 ( .A(REGFILE_SIM_reg_bank_reg_r5_3_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3923_));
INVX1 INVX1_1317 ( .A(REGFILE_SIM_reg_bank_reg_r5_4_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3925_));
INVX1 INVX1_1318 ( .A(REGFILE_SIM_reg_bank_reg_r5_5_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3927_));
INVX1 INVX1_1319 ( .A(REGFILE_SIM_reg_bank_reg_r5_6_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3929_));
INVX1 INVX1_132 ( .A(_abc_40298_new_n885_), .Y(_abc_40298_new_n1070_));
INVX1 INVX1_1320 ( .A(REGFILE_SIM_reg_bank_reg_r5_7_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3931_));
INVX1 INVX1_1321 ( .A(REGFILE_SIM_reg_bank_reg_r5_8_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3933_));
INVX1 INVX1_1322 ( .A(REGFILE_SIM_reg_bank_reg_r5_9_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3935_));
INVX1 INVX1_1323 ( .A(REGFILE_SIM_reg_bank_reg_r5_10_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3937_));
INVX1 INVX1_1324 ( .A(REGFILE_SIM_reg_bank_reg_r5_11_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3939_));
INVX1 INVX1_1325 ( .A(REGFILE_SIM_reg_bank_reg_r5_12_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3941_));
INVX1 INVX1_1326 ( .A(REGFILE_SIM_reg_bank_reg_r5_13_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3943_));
INVX1 INVX1_1327 ( .A(REGFILE_SIM_reg_bank_reg_r5_14_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3945_));
INVX1 INVX1_1328 ( .A(REGFILE_SIM_reg_bank_reg_r5_15_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3947_));
INVX1 INVX1_1329 ( .A(REGFILE_SIM_reg_bank_reg_r5_16_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3949_));
INVX1 INVX1_133 ( .A(_abc_40298_new_n1028_), .Y(_abc_40298_new_n1071_));
INVX1 INVX1_1330 ( .A(REGFILE_SIM_reg_bank_reg_r5_17_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3951_));
INVX1 INVX1_1331 ( .A(REGFILE_SIM_reg_bank_reg_r5_18_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3953_));
INVX1 INVX1_1332 ( .A(REGFILE_SIM_reg_bank_reg_r5_19_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3955_));
INVX1 INVX1_1333 ( .A(REGFILE_SIM_reg_bank_reg_r5_20_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3957_));
INVX1 INVX1_1334 ( .A(REGFILE_SIM_reg_bank_reg_r5_21_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3959_));
INVX1 INVX1_1335 ( .A(REGFILE_SIM_reg_bank_reg_r5_22_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3961_));
INVX1 INVX1_1336 ( .A(REGFILE_SIM_reg_bank_reg_r5_23_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3963_));
INVX1 INVX1_1337 ( .A(REGFILE_SIM_reg_bank_reg_r5_24_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3965_));
INVX1 INVX1_1338 ( .A(REGFILE_SIM_reg_bank_reg_r5_25_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3967_));
INVX1 INVX1_1339 ( .A(REGFILE_SIM_reg_bank_reg_r5_26_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3969_));
INVX1 INVX1_134 ( .A(intr_i), .Y(_abc_40298_new_n1073_));
INVX1 INVX1_1340 ( .A(REGFILE_SIM_reg_bank_reg_r5_27_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3971_));
INVX1 INVX1_1341 ( .A(REGFILE_SIM_reg_bank_reg_r5_28_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3973_));
INVX1 INVX1_1342 ( .A(REGFILE_SIM_reg_bank_reg_r5_29_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3975_));
INVX1 INVX1_1343 ( .A(REGFILE_SIM_reg_bank_reg_r5_30_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3977_));
INVX1 INVX1_1344 ( .A(REGFILE_SIM_reg_bank_reg_r5_31_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3979_));
INVX1 INVX1_1345 ( .A(REGFILE_SIM_reg_bank_reg_r4_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3981_));
INVX1 INVX1_1346 ( .A(REGFILE_SIM_reg_bank_reg_r4_1_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3984_));
INVX1 INVX1_1347 ( .A(REGFILE_SIM_reg_bank_reg_r4_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3986_));
INVX1 INVX1_1348 ( .A(REGFILE_SIM_reg_bank_reg_r4_3_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3988_));
INVX1 INVX1_1349 ( .A(REGFILE_SIM_reg_bank_reg_r4_4_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3990_));
INVX1 INVX1_135 ( .A(_abc_40298_new_n1043_), .Y(_abc_40298_new_n1074_));
INVX1 INVX1_1350 ( .A(REGFILE_SIM_reg_bank_reg_r4_5_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3992_));
INVX1 INVX1_1351 ( .A(REGFILE_SIM_reg_bank_reg_r4_6_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3994_));
INVX1 INVX1_1352 ( .A(REGFILE_SIM_reg_bank_reg_r4_7_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3996_));
INVX1 INVX1_1353 ( .A(REGFILE_SIM_reg_bank_reg_r4_8_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3998_));
INVX1 INVX1_1354 ( .A(REGFILE_SIM_reg_bank_reg_r4_9_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4000_));
INVX1 INVX1_1355 ( .A(REGFILE_SIM_reg_bank_reg_r4_10_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4002_));
INVX1 INVX1_1356 ( .A(REGFILE_SIM_reg_bank_reg_r4_11_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4004_));
INVX1 INVX1_1357 ( .A(REGFILE_SIM_reg_bank_reg_r4_12_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4006_));
INVX1 INVX1_1358 ( .A(REGFILE_SIM_reg_bank_reg_r4_13_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4008_));
INVX1 INVX1_1359 ( .A(REGFILE_SIM_reg_bank_reg_r4_14_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4010_));
INVX1 INVX1_136 ( .A(_abc_40298_new_n1080_), .Y(_abc_40298_new_n1081_));
INVX1 INVX1_1360 ( .A(REGFILE_SIM_reg_bank_reg_r4_15_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4012_));
INVX1 INVX1_1361 ( .A(REGFILE_SIM_reg_bank_reg_r4_16_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4014_));
INVX1 INVX1_1362 ( .A(REGFILE_SIM_reg_bank_reg_r4_17_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4016_));
INVX1 INVX1_1363 ( .A(REGFILE_SIM_reg_bank_reg_r4_18_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4018_));
INVX1 INVX1_1364 ( .A(REGFILE_SIM_reg_bank_reg_r4_19_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4020_));
INVX1 INVX1_1365 ( .A(REGFILE_SIM_reg_bank_reg_r4_20_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4022_));
INVX1 INVX1_1366 ( .A(REGFILE_SIM_reg_bank_reg_r4_21_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4024_));
INVX1 INVX1_1367 ( .A(REGFILE_SIM_reg_bank_reg_r4_22_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4026_));
INVX1 INVX1_1368 ( .A(REGFILE_SIM_reg_bank_reg_r4_23_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4028_));
INVX1 INVX1_1369 ( .A(REGFILE_SIM_reg_bank_reg_r4_24_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4030_));
INVX1 INVX1_137 ( .A(sr_q_9_), .Y(_abc_40298_new_n1089_));
INVX1 INVX1_1370 ( .A(REGFILE_SIM_reg_bank_reg_r4_25_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4032_));
INVX1 INVX1_1371 ( .A(REGFILE_SIM_reg_bank_reg_r4_26_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4034_));
INVX1 INVX1_1372 ( .A(REGFILE_SIM_reg_bank_reg_r4_27_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4036_));
INVX1 INVX1_1373 ( .A(REGFILE_SIM_reg_bank_reg_r4_28_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4038_));
INVX1 INVX1_1374 ( .A(REGFILE_SIM_reg_bank_reg_r4_29_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4040_));
INVX1 INVX1_1375 ( .A(REGFILE_SIM_reg_bank_reg_r4_30_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4042_));
INVX1 INVX1_1376 ( .A(REGFILE_SIM_reg_bank_reg_r4_31_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4044_));
INVX1 INVX1_1377 ( .A(REGFILE_SIM_reg_bank_reg_r3_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4046_));
INVX1 INVX1_1378 ( .A(REGFILE_SIM_reg_bank_reg_r3_1_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4049_));
INVX1 INVX1_1379 ( .A(REGFILE_SIM_reg_bank_reg_r3_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4051_));
INVX1 INVX1_138 ( .A(alu_equal_o), .Y(_abc_40298_new_n1092_));
INVX1 INVX1_1380 ( .A(REGFILE_SIM_reg_bank_reg_r3_3_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4053_));
INVX1 INVX1_1381 ( .A(REGFILE_SIM_reg_bank_reg_r3_4_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4055_));
INVX1 INVX1_1382 ( .A(REGFILE_SIM_reg_bank_reg_r3_5_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4057_));
INVX1 INVX1_1383 ( .A(REGFILE_SIM_reg_bank_reg_r3_6_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4059_));
INVX1 INVX1_1384 ( .A(REGFILE_SIM_reg_bank_reg_r3_7_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4061_));
INVX1 INVX1_1385 ( .A(REGFILE_SIM_reg_bank_reg_r3_8_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4063_));
INVX1 INVX1_1386 ( .A(REGFILE_SIM_reg_bank_reg_r3_9_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4065_));
INVX1 INVX1_1387 ( .A(REGFILE_SIM_reg_bank_reg_r3_10_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4067_));
INVX1 INVX1_1388 ( .A(REGFILE_SIM_reg_bank_reg_r3_11_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4069_));
INVX1 INVX1_1389 ( .A(REGFILE_SIM_reg_bank_reg_r3_12_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4071_));
INVX1 INVX1_139 ( .A(alu_less_than_o), .Y(_abc_40298_new_n1095_));
INVX1 INVX1_1390 ( .A(REGFILE_SIM_reg_bank_reg_r3_13_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4073_));
INVX1 INVX1_1391 ( .A(REGFILE_SIM_reg_bank_reg_r3_14_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4075_));
INVX1 INVX1_1392 ( .A(REGFILE_SIM_reg_bank_reg_r3_15_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4077_));
INVX1 INVX1_1393 ( .A(REGFILE_SIM_reg_bank_reg_r3_16_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4079_));
INVX1 INVX1_1394 ( .A(REGFILE_SIM_reg_bank_reg_r3_17_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4081_));
INVX1 INVX1_1395 ( .A(REGFILE_SIM_reg_bank_reg_r3_18_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4083_));
INVX1 INVX1_1396 ( .A(REGFILE_SIM_reg_bank_reg_r3_19_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4085_));
INVX1 INVX1_1397 ( .A(REGFILE_SIM_reg_bank_reg_r3_20_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4087_));
INVX1 INVX1_1398 ( .A(REGFILE_SIM_reg_bank_reg_r3_21_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4089_));
INVX1 INVX1_1399 ( .A(REGFILE_SIM_reg_bank_reg_r3_22_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4091_));
INVX1 INVX1_14 ( .A(_abc_40298_new_n642_), .Y(_abc_40298_new_n643_));
INVX1 INVX1_140 ( .A(alu_less_than_signed_o), .Y(_abc_40298_new_n1098_));
INVX1 INVX1_1400 ( .A(REGFILE_SIM_reg_bank_reg_r3_23_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4093_));
INVX1 INVX1_1401 ( .A(REGFILE_SIM_reg_bank_reg_r3_24_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4095_));
INVX1 INVX1_1402 ( .A(REGFILE_SIM_reg_bank_reg_r3_25_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4097_));
INVX1 INVX1_1403 ( .A(REGFILE_SIM_reg_bank_reg_r3_26_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4099_));
INVX1 INVX1_1404 ( .A(REGFILE_SIM_reg_bank_reg_r3_27_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4101_));
INVX1 INVX1_1405 ( .A(REGFILE_SIM_reg_bank_reg_r3_28_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4103_));
INVX1 INVX1_1406 ( .A(REGFILE_SIM_reg_bank_reg_r3_29_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4105_));
INVX1 INVX1_1407 ( .A(REGFILE_SIM_reg_bank_reg_r3_30_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4107_));
INVX1 INVX1_1408 ( .A(REGFILE_SIM_reg_bank_reg_r3_31_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4109_));
INVX1 INVX1_1409 ( .A(REGFILE_SIM_reg_bank_reg_r2_fp_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4111_));
INVX1 INVX1_141 ( .A(_abc_40298_new_n1106_), .Y(_abc_40298_new_n1107_));
INVX1 INVX1_1410 ( .A(REGFILE_SIM_reg_bank_reg_r2_fp_1_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4114_));
INVX1 INVX1_1411 ( .A(REGFILE_SIM_reg_bank_reg_r2_fp_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4116_));
INVX1 INVX1_1412 ( .A(REGFILE_SIM_reg_bank_reg_r2_fp_3_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4118_));
INVX1 INVX1_1413 ( .A(REGFILE_SIM_reg_bank_reg_r2_fp_4_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4120_));
INVX1 INVX1_1414 ( .A(REGFILE_SIM_reg_bank_reg_r2_fp_5_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4122_));
INVX1 INVX1_1415 ( .A(REGFILE_SIM_reg_bank_reg_r2_fp_6_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4124_));
INVX1 INVX1_1416 ( .A(REGFILE_SIM_reg_bank_reg_r2_fp_7_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4126_));
INVX1 INVX1_1417 ( .A(REGFILE_SIM_reg_bank_reg_r2_fp_8_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4128_));
INVX1 INVX1_1418 ( .A(REGFILE_SIM_reg_bank_reg_r2_fp_9_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4130_));
INVX1 INVX1_1419 ( .A(REGFILE_SIM_reg_bank_reg_r2_fp_10_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4132_));
INVX1 INVX1_142 ( .A(_abc_40298_new_n1114_), .Y(_abc_40298_new_n1115_));
INVX1 INVX1_1420 ( .A(REGFILE_SIM_reg_bank_reg_r2_fp_11_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4134_));
INVX1 INVX1_1421 ( .A(REGFILE_SIM_reg_bank_reg_r2_fp_12_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4136_));
INVX1 INVX1_1422 ( .A(REGFILE_SIM_reg_bank_reg_r2_fp_13_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4138_));
INVX1 INVX1_1423 ( .A(REGFILE_SIM_reg_bank_reg_r2_fp_14_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4140_));
INVX1 INVX1_1424 ( .A(REGFILE_SIM_reg_bank_reg_r2_fp_15_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4142_));
INVX1 INVX1_1425 ( .A(REGFILE_SIM_reg_bank_reg_r2_fp_16_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4144_));
INVX1 INVX1_1426 ( .A(REGFILE_SIM_reg_bank_reg_r2_fp_17_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4146_));
INVX1 INVX1_1427 ( .A(REGFILE_SIM_reg_bank_reg_r2_fp_18_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4148_));
INVX1 INVX1_1428 ( .A(REGFILE_SIM_reg_bank_reg_r2_fp_19_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4150_));
INVX1 INVX1_1429 ( .A(REGFILE_SIM_reg_bank_reg_r2_fp_20_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4152_));
INVX1 INVX1_143 ( .A(alu_greater_than_signed_o), .Y(_abc_40298_new_n1118_));
INVX1 INVX1_1430 ( .A(REGFILE_SIM_reg_bank_reg_r2_fp_21_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4154_));
INVX1 INVX1_1431 ( .A(REGFILE_SIM_reg_bank_reg_r2_fp_22_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4156_));
INVX1 INVX1_1432 ( .A(REGFILE_SIM_reg_bank_reg_r2_fp_23_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4158_));
INVX1 INVX1_1433 ( .A(REGFILE_SIM_reg_bank_reg_r2_fp_24_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4160_));
INVX1 INVX1_1434 ( .A(REGFILE_SIM_reg_bank_reg_r2_fp_25_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4162_));
INVX1 INVX1_1435 ( .A(REGFILE_SIM_reg_bank_reg_r2_fp_26_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4164_));
INVX1 INVX1_1436 ( .A(REGFILE_SIM_reg_bank_reg_r2_fp_27_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4166_));
INVX1 INVX1_1437 ( .A(REGFILE_SIM_reg_bank_reg_r2_fp_28_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4168_));
INVX1 INVX1_1438 ( .A(REGFILE_SIM_reg_bank_reg_r2_fp_29_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4170_));
INVX1 INVX1_1439 ( .A(REGFILE_SIM_reg_bank_reg_r2_fp_30_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4172_));
INVX1 INVX1_144 ( .A(_abc_40298_new_n1122_), .Y(_abc_40298_new_n1123_));
INVX1 INVX1_1440 ( .A(REGFILE_SIM_reg_bank_reg_r2_fp_31_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4174_));
INVX1 INVX1_1441 ( .A(REGFILE_SIM_reg_bank_rb_i_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4176_));
INVX1 INVX1_1442 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4178_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4179_));
INVX1 INVX1_1443 ( .A(REGFILE_SIM_reg_bank_rb_i_3_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4181_));
INVX1 INVX1_1444 ( .A(REGFILE_SIM_reg_bank_rb_i_4_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4183_));
INVX1 INVX1_1445 ( .A(REGFILE_SIM_reg_bank_rb_i_1_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4188_));
INVX1 INVX1_1446 ( .A(REGFILE_SIM_reg_bank_rb_i_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4193_));
INVX1 INVX1_1447 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4196_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4197_));
INVX1 INVX1_1448 ( .A(REGFILE_SIM_reg_bank_ra_i_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5248_));
INVX1 INVX1_1449 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5250_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5251_));
INVX1 INVX1_145 ( .A(_abc_40298_new_n1124_), .Y(_abc_40298_new_n1125_));
INVX1 INVX1_1450 ( .A(REGFILE_SIM_reg_bank_ra_i_3_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5253_));
INVX1 INVX1_1451 ( .A(REGFILE_SIM_reg_bank_ra_i_4_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5255_));
INVX1 INVX1_1452 ( .A(REGFILE_SIM_reg_bank_ra_i_1_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5260_));
INVX1 INVX1_1453 ( .A(REGFILE_SIM_reg_bank_ra_i_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5265_));
INVX1 INVX1_1454 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5268_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5269_));
INVX1 INVX1_1455 ( .A(rst_i), .Y(REGFILE_SIM_reg_bank__abc_34451_auto_rtlil_cc_1942_NotGate_31954));
INVX1 INVX1_1456 ( .A(alu_b_i_22_), .Y(alu__abc_38674_new_n110_));
INVX1 INVX1_1457 ( .A(alu_a_i_22_), .Y(alu__abc_38674_new_n111_));
INVX1 INVX1_1458 ( .A(alu__abc_38674_new_n114_), .Y(alu__abc_38674_new_n115_));
INVX1 INVX1_1459 ( .A(alu_b_i_23_), .Y(alu__abc_38674_new_n116_));
INVX1 INVX1_146 ( .A(_abc_40298_new_n1130_), .Y(_abc_40298_new_n1131_));
INVX1 INVX1_1460 ( .A(alu_a_i_23_), .Y(alu__abc_38674_new_n117_));
INVX1 INVX1_1461 ( .A(alu_b_i_20_), .Y(alu__abc_38674_new_n121_));
INVX1 INVX1_1462 ( .A(alu_a_i_20_), .Y(alu__abc_38674_new_n122_));
INVX1 INVX1_1463 ( .A(alu__abc_38674_new_n125_), .Y(alu__abc_38674_new_n126_));
INVX1 INVX1_1464 ( .A(alu_b_i_21_), .Y(alu__abc_38674_new_n127_));
INVX1 INVX1_1465 ( .A(alu_a_i_21_), .Y(alu__abc_38674_new_n128_));
INVX1 INVX1_1466 ( .A(alu__abc_38674_new_n132_), .Y(alu__abc_38674_new_n133_));
INVX1 INVX1_1467 ( .A(alu_b_i_16_), .Y(alu__abc_38674_new_n134_));
INVX1 INVX1_1468 ( .A(alu_a_i_16_), .Y(alu__abc_38674_new_n135_));
INVX1 INVX1_1469 ( .A(alu__abc_38674_new_n140_), .Y(alu__abc_38674_new_n141_));
INVX1 INVX1_147 ( .A(_abc_40298_new_n1132_), .Y(_abc_40298_new_n1133_));
INVX1 INVX1_1470 ( .A(alu_b_i_18_), .Y(alu__abc_38674_new_n143_));
INVX1 INVX1_1471 ( .A(alu_a_i_18_), .Y(alu__abc_38674_new_n144_));
INVX1 INVX1_1472 ( .A(alu__abc_38674_new_n149_), .Y(alu__abc_38674_new_n150_));
INVX1 INVX1_1473 ( .A(alu__abc_38674_new_n152_), .Y(alu__abc_38674_new_n153_));
INVX1 INVX1_1474 ( .A(alu_b_i_30_), .Y(alu__abc_38674_new_n155_));
INVX1 INVX1_1475 ( .A(alu_a_i_30_), .Y(alu__abc_38674_new_n156_));
INVX1 INVX1_1476 ( .A(alu_b_i_29_), .Y(alu__abc_38674_new_n164_));
INVX1 INVX1_1477 ( .A(alu_a_i_29_), .Y(alu__abc_38674_new_n165_));
INVX1 INVX1_1478 ( .A(alu__abc_38674_new_n168_), .Y(alu__abc_38674_new_n169_));
INVX1 INVX1_1479 ( .A(alu_b_i_28_), .Y(alu__abc_38674_new_n170_));
INVX1 INVX1_148 ( .A(_abc_40298_new_n1135_), .Y(_abc_40298_new_n1136_));
INVX1 INVX1_1480 ( .A(alu_a_i_28_), .Y(alu__abc_38674_new_n171_));
INVX1 INVX1_1481 ( .A(alu__abc_38674_new_n174_), .Y(alu__abc_38674_new_n175_));
INVX1 INVX1_1482 ( .A(alu_b_i_24_), .Y(alu__abc_38674_new_n177_));
INVX1 INVX1_1483 ( .A(alu_a_i_24_), .Y(alu__abc_38674_new_n178_));
INVX1 INVX1_1484 ( .A(alu__abc_38674_new_n183_), .Y(alu__abc_38674_new_n184_));
INVX1 INVX1_1485 ( .A(alu_b_i_26_), .Y(alu__abc_38674_new_n186_));
INVX1 INVX1_1486 ( .A(alu_a_i_26_), .Y(alu__abc_38674_new_n187_));
INVX1 INVX1_1487 ( .A(alu__abc_38674_new_n190_), .Y(alu__abc_38674_new_n191_));
INVX1 INVX1_1488 ( .A(alu_b_i_27_), .Y(alu__abc_38674_new_n192_));
INVX1 INVX1_1489 ( .A(alu_a_i_27_), .Y(alu__abc_38674_new_n193_));
INVX1 INVX1_149 ( .A(REGFILE_SIM_reg_bank_wr_i), .Y(_abc_40298_new_n1138_));
INVX1 INVX1_1490 ( .A(alu__abc_38674_new_n197_), .Y(alu__abc_38674_new_n198_));
INVX1 INVX1_1491 ( .A(alu_b_i_14_), .Y(alu__abc_38674_new_n201_));
INVX1 INVX1_1492 ( .A(alu_a_i_14_), .Y(alu__abc_38674_new_n202_));
INVX1 INVX1_1493 ( .A(alu__abc_38674_new_n207_), .Y(alu__abc_38674_new_n208_));
INVX1 INVX1_1494 ( .A(alu_b_i_12_), .Y(alu__abc_38674_new_n210_));
INVX1 INVX1_1495 ( .A(alu_a_i_12_), .Y(alu__abc_38674_new_n211_));
INVX1 INVX1_1496 ( .A(alu__abc_38674_new_n214_), .Y(alu__abc_38674_new_n215_));
INVX1 INVX1_1497 ( .A(alu_b_i_13_), .Y(alu__abc_38674_new_n216_));
INVX1 INVX1_1498 ( .A(alu_a_i_13_), .Y(alu__abc_38674_new_n217_));
INVX1 INVX1_1499 ( .A(alu__abc_38674_new_n221_), .Y(alu__abc_38674_new_n222_));
INVX1 INVX1_15 ( .A(_abc_40298_new_n644_), .Y(_abc_40298_new_n645_));
INVX1 INVX1_150 ( .A(esr_q_9_), .Y(_abc_40298_new_n1139_));
INVX1 INVX1_1500 ( .A(alu_b_i_9_), .Y(alu__abc_38674_new_n227_));
INVX1 INVX1_1501 ( .A(alu_a_i_9_), .Y(alu__abc_38674_new_n228_));
INVX1 INVX1_1502 ( .A(alu_b_i_10_), .Y(alu__abc_38674_new_n232_));
INVX1 INVX1_1503 ( .A(alu_a_i_10_), .Y(alu__abc_38674_new_n233_));
INVX1 INVX1_1504 ( .A(alu__abc_38674_new_n235_), .Y(alu__abc_38674_new_n236_));
INVX1 INVX1_1505 ( .A(alu__abc_38674_new_n239_), .Y(alu__abc_38674_new_n240_));
INVX1 INVX1_1506 ( .A(alu__abc_38674_new_n243_), .Y(alu__abc_38674_new_n244_));
INVX1 INVX1_1507 ( .A(alu_a_i_0_), .Y(alu__abc_38674_new_n258_));
INVX1 INVX1_1508 ( .A(alu__abc_38674_new_n260_), .Y(alu__abc_38674_new_n261_));
INVX1 INVX1_1509 ( .A(alu__abc_38674_new_n264_), .Y(alu__abc_38674_new_n265_));
INVX1 INVX1_151 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_9_), .Y(_abc_40298_new_n1140_));
INVX1 INVX1_1510 ( .A(alu_op_i_2_), .Y(alu__abc_38674_new_n277_));
INVX1 INVX1_1511 ( .A(alu__abc_38674_new_n278_), .Y(alu__abc_38674_new_n279_));
INVX1 INVX1_1512 ( .A(alu__abc_38674_new_n280_), .Y(alu__abc_38674_new_n281_));
INVX1 INVX1_1513 ( .A(alu__abc_38674_new_n282_), .Y(alu__abc_38674_new_n283_));
INVX1 INVX1_1514 ( .A(alu_op_i_0_), .Y(alu__abc_38674_new_n284_));
INVX1 INVX1_1515 ( .A(alu__abc_38674_new_n285_), .Y(alu__abc_38674_new_n286_));
INVX1 INVX1_1516 ( .A(alu_op_i_1_), .Y(alu__abc_38674_new_n288_));
INVX1 INVX1_1517 ( .A(alu__abc_38674_new_n289_), .Y(alu__abc_38674_new_n290_));
INVX1 INVX1_1518 ( .A(alu__abc_38674_new_n291_), .Y(alu__abc_38674_new_n292_));
INVX1 INVX1_1519 ( .A(alu_a_i_31_), .Y(alu__abc_38674_new_n294_));
INVX1 INVX1_152 ( .A(esr_q_10_), .Y(_abc_40298_new_n1153_));
INVX1 INVX1_1520 ( .A(alu_a_i_25_), .Y(alu__abc_38674_new_n295_));
INVX1 INVX1_1521 ( .A(alu__abc_38674_new_n298_), .Y(alu__abc_38674_new_n299_));
INVX1 INVX1_1522 ( .A(alu__abc_38674_new_n304_), .Y(alu__abc_38674_new_n305_));
INVX1 INVX1_1523 ( .A(alu__abc_38674_new_n306_), .Y(alu__abc_38674_new_n307_));
INVX1 INVX1_1524 ( .A(alu_a_i_17_), .Y(alu__abc_38674_new_n308_));
INVX1 INVX1_1525 ( .A(alu_a_i_19_), .Y(alu__abc_38674_new_n312_));
INVX1 INVX1_1526 ( .A(alu__abc_38674_new_n319_), .Y(alu__abc_38674_new_n320_));
INVX1 INVX1_1527 ( .A(alu__abc_38674_new_n321_), .Y(alu__abc_38674_new_n322_));
INVX1 INVX1_1528 ( .A(alu__abc_38674_new_n250_), .Y(alu__abc_38674_new_n328_));
INVX1 INVX1_1529 ( .A(alu_a_i_7_), .Y(alu__abc_38674_new_n329_));
INVX1 INVX1_153 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_10_), .Y(_abc_40298_new_n1154_));
INVX1 INVX1_1530 ( .A(alu_a_i_6_), .Y(alu__abc_38674_new_n330_));
INVX1 INVX1_1531 ( .A(alu_a_i_5_), .Y(alu__abc_38674_new_n334_));
INVX1 INVX1_1532 ( .A(alu_a_i_1_), .Y(alu__abc_38674_new_n336_));
INVX1 INVX1_1533 ( .A(alu_b_i_2_), .Y(alu__abc_38674_new_n338_));
INVX1 INVX1_1534 ( .A(alu_b_i_3_), .Y(alu__abc_38674_new_n340_));
INVX1 INVX1_1535 ( .A(alu_a_i_4_), .Y(alu__abc_38674_new_n345_));
INVX1 INVX1_1536 ( .A(alu_a_i_8_), .Y(alu__abc_38674_new_n351_));
INVX1 INVX1_1537 ( .A(alu_a_i_11_), .Y(alu__abc_38674_new_n356_));
INVX1 INVX1_1538 ( .A(alu__abc_38674_new_n209_), .Y(alu__abc_38674_new_n360_));
INVX1 INVX1_1539 ( .A(alu_a_i_15_), .Y(alu__abc_38674_new_n364_));
INVX1 INVX1_154 ( .A(enable_i), .Y(_abc_40298_new_n1166_));
INVX1 INVX1_1540 ( .A(alu__abc_38674_new_n381_), .Y(alu__abc_38674_new_n382_));
INVX1 INVX1_1541 ( .A(alu__abc_38674_new_n159_), .Y(alu__abc_38674_new_n383_));
INVX1 INVX1_1542 ( .A(alu__abc_38674_new_n162_), .Y(alu__abc_38674_new_n384_));
INVX1 INVX1_1543 ( .A(alu__abc_38674_new_n166_), .Y(alu__abc_38674_new_n386_));
INVX1 INVX1_1544 ( .A(alu__abc_38674_new_n172_), .Y(alu__abc_38674_new_n387_));
INVX1 INVX1_1545 ( .A(alu__abc_38674_new_n389_), .Y(alu__abc_38674_new_n390_));
INVX1 INVX1_1546 ( .A(alu__abc_38674_new_n188_), .Y(alu__abc_38674_new_n393_));
INVX1 INVX1_1547 ( .A(alu__abc_38674_new_n194_), .Y(alu__abc_38674_new_n394_));
INVX1 INVX1_1548 ( .A(alu__abc_38674_new_n395_), .Y(alu__abc_38674_new_n396_));
INVX1 INVX1_1549 ( .A(alu__abc_38674_new_n399_), .Y(alu__abc_38674_new_n400_));
INVX1 INVX1_155 ( .A(_abc_40298_new_n1134_), .Y(_abc_40298_new_n1168_));
INVX1 INVX1_1550 ( .A(alu__abc_38674_new_n405_), .Y(alu__abc_38674_new_n406_));
INVX1 INVX1_1551 ( .A(alu__abc_38674_new_n123_), .Y(alu__abc_38674_new_n407_));
INVX1 INVX1_1552 ( .A(alu__abc_38674_new_n129_), .Y(alu__abc_38674_new_n408_));
INVX1 INVX1_1553 ( .A(alu__abc_38674_new_n148_), .Y(alu__abc_38674_new_n415_));
INVX1 INVX1_1554 ( .A(alu__abc_38674_new_n270_), .Y(alu__abc_38674_new_n423_));
INVX1 INVX1_1555 ( .A(alu__abc_38674_new_n437_), .Y(alu__abc_38674_new_n438_));
INVX1 INVX1_1556 ( .A(alu__abc_38674_new_n231_), .Y(alu__abc_38674_new_n446_));
INVX1 INVX1_1557 ( .A(alu__abc_38674_new_n461_), .Y(alu__abc_38674_new_n462_));
INVX1 INVX1_1558 ( .A(alu__abc_38674_new_n471_), .Y(alu__abc_38674_new_n472_));
INVX1 INVX1_1559 ( .A(alu__abc_38674_new_n473_), .Y(alu__abc_38674_new_n474_));
INVX1 INVX1_156 ( .A(_abc_40298_new_n1169_), .Y(_abc_40298_new_n1170_));
INVX1 INVX1_1560 ( .A(alu__abc_38674_new_n145_), .Y(alu__abc_38674_new_n485_));
INVX1 INVX1_1561 ( .A(alu__abc_38674_new_n414_), .Y(alu__abc_38674_new_n486_));
INVX1 INVX1_1562 ( .A(alu__abc_38674_new_n466_), .Y(alu__abc_38674_new_n487_));
INVX1 INVX1_1563 ( .A(alu__abc_38674_new_n409_), .Y(alu__abc_38674_new_n494_));
INVX1 INVX1_1564 ( .A(alu__abc_38674_new_n179_), .Y(alu__abc_38674_new_n501_));
INVX1 INVX1_1565 ( .A(alu__abc_38674_new_n503_), .Y(alu__abc_38674_new_n504_));
INVX1 INVX1_1566 ( .A(alu__abc_38674_new_n507_), .Y(alu__abc_38674_new_n508_));
INVX1 INVX1_1567 ( .A(alu__abc_38674_new_n465_), .Y(alu__abc_38674_new_n509_));
INVX1 INVX1_1568 ( .A(alu__abc_38674_new_n510_), .Y(alu__abc_38674_new_n511_));
INVX1 INVX1_1569 ( .A(alu__abc_38674_new_n203_), .Y(alu__abc_38674_new_n512_));
INVX1 INVX1_157 ( .A(_abc_40298_new_n1175_), .Y(_abc_40298_new_n1176_));
INVX1 INVX1_1570 ( .A(alu__abc_38674_new_n452_), .Y(alu__abc_38674_new_n513_));
INVX1 INVX1_1571 ( .A(alu_b_i_4_), .Y(alu__abc_38674_new_n519_));
INVX1 INVX1_1572 ( .A(alu__abc_38674_new_n453_), .Y(alu__abc_38674_new_n529_));
INVX1 INVX1_1573 ( .A(alu__abc_38674_new_n456_), .Y(alu__abc_38674_new_n530_));
INVX1 INVX1_1574 ( .A(alu__abc_38674_new_n537_), .Y(alu__abc_38674_new_n538_));
INVX1 INVX1_1575 ( .A(alu__abc_38674_new_n225_), .Y(alu__abc_38674_new_n539_));
INVX1 INVX1_1576 ( .A(alu__abc_38674_new_n271_), .Y(alu__abc_38674_new_n555_));
INVX1 INVX1_1577 ( .A(alu_b_i_1_), .Y(alu__abc_38674_new_n559_));
INVX1 INVX1_1578 ( .A(alu_b_i_0_), .Y(alu__abc_38674_new_n562_));
INVX1 INVX1_1579 ( .A(alu__abc_38674_new_n565_), .Y(alu__abc_38674_new_n566_));
INVX1 INVX1_158 ( .A(_abc_40298_new_n1011_), .Y(_abc_40298_new_n1177_));
INVX1 INVX1_1580 ( .A(alu__abc_38674_new_n212_), .Y(alu__abc_38674_new_n578_));
INVX1 INVX1_1581 ( .A(alu__abc_38674_new_n451_), .Y(alu__abc_38674_new_n579_));
INVX1 INVX1_1582 ( .A(alu__abc_38674_new_n460_), .Y(alu__abc_38674_new_n585_));
INVX1 INVX1_1583 ( .A(alu__abc_38674_new_n157_), .Y(alu__abc_38674_new_n610_));
INVX1 INVX1_1584 ( .A(alu__abc_38674_new_n619_), .Y(alu__abc_38674_new_n620_));
INVX1 INVX1_1585 ( .A(alu__abc_38674_new_n623_), .Y(alu__abc_38674_new_n624_));
INVX1 INVX1_1586 ( .A(alu_a_i_3_), .Y(alu__abc_38674_new_n641_));
INVX1 INVX1_1587 ( .A(alu__abc_38674_new_n644_), .Y(alu__abc_38674_new_n645_));
INVX1 INVX1_1588 ( .A(alu__abc_38674_new_n660_), .Y(alu__abc_38674_new_n661_));
INVX1 INVX1_1589 ( .A(alu__abc_38674_new_n666_), .Y(alu__abc_38674_new_n667_));
INVX1 INVX1_159 ( .A(_abc_40298_new_n1076_), .Y(_abc_40298_new_n1181_));
INVX1 INVX1_1590 ( .A(alu__abc_38674_new_n673_), .Y(alu__abc_38674_new_n674_));
INVX1 INVX1_1591 ( .A(alu__abc_38674_new_n679_), .Y(alu__abc_38674_new_n680_));
INVX1 INVX1_1592 ( .A(alu__abc_38674_new_n259_), .Y(alu__abc_38674_new_n695_));
INVX1 INVX1_1593 ( .A(alu__abc_38674_new_n656_), .Y(alu__abc_38674_new_n698_));
INVX1 INVX1_1594 ( .A(alu__abc_38674_new_n699_), .Y(alu__abc_38674_new_n700_));
INVX1 INVX1_1595 ( .A(alu__abc_38674_new_n701_), .Y(alu__abc_38674_new_n702_));
INVX1 INVX1_1596 ( .A(alu__abc_38674_new_n712_), .Y(alu__abc_38674_new_n713_));
INVX1 INVX1_1597 ( .A(alu__abc_38674_new_n728_), .Y(alu__abc_38674_new_n729_));
INVX1 INVX1_1598 ( .A(alu__abc_38674_new_n743_), .Y(alu__abc_38674_new_n744_));
INVX1 INVX1_1599 ( .A(alu__abc_38674_new_n753_), .Y(alu__abc_38674_new_n754_));
INVX1 INVX1_16 ( .A(_abc_40298_new_n647_), .Y(_abc_40298_new_n648_));
INVX1 INVX1_160 ( .A(_abc_40298_new_n1054_), .Y(_abc_40298_new_n1182_));
INVX1 INVX1_1600 ( .A(alu__abc_38674_new_n758_), .Y(alu__abc_38674_new_n759_));
INVX1 INVX1_1601 ( .A(alu__abc_38674_new_n763_), .Y(alu__abc_38674_new_n764_));
INVX1 INVX1_1602 ( .A(alu__abc_38674_new_n706_), .Y(alu__abc_38674_new_n782_));
INVX1 INVX1_1603 ( .A(alu__abc_38674_new_n703_), .Y(alu__abc_38674_new_n787_));
INVX1 INVX1_1604 ( .A(alu__abc_38674_new_n705_), .Y(alu__abc_38674_new_n788_));
INVX1 INVX1_1605 ( .A(alu__abc_38674_new_n799_), .Y(alu__abc_38674_new_n800_));
INVX1 INVX1_1606 ( .A(alu__abc_38674_new_n677_), .Y(alu__abc_38674_new_n805_));
INVX1 INVX1_1607 ( .A(alu__abc_38674_new_n807_), .Y(alu__abc_38674_new_n808_));
INVX1 INVX1_1608 ( .A(alu__abc_38674_new_n814_), .Y(alu__abc_38674_new_n815_));
INVX1 INVX1_1609 ( .A(alu__abc_38674_new_n817_), .Y(alu__abc_38674_new_n818_));
INVX1 INVX1_161 ( .A(_abc_40298_new_n1185_), .Y(_abc_40298_new_n1186_));
INVX1 INVX1_1610 ( .A(alu__abc_38674_new_n650_), .Y(alu__abc_38674_new_n819_));
INVX1 INVX1_1611 ( .A(alu__abc_38674_new_n636_), .Y(alu__abc_38674_new_n825_));
INVX1 INVX1_1612 ( .A(alu__abc_38674_new_n268_), .Y(alu__abc_38674_new_n834_));
INVX1 INVX1_1613 ( .A(alu__abc_38674_new_n710_), .Y(alu__abc_38674_new_n844_));
INVX1 INVX1_1614 ( .A(alu__abc_38674_new_n855_), .Y(alu__abc_38674_new_n856_));
INVX1 INVX1_1615 ( .A(alu__abc_38674_new_n751_), .Y(alu__abc_38674_new_n860_));
INVX1 INVX1_1616 ( .A(alu__abc_38674_new_n870_), .Y(alu__abc_38674_new_n871_));
INVX1 INVX1_1617 ( .A(alu__abc_38674_new_n731_), .Y(alu__abc_38674_new_n872_));
INVX1 INVX1_1618 ( .A(alu__abc_38674_new_n558_), .Y(alu__abc_38674_new_n883_));
INVX1 INVX1_1619 ( .A(alu__abc_38674_new_n778_), .Y(alu__abc_38674_new_n884_));
INVX1 INVX1_162 ( .A(epc_q_0_), .Y(_abc_40298_new_n1188_));
INVX1 INVX1_1620 ( .A(alu__abc_38674_new_n337_), .Y(alu__abc_38674_new_n895_));
INVX1 INVX1_1621 ( .A(alu__abc_38674_new_n658_), .Y(alu__abc_38674_new_n908_));
INVX1 INVX1_1622 ( .A(alu__abc_38674_new_n685_), .Y(alu__abc_38674_new_n912_));
INVX1 INVX1_1623 ( .A(alu__abc_38674_new_n918_), .Y(alu__abc_38674_new_n919_));
INVX1 INVX1_1624 ( .A(alu__abc_38674_new_n926_), .Y(alu__abc_38674_new_n927_));
INVX1 INVX1_1625 ( .A(alu__abc_38674_new_n929_), .Y(alu__abc_38674_new_n930_));
INVX1 INVX1_1626 ( .A(alu__abc_38674_new_n917_), .Y(alu__abc_38674_new_n941_));
INVX1 INVX1_1627 ( .A(alu__abc_38674_new_n957_), .Y(alu__abc_38674_new_n958_));
INVX1 INVX1_1628 ( .A(alu__abc_38674_new_n552_), .Y(alu__abc_38674_new_n967_));
INVX1 INVX1_1629 ( .A(alu__abc_38674_new_n348_), .Y(alu__abc_38674_new_n976_));
INVX1 INVX1_163 ( .A(epc_q_1_), .Y(_abc_40298_new_n1200_));
INVX1 INVX1_1630 ( .A(alu__abc_38674_new_n995_), .Y(alu__abc_38674_new_n996_));
INVX1 INVX1_1631 ( .A(alu__abc_38674_new_n1019_), .Y(alu__abc_38674_new_n1020_));
INVX1 INVX1_1632 ( .A(alu__abc_38674_new_n955_), .Y(alu__abc_38674_new_n1026_));
INVX1 INVX1_1633 ( .A(alu__abc_38674_new_n540_), .Y(alu__abc_38674_new_n1043_));
INVX1 INVX1_1634 ( .A(alu__abc_38674_new_n687_), .Y(alu__abc_38674_new_n1050_));
INVX1 INVX1_1635 ( .A(alu__abc_38674_new_n696_), .Y(alu__abc_38674_new_n1057_));
INVX1 INVX1_1636 ( .A(alu__abc_38674_new_n993_), .Y(alu__abc_38674_new_n1059_));
INVX1 INVX1_1637 ( .A(alu__abc_38674_new_n1063_), .Y(alu__abc_38674_new_n1064_));
INVX1 INVX1_1638 ( .A(alu__abc_38674_new_n1053_), .Y(alu__abc_38674_new_n1079_));
INVX1 INVX1_1639 ( .A(alu__abc_38674_new_n1028_), .Y(alu__abc_38674_new_n1086_));
INVX1 INVX1_164 ( .A(pc_q_2_), .Y(_abc_40298_new_n1215_));
INVX1 INVX1_1640 ( .A(alu__abc_38674_new_n352_), .Y(alu__abc_38674_new_n1098_));
INVX1 INVX1_1641 ( .A(alu__abc_38674_new_n1112_), .Y(alu__abc_38674_new_n1113_));
INVX1 INVX1_1642 ( .A(alu__abc_38674_new_n1123_), .Y(alu__abc_38674_new_n1124_));
INVX1 INVX1_1643 ( .A(alu__abc_38674_new_n1147_), .Y(alu__abc_38674_new_n1148_));
INVX1 INVX1_1644 ( .A(alu__abc_38674_new_n1030_), .Y(alu__abc_38674_new_n1151_));
INVX1 INVX1_1645 ( .A(alu__abc_38674_new_n1153_), .Y(alu__abc_38674_new_n1154_));
INVX1 INVX1_1646 ( .A(alu__abc_38674_new_n1158_), .Y(alu__abc_38674_new_n1159_));
INVX1 INVX1_1647 ( .A(alu__abc_38674_new_n1161_), .Y(alu__abc_38674_new_n1162_));
INVX1 INVX1_1648 ( .A(alu__abc_38674_new_n1174_), .Y(alu__abc_38674_new_n1175_));
INVX1 INVX1_1649 ( .A(alu__abc_38674_new_n1184_), .Y(alu__abc_38674_new_n1185_));
INVX1 INVX1_165 ( .A(epc_q_3_), .Y(_abc_40298_new_n1229_));
INVX1 INVX1_1650 ( .A(alu__abc_38674_new_n1191_), .Y(alu__abc_38674_new_n1192_));
INVX1 INVX1_1651 ( .A(alu__abc_38674_new_n361_), .Y(alu__abc_38674_new_n1209_));
INVX1 INVX1_1652 ( .A(alu__abc_38674_new_n1219_), .Y(alu__abc_38674_new_n1220_));
INVX1 INVX1_1653 ( .A(alu__abc_38674_new_n1222_), .Y(alu__abc_38674_new_n1223_));
INVX1 INVX1_1654 ( .A(alu__abc_38674_new_n1126_), .Y(alu__abc_38674_new_n1246_));
INVX1 INVX1_1655 ( .A(alu__abc_38674_new_n1180_), .Y(alu__abc_38674_new_n1247_));
INVX1 INVX1_1656 ( .A(alu__abc_38674_new_n1254_), .Y(alu__abc_38674_new_n1255_));
INVX1 INVX1_1657 ( .A(alu__abc_38674_new_n1021_), .Y(alu__abc_38674_new_n1276_));
INVX1 INVX1_1658 ( .A(alu__abc_38674_new_n1282_), .Y(alu__abc_38674_new_n1283_));
INVX1 INVX1_1659 ( .A(alu__abc_38674_new_n1305_), .Y(alu__abc_38674_new_n1306_));
INVX1 INVX1_166 ( .A(_abc_40298_new_n1213_), .Y(_abc_40298_new_n1232_));
INVX1 INVX1_1660 ( .A(alu__abc_38674_new_n1309_), .Y(alu__abc_38674_new_n1310_));
INVX1 INVX1_1661 ( .A(alu__abc_38674_new_n1312_), .Y(alu__abc_38674_new_n1313_));
INVX1 INVX1_1662 ( .A(alu__abc_38674_new_n1317_), .Y(alu__abc_38674_new_n1318_));
INVX1 INVX1_1663 ( .A(alu__abc_38674_new_n1336_), .Y(alu__abc_38674_new_n1337_));
INVX1 INVX1_1664 ( .A(alu__abc_38674_new_n138_), .Y(alu__abc_38674_new_n1350_));
INVX1 INVX1_1665 ( .A(alu__abc_38674_new_n139_), .Y(alu__abc_38674_new_n1351_));
INVX1 INVX1_1666 ( .A(alu__abc_38674_new_n1371_), .Y(alu__abc_38674_new_n1372_));
INVX1 INVX1_1667 ( .A(alu__abc_38674_new_n1128_), .Y(alu__abc_38674_new_n1375_));
INVX1 INVX1_1668 ( .A(alu__abc_38674_new_n490_), .Y(alu__abc_38674_new_n1384_));
INVX1 INVX1_1669 ( .A(alu__abc_38674_new_n1385_), .Y(alu__abc_38674_new_n1411_));
INVX1 INVX1_167 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_3_), .Y(_abc_40298_new_n1233_));
INVX1 INVX1_1670 ( .A(alu__abc_38674_new_n1425_), .Y(alu__abc_38674_new_n1426_));
INVX1 INVX1_1671 ( .A(alu__abc_38674_new_n923_), .Y(alu__abc_38674_new_n1437_));
INVX1 INVX1_1672 ( .A(alu__abc_38674_new_n1417_), .Y(alu__abc_38674_new_n1445_));
INVX1 INVX1_1673 ( .A(alu__abc_38674_new_n1453_), .Y(alu__abc_38674_new_n1454_));
INVX1 INVX1_1674 ( .A(alu__abc_38674_new_n410_), .Y(alu__abc_38674_new_n1461_));
INVX1 INVX1_1675 ( .A(alu__abc_38674_new_n1252_), .Y(alu__abc_38674_new_n1474_));
INVX1 INVX1_1676 ( .A(alu__abc_38674_new_n113_), .Y(alu__abc_38674_new_n1492_));
INVX1 INVX1_1677 ( .A(alu__abc_38674_new_n1392_), .Y(alu__abc_38674_new_n1506_));
INVX1 INVX1_1678 ( .A(alu__abc_38674_new_n1285_), .Y(alu__abc_38674_new_n1512_));
INVX1 INVX1_1679 ( .A(alu__abc_38674_new_n1500_), .Y(alu__abc_38674_new_n1524_));
INVX1 INVX1_168 ( .A(_abc_40298_new_n1246_), .Y(_abc_40298_new_n1247_));
INVX1 INVX1_1680 ( .A(alu__abc_38674_new_n1528_), .Y(alu__abc_38674_new_n1529_));
INVX1 INVX1_1681 ( .A(alu__abc_38674_new_n1507_), .Y(alu__abc_38674_new_n1551_));
INVX1 INVX1_1682 ( .A(alu__abc_38674_new_n1558_), .Y(alu__abc_38674_new_n1559_));
INVX1 INVX1_1683 ( .A(alu__abc_38674_new_n499_), .Y(alu__abc_38674_new_n1573_));
INVX1 INVX1_1684 ( .A(alu__abc_38674_new_n1477_), .Y(alu__abc_38674_new_n1584_));
INVX1 INVX1_1685 ( .A(alu__abc_38674_new_n1585_), .Y(alu__abc_38674_new_n1586_));
INVX1 INVX1_1686 ( .A(alu__abc_38674_new_n1607_), .Y(alu__abc_38674_new_n1608_));
INVX1 INVX1_1687 ( .A(alu__abc_38674_new_n484_), .Y(alu__abc_38674_new_n1624_));
INVX1 INVX1_1688 ( .A(alu__abc_38674_new_n173_), .Y(alu__abc_38674_new_n1639_));
INVX1 INVX1_1689 ( .A(alu__abc_38674_new_n1646_), .Y(alu__abc_38674_new_n1647_));
INVX1 INVX1_169 ( .A(epc_q_4_), .Y(_abc_40298_new_n1252_));
INVX1 INVX1_1690 ( .A(alu__abc_38674_new_n483_), .Y(alu__abc_38674_new_n1649_));
INVX1 INVX1_1691 ( .A(alu__abc_38674_new_n1225_), .Y(alu__abc_38674_new_n1655_));
INVX1 INVX1_1692 ( .A(alu__abc_38674_new_n616_), .Y(alu__abc_38674_new_n1671_));
INVX1 INVX1_1693 ( .A(alu__abc_38674_new_n1692_), .Y(alu__abc_38674_new_n1693_));
INVX1 INVX1_1694 ( .A(alu__abc_38674_new_n1699_), .Y(alu__abc_38674_new_n1700_));
INVX1 INVX1_1695 ( .A(alu__abc_38674_new_n1511_), .Y(alu__abc_38674_new_n1705_));
INVX1 INVX1_1696 ( .A(alu__abc_38674_new_n375_), .Y(alu__abc_38674_new_n1726_));
INVX1 INVX1_17 ( .A(_abc_40298_new_n649_), .Y(_abc_40298_new_n650_));
INVX1 INVX1_170 ( .A(pc_q_3_), .Y(_abc_40298_new_n1255_));
INVX1 INVX1_171 ( .A(pc_q_4_), .Y(_abc_40298_new_n1256_));
INVX1 INVX1_172 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_4_), .Y(_abc_40298_new_n1260_));
INVX1 INVX1_173 ( .A(_abc_40298_new_n1279_), .Y(_abc_40298_new_n1280_));
INVX1 INVX1_174 ( .A(pc_q_5_), .Y(_abc_40298_new_n1287_));
INVX1 INVX1_175 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_5_), .Y(_abc_40298_new_n1293_));
INVX1 INVX1_176 ( .A(pc_q_6_), .Y(_abc_40298_new_n1302_));
INVX1 INVX1_177 ( .A(_abc_40298_new_n1304_), .Y(_abc_40298_new_n1305_));
INVX1 INVX1_178 ( .A(_abc_40298_new_n1306_), .Y(_abc_40298_new_n1308_));
INVX1 INVX1_179 ( .A(epc_q_6_), .Y(_abc_40298_new_n1309_));
INVX1 INVX1_18 ( .A(_abc_40298_new_n625_), .Y(_abc_40298_new_n651_));
INVX1 INVX1_180 ( .A(int32_r_4_), .Y(_abc_40298_new_n1315_));
INVX1 INVX1_181 ( .A(_abc_40298_new_n1317_), .Y(_abc_40298_new_n1318_));
INVX1 INVX1_182 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_6_), .Y(_abc_40298_new_n1322_));
INVX1 INVX1_183 ( .A(pc_q_7_), .Y(_abc_40298_new_n1332_));
INVX1 INVX1_184 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_7_), .Y(_abc_40298_new_n1338_));
INVX1 INVX1_185 ( .A(epc_q_7_), .Y(_abc_40298_new_n1339_));
INVX1 INVX1_186 ( .A(int32_r_5_), .Y(_abc_40298_new_n1341_));
INVX1 INVX1_187 ( .A(_abc_40298_new_n1313_), .Y(_abc_40298_new_n1344_));
INVX1 INVX1_188 ( .A(_abc_40298_new_n1316_), .Y(_abc_40298_new_n1345_));
INVX1 INVX1_189 ( .A(_abc_40298_new_n1343_), .Y(_abc_40298_new_n1348_));
INVX1 INVX1_19 ( .A(_abc_40298_new_n654_), .Y(_abc_40298_new_n655_));
INVX1 INVX1_190 ( .A(_abc_40298_new_n1349_), .Y(_abc_40298_new_n1350_));
INVX1 INVX1_191 ( .A(pc_q_8_), .Y(_abc_40298_new_n1362_));
INVX1 INVX1_192 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_8_), .Y(_abc_40298_new_n1368_));
INVX1 INVX1_193 ( .A(epc_q_8_), .Y(_abc_40298_new_n1369_));
INVX1 INVX1_194 ( .A(_abc_40298_new_n1342_), .Y(_abc_40298_new_n1370_));
INVX1 INVX1_195 ( .A(_abc_40298_new_n1372_), .Y(_abc_40298_new_n1373_));
INVX1 INVX1_196 ( .A(_abc_40298_new_n1384_), .Y(_abc_40298_new_n1385_));
INVX1 INVX1_197 ( .A(epc_q_9_), .Y(_abc_40298_new_n1395_));
INVX1 INVX1_198 ( .A(_abc_40298_new_n886_), .Y(_abc_40298_new_n1396_));
INVX1 INVX1_199 ( .A(pc_q_9_), .Y(_abc_40298_new_n1399_));
INVX1 INVX1_2 ( .A(inst_r_3_), .Y(_abc_40298_new_n619_));
INVX1 INVX1_20 ( .A(inst_r_1_), .Y(_abc_40298_new_n656_));
INVX1 INVX1_200 ( .A(pc_q_10_), .Y(_abc_40298_new_n1414_));
INVX1 INVX1_201 ( .A(_abc_40298_new_n1416_), .Y(_abc_40298_new_n1417_));
INVX1 INVX1_202 ( .A(_abc_40298_new_n1418_), .Y(_abc_40298_new_n1419_));
INVX1 INVX1_203 ( .A(_abc_40298_new_n1428_), .Y(_abc_40298_new_n1429_));
INVX1 INVX1_204 ( .A(_abc_40298_new_n1431_), .Y(_abc_40298_new_n1432_));
INVX1 INVX1_205 ( .A(_abc_40298_new_n1430_), .Y(_abc_40298_new_n1434_));
INVX1 INVX1_206 ( .A(epc_q_10_), .Y(_abc_40298_new_n1437_));
INVX1 INVX1_207 ( .A(pc_q_11_), .Y(_abc_40298_new_n1447_));
INVX1 INVX1_208 ( .A(epc_q_11_), .Y(_abc_40298_new_n1454_));
INVX1 INVX1_209 ( .A(alu_op_r_6_), .Y(_abc_40298_new_n1455_));
INVX1 INVX1_21 ( .A(_abc_40298_new_n658_), .Y(_abc_40298_new_n659_));
INVX1 INVX1_210 ( .A(alu_op_r_7_), .Y(_abc_40298_new_n1457_));
INVX1 INVX1_211 ( .A(_abc_40298_new_n1460_), .Y(_abc_40298_new_n1461_));
INVX1 INVX1_212 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_11_), .Y(_abc_40298_new_n1466_));
INVX1 INVX1_213 ( .A(pc_q_12_), .Y(_abc_40298_new_n1473_));
INVX1 INVX1_214 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_12_), .Y(_abc_40298_new_n1478_));
INVX1 INVX1_215 ( .A(epc_q_12_), .Y(_abc_40298_new_n1479_));
INVX1 INVX1_216 ( .A(_abc_40298_new_n1459_), .Y(_abc_40298_new_n1482_));
INVX1 INVX1_217 ( .A(_abc_40298_new_n1480_), .Y(_abc_40298_new_n1485_));
INVX1 INVX1_218 ( .A(_abc_40298_new_n1486_), .Y(_abc_40298_new_n1487_));
INVX1 INVX1_219 ( .A(_abc_40298_new_n1491_), .Y(_abc_40298_new_n1492_));
INVX1 INVX1_22 ( .A(_abc_40298_new_n663_), .Y(_abc_40298_new_n664_));
INVX1 INVX1_220 ( .A(_abc_40298_new_n1494_), .Y(_abc_40298_new_n1495_));
INVX1 INVX1_221 ( .A(_abc_40298_new_n1502_), .Y(_abc_40298_new_n1503_));
INVX1 INVX1_222 ( .A(pc_q_13_), .Y(_abc_40298_new_n1512_));
INVX1 INVX1_223 ( .A(REGFILE_SIM_reg_bank_rb_i_0_), .Y(_abc_40298_new_n1513_));
INVX1 INVX1_224 ( .A(_abc_40298_new_n1515_), .Y(_abc_40298_new_n1519_));
INVX1 INVX1_225 ( .A(pc_q_14_), .Y(_abc_40298_new_n1532_));
INVX1 INVX1_226 ( .A(_abc_40298_new_n1534_), .Y(_abc_40298_new_n1535_));
INVX1 INVX1_227 ( .A(_abc_40298_new_n1536_), .Y(_abc_40298_new_n1537_));
INVX1 INVX1_228 ( .A(_abc_40298_new_n1517_), .Y(_abc_40298_new_n1540_));
INVX1 INVX1_229 ( .A(_abc_40298_new_n1544_), .Y(_abc_40298_new_n1545_));
INVX1 INVX1_23 ( .A(state_q_2_), .Y(_abc_40298_new_n666_));
INVX1 INVX1_230 ( .A(_abc_40298_new_n1547_), .Y(_abc_40298_new_n1548_));
INVX1 INVX1_231 ( .A(_abc_40298_new_n1542_), .Y(_abc_40298_new_n1549_));
INVX1 INVX1_232 ( .A(pc_q_15_), .Y(_abc_40298_new_n1561_));
INVX1 INVX1_233 ( .A(_abc_40298_new_n1564_), .Y(_abc_40298_new_n1565_));
INVX1 INVX1_234 ( .A(_abc_40298_new_n1566_), .Y(_abc_40298_new_n1568_));
INVX1 INVX1_235 ( .A(epc_q_15_), .Y(_abc_40298_new_n1569_));
INVX1 INVX1_236 ( .A(_abc_40298_new_n1571_), .Y(_abc_40298_new_n1572_));
INVX1 INVX1_237 ( .A(_abc_40298_new_n1573_), .Y(_abc_40298_new_n1574_));
INVX1 INVX1_238 ( .A(pc_q_16_), .Y(_abc_40298_new_n1587_));
INVX1 INVX1_239 ( .A(REGFILE_SIM_reg_bank_rb_i_3_), .Y(_abc_40298_new_n1604_));
INVX1 INVX1_24 ( .A(state_q_3_), .Y(_abc_40298_new_n667_));
INVX1 INVX1_240 ( .A(_abc_40298_new_n1606_), .Y(_abc_40298_new_n1607_));
INVX1 INVX1_241 ( .A(_abc_40298_new_n1613_), .Y(_abc_40298_new_n1614_));
INVX1 INVX1_242 ( .A(pc_q_17_), .Y(_abc_40298_new_n1620_));
INVX1 INVX1_243 ( .A(_abc_40298_new_n1623_), .Y(_abc_40298_new_n1625_));
INVX1 INVX1_244 ( .A(REGFILE_SIM_reg_bank_rb_i_4_), .Y(_abc_40298_new_n1628_));
INVX1 INVX1_245 ( .A(_abc_40298_new_n1630_), .Y(_abc_40298_new_n1631_));
INVX1 INVX1_246 ( .A(pc_q_18_), .Y(_abc_40298_new_n1644_));
INVX1 INVX1_247 ( .A(_abc_40298_new_n1646_), .Y(_abc_40298_new_n1647_));
INVX1 INVX1_248 ( .A(_abc_40298_new_n1648_), .Y(_abc_40298_new_n1649_));
INVX1 INVX1_249 ( .A(_abc_40298_new_n1602_), .Y(_abc_40298_new_n1652_));
INVX1 INVX1_25 ( .A(alu_p_o_0_), .Y(_abc_40298_new_n671_));
INVX1 INVX1_250 ( .A(_abc_40298_new_n1654_), .Y(_abc_40298_new_n1655_));
INVX1 INVX1_251 ( .A(REGFILE_SIM_reg_bank_ra_i_0_), .Y(_abc_40298_new_n1658_));
INVX1 INVX1_252 ( .A(_abc_40298_new_n1660_), .Y(_abc_40298_new_n1661_));
INVX1 INVX1_253 ( .A(_abc_40298_new_n1656_), .Y(_abc_40298_new_n1663_));
INVX1 INVX1_254 ( .A(pc_q_19_), .Y(_abc_40298_new_n1675_));
INVX1 INVX1_255 ( .A(_abc_40298_new_n1677_), .Y(_abc_40298_new_n1679_));
INVX1 INVX1_256 ( .A(REGFILE_SIM_reg_bank_ra_i_1_), .Y(_abc_40298_new_n1683_));
INVX1 INVX1_257 ( .A(pc_q_20_), .Y(_abc_40298_new_n1697_));
INVX1 INVX1_258 ( .A(_abc_40298_new_n1700_), .Y(_abc_40298_new_n1701_));
INVX1 INVX1_259 ( .A(_abc_40298_new_n1706_), .Y(_abc_40298_new_n1707_));
INVX1 INVX1_26 ( .A(mem_offset_q_1_), .Y(_abc_40298_new_n672_));
INVX1 INVX1_260 ( .A(_abc_40298_new_n1653_), .Y(_abc_40298_new_n1708_));
INVX1 INVX1_261 ( .A(REGFILE_SIM_reg_bank_ra_i_2_), .Y(_abc_40298_new_n1712_));
INVX1 INVX1_262 ( .A(pc_q_21_), .Y(_abc_40298_new_n1726_));
INVX1 INVX1_263 ( .A(_abc_40298_new_n1729_), .Y(_abc_40298_new_n1731_));
INVX1 INVX1_264 ( .A(_abc_40298_new_n1713_), .Y(_abc_40298_new_n1733_));
INVX1 INVX1_265 ( .A(REGFILE_SIM_reg_bank_ra_i_3_), .Y(_abc_40298_new_n1735_));
INVX1 INVX1_266 ( .A(_abc_40298_new_n1710_), .Y(_abc_40298_new_n1739_));
INVX1 INVX1_267 ( .A(pc_q_22_), .Y(_abc_40298_new_n1753_));
INVX1 INVX1_268 ( .A(_abc_40298_new_n1755_), .Y(_abc_40298_new_n1756_));
INVX1 INVX1_269 ( .A(_abc_40298_new_n1757_), .Y(_abc_40298_new_n1758_));
INVX1 INVX1_27 ( .A(mem_offset_q_0_), .Y(_abc_40298_new_n676_));
INVX1 INVX1_270 ( .A(_abc_40298_new_n1741_), .Y(_abc_40298_new_n1761_));
INVX1 INVX1_271 ( .A(REGFILE_SIM_reg_bank_ra_i_4_), .Y(_abc_40298_new_n1766_));
INVX1 INVX1_272 ( .A(_abc_40298_new_n1768_), .Y(_abc_40298_new_n1769_));
INVX1 INVX1_273 ( .A(_abc_40298_new_n1764_), .Y(_abc_40298_new_n1771_));
INVX1 INVX1_274 ( .A(pc_q_23_), .Y(_abc_40298_new_n1783_));
INVX1 INVX1_275 ( .A(_abc_40298_new_n1785_), .Y(_abc_40298_new_n1787_));
INVX1 INVX1_276 ( .A(_abc_40298_new_n1792_), .Y(_abc_40298_new_n1793_));
INVX1 INVX1_277 ( .A(pc_q_24_), .Y(_abc_40298_new_n1805_));
INVX1 INVX1_278 ( .A(_abc_40298_new_n1808_), .Y(_abc_40298_new_n1809_));
INVX1 INVX1_279 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_24_), .Y(_abc_40298_new_n1811_));
INVX1 INVX1_28 ( .A(_abc_40298_new_n682_), .Y(_abc_40298_new_n683_));
INVX1 INVX1_280 ( .A(_abc_40298_new_n1763_), .Y(_abc_40298_new_n1814_));
INVX1 INVX1_281 ( .A(_abc_40298_new_n1813_), .Y(_abc_40298_new_n1818_));
INVX1 INVX1_282 ( .A(_abc_40298_new_n1824_), .Y(_abc_40298_new_n1827_));
INVX1 INVX1_283 ( .A(_abc_40298_new_n1834_), .Y(_abc_40298_new_n1835_));
INVX1 INVX1_284 ( .A(pc_q_25_), .Y(_abc_40298_new_n1844_));
INVX1 INVX1_285 ( .A(_abc_40298_new_n1823_), .Y(_abc_40298_new_n1847_));
INVX1 INVX1_286 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_25_), .Y(_abc_40298_new_n1853_));
INVX1 INVX1_287 ( .A(pc_q_26_), .Y(_abc_40298_new_n1862_));
INVX1 INVX1_288 ( .A(_abc_40298_new_n1864_), .Y(_abc_40298_new_n1865_));
INVX1 INVX1_289 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_26_), .Y(_abc_40298_new_n1868_));
INVX1 INVX1_29 ( .A(\mem_dat_i[1] ), .Y(_abc_40298_new_n694_));
INVX1 INVX1_290 ( .A(_abc_40298_new_n1846_), .Y(_abc_40298_new_n1869_));
INVX1 INVX1_291 ( .A(_abc_40298_new_n1872_), .Y(_abc_40298_new_n1873_));
INVX1 INVX1_292 ( .A(_abc_40298_new_n1877_), .Y(_abc_40298_new_n1878_));
INVX1 INVX1_293 ( .A(_abc_40298_new_n1891_), .Y(_abc_40298_new_n1892_));
INVX1 INVX1_294 ( .A(pc_q_27_), .Y(_abc_40298_new_n1895_));
INVX1 INVX1_295 ( .A(_abc_40298_new_n1876_), .Y(_abc_40298_new_n1898_));
INVX1 INVX1_296 ( .A(pc_q_28_), .Y(_abc_40298_new_n1911_));
INVX1 INVX1_297 ( .A(epc_q_28_), .Y(_abc_40298_new_n1916_));
INVX1 INVX1_298 ( .A(_abc_40298_new_n1897_), .Y(_abc_40298_new_n1917_));
INVX1 INVX1_299 ( .A(_abc_40298_new_n1919_), .Y(_abc_40298_new_n1920_));
INVX1 INVX1_3 ( .A(_abc_40298_new_n620_), .Y(_abc_40298_new_n621_));
INVX1 INVX1_30 ( .A(_abc_40298_new_n687_), .Y(_abc_40298_new_n695_));
INVX1 INVX1_300 ( .A(_abc_40298_new_n1918_), .Y(_abc_40298_new_n1922_));
INVX1 INVX1_301 ( .A(_abc_40298_new_n1944_), .Y(_abc_40298_new_n1945_));
INVX1 INVX1_302 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_29_), .Y(_abc_40298_new_n1950_));
INVX1 INVX1_303 ( .A(pc_q_29_), .Y(_abc_40298_new_n1960_));
INVX1 INVX1_304 ( .A(pc_q_30_), .Y(_abc_40298_new_n1961_));
INVX1 INVX1_305 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_30_), .Y(_abc_40298_new_n1967_));
INVX1 INVX1_306 ( .A(_abc_40298_new_n1974_), .Y(_abc_40298_new_n1975_));
INVX1 INVX1_307 ( .A(_abc_40298_new_n1972_), .Y(_abc_40298_new_n1989_));
INVX1 INVX1_308 ( .A(_abc_40298_new_n1973_), .Y(_abc_40298_new_n1990_));
INVX1 INVX1_309 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_31_), .Y(_abc_40298_new_n1996_));
INVX1 INVX1_31 ( .A(_abc_40298_new_n679_), .Y(_abc_40298_new_n699_));
INVX1 INVX1_310 ( .A(pc_q_31_), .Y(_abc_40298_new_n1999_));
INVX1 INVX1_311 ( .A(_abc_40298_new_n2014_), .Y(_abc_40298_new_n2024_));
INVX1 INVX1_312 ( .A(_abc_40298_new_n1027_), .Y(_abc_40298_new_n2043_));
INVX1 INVX1_313 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_0_), .Y(_abc_40298_new_n2139_));
INVX1 INVX1_314 ( .A(_abc_40298_new_n2140_), .Y(_abc_40298_new_n2141_));
INVX1 INVX1_315 ( .A(_abc_40298_new_n931_), .Y(_abc_40298_new_n2147_));
INVX1 INVX1_316 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_1_), .Y(_abc_40298_new_n2153_));
INVX1 INVX1_317 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_13_), .Y(_abc_40298_new_n2190_));
INVX1 INVX1_318 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_14_), .Y(_abc_40298_new_n2193_));
INVX1 INVX1_319 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_15_), .Y(_abc_40298_new_n2196_));
INVX1 INVX1_32 ( .A(_abc_40298_new_n701_), .Y(_abc_40298_new_n702_));
INVX1 INVX1_320 ( .A(_abc_40298_new_n980_), .Y(_abc_40298_new_n2203_));
INVX1 INVX1_321 ( .A(_abc_40298_new_n930_), .Y(_abc_40298_new_n2205_));
INVX1 INVX1_322 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_0_), .Y(_abc_40298_new_n2280_));
INVX1 INVX1_323 ( .A(next_pc_r_0_), .Y(_abc_40298_new_n2281_));
INVX1 INVX1_324 ( .A(_abc_40298_new_n2282_), .Y(_abc_40298_new_n2283_));
INVX1 INVX1_325 ( .A(_abc_40298_new_n2289_), .Y(_abc_40298_new_n2290_));
INVX1 INVX1_326 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_1_), .Y(_abc_40298_new_n2292_));
INVX1 INVX1_327 ( .A(next_pc_r_1_), .Y(_abc_40298_new_n2293_));
INVX1 INVX1_328 ( .A(_abc_40298_new_n2296_), .Y(_abc_40298_new_n2297_));
INVX1 INVX1_329 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_2_), .Y(_abc_40298_new_n2299_));
INVX1 INVX1_33 ( .A(\mem_dat_i[2] ), .Y(_abc_40298_new_n707_));
INVX1 INVX1_330 ( .A(_abc_40298_new_n2286_), .Y(_abc_40298_new_n2302_));
INVX1 INVX1_331 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_3_), .Y(_abc_40298_new_n2307_));
INVX1 INVX1_332 ( .A(_abc_40298_new_n2311_), .Y(_abc_40298_new_n2312_));
INVX1 INVX1_333 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_4_), .Y(_abc_40298_new_n2314_));
INVX1 INVX1_334 ( .A(_abc_40298_new_n2318_), .Y(_abc_40298_new_n2319_));
INVX1 INVX1_335 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_5_), .Y(_abc_40298_new_n2321_));
INVX1 INVX1_336 ( .A(_abc_40298_new_n2324_), .Y(_abc_40298_new_n2325_));
INVX1 INVX1_337 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_6_), .Y(_abc_40298_new_n2327_));
INVX1 INVX1_338 ( .A(_abc_40298_new_n2331_), .Y(_abc_40298_new_n2332_));
INVX1 INVX1_339 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_7_), .Y(_abc_40298_new_n2334_));
INVX1 INVX1_34 ( .A(_abc_40298_new_n712_), .Y(_abc_40298_new_n713_));
INVX1 INVX1_340 ( .A(_abc_40298_new_n1334_), .Y(_abc_40298_new_n2335_));
INVX1 INVX1_341 ( .A(_abc_40298_new_n2339_), .Y(_abc_40298_new_n2340_));
INVX1 INVX1_342 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_8_), .Y(_abc_40298_new_n2342_));
INVX1 INVX1_343 ( .A(_abc_40298_new_n2346_), .Y(_abc_40298_new_n2347_));
INVX1 INVX1_344 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_9_), .Y(_abc_40298_new_n2352_));
INVX1 INVX1_345 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_10_), .Y(_abc_40298_new_n2358_));
INVX1 INVX1_346 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_16_), .Y(_abc_40298_new_n2385_));
INVX1 INVX1_347 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_17_), .Y(_abc_40298_new_n2392_));
INVX1 INVX1_348 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_18_), .Y(_abc_40298_new_n2399_));
INVX1 INVX1_349 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_19_), .Y(_abc_40298_new_n2406_));
INVX1 INVX1_35 ( .A(\mem_dat_i[3] ), .Y(_abc_40298_new_n718_));
INVX1 INVX1_350 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_20_), .Y(_abc_40298_new_n2413_));
INVX1 INVX1_351 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_21_), .Y(_abc_40298_new_n2420_));
INVX1 INVX1_352 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_22_), .Y(_abc_40298_new_n2427_));
INVX1 INVX1_353 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_23_), .Y(_abc_40298_new_n2434_));
INVX1 INVX1_354 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_24_), .Y(_abc_40298_new_n2441_));
INVX1 INVX1_355 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_25_), .Y(_abc_40298_new_n2448_));
INVX1 INVX1_356 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_26_), .Y(_abc_40298_new_n2455_));
INVX1 INVX1_357 ( .A(int32_r_10_), .Y(_abc_40298_new_n2456_));
INVX1 INVX1_358 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_27_), .Y(_abc_40298_new_n2463_));
INVX1 INVX1_359 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_28_), .Y(_abc_40298_new_n2470_));
INVX1 INVX1_36 ( .A(_abc_40298_new_n723_), .Y(_abc_40298_new_n724_));
INVX1 INVX1_360 ( .A(REGFILE_SIM_reg_bank_rb_i_1_), .Y(_abc_40298_new_n2471_));
INVX1 INVX1_361 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_29_), .Y(_abc_40298_new_n2478_));
INVX1 INVX1_362 ( .A(REGFILE_SIM_reg_bank_rb_i_2_), .Y(_abc_40298_new_n2479_));
INVX1 INVX1_363 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_30_), .Y(_abc_40298_new_n2486_));
INVX1 INVX1_364 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_31_), .Y(_abc_40298_new_n2493_));
INVX1 INVX1_365 ( .A(_abc_40298_new_n2284_), .Y(_abc_40298_new_n2510_));
INVX1 INVX1_366 ( .A(_abc_40298_new_n2513_), .Y(_abc_40298_new_n2514_));
INVX1 INVX1_367 ( .A(_abc_40298_new_n2515_), .Y(_abc_40298_new_n2516_));
INVX1 INVX1_368 ( .A(_abc_40298_new_n2518_), .Y(_abc_40298_new_n2519_));
INVX1 INVX1_369 ( .A(_abc_40298_new_n2521_), .Y(_abc_40298_new_n2522_));
INVX1 INVX1_37 ( .A(alu_p_o_4_), .Y(_abc_40298_new_n728_));
INVX1 INVX1_370 ( .A(\mem_dat_i[0] ), .Y(_abc_40298_new_n2524_));
INVX1 INVX1_371 ( .A(\mem_dat_i[4] ), .Y(_abc_40298_new_n2530_));
INVX1 INVX1_372 ( .A(\mem_dat_i[5] ), .Y(_abc_40298_new_n2532_));
INVX1 INVX1_373 ( .A(\mem_dat_i[7] ), .Y(_abc_40298_new_n2535_));
INVX1 INVX1_374 ( .A(\mem_dat_i[8] ), .Y(_abc_40298_new_n2537_));
INVX1 INVX1_375 ( .A(\mem_dat_i[12] ), .Y(_abc_40298_new_n2542_));
INVX1 INVX1_376 ( .A(\mem_dat_i[13] ), .Y(_abc_40298_new_n2544_));
INVX1 INVX1_377 ( .A(\mem_dat_i[15] ), .Y(_abc_40298_new_n2547_));
INVX1 INVX1_378 ( .A(\mem_sel_o[0] ), .Y(_abc_40298_new_n2567_));
INVX1 INVX1_379 ( .A(_abc_40298_new_n641_), .Y(_abc_40298_new_n2568_));
INVX1 INVX1_38 ( .A(alu_p_o_5_), .Y(_abc_40298_new_n737_));
INVX1 INVX1_380 ( .A(_abc_40298_new_n2569_), .Y(_abc_40298_new_n2570_));
INVX1 INVX1_381 ( .A(_abc_40298_new_n2576_), .Y(_abc_40298_new_n2577_));
INVX1 INVX1_382 ( .A(_abc_40298_new_n2520_), .Y(_abc_40298_new_n2580_));
INVX1 INVX1_383 ( .A(\mem_sel_o[1] ), .Y(_abc_40298_new_n2584_));
INVX1 INVX1_384 ( .A(_abc_40298_new_n2585_), .Y(_abc_40298_new_n2586_));
INVX1 INVX1_385 ( .A(_abc_40298_new_n2572_), .Y(_abc_40298_new_n2587_));
INVX1 INVX1_386 ( .A(\mem_sel_o[2] ), .Y(_abc_40298_new_n2592_));
INVX1 INVX1_387 ( .A(\mem_sel_o[3] ), .Y(_abc_40298_new_n2600_));
INVX1 INVX1_388 ( .A(_abc_40298_new_n2601_), .Y(_abc_40298_new_n2602_));
INVX1 INVX1_389 ( .A(_abc_40298_new_n2593_), .Y(_abc_40298_new_n2603_));
INVX1 INVX1_39 ( .A(\mem_dat_i[6] ), .Y(_abc_40298_new_n747_));
INVX1 INVX1_390 ( .A(\mem_dat_o[0] ), .Y(_abc_40298_new_n2607_));
INVX1 INVX1_391 ( .A(_abc_40298_new_n2571_), .Y(_abc_40298_new_n2608_));
INVX1 INVX1_392 ( .A(_abc_40298_new_n2611_), .Y(_abc_40298_new_n2612_));
INVX1 INVX1_393 ( .A(\mem_dat_o[1] ), .Y(_abc_40298_new_n2618_));
INVX1 INVX1_394 ( .A(\mem_dat_o[2] ), .Y(_abc_40298_new_n2626_));
INVX1 INVX1_395 ( .A(\mem_dat_o[3] ), .Y(_abc_40298_new_n2634_));
INVX1 INVX1_396 ( .A(\mem_dat_o[4] ), .Y(_abc_40298_new_n2642_));
INVX1 INVX1_397 ( .A(\mem_dat_o[5] ), .Y(_abc_40298_new_n2650_));
INVX1 INVX1_398 ( .A(\mem_dat_o[6] ), .Y(_abc_40298_new_n2658_));
INVX1 INVX1_399 ( .A(\mem_dat_o[7] ), .Y(_abc_40298_new_n2666_));
INVX1 INVX1_4 ( .A(opcode_q_24_), .Y(_abc_40298_new_n623_));
INVX1 INVX1_40 ( .A(alu_p_o_8_), .Y(_abc_40298_new_n763_));
INVX1 INVX1_400 ( .A(\mem_dat_o[8] ), .Y(_abc_40298_new_n2674_));
INVX1 INVX1_401 ( .A(\mem_dat_o[9] ), .Y(_abc_40298_new_n2683_));
INVX1 INVX1_402 ( .A(\mem_dat_o[10] ), .Y(_abc_40298_new_n2692_));
INVX1 INVX1_403 ( .A(\mem_dat_o[11] ), .Y(_abc_40298_new_n2701_));
INVX1 INVX1_404 ( .A(\mem_dat_o[12] ), .Y(_abc_40298_new_n2710_));
INVX1 INVX1_405 ( .A(\mem_dat_o[13] ), .Y(_abc_40298_new_n2719_));
INVX1 INVX1_406 ( .A(\mem_dat_o[14] ), .Y(_abc_40298_new_n2728_));
INVX1 INVX1_407 ( .A(\mem_dat_o[15] ), .Y(_abc_40298_new_n2737_));
INVX1 INVX1_408 ( .A(\mem_dat_o[16] ), .Y(_abc_40298_new_n2746_));
INVX1 INVX1_409 ( .A(\mem_dat_o[17] ), .Y(_abc_40298_new_n2754_));
INVX1 INVX1_41 ( .A(_abc_40298_new_n653_), .Y(_abc_40298_new_n766_));
INVX1 INVX1_410 ( .A(\mem_dat_o[18] ), .Y(_abc_40298_new_n2762_));
INVX1 INVX1_411 ( .A(\mem_dat_o[19] ), .Y(_abc_40298_new_n2770_));
INVX1 INVX1_412 ( .A(\mem_dat_o[20] ), .Y(_abc_40298_new_n2778_));
INVX1 INVX1_413 ( .A(\mem_dat_o[21] ), .Y(_abc_40298_new_n2786_));
INVX1 INVX1_414 ( .A(\mem_dat_o[22] ), .Y(_abc_40298_new_n2794_));
INVX1 INVX1_415 ( .A(\mem_dat_o[23] ), .Y(_abc_40298_new_n2802_));
INVX1 INVX1_416 ( .A(\mem_dat_o[24] ), .Y(_abc_40298_new_n2810_));
INVX1 INVX1_417 ( .A(\mem_dat_o[25] ), .Y(_abc_40298_new_n2819_));
INVX1 INVX1_418 ( .A(\mem_dat_o[26] ), .Y(_abc_40298_new_n2828_));
INVX1 INVX1_419 ( .A(\mem_dat_o[27] ), .Y(_abc_40298_new_n2837_));
INVX1 INVX1_42 ( .A(alu_p_o_9_), .Y(_abc_40298_new_n769_));
INVX1 INVX1_420 ( .A(\mem_dat_o[28] ), .Y(_abc_40298_new_n2846_));
INVX1 INVX1_421 ( .A(\mem_dat_o[29] ), .Y(_abc_40298_new_n2855_));
INVX1 INVX1_422 ( .A(\mem_dat_o[30] ), .Y(_abc_40298_new_n2864_));
INVX1 INVX1_423 ( .A(\mem_dat_o[31] ), .Y(_abc_40298_new_n2873_));
INVX1 INVX1_424 ( .A(mem_we_o), .Y(_abc_40298_new_n2882_));
INVX1 INVX1_425 ( .A(_abc_40298_new_n2883_), .Y(_abc_40298_new_n2884_));
INVX1 INVX1_426 ( .A(_abc_40298_new_n669_), .Y(_abc_40298_new_n2902_));
INVX1 INVX1_427 ( .A(_abc_40298_new_n2907_), .Y(_abc_40298_new_n2908_));
INVX1 INVX1_428 ( .A(_abc_40298_new_n2912_), .Y(_abc_40298_new_n2922_));
INVX1 INVX1_429 ( .A(_abc_40298_new_n2920_), .Y(_abc_40298_new_n2932_));
INVX1 INVX1_43 ( .A(\mem_dat_i[9] ), .Y(_abc_40298_new_n770_));
INVX1 INVX1_430 ( .A(_abc_40298_new_n2930_), .Y(_abc_40298_new_n2933_));
INVX1 INVX1_431 ( .A(_abc_40298_new_n2944_), .Y(_abc_40298_new_n2951_));
INVX1 INVX1_432 ( .A(_abc_40298_new_n3023_), .Y(_abc_40298_new_n3032_));
INVX1 INVX1_433 ( .A(_abc_40298_new_n3054_), .Y(_abc_40298_new_n3055_));
INVX1 INVX1_434 ( .A(_abc_40298_new_n3051_), .Y(_abc_40298_new_n3057_));
INVX1 INVX1_435 ( .A(_abc_40298_new_n3087_), .Y(_abc_40298_new_n3088_));
INVX1 INVX1_436 ( .A(_abc_40298_new_n3106_), .Y(_abc_40298_new_n3107_));
INVX1 INVX1_437 ( .A(_abc_40298_new_n3115_), .Y(_abc_40298_new_n3116_));
INVX1 INVX1_438 ( .A(_abc_40298_new_n3129_), .Y(_abc_40298_new_n3130_));
INVX1 INVX1_439 ( .A(_abc_40298_new_n3137_), .Y(_abc_40298_new_n3138_));
INVX1 INVX1_44 ( .A(_abc_40298_new_n686_), .Y(_abc_40298_new_n771_));
INVX1 INVX1_440 ( .A(_abc_40298_new_n3145_), .Y(_abc_40298_new_n3146_));
INVX1 INVX1_441 ( .A(_abc_40298_new_n3166_), .Y(_abc_40298_new_n3181_));
INVX1 INVX1_442 ( .A(rst_i), .Y(_abc_40298_auto_rtlil_cc_1942_NotGate_33938));
INVX1 INVX1_443 ( .A(REGFILE_SIM_reg_bank_reg_r31_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2099_));
INVX1 INVX1_444 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2100_));
INVX1 INVX1_445 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2104_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2105_));
INVX1 INVX1_446 ( .A(REGFILE_SIM_reg_bank_reg_r31_1_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2108_));
INVX1 INVX1_447 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_1_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2109_));
INVX1 INVX1_448 ( .A(REGFILE_SIM_reg_bank_reg_r31_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2111_));
INVX1 INVX1_449 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2112_));
INVX1 INVX1_45 ( .A(alu_p_o_10_), .Y(_abc_40298_new_n775_));
INVX1 INVX1_450 ( .A(REGFILE_SIM_reg_bank_reg_r31_3_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2114_));
INVX1 INVX1_451 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_3_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2115_));
INVX1 INVX1_452 ( .A(REGFILE_SIM_reg_bank_reg_r31_4_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2117_));
INVX1 INVX1_453 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_4_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2118_));
INVX1 INVX1_454 ( .A(REGFILE_SIM_reg_bank_reg_r31_5_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2120_));
INVX1 INVX1_455 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_5_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2121_));
INVX1 INVX1_456 ( .A(REGFILE_SIM_reg_bank_reg_r31_6_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2123_));
INVX1 INVX1_457 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_6_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2124_));
INVX1 INVX1_458 ( .A(REGFILE_SIM_reg_bank_reg_r31_7_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2126_));
INVX1 INVX1_459 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_7_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2127_));
INVX1 INVX1_46 ( .A(\mem_dat_i[10] ), .Y(_abc_40298_new_n776_));
INVX1 INVX1_460 ( .A(REGFILE_SIM_reg_bank_reg_r31_8_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2129_));
INVX1 INVX1_461 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_8_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2130_));
INVX1 INVX1_462 ( .A(REGFILE_SIM_reg_bank_reg_r31_9_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2132_));
INVX1 INVX1_463 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_9_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2133_));
INVX1 INVX1_464 ( .A(REGFILE_SIM_reg_bank_reg_r31_10_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2135_));
INVX1 INVX1_465 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_10_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2136_));
INVX1 INVX1_466 ( .A(REGFILE_SIM_reg_bank_reg_r31_11_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2138_));
INVX1 INVX1_467 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_11_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2139_));
INVX1 INVX1_468 ( .A(REGFILE_SIM_reg_bank_reg_r31_12_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2141_));
INVX1 INVX1_469 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_12_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2142_));
INVX1 INVX1_47 ( .A(alu_p_o_11_), .Y(_abc_40298_new_n780_));
INVX1 INVX1_470 ( .A(REGFILE_SIM_reg_bank_reg_r31_13_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2144_));
INVX1 INVX1_471 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_13_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2145_));
INVX1 INVX1_472 ( .A(REGFILE_SIM_reg_bank_reg_r31_14_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2147_));
INVX1 INVX1_473 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_14_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2148_));
INVX1 INVX1_474 ( .A(REGFILE_SIM_reg_bank_reg_r31_15_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2150_));
INVX1 INVX1_475 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_15_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2151_));
INVX1 INVX1_476 ( .A(REGFILE_SIM_reg_bank_reg_r31_16_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2153_));
INVX1 INVX1_477 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_16_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2154_));
INVX1 INVX1_478 ( .A(REGFILE_SIM_reg_bank_reg_r31_17_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2156_));
INVX1 INVX1_479 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_17_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2157_));
INVX1 INVX1_48 ( .A(\mem_dat_i[11] ), .Y(_abc_40298_new_n781_));
INVX1 INVX1_480 ( .A(REGFILE_SIM_reg_bank_reg_r31_18_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2159_));
INVX1 INVX1_481 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_18_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2160_));
INVX1 INVX1_482 ( .A(REGFILE_SIM_reg_bank_reg_r31_19_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2162_));
INVX1 INVX1_483 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_19_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2163_));
INVX1 INVX1_484 ( .A(REGFILE_SIM_reg_bank_reg_r31_20_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2165_));
INVX1 INVX1_485 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_20_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2166_));
INVX1 INVX1_486 ( .A(REGFILE_SIM_reg_bank_reg_r31_21_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2168_));
INVX1 INVX1_487 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_21_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2169_));
INVX1 INVX1_488 ( .A(REGFILE_SIM_reg_bank_reg_r31_22_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2171_));
INVX1 INVX1_489 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_22_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2172_));
INVX1 INVX1_49 ( .A(alu_p_o_12_), .Y(_abc_40298_new_n785_));
INVX1 INVX1_490 ( .A(REGFILE_SIM_reg_bank_reg_r31_23_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2174_));
INVX1 INVX1_491 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_23_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2175_));
INVX1 INVX1_492 ( .A(REGFILE_SIM_reg_bank_reg_r31_24_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2177_));
INVX1 INVX1_493 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_24_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2178_));
INVX1 INVX1_494 ( .A(REGFILE_SIM_reg_bank_reg_r31_25_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2180_));
INVX1 INVX1_495 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_25_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2181_));
INVX1 INVX1_496 ( .A(REGFILE_SIM_reg_bank_reg_r31_26_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2183_));
INVX1 INVX1_497 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_26_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2184_));
INVX1 INVX1_498 ( .A(REGFILE_SIM_reg_bank_reg_r31_27_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2186_));
INVX1 INVX1_499 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_27_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2187_));
INVX1 INVX1_5 ( .A(opcode_q_25_), .Y(_abc_40298_new_n624_));
INVX1 INVX1_50 ( .A(alu_p_o_13_), .Y(_abc_40298_new_n789_));
INVX1 INVX1_500 ( .A(REGFILE_SIM_reg_bank_reg_r31_28_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2189_));
INVX1 INVX1_501 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_28_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2190_));
INVX1 INVX1_502 ( .A(REGFILE_SIM_reg_bank_reg_r31_29_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2192_));
INVX1 INVX1_503 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_29_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2193_));
INVX1 INVX1_504 ( .A(REGFILE_SIM_reg_bank_reg_r31_30_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2195_));
INVX1 INVX1_505 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_30_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2196_));
INVX1 INVX1_506 ( .A(REGFILE_SIM_reg_bank_reg_r31_31_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2198_));
INVX1 INVX1_507 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_31_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2199_));
INVX1 INVX1_508 ( .A(REGFILE_SIM_reg_bank_reg_r30_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2201_));
INVX1 INVX1_509 ( .A(REGFILE_SIM_reg_bank_rd_i_1_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2202_));
INVX1 INVX1_51 ( .A(alu_p_o_14_), .Y(_abc_40298_new_n793_));
INVX1 INVX1_510 ( .A(REGFILE_SIM_reg_bank_reg_r30_1_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2207_));
INVX1 INVX1_511 ( .A(REGFILE_SIM_reg_bank_reg_r30_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2209_));
INVX1 INVX1_512 ( .A(REGFILE_SIM_reg_bank_reg_r30_3_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2211_));
INVX1 INVX1_513 ( .A(REGFILE_SIM_reg_bank_reg_r30_4_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2213_));
INVX1 INVX1_514 ( .A(REGFILE_SIM_reg_bank_reg_r30_5_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2215_));
INVX1 INVX1_515 ( .A(REGFILE_SIM_reg_bank_reg_r30_6_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2217_));
INVX1 INVX1_516 ( .A(REGFILE_SIM_reg_bank_reg_r30_7_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2219_));
INVX1 INVX1_517 ( .A(REGFILE_SIM_reg_bank_reg_r30_8_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2221_));
INVX1 INVX1_518 ( .A(REGFILE_SIM_reg_bank_reg_r30_9_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2223_));
INVX1 INVX1_519 ( .A(REGFILE_SIM_reg_bank_reg_r30_10_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2225_));
INVX1 INVX1_52 ( .A(\mem_dat_i[14] ), .Y(_abc_40298_new_n794_));
INVX1 INVX1_520 ( .A(REGFILE_SIM_reg_bank_reg_r30_11_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2227_));
INVX1 INVX1_521 ( .A(REGFILE_SIM_reg_bank_reg_r30_12_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2229_));
INVX1 INVX1_522 ( .A(REGFILE_SIM_reg_bank_reg_r30_13_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2231_));
INVX1 INVX1_523 ( .A(REGFILE_SIM_reg_bank_reg_r30_14_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2233_));
INVX1 INVX1_524 ( .A(REGFILE_SIM_reg_bank_reg_r30_15_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2235_));
INVX1 INVX1_525 ( .A(REGFILE_SIM_reg_bank_reg_r30_16_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2237_));
INVX1 INVX1_526 ( .A(REGFILE_SIM_reg_bank_reg_r30_17_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2239_));
INVX1 INVX1_527 ( .A(REGFILE_SIM_reg_bank_reg_r30_18_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2241_));
INVX1 INVX1_528 ( .A(REGFILE_SIM_reg_bank_reg_r30_19_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2243_));
INVX1 INVX1_529 ( .A(REGFILE_SIM_reg_bank_reg_r30_20_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2245_));
INVX1 INVX1_53 ( .A(alu_p_o_15_), .Y(_abc_40298_new_n799_));
INVX1 INVX1_530 ( .A(REGFILE_SIM_reg_bank_reg_r30_21_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2247_));
INVX1 INVX1_531 ( .A(REGFILE_SIM_reg_bank_reg_r30_22_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2249_));
INVX1 INVX1_532 ( .A(REGFILE_SIM_reg_bank_reg_r30_23_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2251_));
INVX1 INVX1_533 ( .A(REGFILE_SIM_reg_bank_reg_r30_24_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2253_));
INVX1 INVX1_534 ( .A(REGFILE_SIM_reg_bank_reg_r30_25_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2255_));
INVX1 INVX1_535 ( .A(REGFILE_SIM_reg_bank_reg_r30_26_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2257_));
INVX1 INVX1_536 ( .A(REGFILE_SIM_reg_bank_reg_r30_27_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2259_));
INVX1 INVX1_537 ( .A(REGFILE_SIM_reg_bank_reg_r30_28_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2261_));
INVX1 INVX1_538 ( .A(REGFILE_SIM_reg_bank_reg_r30_29_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2263_));
INVX1 INVX1_539 ( .A(REGFILE_SIM_reg_bank_reg_r30_30_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2265_));
INVX1 INVX1_54 ( .A(alu_p_o_16_), .Y(_abc_40298_new_n803_));
INVX1 INVX1_540 ( .A(REGFILE_SIM_reg_bank_reg_r30_31_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2267_));
INVX1 INVX1_541 ( .A(REGFILE_SIM_reg_bank_reg_r29_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2269_));
INVX1 INVX1_542 ( .A(REGFILE_SIM_reg_bank_reg_r29_1_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2274_));
INVX1 INVX1_543 ( .A(REGFILE_SIM_reg_bank_reg_r29_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2276_));
INVX1 INVX1_544 ( .A(REGFILE_SIM_reg_bank_reg_r29_3_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2278_));
INVX1 INVX1_545 ( .A(REGFILE_SIM_reg_bank_reg_r29_4_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2280_));
INVX1 INVX1_546 ( .A(REGFILE_SIM_reg_bank_reg_r29_5_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2282_));
INVX1 INVX1_547 ( .A(REGFILE_SIM_reg_bank_reg_r29_6_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2284_));
INVX1 INVX1_548 ( .A(REGFILE_SIM_reg_bank_reg_r29_7_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2286_));
INVX1 INVX1_549 ( .A(REGFILE_SIM_reg_bank_reg_r29_8_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2288_));
INVX1 INVX1_55 ( .A(\mem_dat_i[16] ), .Y(_abc_40298_new_n805_));
INVX1 INVX1_550 ( .A(REGFILE_SIM_reg_bank_reg_r29_9_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2290_));
INVX1 INVX1_551 ( .A(REGFILE_SIM_reg_bank_reg_r29_10_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2292_));
INVX1 INVX1_552 ( .A(REGFILE_SIM_reg_bank_reg_r29_11_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2294_));
INVX1 INVX1_553 ( .A(REGFILE_SIM_reg_bank_reg_r29_12_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2296_));
INVX1 INVX1_554 ( .A(REGFILE_SIM_reg_bank_reg_r29_13_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2298_));
INVX1 INVX1_555 ( .A(REGFILE_SIM_reg_bank_reg_r29_14_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2300_));
INVX1 INVX1_556 ( .A(REGFILE_SIM_reg_bank_reg_r29_15_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2302_));
INVX1 INVX1_557 ( .A(REGFILE_SIM_reg_bank_reg_r29_16_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2304_));
INVX1 INVX1_558 ( .A(REGFILE_SIM_reg_bank_reg_r29_17_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2306_));
INVX1 INVX1_559 ( .A(REGFILE_SIM_reg_bank_reg_r29_18_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2308_));
INVX1 INVX1_56 ( .A(alu_p_o_17_), .Y(_abc_40298_new_n809_));
INVX1 INVX1_560 ( .A(REGFILE_SIM_reg_bank_reg_r29_19_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2310_));
INVX1 INVX1_561 ( .A(REGFILE_SIM_reg_bank_reg_r29_20_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2312_));
INVX1 INVX1_562 ( .A(REGFILE_SIM_reg_bank_reg_r29_21_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2314_));
INVX1 INVX1_563 ( .A(REGFILE_SIM_reg_bank_reg_r29_22_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2316_));
INVX1 INVX1_564 ( .A(REGFILE_SIM_reg_bank_reg_r29_23_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2318_));
INVX1 INVX1_565 ( .A(REGFILE_SIM_reg_bank_reg_r29_24_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2320_));
INVX1 INVX1_566 ( .A(REGFILE_SIM_reg_bank_reg_r29_25_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2322_));
INVX1 INVX1_567 ( .A(REGFILE_SIM_reg_bank_reg_r29_26_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2324_));
INVX1 INVX1_568 ( .A(REGFILE_SIM_reg_bank_reg_r29_27_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2326_));
INVX1 INVX1_569 ( .A(REGFILE_SIM_reg_bank_reg_r29_28_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2328_));
INVX1 INVX1_57 ( .A(\mem_dat_i[17] ), .Y(_abc_40298_new_n810_));
INVX1 INVX1_570 ( .A(REGFILE_SIM_reg_bank_reg_r29_29_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2330_));
INVX1 INVX1_571 ( .A(REGFILE_SIM_reg_bank_reg_r29_30_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2332_));
INVX1 INVX1_572 ( .A(REGFILE_SIM_reg_bank_reg_r29_31_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2334_));
INVX1 INVX1_573 ( .A(REGFILE_SIM_reg_bank_reg_r28_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2336_));
INVX1 INVX1_574 ( .A(REGFILE_SIM_reg_bank_reg_r28_1_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2341_));
INVX1 INVX1_575 ( .A(REGFILE_SIM_reg_bank_reg_r28_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2343_));
INVX1 INVX1_576 ( .A(REGFILE_SIM_reg_bank_reg_r28_3_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2345_));
INVX1 INVX1_577 ( .A(REGFILE_SIM_reg_bank_reg_r28_4_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2347_));
INVX1 INVX1_578 ( .A(REGFILE_SIM_reg_bank_reg_r28_5_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2349_));
INVX1 INVX1_579 ( .A(REGFILE_SIM_reg_bank_reg_r28_6_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2351_));
INVX1 INVX1_58 ( .A(alu_p_o_18_), .Y(_abc_40298_new_n814_));
INVX1 INVX1_580 ( .A(REGFILE_SIM_reg_bank_reg_r28_7_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2353_));
INVX1 INVX1_581 ( .A(REGFILE_SIM_reg_bank_reg_r28_8_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2355_));
INVX1 INVX1_582 ( .A(REGFILE_SIM_reg_bank_reg_r28_9_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2357_));
INVX1 INVX1_583 ( .A(REGFILE_SIM_reg_bank_reg_r28_10_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2359_));
INVX1 INVX1_584 ( .A(REGFILE_SIM_reg_bank_reg_r28_11_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2361_));
INVX1 INVX1_585 ( .A(REGFILE_SIM_reg_bank_reg_r28_12_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2363_));
INVX1 INVX1_586 ( .A(REGFILE_SIM_reg_bank_reg_r28_13_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2365_));
INVX1 INVX1_587 ( .A(REGFILE_SIM_reg_bank_reg_r28_14_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2367_));
INVX1 INVX1_588 ( .A(REGFILE_SIM_reg_bank_reg_r28_15_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2369_));
INVX1 INVX1_589 ( .A(REGFILE_SIM_reg_bank_reg_r28_16_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2371_));
INVX1 INVX1_59 ( .A(\mem_dat_i[18] ), .Y(_abc_40298_new_n815_));
INVX1 INVX1_590 ( .A(REGFILE_SIM_reg_bank_reg_r28_17_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2373_));
INVX1 INVX1_591 ( .A(REGFILE_SIM_reg_bank_reg_r28_18_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2375_));
INVX1 INVX1_592 ( .A(REGFILE_SIM_reg_bank_reg_r28_19_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2377_));
INVX1 INVX1_593 ( .A(REGFILE_SIM_reg_bank_reg_r28_20_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2379_));
INVX1 INVX1_594 ( .A(REGFILE_SIM_reg_bank_reg_r28_21_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2381_));
INVX1 INVX1_595 ( .A(REGFILE_SIM_reg_bank_reg_r28_22_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2383_));
INVX1 INVX1_596 ( .A(REGFILE_SIM_reg_bank_reg_r28_23_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2385_));
INVX1 INVX1_597 ( .A(REGFILE_SIM_reg_bank_reg_r28_24_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2387_));
INVX1 INVX1_598 ( .A(REGFILE_SIM_reg_bank_reg_r28_25_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2389_));
INVX1 INVX1_599 ( .A(REGFILE_SIM_reg_bank_reg_r28_26_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2391_));
INVX1 INVX1_6 ( .A(_abc_40298_new_n628_), .Y(inst_trap_w));
INVX1 INVX1_60 ( .A(alu_p_o_19_), .Y(_abc_40298_new_n819_));
INVX1 INVX1_600 ( .A(REGFILE_SIM_reg_bank_reg_r28_27_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2393_));
INVX1 INVX1_601 ( .A(REGFILE_SIM_reg_bank_reg_r28_28_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2395_));
INVX1 INVX1_602 ( .A(REGFILE_SIM_reg_bank_reg_r28_29_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2397_));
INVX1 INVX1_603 ( .A(REGFILE_SIM_reg_bank_reg_r28_30_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2399_));
INVX1 INVX1_604 ( .A(REGFILE_SIM_reg_bank_reg_r28_31_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2401_));
INVX1 INVX1_605 ( .A(REGFILE_SIM_reg_bank_reg_r27_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2403_));
INVX1 INVX1_606 ( .A(REGFILE_SIM_reg_bank_rd_i_3_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2404_));
INVX1 INVX1_607 ( .A(REGFILE_SIM_reg_bank_reg_r27_1_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2409_));
INVX1 INVX1_608 ( .A(REGFILE_SIM_reg_bank_reg_r27_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2411_));
INVX1 INVX1_609 ( .A(REGFILE_SIM_reg_bank_reg_r27_3_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2413_));
INVX1 INVX1_61 ( .A(\mem_dat_i[19] ), .Y(_abc_40298_new_n820_));
INVX1 INVX1_610 ( .A(REGFILE_SIM_reg_bank_reg_r27_4_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2415_));
INVX1 INVX1_611 ( .A(REGFILE_SIM_reg_bank_reg_r27_5_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2417_));
INVX1 INVX1_612 ( .A(REGFILE_SIM_reg_bank_reg_r27_6_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2419_));
INVX1 INVX1_613 ( .A(REGFILE_SIM_reg_bank_reg_r27_7_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2421_));
INVX1 INVX1_614 ( .A(REGFILE_SIM_reg_bank_reg_r27_8_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2423_));
INVX1 INVX1_615 ( .A(REGFILE_SIM_reg_bank_reg_r27_9_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2425_));
INVX1 INVX1_616 ( .A(REGFILE_SIM_reg_bank_reg_r27_10_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2427_));
INVX1 INVX1_617 ( .A(REGFILE_SIM_reg_bank_reg_r27_11_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2429_));
INVX1 INVX1_618 ( .A(REGFILE_SIM_reg_bank_reg_r27_12_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2431_));
INVX1 INVX1_619 ( .A(REGFILE_SIM_reg_bank_reg_r27_13_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2433_));
INVX1 INVX1_62 ( .A(alu_p_o_20_), .Y(_abc_40298_new_n824_));
INVX1 INVX1_620 ( .A(REGFILE_SIM_reg_bank_reg_r27_14_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2435_));
INVX1 INVX1_621 ( .A(REGFILE_SIM_reg_bank_reg_r27_15_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2437_));
INVX1 INVX1_622 ( .A(REGFILE_SIM_reg_bank_reg_r27_16_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2439_));
INVX1 INVX1_623 ( .A(REGFILE_SIM_reg_bank_reg_r27_17_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2441_));
INVX1 INVX1_624 ( .A(REGFILE_SIM_reg_bank_reg_r27_18_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2443_));
INVX1 INVX1_625 ( .A(REGFILE_SIM_reg_bank_reg_r27_19_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2445_));
INVX1 INVX1_626 ( .A(REGFILE_SIM_reg_bank_reg_r27_20_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2447_));
INVX1 INVX1_627 ( .A(REGFILE_SIM_reg_bank_reg_r27_21_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2449_));
INVX1 INVX1_628 ( .A(REGFILE_SIM_reg_bank_reg_r27_22_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2451_));
INVX1 INVX1_629 ( .A(REGFILE_SIM_reg_bank_reg_r27_23_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2453_));
INVX1 INVX1_63 ( .A(\mem_dat_i[20] ), .Y(_abc_40298_new_n825_));
INVX1 INVX1_630 ( .A(REGFILE_SIM_reg_bank_reg_r27_24_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2455_));
INVX1 INVX1_631 ( .A(REGFILE_SIM_reg_bank_reg_r27_25_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2457_));
INVX1 INVX1_632 ( .A(REGFILE_SIM_reg_bank_reg_r27_26_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2459_));
INVX1 INVX1_633 ( .A(REGFILE_SIM_reg_bank_reg_r27_27_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2461_));
INVX1 INVX1_634 ( .A(REGFILE_SIM_reg_bank_reg_r27_28_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2463_));
INVX1 INVX1_635 ( .A(REGFILE_SIM_reg_bank_reg_r27_29_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2465_));
INVX1 INVX1_636 ( .A(REGFILE_SIM_reg_bank_reg_r27_30_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2467_));
INVX1 INVX1_637 ( .A(REGFILE_SIM_reg_bank_reg_r27_31_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2469_));
INVX1 INVX1_638 ( .A(REGFILE_SIM_reg_bank_reg_r26_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2471_));
INVX1 INVX1_639 ( .A(REGFILE_SIM_reg_bank_reg_r26_1_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2475_));
INVX1 INVX1_64 ( .A(alu_p_o_21_), .Y(_abc_40298_new_n829_));
INVX1 INVX1_640 ( .A(REGFILE_SIM_reg_bank_reg_r26_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2477_));
INVX1 INVX1_641 ( .A(REGFILE_SIM_reg_bank_reg_r26_3_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2479_));
INVX1 INVX1_642 ( .A(REGFILE_SIM_reg_bank_reg_r26_4_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2481_));
INVX1 INVX1_643 ( .A(REGFILE_SIM_reg_bank_reg_r26_5_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2483_));
INVX1 INVX1_644 ( .A(REGFILE_SIM_reg_bank_reg_r26_6_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2485_));
INVX1 INVX1_645 ( .A(REGFILE_SIM_reg_bank_reg_r26_7_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2487_));
INVX1 INVX1_646 ( .A(REGFILE_SIM_reg_bank_reg_r26_8_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2489_));
INVX1 INVX1_647 ( .A(REGFILE_SIM_reg_bank_reg_r26_9_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2491_));
INVX1 INVX1_648 ( .A(REGFILE_SIM_reg_bank_reg_r26_10_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2493_));
INVX1 INVX1_649 ( .A(REGFILE_SIM_reg_bank_reg_r26_11_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2495_));
INVX1 INVX1_65 ( .A(\mem_dat_i[21] ), .Y(_abc_40298_new_n830_));
INVX1 INVX1_650 ( .A(REGFILE_SIM_reg_bank_reg_r26_12_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2497_));
INVX1 INVX1_651 ( .A(REGFILE_SIM_reg_bank_reg_r26_13_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2499_));
INVX1 INVX1_652 ( .A(REGFILE_SIM_reg_bank_reg_r26_14_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2501_));
INVX1 INVX1_653 ( .A(REGFILE_SIM_reg_bank_reg_r26_15_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2503_));
INVX1 INVX1_654 ( .A(REGFILE_SIM_reg_bank_reg_r26_16_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2505_));
INVX1 INVX1_655 ( .A(REGFILE_SIM_reg_bank_reg_r26_17_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2507_));
INVX1 INVX1_656 ( .A(REGFILE_SIM_reg_bank_reg_r26_18_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2509_));
INVX1 INVX1_657 ( .A(REGFILE_SIM_reg_bank_reg_r26_19_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2511_));
INVX1 INVX1_658 ( .A(REGFILE_SIM_reg_bank_reg_r26_20_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2513_));
INVX1 INVX1_659 ( .A(REGFILE_SIM_reg_bank_reg_r26_21_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2515_));
INVX1 INVX1_66 ( .A(alu_p_o_22_), .Y(_abc_40298_new_n834_));
INVX1 INVX1_660 ( .A(REGFILE_SIM_reg_bank_reg_r26_22_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2517_));
INVX1 INVX1_661 ( .A(REGFILE_SIM_reg_bank_reg_r26_23_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2519_));
INVX1 INVX1_662 ( .A(REGFILE_SIM_reg_bank_reg_r26_24_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2521_));
INVX1 INVX1_663 ( .A(REGFILE_SIM_reg_bank_reg_r26_25_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2523_));
INVX1 INVX1_664 ( .A(REGFILE_SIM_reg_bank_reg_r26_26_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2525_));
INVX1 INVX1_665 ( .A(REGFILE_SIM_reg_bank_reg_r26_27_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2527_));
INVX1 INVX1_666 ( .A(REGFILE_SIM_reg_bank_reg_r26_28_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2529_));
INVX1 INVX1_667 ( .A(REGFILE_SIM_reg_bank_reg_r26_29_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2531_));
INVX1 INVX1_668 ( .A(REGFILE_SIM_reg_bank_reg_r26_30_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2533_));
INVX1 INVX1_669 ( .A(REGFILE_SIM_reg_bank_reg_r26_31_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2535_));
INVX1 INVX1_67 ( .A(\mem_dat_i[22] ), .Y(_abc_40298_new_n835_));
INVX1 INVX1_670 ( .A(REGFILE_SIM_reg_bank_reg_r25_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2537_));
INVX1 INVX1_671 ( .A(REGFILE_SIM_reg_bank_reg_r25_1_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2541_));
INVX1 INVX1_672 ( .A(REGFILE_SIM_reg_bank_reg_r25_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2543_));
INVX1 INVX1_673 ( .A(REGFILE_SIM_reg_bank_reg_r25_3_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2545_));
INVX1 INVX1_674 ( .A(REGFILE_SIM_reg_bank_reg_r25_4_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2547_));
INVX1 INVX1_675 ( .A(REGFILE_SIM_reg_bank_reg_r25_5_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2549_));
INVX1 INVX1_676 ( .A(REGFILE_SIM_reg_bank_reg_r25_6_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2551_));
INVX1 INVX1_677 ( .A(REGFILE_SIM_reg_bank_reg_r25_7_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2553_));
INVX1 INVX1_678 ( .A(REGFILE_SIM_reg_bank_reg_r25_8_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2555_));
INVX1 INVX1_679 ( .A(REGFILE_SIM_reg_bank_reg_r25_9_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2557_));
INVX1 INVX1_68 ( .A(alu_p_o_23_), .Y(_abc_40298_new_n839_));
INVX1 INVX1_680 ( .A(REGFILE_SIM_reg_bank_reg_r25_10_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2559_));
INVX1 INVX1_681 ( .A(REGFILE_SIM_reg_bank_reg_r25_11_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2561_));
INVX1 INVX1_682 ( .A(REGFILE_SIM_reg_bank_reg_r25_12_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2563_));
INVX1 INVX1_683 ( .A(REGFILE_SIM_reg_bank_reg_r25_13_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2565_));
INVX1 INVX1_684 ( .A(REGFILE_SIM_reg_bank_reg_r25_14_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2567_));
INVX1 INVX1_685 ( .A(REGFILE_SIM_reg_bank_reg_r25_15_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2569_));
INVX1 INVX1_686 ( .A(REGFILE_SIM_reg_bank_reg_r25_16_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2571_));
INVX1 INVX1_687 ( .A(REGFILE_SIM_reg_bank_reg_r25_17_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2573_));
INVX1 INVX1_688 ( .A(REGFILE_SIM_reg_bank_reg_r25_18_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2575_));
INVX1 INVX1_689 ( .A(REGFILE_SIM_reg_bank_reg_r25_19_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2577_));
INVX1 INVX1_69 ( .A(\mem_dat_i[23] ), .Y(_abc_40298_new_n840_));
INVX1 INVX1_690 ( .A(REGFILE_SIM_reg_bank_reg_r25_20_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2579_));
INVX1 INVX1_691 ( .A(REGFILE_SIM_reg_bank_reg_r25_21_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2581_));
INVX1 INVX1_692 ( .A(REGFILE_SIM_reg_bank_reg_r25_22_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2583_));
INVX1 INVX1_693 ( .A(REGFILE_SIM_reg_bank_reg_r25_23_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2585_));
INVX1 INVX1_694 ( .A(REGFILE_SIM_reg_bank_reg_r25_24_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2587_));
INVX1 INVX1_695 ( .A(REGFILE_SIM_reg_bank_reg_r25_25_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2589_));
INVX1 INVX1_696 ( .A(REGFILE_SIM_reg_bank_reg_r25_26_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2591_));
INVX1 INVX1_697 ( .A(REGFILE_SIM_reg_bank_reg_r25_27_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2593_));
INVX1 INVX1_698 ( .A(REGFILE_SIM_reg_bank_reg_r25_28_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2595_));
INVX1 INVX1_699 ( .A(REGFILE_SIM_reg_bank_reg_r25_29_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2597_));
INVX1 INVX1_7 ( .A(mem_ack_i), .Y(_abc_40298_new_n630_));
INVX1 INVX1_70 ( .A(alu_p_o_24_), .Y(_abc_40298_new_n844_));
INVX1 INVX1_700 ( .A(REGFILE_SIM_reg_bank_reg_r25_30_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2599_));
INVX1 INVX1_701 ( .A(REGFILE_SIM_reg_bank_reg_r25_31_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2601_));
INVX1 INVX1_702 ( .A(REGFILE_SIM_reg_bank_reg_r23_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2668_));
INVX1 INVX1_703 ( .A(REGFILE_SIM_reg_bank_reg_r23_1_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2673_));
INVX1 INVX1_704 ( .A(REGFILE_SIM_reg_bank_reg_r23_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2675_));
INVX1 INVX1_705 ( .A(REGFILE_SIM_reg_bank_reg_r23_3_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2677_));
INVX1 INVX1_706 ( .A(REGFILE_SIM_reg_bank_reg_r23_4_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2679_));
INVX1 INVX1_707 ( .A(REGFILE_SIM_reg_bank_reg_r23_5_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2681_));
INVX1 INVX1_708 ( .A(REGFILE_SIM_reg_bank_reg_r23_6_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2683_));
INVX1 INVX1_709 ( .A(REGFILE_SIM_reg_bank_reg_r23_7_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2685_));
INVX1 INVX1_71 ( .A(\mem_dat_i[24] ), .Y(_abc_40298_new_n845_));
INVX1 INVX1_710 ( .A(REGFILE_SIM_reg_bank_reg_r23_8_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2687_));
INVX1 INVX1_711 ( .A(REGFILE_SIM_reg_bank_reg_r23_9_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2689_));
INVX1 INVX1_712 ( .A(REGFILE_SIM_reg_bank_reg_r23_10_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2691_));
INVX1 INVX1_713 ( .A(REGFILE_SIM_reg_bank_reg_r23_11_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2693_));
INVX1 INVX1_714 ( .A(REGFILE_SIM_reg_bank_reg_r23_12_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2695_));
INVX1 INVX1_715 ( .A(REGFILE_SIM_reg_bank_reg_r23_13_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2697_));
INVX1 INVX1_716 ( .A(REGFILE_SIM_reg_bank_reg_r23_14_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2699_));
INVX1 INVX1_717 ( .A(REGFILE_SIM_reg_bank_reg_r23_15_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2701_));
INVX1 INVX1_718 ( .A(REGFILE_SIM_reg_bank_reg_r23_16_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2703_));
INVX1 INVX1_719 ( .A(REGFILE_SIM_reg_bank_reg_r23_17_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2705_));
INVX1 INVX1_72 ( .A(alu_p_o_25_), .Y(_abc_40298_new_n849_));
INVX1 INVX1_720 ( .A(REGFILE_SIM_reg_bank_reg_r23_18_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2707_));
INVX1 INVX1_721 ( .A(REGFILE_SIM_reg_bank_reg_r23_19_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2709_));
INVX1 INVX1_722 ( .A(REGFILE_SIM_reg_bank_reg_r23_20_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2711_));
INVX1 INVX1_723 ( .A(REGFILE_SIM_reg_bank_reg_r23_21_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2713_));
INVX1 INVX1_724 ( .A(REGFILE_SIM_reg_bank_reg_r23_22_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2715_));
INVX1 INVX1_725 ( .A(REGFILE_SIM_reg_bank_reg_r23_23_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2717_));
INVX1 INVX1_726 ( .A(REGFILE_SIM_reg_bank_reg_r23_24_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2719_));
INVX1 INVX1_727 ( .A(REGFILE_SIM_reg_bank_reg_r23_25_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2721_));
INVX1 INVX1_728 ( .A(REGFILE_SIM_reg_bank_reg_r23_26_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2723_));
INVX1 INVX1_729 ( .A(REGFILE_SIM_reg_bank_reg_r23_27_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2725_));
INVX1 INVX1_73 ( .A(\mem_dat_i[25] ), .Y(_abc_40298_new_n850_));
INVX1 INVX1_730 ( .A(REGFILE_SIM_reg_bank_reg_r23_28_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2727_));
INVX1 INVX1_731 ( .A(REGFILE_SIM_reg_bank_reg_r23_29_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2729_));
INVX1 INVX1_732 ( .A(REGFILE_SIM_reg_bank_reg_r23_30_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2731_));
INVX1 INVX1_733 ( .A(REGFILE_SIM_reg_bank_reg_r23_31_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2733_));
INVX1 INVX1_734 ( .A(REGFILE_SIM_reg_bank_reg_r22_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2735_));
INVX1 INVX1_735 ( .A(REGFILE_SIM_reg_bank_reg_r22_1_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2739_));
INVX1 INVX1_736 ( .A(REGFILE_SIM_reg_bank_reg_r22_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2741_));
INVX1 INVX1_737 ( .A(REGFILE_SIM_reg_bank_reg_r22_3_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2743_));
INVX1 INVX1_738 ( .A(REGFILE_SIM_reg_bank_reg_r22_4_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2745_));
INVX1 INVX1_739 ( .A(REGFILE_SIM_reg_bank_reg_r22_5_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2747_));
INVX1 INVX1_74 ( .A(alu_p_o_26_), .Y(_abc_40298_new_n854_));
INVX1 INVX1_740 ( .A(REGFILE_SIM_reg_bank_reg_r22_6_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2749_));
INVX1 INVX1_741 ( .A(REGFILE_SIM_reg_bank_reg_r22_7_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2751_));
INVX1 INVX1_742 ( .A(REGFILE_SIM_reg_bank_reg_r22_8_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2753_));
INVX1 INVX1_743 ( .A(REGFILE_SIM_reg_bank_reg_r22_9_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2755_));
INVX1 INVX1_744 ( .A(REGFILE_SIM_reg_bank_reg_r22_10_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2757_));
INVX1 INVX1_745 ( .A(REGFILE_SIM_reg_bank_reg_r22_11_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2759_));
INVX1 INVX1_746 ( .A(REGFILE_SIM_reg_bank_reg_r22_12_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2761_));
INVX1 INVX1_747 ( .A(REGFILE_SIM_reg_bank_reg_r22_13_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2763_));
INVX1 INVX1_748 ( .A(REGFILE_SIM_reg_bank_reg_r22_14_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2765_));
INVX1 INVX1_749 ( .A(REGFILE_SIM_reg_bank_reg_r22_15_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2767_));
INVX1 INVX1_75 ( .A(\mem_dat_i[26] ), .Y(_abc_40298_new_n855_));
INVX1 INVX1_750 ( .A(REGFILE_SIM_reg_bank_reg_r22_16_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2769_));
INVX1 INVX1_751 ( .A(REGFILE_SIM_reg_bank_reg_r22_17_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2771_));
INVX1 INVX1_752 ( .A(REGFILE_SIM_reg_bank_reg_r22_18_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2773_));
INVX1 INVX1_753 ( .A(REGFILE_SIM_reg_bank_reg_r22_19_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2775_));
INVX1 INVX1_754 ( .A(REGFILE_SIM_reg_bank_reg_r22_20_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2777_));
INVX1 INVX1_755 ( .A(REGFILE_SIM_reg_bank_reg_r22_21_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2779_));
INVX1 INVX1_756 ( .A(REGFILE_SIM_reg_bank_reg_r22_22_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2781_));
INVX1 INVX1_757 ( .A(REGFILE_SIM_reg_bank_reg_r22_23_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2783_));
INVX1 INVX1_758 ( .A(REGFILE_SIM_reg_bank_reg_r22_24_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2785_));
INVX1 INVX1_759 ( .A(REGFILE_SIM_reg_bank_reg_r22_25_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2787_));
INVX1 INVX1_76 ( .A(alu_p_o_27_), .Y(_abc_40298_new_n859_));
INVX1 INVX1_760 ( .A(REGFILE_SIM_reg_bank_reg_r22_26_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2789_));
INVX1 INVX1_761 ( .A(REGFILE_SIM_reg_bank_reg_r22_27_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2791_));
INVX1 INVX1_762 ( .A(REGFILE_SIM_reg_bank_reg_r22_28_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2793_));
INVX1 INVX1_763 ( .A(REGFILE_SIM_reg_bank_reg_r22_29_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2795_));
INVX1 INVX1_764 ( .A(REGFILE_SIM_reg_bank_reg_r22_30_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2797_));
INVX1 INVX1_765 ( .A(REGFILE_SIM_reg_bank_reg_r22_31_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2799_));
INVX1 INVX1_766 ( .A(REGFILE_SIM_reg_bank_reg_r21_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2801_));
INVX1 INVX1_767 ( .A(REGFILE_SIM_reg_bank_reg_r21_1_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2805_));
INVX1 INVX1_768 ( .A(REGFILE_SIM_reg_bank_reg_r21_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2807_));
INVX1 INVX1_769 ( .A(REGFILE_SIM_reg_bank_reg_r21_3_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2809_));
INVX1 INVX1_77 ( .A(\mem_dat_i[27] ), .Y(_abc_40298_new_n860_));
INVX1 INVX1_770 ( .A(REGFILE_SIM_reg_bank_reg_r21_4_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2811_));
INVX1 INVX1_771 ( .A(REGFILE_SIM_reg_bank_reg_r21_5_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2813_));
INVX1 INVX1_772 ( .A(REGFILE_SIM_reg_bank_reg_r21_6_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2815_));
INVX1 INVX1_773 ( .A(REGFILE_SIM_reg_bank_reg_r21_7_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2817_));
INVX1 INVX1_774 ( .A(REGFILE_SIM_reg_bank_reg_r21_8_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2819_));
INVX1 INVX1_775 ( .A(REGFILE_SIM_reg_bank_reg_r21_9_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2821_));
INVX1 INVX1_776 ( .A(REGFILE_SIM_reg_bank_reg_r21_10_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2823_));
INVX1 INVX1_777 ( .A(REGFILE_SIM_reg_bank_reg_r21_11_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2825_));
INVX1 INVX1_778 ( .A(REGFILE_SIM_reg_bank_reg_r21_12_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2827_));
INVX1 INVX1_779 ( .A(REGFILE_SIM_reg_bank_reg_r21_13_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2829_));
INVX1 INVX1_78 ( .A(alu_p_o_28_), .Y(_abc_40298_new_n864_));
INVX1 INVX1_780 ( .A(REGFILE_SIM_reg_bank_reg_r21_14_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2831_));
INVX1 INVX1_781 ( .A(REGFILE_SIM_reg_bank_reg_r21_15_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2833_));
INVX1 INVX1_782 ( .A(REGFILE_SIM_reg_bank_reg_r21_16_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2835_));
INVX1 INVX1_783 ( .A(REGFILE_SIM_reg_bank_reg_r21_17_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2837_));
INVX1 INVX1_784 ( .A(REGFILE_SIM_reg_bank_reg_r21_18_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2839_));
INVX1 INVX1_785 ( .A(REGFILE_SIM_reg_bank_reg_r21_19_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2841_));
INVX1 INVX1_786 ( .A(REGFILE_SIM_reg_bank_reg_r21_20_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2843_));
INVX1 INVX1_787 ( .A(REGFILE_SIM_reg_bank_reg_r21_21_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2845_));
INVX1 INVX1_788 ( .A(REGFILE_SIM_reg_bank_reg_r21_22_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2847_));
INVX1 INVX1_789 ( .A(REGFILE_SIM_reg_bank_reg_r21_23_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2849_));
INVX1 INVX1_79 ( .A(\mem_dat_i[28] ), .Y(_abc_40298_new_n865_));
INVX1 INVX1_790 ( .A(REGFILE_SIM_reg_bank_reg_r21_24_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2851_));
INVX1 INVX1_791 ( .A(REGFILE_SIM_reg_bank_reg_r21_25_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2853_));
INVX1 INVX1_792 ( .A(REGFILE_SIM_reg_bank_reg_r21_26_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2855_));
INVX1 INVX1_793 ( .A(REGFILE_SIM_reg_bank_reg_r21_27_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2857_));
INVX1 INVX1_794 ( .A(REGFILE_SIM_reg_bank_reg_r21_28_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2859_));
INVX1 INVX1_795 ( .A(REGFILE_SIM_reg_bank_reg_r21_29_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2861_));
INVX1 INVX1_796 ( .A(REGFILE_SIM_reg_bank_reg_r21_30_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2863_));
INVX1 INVX1_797 ( .A(REGFILE_SIM_reg_bank_reg_r21_31_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2865_));
INVX1 INVX1_798 ( .A(REGFILE_SIM_reg_bank_reg_r20_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2867_));
INVX1 INVX1_799 ( .A(REGFILE_SIM_reg_bank_reg_r20_1_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2870_));
INVX1 INVX1_8 ( .A(state_q_1_), .Y(_abc_40298_new_n631_));
INVX1 INVX1_80 ( .A(alu_p_o_29_), .Y(_abc_40298_new_n869_));
INVX1 INVX1_800 ( .A(REGFILE_SIM_reg_bank_reg_r20_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2872_));
INVX1 INVX1_801 ( .A(REGFILE_SIM_reg_bank_reg_r20_3_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2874_));
INVX1 INVX1_802 ( .A(REGFILE_SIM_reg_bank_reg_r20_4_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2876_));
INVX1 INVX1_803 ( .A(REGFILE_SIM_reg_bank_reg_r20_5_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2878_));
INVX1 INVX1_804 ( .A(REGFILE_SIM_reg_bank_reg_r20_6_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2880_));
INVX1 INVX1_805 ( .A(REGFILE_SIM_reg_bank_reg_r20_7_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2882_));
INVX1 INVX1_806 ( .A(REGFILE_SIM_reg_bank_reg_r20_8_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2884_));
INVX1 INVX1_807 ( .A(REGFILE_SIM_reg_bank_reg_r20_9_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2886_));
INVX1 INVX1_808 ( .A(REGFILE_SIM_reg_bank_reg_r20_10_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2888_));
INVX1 INVX1_809 ( .A(REGFILE_SIM_reg_bank_reg_r20_11_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2890_));
INVX1 INVX1_81 ( .A(\mem_dat_i[29] ), .Y(_abc_40298_new_n870_));
INVX1 INVX1_810 ( .A(REGFILE_SIM_reg_bank_reg_r20_12_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2892_));
INVX1 INVX1_811 ( .A(REGFILE_SIM_reg_bank_reg_r20_13_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2894_));
INVX1 INVX1_812 ( .A(REGFILE_SIM_reg_bank_reg_r20_14_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2896_));
INVX1 INVX1_813 ( .A(REGFILE_SIM_reg_bank_reg_r20_15_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2898_));
INVX1 INVX1_814 ( .A(REGFILE_SIM_reg_bank_reg_r20_16_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2900_));
INVX1 INVX1_815 ( .A(REGFILE_SIM_reg_bank_reg_r20_17_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2902_));
INVX1 INVX1_816 ( .A(REGFILE_SIM_reg_bank_reg_r20_18_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2904_));
INVX1 INVX1_817 ( .A(REGFILE_SIM_reg_bank_reg_r20_19_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2906_));
INVX1 INVX1_818 ( .A(REGFILE_SIM_reg_bank_reg_r20_20_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2908_));
INVX1 INVX1_819 ( .A(REGFILE_SIM_reg_bank_reg_r20_21_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2910_));
INVX1 INVX1_82 ( .A(alu_p_o_30_), .Y(_abc_40298_new_n874_));
INVX1 INVX1_820 ( .A(REGFILE_SIM_reg_bank_reg_r20_22_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2912_));
INVX1 INVX1_821 ( .A(REGFILE_SIM_reg_bank_reg_r20_23_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2914_));
INVX1 INVX1_822 ( .A(REGFILE_SIM_reg_bank_reg_r20_24_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2916_));
INVX1 INVX1_823 ( .A(REGFILE_SIM_reg_bank_reg_r20_25_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2918_));
INVX1 INVX1_824 ( .A(REGFILE_SIM_reg_bank_reg_r20_26_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2920_));
INVX1 INVX1_825 ( .A(REGFILE_SIM_reg_bank_reg_r20_27_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2922_));
INVX1 INVX1_826 ( .A(REGFILE_SIM_reg_bank_reg_r20_28_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2924_));
INVX1 INVX1_827 ( .A(REGFILE_SIM_reg_bank_reg_r20_29_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2926_));
INVX1 INVX1_828 ( .A(REGFILE_SIM_reg_bank_reg_r20_30_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2928_));
INVX1 INVX1_829 ( .A(REGFILE_SIM_reg_bank_reg_r20_31_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2930_));
INVX1 INVX1_83 ( .A(\mem_dat_i[30] ), .Y(_abc_40298_new_n875_));
INVX1 INVX1_830 ( .A(REGFILE_SIM_reg_bank_reg_r19_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2932_));
INVX1 INVX1_831 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2933_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2934_));
INVX1 INVX1_832 ( .A(REGFILE_SIM_reg_bank_reg_r19_1_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2938_));
INVX1 INVX1_833 ( .A(REGFILE_SIM_reg_bank_reg_r19_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2940_));
INVX1 INVX1_834 ( .A(REGFILE_SIM_reg_bank_reg_r19_3_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2942_));
INVX1 INVX1_835 ( .A(REGFILE_SIM_reg_bank_reg_r19_4_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2944_));
INVX1 INVX1_836 ( .A(REGFILE_SIM_reg_bank_reg_r19_5_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2946_));
INVX1 INVX1_837 ( .A(REGFILE_SIM_reg_bank_reg_r19_6_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2948_));
INVX1 INVX1_838 ( .A(REGFILE_SIM_reg_bank_reg_r19_7_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2950_));
INVX1 INVX1_839 ( .A(REGFILE_SIM_reg_bank_reg_r19_8_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2952_));
INVX1 INVX1_84 ( .A(alu_p_o_31_), .Y(_abc_40298_new_n879_));
INVX1 INVX1_840 ( .A(REGFILE_SIM_reg_bank_reg_r19_9_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2954_));
INVX1 INVX1_841 ( .A(REGFILE_SIM_reg_bank_reg_r19_10_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2956_));
INVX1 INVX1_842 ( .A(REGFILE_SIM_reg_bank_reg_r19_11_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2958_));
INVX1 INVX1_843 ( .A(REGFILE_SIM_reg_bank_reg_r19_12_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2960_));
INVX1 INVX1_844 ( .A(REGFILE_SIM_reg_bank_reg_r19_13_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2962_));
INVX1 INVX1_845 ( .A(REGFILE_SIM_reg_bank_reg_r19_14_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2964_));
INVX1 INVX1_846 ( .A(REGFILE_SIM_reg_bank_reg_r19_15_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2966_));
INVX1 INVX1_847 ( .A(REGFILE_SIM_reg_bank_reg_r19_16_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2968_));
INVX1 INVX1_848 ( .A(REGFILE_SIM_reg_bank_reg_r19_17_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2970_));
INVX1 INVX1_849 ( .A(REGFILE_SIM_reg_bank_reg_r19_18_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2972_));
INVX1 INVX1_85 ( .A(\mem_dat_i[31] ), .Y(_abc_40298_new_n880_));
INVX1 INVX1_850 ( .A(REGFILE_SIM_reg_bank_reg_r19_19_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2974_));
INVX1 INVX1_851 ( .A(REGFILE_SIM_reg_bank_reg_r19_20_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2976_));
INVX1 INVX1_852 ( .A(REGFILE_SIM_reg_bank_reg_r19_21_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2978_));
INVX1 INVX1_853 ( .A(REGFILE_SIM_reg_bank_reg_r19_22_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2980_));
INVX1 INVX1_854 ( .A(REGFILE_SIM_reg_bank_reg_r19_23_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2982_));
INVX1 INVX1_855 ( .A(REGFILE_SIM_reg_bank_reg_r19_24_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2984_));
INVX1 INVX1_856 ( .A(REGFILE_SIM_reg_bank_reg_r19_25_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2986_));
INVX1 INVX1_857 ( .A(REGFILE_SIM_reg_bank_reg_r19_26_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2988_));
INVX1 INVX1_858 ( .A(REGFILE_SIM_reg_bank_reg_r19_27_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2990_));
INVX1 INVX1_859 ( .A(REGFILE_SIM_reg_bank_reg_r19_28_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2992_));
INVX1 INVX1_86 ( .A(_abc_40298_new_n887_), .Y(_abc_40298_new_n888_));
INVX1 INVX1_860 ( .A(REGFILE_SIM_reg_bank_reg_r19_29_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2994_));
INVX1 INVX1_861 ( .A(REGFILE_SIM_reg_bank_reg_r19_30_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2996_));
INVX1 INVX1_862 ( .A(REGFILE_SIM_reg_bank_reg_r19_31_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2998_));
INVX1 INVX1_863 ( .A(REGFILE_SIM_reg_bank_reg_r18_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3000_));
INVX1 INVX1_864 ( .A(REGFILE_SIM_reg_bank_reg_r18_1_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3004_));
INVX1 INVX1_865 ( .A(REGFILE_SIM_reg_bank_reg_r18_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3006_));
INVX1 INVX1_866 ( .A(REGFILE_SIM_reg_bank_reg_r18_3_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3008_));
INVX1 INVX1_867 ( .A(REGFILE_SIM_reg_bank_reg_r18_4_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3010_));
INVX1 INVX1_868 ( .A(REGFILE_SIM_reg_bank_reg_r18_5_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3012_));
INVX1 INVX1_869 ( .A(REGFILE_SIM_reg_bank_reg_r18_6_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3014_));
INVX1 INVX1_87 ( .A(_abc_40298_new_n891_), .Y(_abc_40298_new_n892_));
INVX1 INVX1_870 ( .A(REGFILE_SIM_reg_bank_reg_r18_7_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3016_));
INVX1 INVX1_871 ( .A(REGFILE_SIM_reg_bank_reg_r18_8_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3018_));
INVX1 INVX1_872 ( .A(REGFILE_SIM_reg_bank_reg_r18_9_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3020_));
INVX1 INVX1_873 ( .A(REGFILE_SIM_reg_bank_reg_r18_10_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3022_));
INVX1 INVX1_874 ( .A(REGFILE_SIM_reg_bank_reg_r18_11_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3024_));
INVX1 INVX1_875 ( .A(REGFILE_SIM_reg_bank_reg_r18_12_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3026_));
INVX1 INVX1_876 ( .A(REGFILE_SIM_reg_bank_reg_r18_13_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3028_));
INVX1 INVX1_877 ( .A(REGFILE_SIM_reg_bank_reg_r18_14_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3030_));
INVX1 INVX1_878 ( .A(REGFILE_SIM_reg_bank_reg_r18_15_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3032_));
INVX1 INVX1_879 ( .A(REGFILE_SIM_reg_bank_reg_r18_16_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3034_));
INVX1 INVX1_88 ( .A(_abc_40298_new_n894_), .Y(_abc_40298_new_n895_));
INVX1 INVX1_880 ( .A(REGFILE_SIM_reg_bank_reg_r18_17_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3036_));
INVX1 INVX1_881 ( .A(REGFILE_SIM_reg_bank_reg_r18_18_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3038_));
INVX1 INVX1_882 ( .A(REGFILE_SIM_reg_bank_reg_r18_19_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3040_));
INVX1 INVX1_883 ( .A(REGFILE_SIM_reg_bank_reg_r18_20_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3042_));
INVX1 INVX1_884 ( .A(REGFILE_SIM_reg_bank_reg_r18_21_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3044_));
INVX1 INVX1_885 ( .A(REGFILE_SIM_reg_bank_reg_r18_22_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3046_));
INVX1 INVX1_886 ( .A(REGFILE_SIM_reg_bank_reg_r18_23_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3048_));
INVX1 INVX1_887 ( .A(REGFILE_SIM_reg_bank_reg_r18_24_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3050_));
INVX1 INVX1_888 ( .A(REGFILE_SIM_reg_bank_reg_r18_25_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3052_));
INVX1 INVX1_889 ( .A(REGFILE_SIM_reg_bank_reg_r18_26_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3054_));
INVX1 INVX1_89 ( .A(alu_op_r_2_), .Y(_abc_40298_new_n898_));
INVX1 INVX1_890 ( .A(REGFILE_SIM_reg_bank_reg_r18_27_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3056_));
INVX1 INVX1_891 ( .A(REGFILE_SIM_reg_bank_reg_r18_28_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3058_));
INVX1 INVX1_892 ( .A(REGFILE_SIM_reg_bank_reg_r18_29_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3060_));
INVX1 INVX1_893 ( .A(REGFILE_SIM_reg_bank_reg_r18_30_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3062_));
INVX1 INVX1_894 ( .A(REGFILE_SIM_reg_bank_reg_r18_31_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3064_));
INVX1 INVX1_895 ( .A(REGFILE_SIM_reg_bank_reg_r17_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3066_));
INVX1 INVX1_896 ( .A(REGFILE_SIM_reg_bank_reg_r17_1_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3070_));
INVX1 INVX1_897 ( .A(REGFILE_SIM_reg_bank_reg_r17_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3072_));
INVX1 INVX1_898 ( .A(REGFILE_SIM_reg_bank_reg_r17_3_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3074_));
INVX1 INVX1_899 ( .A(REGFILE_SIM_reg_bank_reg_r17_4_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3076_));
INVX1 INVX1_9 ( .A(state_q_4_), .Y(_abc_40298_new_n634_));
INVX1 INVX1_90 ( .A(alu_op_r_3_), .Y(_abc_40298_new_n903_));
INVX1 INVX1_900 ( .A(REGFILE_SIM_reg_bank_reg_r17_5_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3078_));
INVX1 INVX1_901 ( .A(REGFILE_SIM_reg_bank_reg_r17_6_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3080_));
INVX1 INVX1_902 ( .A(REGFILE_SIM_reg_bank_reg_r17_7_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3082_));
INVX1 INVX1_903 ( .A(REGFILE_SIM_reg_bank_reg_r17_8_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3084_));
INVX1 INVX1_904 ( .A(REGFILE_SIM_reg_bank_reg_r17_9_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3086_));
INVX1 INVX1_905 ( .A(REGFILE_SIM_reg_bank_reg_r17_10_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3088_));
INVX1 INVX1_906 ( .A(REGFILE_SIM_reg_bank_reg_r17_11_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3090_));
INVX1 INVX1_907 ( .A(REGFILE_SIM_reg_bank_reg_r17_12_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3092_));
INVX1 INVX1_908 ( .A(REGFILE_SIM_reg_bank_reg_r17_13_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3094_));
INVX1 INVX1_909 ( .A(REGFILE_SIM_reg_bank_reg_r17_14_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3096_));
INVX1 INVX1_91 ( .A(_abc_40298_new_n897_), .Y(_abc_40298_new_n906_));
INVX1 INVX1_910 ( .A(REGFILE_SIM_reg_bank_reg_r17_15_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3098_));
INVX1 INVX1_911 ( .A(REGFILE_SIM_reg_bank_reg_r17_16_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3100_));
INVX1 INVX1_912 ( .A(REGFILE_SIM_reg_bank_reg_r17_17_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3102_));
INVX1 INVX1_913 ( .A(REGFILE_SIM_reg_bank_reg_r17_18_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3104_));
INVX1 INVX1_914 ( .A(REGFILE_SIM_reg_bank_reg_r17_19_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3106_));
INVX1 INVX1_915 ( .A(REGFILE_SIM_reg_bank_reg_r17_20_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3108_));
INVX1 INVX1_916 ( .A(REGFILE_SIM_reg_bank_reg_r17_21_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3110_));
INVX1 INVX1_917 ( .A(REGFILE_SIM_reg_bank_reg_r17_22_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3112_));
INVX1 INVX1_918 ( .A(REGFILE_SIM_reg_bank_reg_r17_23_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3114_));
INVX1 INVX1_919 ( .A(REGFILE_SIM_reg_bank_reg_r17_24_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3116_));
INVX1 INVX1_92 ( .A(_abc_40298_new_n901_), .Y(_abc_40298_new_n908_));
INVX1 INVX1_920 ( .A(REGFILE_SIM_reg_bank_reg_r17_25_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3118_));
INVX1 INVX1_921 ( .A(REGFILE_SIM_reg_bank_reg_r17_26_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3120_));
INVX1 INVX1_922 ( .A(REGFILE_SIM_reg_bank_reg_r17_27_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3122_));
INVX1 INVX1_923 ( .A(REGFILE_SIM_reg_bank_reg_r17_28_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3124_));
INVX1 INVX1_924 ( .A(REGFILE_SIM_reg_bank_reg_r17_29_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3126_));
INVX1 INVX1_925 ( .A(REGFILE_SIM_reg_bank_reg_r17_30_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3128_));
INVX1 INVX1_926 ( .A(REGFILE_SIM_reg_bank_reg_r17_31_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3130_));
INVX1 INVX1_927 ( .A(REGFILE_SIM_reg_bank_reg_r16_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3132_));
INVX1 INVX1_928 ( .A(REGFILE_SIM_reg_bank_reg_r16_1_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3135_));
INVX1 INVX1_929 ( .A(REGFILE_SIM_reg_bank_reg_r16_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3137_));
INVX1 INVX1_93 ( .A(alu_op_r_1_), .Y(_abc_40298_new_n909_));
INVX1 INVX1_930 ( .A(REGFILE_SIM_reg_bank_reg_r16_3_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3139_));
INVX1 INVX1_931 ( .A(REGFILE_SIM_reg_bank_reg_r16_4_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3141_));
INVX1 INVX1_932 ( .A(REGFILE_SIM_reg_bank_reg_r16_5_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3143_));
INVX1 INVX1_933 ( .A(REGFILE_SIM_reg_bank_reg_r16_6_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3145_));
INVX1 INVX1_934 ( .A(REGFILE_SIM_reg_bank_reg_r16_7_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3147_));
INVX1 INVX1_935 ( .A(REGFILE_SIM_reg_bank_reg_r16_8_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3149_));
INVX1 INVX1_936 ( .A(REGFILE_SIM_reg_bank_reg_r16_9_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3151_));
INVX1 INVX1_937 ( .A(REGFILE_SIM_reg_bank_reg_r16_10_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3153_));
INVX1 INVX1_938 ( .A(REGFILE_SIM_reg_bank_reg_r16_11_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3155_));
INVX1 INVX1_939 ( .A(REGFILE_SIM_reg_bank_reg_r16_12_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3157_));
INVX1 INVX1_94 ( .A(alu_op_r_0_), .Y(_abc_40298_new_n911_));
INVX1 INVX1_940 ( .A(REGFILE_SIM_reg_bank_reg_r16_13_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3159_));
INVX1 INVX1_941 ( .A(REGFILE_SIM_reg_bank_reg_r16_14_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3161_));
INVX1 INVX1_942 ( .A(REGFILE_SIM_reg_bank_reg_r16_15_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3163_));
INVX1 INVX1_943 ( .A(REGFILE_SIM_reg_bank_reg_r16_16_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3165_));
INVX1 INVX1_944 ( .A(REGFILE_SIM_reg_bank_reg_r16_17_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3167_));
INVX1 INVX1_945 ( .A(REGFILE_SIM_reg_bank_reg_r16_18_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3169_));
INVX1 INVX1_946 ( .A(REGFILE_SIM_reg_bank_reg_r16_19_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3171_));
INVX1 INVX1_947 ( .A(REGFILE_SIM_reg_bank_reg_r16_20_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3173_));
INVX1 INVX1_948 ( .A(REGFILE_SIM_reg_bank_reg_r16_21_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3175_));
INVX1 INVX1_949 ( .A(REGFILE_SIM_reg_bank_reg_r16_22_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3177_));
INVX1 INVX1_95 ( .A(alu_op_r_4_), .Y(_abc_40298_new_n917_));
INVX1 INVX1_950 ( .A(REGFILE_SIM_reg_bank_reg_r16_23_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3179_));
INVX1 INVX1_951 ( .A(REGFILE_SIM_reg_bank_reg_r16_24_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3181_));
INVX1 INVX1_952 ( .A(REGFILE_SIM_reg_bank_reg_r16_25_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3183_));
INVX1 INVX1_953 ( .A(REGFILE_SIM_reg_bank_reg_r16_26_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3185_));
INVX1 INVX1_954 ( .A(REGFILE_SIM_reg_bank_reg_r16_27_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3187_));
INVX1 INVX1_955 ( .A(REGFILE_SIM_reg_bank_reg_r16_28_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3189_));
INVX1 INVX1_956 ( .A(REGFILE_SIM_reg_bank_reg_r16_29_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3191_));
INVX1 INVX1_957 ( .A(REGFILE_SIM_reg_bank_reg_r16_30_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3193_));
INVX1 INVX1_958 ( .A(REGFILE_SIM_reg_bank_reg_r16_31_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3195_));
INVX1 INVX1_959 ( .A(REGFILE_SIM_reg_bank_reg_r15_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3197_));
INVX1 INVX1_96 ( .A(_abc_40298_new_n918_), .Y(_abc_40298_new_n919_));
INVX1 INVX1_960 ( .A(REGFILE_SIM_reg_bank_wr_i), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3198_));
INVX1 INVX1_961 ( .A(REGFILE_SIM_reg_bank_reg_r15_1_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3202_));
INVX1 INVX1_962 ( .A(REGFILE_SIM_reg_bank_reg_r15_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3204_));
INVX1 INVX1_963 ( .A(REGFILE_SIM_reg_bank_reg_r15_3_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3206_));
INVX1 INVX1_964 ( .A(REGFILE_SIM_reg_bank_reg_r15_4_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3208_));
INVX1 INVX1_965 ( .A(REGFILE_SIM_reg_bank_reg_r15_5_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3210_));
INVX1 INVX1_966 ( .A(REGFILE_SIM_reg_bank_reg_r15_6_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3212_));
INVX1 INVX1_967 ( .A(REGFILE_SIM_reg_bank_reg_r15_7_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3214_));
INVX1 INVX1_968 ( .A(REGFILE_SIM_reg_bank_reg_r15_8_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3216_));
INVX1 INVX1_969 ( .A(REGFILE_SIM_reg_bank_reg_r15_9_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3218_));
INVX1 INVX1_97 ( .A(_abc_40298_new_n899_), .Y(_abc_40298_new_n925_));
INVX1 INVX1_970 ( .A(REGFILE_SIM_reg_bank_reg_r15_10_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3220_));
INVX1 INVX1_971 ( .A(REGFILE_SIM_reg_bank_reg_r15_11_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3222_));
INVX1 INVX1_972 ( .A(REGFILE_SIM_reg_bank_reg_r15_12_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3224_));
INVX1 INVX1_973 ( .A(REGFILE_SIM_reg_bank_reg_r15_13_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3226_));
INVX1 INVX1_974 ( .A(REGFILE_SIM_reg_bank_reg_r15_14_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3228_));
INVX1 INVX1_975 ( .A(REGFILE_SIM_reg_bank_reg_r15_15_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3230_));
INVX1 INVX1_976 ( .A(REGFILE_SIM_reg_bank_reg_r15_16_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3232_));
INVX1 INVX1_977 ( .A(REGFILE_SIM_reg_bank_reg_r15_17_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3234_));
INVX1 INVX1_978 ( .A(REGFILE_SIM_reg_bank_reg_r15_18_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3236_));
INVX1 INVX1_979 ( .A(REGFILE_SIM_reg_bank_reg_r15_19_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3238_));
INVX1 INVX1_98 ( .A(_abc_40298_new_n932_), .Y(_abc_40298_new_n933_));
INVX1 INVX1_980 ( .A(REGFILE_SIM_reg_bank_reg_r15_20_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3240_));
INVX1 INVX1_981 ( .A(REGFILE_SIM_reg_bank_reg_r15_21_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3242_));
INVX1 INVX1_982 ( .A(REGFILE_SIM_reg_bank_reg_r15_22_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3244_));
INVX1 INVX1_983 ( .A(REGFILE_SIM_reg_bank_reg_r15_23_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3246_));
INVX1 INVX1_984 ( .A(REGFILE_SIM_reg_bank_reg_r15_24_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3248_));
INVX1 INVX1_985 ( .A(REGFILE_SIM_reg_bank_reg_r15_25_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3250_));
INVX1 INVX1_986 ( .A(REGFILE_SIM_reg_bank_reg_r15_26_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3252_));
INVX1 INVX1_987 ( .A(REGFILE_SIM_reg_bank_reg_r15_27_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3254_));
INVX1 INVX1_988 ( .A(REGFILE_SIM_reg_bank_reg_r15_28_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3256_));
INVX1 INVX1_989 ( .A(REGFILE_SIM_reg_bank_reg_r15_29_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3258_));
INVX1 INVX1_99 ( .A(opcode_q_23_), .Y(_abc_40298_new_n938_));
INVX1 INVX1_990 ( .A(REGFILE_SIM_reg_bank_reg_r15_30_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3260_));
INVX1 INVX1_991 ( .A(REGFILE_SIM_reg_bank_reg_r15_31_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3262_));
INVX1 INVX1_992 ( .A(REGFILE_SIM_reg_bank_reg_r14_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3264_));
INVX1 INVX1_993 ( .A(REGFILE_SIM_reg_bank_reg_r14_1_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3267_));
INVX1 INVX1_994 ( .A(REGFILE_SIM_reg_bank_reg_r14_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3269_));
INVX1 INVX1_995 ( .A(REGFILE_SIM_reg_bank_reg_r14_3_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3271_));
INVX1 INVX1_996 ( .A(REGFILE_SIM_reg_bank_reg_r14_4_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3273_));
INVX1 INVX1_997 ( .A(REGFILE_SIM_reg_bank_reg_r14_5_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3275_));
INVX1 INVX1_998 ( .A(REGFILE_SIM_reg_bank_reg_r14_6_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3277_));
INVX1 INVX1_999 ( .A(REGFILE_SIM_reg_bank_reg_r14_7_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3279_));
MUX2X1 MUX2X1_1 ( .A(_abc_40298_new_n1139_), .B(_abc_40298_new_n1140_), .S(_abc_40298_new_n1082_), .Y(_abc_40298_new_n1141_));
MUX2X1 MUX2X1_10 ( .A(epc_q_9_), .B(REGFILE_SIM_reg_bank_reg_rb_o_9_), .S(_abc_40298_new_n1187_), .Y(_abc_40298_new_n1393_));
MUX2X1 MUX2X1_100 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2198_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2199_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2106_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__31_));
MUX2X1 MUX2X1_1000 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2115_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4118_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4112_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__3_));
MUX2X1 MUX2X1_1001 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2118_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4120_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4112_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__4_));
MUX2X1 MUX2X1_1002 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2121_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4122_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4112_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__5_));
MUX2X1 MUX2X1_1003 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2124_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4124_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4112_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__6_));
MUX2X1 MUX2X1_1004 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2127_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4126_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4112_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__7_));
MUX2X1 MUX2X1_1005 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2130_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4128_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4112_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__8_));
MUX2X1 MUX2X1_1006 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2133_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4130_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4112_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__9_));
MUX2X1 MUX2X1_1007 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2136_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4132_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4112_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__10_));
MUX2X1 MUX2X1_1008 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2139_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4134_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4112_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__11_));
MUX2X1 MUX2X1_1009 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2142_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4136_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4112_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__12_));
MUX2X1 MUX2X1_101 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2201_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2100_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2205_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__0_));
MUX2X1 MUX2X1_1010 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2145_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4138_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4112_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__13_));
MUX2X1 MUX2X1_1011 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2148_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4140_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4112_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__14_));
MUX2X1 MUX2X1_1012 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2151_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4142_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4112_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__15_));
MUX2X1 MUX2X1_1013 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2154_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4144_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4112_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__16_));
MUX2X1 MUX2X1_1014 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2157_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4146_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4112_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__17_));
MUX2X1 MUX2X1_1015 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2160_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4148_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4112_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__18_));
MUX2X1 MUX2X1_1016 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2163_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4150_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4112_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__19_));
MUX2X1 MUX2X1_1017 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2166_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4152_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4112_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__20_));
MUX2X1 MUX2X1_1018 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2169_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4154_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4112_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__21_));
MUX2X1 MUX2X1_1019 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2172_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4156_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4112_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__22_));
MUX2X1 MUX2X1_102 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2207_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2109_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2205_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__1_));
MUX2X1 MUX2X1_1020 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2175_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4158_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4112_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__23_));
MUX2X1 MUX2X1_1021 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2178_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4160_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4112_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__24_));
MUX2X1 MUX2X1_1022 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2181_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4162_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4112_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__25_));
MUX2X1 MUX2X1_1023 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2184_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4164_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4112_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__26_));
MUX2X1 MUX2X1_1024 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2187_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4166_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4112_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__27_));
MUX2X1 MUX2X1_1025 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2190_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4168_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4112_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__28_));
MUX2X1 MUX2X1_1026 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2193_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4170_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4112_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__29_));
MUX2X1 MUX2X1_1027 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2196_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4172_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4112_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__30_));
MUX2X1 MUX2X1_1028 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2199_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4174_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4112_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__31_));
MUX2X1 MUX2X1_1029 ( .A(alu__abc_38674_new_n632_), .B(alu__abc_38674_new_n630_), .S(alu__abc_38674_new_n559_), .Y(alu__abc_38674_new_n633_));
MUX2X1 MUX2X1_103 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2209_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2112_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2205_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__2_));
MUX2X1 MUX2X1_1030 ( .A(alu__abc_38674_new_n364_), .B(alu__abc_38674_new_n202_), .S(alu_b_i_0_), .Y(alu__abc_38674_new_n634_));
MUX2X1 MUX2X1_1031 ( .A(alu__abc_38674_new_n329_), .B(alu__abc_38674_new_n330_), .S(alu_b_i_0_), .Y(alu__abc_38674_new_n648_));
MUX2X1 MUX2X1_1032 ( .A(alu__abc_38674_new_n165_), .B(alu__abc_38674_new_n171_), .S(alu_b_i_0_), .Y(alu__abc_38674_new_n662_));
MUX2X1 MUX2X1_1033 ( .A(alu__abc_38674_new_n117_), .B(alu__abc_38674_new_n111_), .S(alu_b_i_0_), .Y(alu__abc_38674_new_n675_));
MUX2X1 MUX2X1_1034 ( .A(alu__abc_38674_new_n308_), .B(alu__abc_38674_new_n135_), .S(alu_b_i_0_), .Y(alu__abc_38674_new_n681_));
MUX2X1 MUX2X1_1035 ( .A(alu__abc_38674_new_n345_), .B(alu__abc_38674_new_n641_), .S(alu_b_i_0_), .Y(alu__abc_38674_new_n717_));
MUX2X1 MUX2X1_1036 ( .A(alu__abc_38674_new_n351_), .B(alu__abc_38674_new_n329_), .S(alu_b_i_0_), .Y(alu__abc_38674_new_n722_));
MUX2X1 MUX2X1_1037 ( .A(alu__abc_38674_new_n330_), .B(alu__abc_38674_new_n334_), .S(alu_b_i_0_), .Y(alu__abc_38674_new_n723_));
MUX2X1 MUX2X1_1038 ( .A(alu__abc_38674_new_n723_), .B(alu__abc_38674_new_n722_), .S(alu__abc_38674_new_n559_), .Y(alu__abc_38674_new_n724_));
MUX2X1 MUX2X1_1039 ( .A(alu__abc_38674_new_n721_), .B(alu__abc_38674_new_n724_), .S(alu__abc_38674_new_n338_), .Y(alu__abc_38674_new_n725_));
MUX2X1 MUX2X1_104 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2211_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2115_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2205_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__3_));
MUX2X1 MUX2X1_1040 ( .A(alu__abc_38674_new_n233_), .B(alu__abc_38674_new_n228_), .S(alu_b_i_0_), .Y(alu__abc_38674_new_n734_));
MUX2X1 MUX2X1_1041 ( .A(alu__abc_38674_new_n733_), .B(alu__abc_38674_new_n738_), .S(alu_b_i_2_), .Y(alu__abc_38674_new_n739_));
MUX2X1 MUX2X1_1042 ( .A(alu__abc_38674_new_n144_), .B(alu__abc_38674_new_n308_), .S(alu_b_i_0_), .Y(alu__abc_38674_new_n749_));
MUX2X1 MUX2X1_1043 ( .A(alu__abc_38674_new_n681_), .B(alu__abc_38674_new_n634_), .S(alu_b_i_1_), .Y(alu__abc_38674_new_n824_));
MUX2X1 MUX2X1_1044 ( .A(alu__abc_38674_new_n827_), .B(alu__abc_38674_new_n824_), .S(alu__abc_38674_new_n338_), .Y(alu__abc_38674_new_n828_));
MUX2X1 MUX2X1_1045 ( .A(alu__abc_38674_new_n723_), .B(alu__abc_38674_new_n717_), .S(alu_b_i_1_), .Y(alu__abc_38674_new_n866_));
MUX2X1 MUX2X1_1046 ( .A(alu__abc_38674_new_n734_), .B(alu__abc_38674_new_n722_), .S(alu_b_i_1_), .Y(alu__abc_38674_new_n867_));
MUX2X1 MUX2X1_1047 ( .A(alu__abc_38674_new_n867_), .B(alu__abc_38674_new_n866_), .S(alu_b_i_2_), .Y(alu__abc_38674_new_n868_));
MUX2X1 MUX2X1_1048 ( .A(alu__abc_38674_new_n738_), .B(alu__abc_38674_new_n724_), .S(alu_b_i_2_), .Y(alu__abc_38674_new_n947_));
MUX2X1 MUX2X1_1049 ( .A(alu__abc_38674_new_n810_), .B(alu__abc_38674_new_n803_), .S(alu__abc_38674_new_n338_), .Y(alu__abc_38674_new_n988_));
MUX2X1 MUX2X1_105 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2213_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2118_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2205_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__4_));
MUX2X1 MUX2X1_1050 ( .A(alu__abc_38674_new_n991_), .B(alu__abc_38674_new_n987_), .S(alu_b_i_4_), .Y(alu__abc_38674_new_n992_));
MUX2X1 MUX2X1_1051 ( .A(alu__abc_38674_new_n874_), .B(alu__abc_38674_new_n867_), .S(alu_b_i_2_), .Y(alu__abc_38674_new_n1013_));
MUX2X1 MUX2X1_1052 ( .A(alu__abc_38674_new_n202_), .B(alu__abc_38674_new_n364_), .S(alu_b_i_0_), .Y(alu__abc_38674_new_n1280_));
MUX2X1 MUX2X1_1053 ( .A(alu__abc_38674_new_n1315_), .B(alu__abc_38674_new_n1066_), .S(alu__abc_38674_new_n340_), .Y(alu__abc_38674_new_n1316_));
MUX2X1 MUX2X1_1054 ( .A(alu__abc_38674_new_n135_), .B(alu__abc_38674_new_n308_), .S(alu_b_i_0_), .Y(alu__abc_38674_new_n1343_));
MUX2X1 MUX2X1_1055 ( .A(alu__abc_38674_new_n1343_), .B(alu__abc_38674_new_n1280_), .S(alu__abc_38674_new_n559_), .Y(alu__abc_38674_new_n1344_));
MUX2X1 MUX2X1_1056 ( .A(alu__abc_38674_new_n1456_), .B(alu__abc_38674_new_n1344_), .S(alu__abc_38674_new_n338_), .Y(alu__abc_38674_new_n1457_));
MUX2X1 MUX2X1_1057 ( .A(alu__abc_38674_new_n1534_), .B(alu__abc_38674_new_n1475_), .S(alu__abc_38674_new_n559_), .Y(alu__abc_38674_new_n1535_));
MUX2X1 MUX2X1_1058 ( .A(alu__abc_38674_new_n1612_), .B(alu__abc_38674_new_n1394_), .S(alu__abc_38674_new_n340_), .Y(alu__abc_38674_new_n1613_));
MUX2X1 MUX2X1_1059 ( .A(alu__abc_38674_new_n1554_), .B(alu__abc_38674_new_n1658_), .S(alu_b_i_2_), .Y(alu__abc_38674_new_n1659_));
MUX2X1 MUX2X1_106 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2215_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2121_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2205_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__5_));
MUX2X1 MUX2X1_1060 ( .A(alu__abc_38674_new_n1659_), .B(alu__abc_38674_new_n1457_), .S(alu__abc_38674_new_n340_), .Y(alu__abc_38674_new_n1660_));
MUX2X1 MUX2X1_1061 ( .A(alu__abc_38674_new_n1588_), .B(alu__abc_38674_new_n1682_), .S(alu_b_i_2_), .Y(alu__abc_38674_new_n1683_));
MUX2X1 MUX2X1_1062 ( .A(alu__abc_38674_new_n1706_), .B(alu__abc_38674_new_n1656_), .S(alu__abc_38674_new_n559_), .Y(alu__abc_38674_new_n1707_));
MUX2X1 MUX2X1_107 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2217_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2124_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2205_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__6_));
MUX2X1 MUX2X1_108 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2219_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2127_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2205_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__7_));
MUX2X1 MUX2X1_109 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2221_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2130_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2205_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__8_));
MUX2X1 MUX2X1_11 ( .A(epc_q_10_), .B(REGFILE_SIM_reg_bank_reg_rb_o_10_), .S(_abc_40298_new_n1187_), .Y(_abc_40298_new_n1421_));
MUX2X1 MUX2X1_110 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2223_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2133_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2205_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__9_));
MUX2X1 MUX2X1_111 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2225_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2136_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2205_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__10_));
MUX2X1 MUX2X1_112 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2227_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2139_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2205_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__11_));
MUX2X1 MUX2X1_113 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2229_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2142_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2205_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__12_));
MUX2X1 MUX2X1_114 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2231_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2145_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2205_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__13_));
MUX2X1 MUX2X1_115 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2233_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2148_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2205_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__14_));
MUX2X1 MUX2X1_116 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2235_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2151_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2205_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__15_));
MUX2X1 MUX2X1_117 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2237_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2154_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2205_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__16_));
MUX2X1 MUX2X1_118 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2239_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2157_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2205_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__17_));
MUX2X1 MUX2X1_119 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2241_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2160_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2205_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__18_));
MUX2X1 MUX2X1_12 ( .A(epc_q_11_), .B(REGFILE_SIM_reg_bank_reg_rb_o_11_), .S(_abc_40298_new_n1187_), .Y(_abc_40298_new_n1452_));
MUX2X1 MUX2X1_120 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2243_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2163_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2205_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__19_));
MUX2X1 MUX2X1_121 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2245_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2166_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2205_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__20_));
MUX2X1 MUX2X1_122 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2247_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2169_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2205_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__21_));
MUX2X1 MUX2X1_123 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2249_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2172_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2205_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__22_));
MUX2X1 MUX2X1_124 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2251_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2175_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2205_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__23_));
MUX2X1 MUX2X1_125 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2253_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2178_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2205_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__24_));
MUX2X1 MUX2X1_126 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2255_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2181_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2205_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__25_));
MUX2X1 MUX2X1_127 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2257_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2184_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2205_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__26_));
MUX2X1 MUX2X1_128 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2259_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2187_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2205_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__27_));
MUX2X1 MUX2X1_129 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2261_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2190_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2205_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__28_));
MUX2X1 MUX2X1_13 ( .A(epc_q_12_), .B(REGFILE_SIM_reg_bank_reg_rb_o_12_), .S(_abc_40298_new_n1187_), .Y(_abc_40298_new_n1504_));
MUX2X1 MUX2X1_130 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2263_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2193_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2205_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__29_));
MUX2X1 MUX2X1_131 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2265_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2196_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2205_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__30_));
MUX2X1 MUX2X1_132 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2267_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2199_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2205_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__31_));
MUX2X1 MUX2X1_133 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2269_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2100_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2272_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__0_));
MUX2X1 MUX2X1_134 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2274_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2109_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2272_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__1_));
MUX2X1 MUX2X1_135 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2276_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2112_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2272_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__2_));
MUX2X1 MUX2X1_136 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2278_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2115_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2272_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__3_));
MUX2X1 MUX2X1_137 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2280_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2118_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2272_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__4_));
MUX2X1 MUX2X1_138 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2282_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2121_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2272_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__5_));
MUX2X1 MUX2X1_139 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2284_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2124_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2272_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__6_));
MUX2X1 MUX2X1_14 ( .A(epc_q_13_), .B(REGFILE_SIM_reg_bank_reg_rb_o_13_), .S(_abc_40298_new_n1187_), .Y(_abc_40298_new_n1527_));
MUX2X1 MUX2X1_140 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2286_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2127_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2272_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__7_));
MUX2X1 MUX2X1_141 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2288_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2130_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2272_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__8_));
MUX2X1 MUX2X1_142 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2290_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2133_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2272_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__9_));
MUX2X1 MUX2X1_143 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2292_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2136_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2272_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__10_));
MUX2X1 MUX2X1_144 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2294_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2139_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2272_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__11_));
MUX2X1 MUX2X1_145 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2296_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2142_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2272_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__12_));
MUX2X1 MUX2X1_146 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2298_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2145_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2272_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__13_));
MUX2X1 MUX2X1_147 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2300_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2148_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2272_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__14_));
MUX2X1 MUX2X1_148 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2302_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2151_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2272_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__15_));
MUX2X1 MUX2X1_149 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2304_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2154_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2272_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__16_));
MUX2X1 MUX2X1_15 ( .A(epc_q_14_), .B(REGFILE_SIM_reg_bank_reg_rb_o_14_), .S(_abc_40298_new_n1187_), .Y(_abc_40298_new_n1556_));
MUX2X1 MUX2X1_150 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2306_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2157_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2272_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__17_));
MUX2X1 MUX2X1_151 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2308_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2160_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2272_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__18_));
MUX2X1 MUX2X1_152 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2310_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2163_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2272_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__19_));
MUX2X1 MUX2X1_153 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2312_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2166_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2272_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__20_));
MUX2X1 MUX2X1_154 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2314_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2169_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2272_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__21_));
MUX2X1 MUX2X1_155 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2316_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2172_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2272_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__22_));
MUX2X1 MUX2X1_156 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2318_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2175_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2272_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__23_));
MUX2X1 MUX2X1_157 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2320_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2178_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2272_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__24_));
MUX2X1 MUX2X1_158 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2322_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2181_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2272_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__25_));
MUX2X1 MUX2X1_159 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2324_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2184_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2272_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__26_));
MUX2X1 MUX2X1_16 ( .A(epc_q_15_), .B(REGFILE_SIM_reg_bank_reg_rb_o_15_), .S(_abc_40298_new_n1187_), .Y(_abc_40298_new_n1582_));
MUX2X1 MUX2X1_160 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2326_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2187_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2272_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__27_));
MUX2X1 MUX2X1_161 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2328_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2190_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2272_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__28_));
MUX2X1 MUX2X1_162 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2330_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2193_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2272_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__29_));
MUX2X1 MUX2X1_163 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2332_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2196_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2272_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__30_));
MUX2X1 MUX2X1_164 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2334_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2199_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2272_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__31_));
MUX2X1 MUX2X1_165 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2336_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2100_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2339_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__0_));
MUX2X1 MUX2X1_166 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2341_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2109_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2339_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__1_));
MUX2X1 MUX2X1_167 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2343_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2112_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2339_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__2_));
MUX2X1 MUX2X1_168 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2345_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2115_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2339_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__3_));
MUX2X1 MUX2X1_169 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2347_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2118_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2339_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__4_));
MUX2X1 MUX2X1_17 ( .A(epc_q_16_), .B(REGFILE_SIM_reg_bank_reg_rb_o_16_), .S(_abc_40298_new_n1187_), .Y(_abc_40298_new_n1615_));
MUX2X1 MUX2X1_170 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2349_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2121_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2339_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__5_));
MUX2X1 MUX2X1_171 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2351_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2124_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2339_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__6_));
MUX2X1 MUX2X1_172 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2353_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2127_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2339_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__7_));
MUX2X1 MUX2X1_173 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2355_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2130_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2339_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__8_));
MUX2X1 MUX2X1_174 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2357_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2133_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2339_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__9_));
MUX2X1 MUX2X1_175 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2359_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2136_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2339_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__10_));
MUX2X1 MUX2X1_176 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2361_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2139_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2339_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__11_));
MUX2X1 MUX2X1_177 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2363_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2142_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2339_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__12_));
MUX2X1 MUX2X1_178 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2365_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2145_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2339_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__13_));
MUX2X1 MUX2X1_179 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2367_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2148_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2339_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__14_));
MUX2X1 MUX2X1_18 ( .A(epc_q_17_), .B(REGFILE_SIM_reg_bank_reg_rb_o_17_), .S(_abc_40298_new_n1187_), .Y(_abc_40298_new_n1639_));
MUX2X1 MUX2X1_180 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2369_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2151_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2339_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__15_));
MUX2X1 MUX2X1_181 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2371_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2154_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2339_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__16_));
MUX2X1 MUX2X1_182 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2373_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2157_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2339_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__17_));
MUX2X1 MUX2X1_183 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2375_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2160_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2339_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__18_));
MUX2X1 MUX2X1_184 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2377_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2163_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2339_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__19_));
MUX2X1 MUX2X1_185 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2379_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2166_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2339_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__20_));
MUX2X1 MUX2X1_186 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2381_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2169_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2339_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__21_));
MUX2X1 MUX2X1_187 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2383_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2172_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2339_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__22_));
MUX2X1 MUX2X1_188 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2385_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2175_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2339_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__23_));
MUX2X1 MUX2X1_189 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2387_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2178_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2339_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__24_));
MUX2X1 MUX2X1_19 ( .A(epc_q_18_), .B(REGFILE_SIM_reg_bank_reg_rb_o_18_), .S(_abc_40298_new_n1187_), .Y(_abc_40298_new_n1669_));
MUX2X1 MUX2X1_190 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2389_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2181_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2339_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__25_));
MUX2X1 MUX2X1_191 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2391_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2184_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2339_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__26_));
MUX2X1 MUX2X1_192 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2393_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2187_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2339_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__27_));
MUX2X1 MUX2X1_193 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2395_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2190_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2339_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__28_));
MUX2X1 MUX2X1_194 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2397_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2193_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2339_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__29_));
MUX2X1 MUX2X1_195 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2399_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2196_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2339_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__30_));
MUX2X1 MUX2X1_196 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2401_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2199_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2339_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__31_));
MUX2X1 MUX2X1_197 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2403_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2100_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2407_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__0_));
MUX2X1 MUX2X1_198 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2409_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2109_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2407_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__1_));
MUX2X1 MUX2X1_199 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2411_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2112_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2407_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__2_));
MUX2X1 MUX2X1_2 ( .A(alu_c_o), .B(alu_c_i), .S(alu_c_update_o), .Y(_abc_40298_new_n1145_));
MUX2X1 MUX2X1_20 ( .A(epc_q_19_), .B(REGFILE_SIM_reg_bank_reg_rb_o_19_), .S(_abc_40298_new_n1187_), .Y(_abc_40298_new_n1692_));
MUX2X1 MUX2X1_200 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2413_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2115_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2407_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__3_));
MUX2X1 MUX2X1_201 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2415_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2118_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2407_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__4_));
MUX2X1 MUX2X1_202 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2417_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2121_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2407_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__5_));
MUX2X1 MUX2X1_203 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2419_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2124_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2407_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__6_));
MUX2X1 MUX2X1_204 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2421_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2127_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2407_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__7_));
MUX2X1 MUX2X1_205 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2423_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2130_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2407_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__8_));
MUX2X1 MUX2X1_206 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2425_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2133_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2407_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__9_));
MUX2X1 MUX2X1_207 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2427_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2136_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2407_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__10_));
MUX2X1 MUX2X1_208 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2429_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2139_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2407_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__11_));
MUX2X1 MUX2X1_209 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2431_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2142_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2407_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__12_));
MUX2X1 MUX2X1_21 ( .A(epc_q_20_), .B(REGFILE_SIM_reg_bank_reg_rb_o_20_), .S(_abc_40298_new_n1187_), .Y(_abc_40298_new_n1721_));
MUX2X1 MUX2X1_210 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2433_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2145_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2407_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__13_));
MUX2X1 MUX2X1_211 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2435_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2148_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2407_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__14_));
MUX2X1 MUX2X1_212 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2437_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2151_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2407_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__15_));
MUX2X1 MUX2X1_213 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2439_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2154_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2407_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__16_));
MUX2X1 MUX2X1_214 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2441_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2157_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2407_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__17_));
MUX2X1 MUX2X1_215 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2443_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2160_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2407_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__18_));
MUX2X1 MUX2X1_216 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2445_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2163_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2407_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__19_));
MUX2X1 MUX2X1_217 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2447_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2166_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2407_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__20_));
MUX2X1 MUX2X1_218 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2449_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2169_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2407_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__21_));
MUX2X1 MUX2X1_219 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2451_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2172_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2407_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__22_));
MUX2X1 MUX2X1_22 ( .A(epc_q_21_), .B(REGFILE_SIM_reg_bank_reg_rb_o_21_), .S(_abc_40298_new_n1187_), .Y(_abc_40298_new_n1748_));
MUX2X1 MUX2X1_220 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2453_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2175_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2407_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__23_));
MUX2X1 MUX2X1_221 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2455_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2178_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2407_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__24_));
MUX2X1 MUX2X1_222 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2457_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2181_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2407_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__25_));
MUX2X1 MUX2X1_223 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2459_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2184_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2407_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__26_));
MUX2X1 MUX2X1_224 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2461_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2187_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2407_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__27_));
MUX2X1 MUX2X1_225 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2463_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2190_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2407_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__28_));
MUX2X1 MUX2X1_226 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2465_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2193_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2407_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__29_));
MUX2X1 MUX2X1_227 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2467_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2196_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2407_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__30_));
MUX2X1 MUX2X1_228 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2469_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2199_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2407_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__31_));
MUX2X1 MUX2X1_229 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2471_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2100_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2473_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__0_));
MUX2X1 MUX2X1_23 ( .A(epc_q_22_), .B(REGFILE_SIM_reg_bank_reg_rb_o_22_), .S(_abc_40298_new_n1187_), .Y(_abc_40298_new_n1777_));
MUX2X1 MUX2X1_230 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2475_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2109_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2473_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__1_));
MUX2X1 MUX2X1_231 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2477_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2112_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2473_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__2_));
MUX2X1 MUX2X1_232 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2479_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2115_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2473_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__3_));
MUX2X1 MUX2X1_233 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2481_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2118_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2473_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__4_));
MUX2X1 MUX2X1_234 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2483_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2121_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2473_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__5_));
MUX2X1 MUX2X1_235 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2485_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2124_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2473_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__6_));
MUX2X1 MUX2X1_236 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2487_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2127_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2473_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__7_));
MUX2X1 MUX2X1_237 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2489_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2130_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2473_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__8_));
MUX2X1 MUX2X1_238 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2491_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2133_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2473_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__9_));
MUX2X1 MUX2X1_239 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2493_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2136_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2473_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__10_));
MUX2X1 MUX2X1_24 ( .A(epc_q_23_), .B(REGFILE_SIM_reg_bank_reg_rb_o_23_), .S(_abc_40298_new_n1187_), .Y(_abc_40298_new_n1800_));
MUX2X1 MUX2X1_240 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2495_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2139_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2473_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__11_));
MUX2X1 MUX2X1_241 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2497_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2142_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2473_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__12_));
MUX2X1 MUX2X1_242 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2499_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2145_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2473_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__13_));
MUX2X1 MUX2X1_243 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2501_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2148_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2473_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__14_));
MUX2X1 MUX2X1_244 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2503_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2151_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2473_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__15_));
MUX2X1 MUX2X1_245 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2505_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2154_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2473_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__16_));
MUX2X1 MUX2X1_246 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2507_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2157_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2473_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__17_));
MUX2X1 MUX2X1_247 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2509_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2160_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2473_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__18_));
MUX2X1 MUX2X1_248 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2511_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2163_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2473_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__19_));
MUX2X1 MUX2X1_249 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2513_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2166_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2473_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__20_));
MUX2X1 MUX2X1_25 ( .A(epc_q_24_), .B(REGFILE_SIM_reg_bank_reg_rb_o_24_), .S(_abc_40298_new_n1187_), .Y(_abc_40298_new_n1836_));
MUX2X1 MUX2X1_250 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2515_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2169_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2473_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__21_));
MUX2X1 MUX2X1_251 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2517_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2172_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2473_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__22_));
MUX2X1 MUX2X1_252 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2519_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2175_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2473_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__23_));
MUX2X1 MUX2X1_253 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2521_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2178_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2473_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__24_));
MUX2X1 MUX2X1_254 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2523_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2181_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2473_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__25_));
MUX2X1 MUX2X1_255 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2525_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2184_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2473_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__26_));
MUX2X1 MUX2X1_256 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2527_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2187_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2473_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__27_));
MUX2X1 MUX2X1_257 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2529_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2190_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2473_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__28_));
MUX2X1 MUX2X1_258 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2531_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2193_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2473_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__29_));
MUX2X1 MUX2X1_259 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2533_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2196_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2473_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__30_));
MUX2X1 MUX2X1_26 ( .A(epc_q_25_), .B(REGFILE_SIM_reg_bank_reg_rb_o_25_), .S(_abc_40298_new_n1187_), .Y(_abc_40298_new_n1857_));
MUX2X1 MUX2X1_260 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2535_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2199_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2473_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__31_));
MUX2X1 MUX2X1_261 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2537_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2100_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2539_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__0_));
MUX2X1 MUX2X1_262 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2541_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2109_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2539_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__1_));
MUX2X1 MUX2X1_263 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2543_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2112_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2539_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__2_));
MUX2X1 MUX2X1_264 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2545_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2115_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2539_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__3_));
MUX2X1 MUX2X1_265 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2547_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2118_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2539_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__4_));
MUX2X1 MUX2X1_266 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2549_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2121_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2539_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__5_));
MUX2X1 MUX2X1_267 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2551_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2124_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2539_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__6_));
MUX2X1 MUX2X1_268 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2553_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2127_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2539_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__7_));
MUX2X1 MUX2X1_269 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2555_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2130_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2539_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__8_));
MUX2X1 MUX2X1_27 ( .A(_abc_40298_new_n1883_), .B(_abc_40298_new_n1866_), .S(_abc_40298_new_n1213_), .Y(_abc_40298_new_n1884_));
MUX2X1 MUX2X1_270 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2557_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2133_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2539_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__9_));
MUX2X1 MUX2X1_271 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2559_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2136_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2539_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__10_));
MUX2X1 MUX2X1_272 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2561_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2139_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2539_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__11_));
MUX2X1 MUX2X1_273 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2563_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2142_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2539_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__12_));
MUX2X1 MUX2X1_274 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2565_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2145_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2539_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__13_));
MUX2X1 MUX2X1_275 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2567_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2148_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2539_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__14_));
MUX2X1 MUX2X1_276 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2569_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2151_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2539_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__15_));
MUX2X1 MUX2X1_277 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2571_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2154_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2539_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__16_));
MUX2X1 MUX2X1_278 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2573_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2157_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2539_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__17_));
MUX2X1 MUX2X1_279 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2575_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2160_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2539_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__18_));
MUX2X1 MUX2X1_28 ( .A(epc_q_26_), .B(REGFILE_SIM_reg_bank_reg_rb_o_26_), .S(_abc_40298_new_n1187_), .Y(_abc_40298_new_n1886_));
MUX2X1 MUX2X1_280 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2577_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2163_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2539_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__19_));
MUX2X1 MUX2X1_281 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2579_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2166_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2539_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__20_));
MUX2X1 MUX2X1_282 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2581_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2169_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2539_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__21_));
MUX2X1 MUX2X1_283 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2583_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2172_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2539_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__22_));
MUX2X1 MUX2X1_284 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2585_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2175_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2539_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__23_));
MUX2X1 MUX2X1_285 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2587_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2178_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2539_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__24_));
MUX2X1 MUX2X1_286 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2589_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2181_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2539_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__25_));
MUX2X1 MUX2X1_287 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2591_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2184_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2539_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__26_));
MUX2X1 MUX2X1_288 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2593_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2187_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2539_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__27_));
MUX2X1 MUX2X1_289 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2595_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2190_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2539_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__28_));
MUX2X1 MUX2X1_29 ( .A(_abc_40298_new_n1902_), .B(REGFILE_SIM_reg_bank_reg_rb_o_27_), .S(_abc_40298_new_n1175_), .Y(_abc_40298_new_n1903_));
MUX2X1 MUX2X1_290 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2597_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2193_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2539_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__29_));
MUX2X1 MUX2X1_291 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2599_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2196_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2539_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__30_));
MUX2X1 MUX2X1_292 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2601_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2199_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2539_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__31_));
MUX2X1 MUX2X1_293 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2668_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2100_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2671_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__0_));
MUX2X1 MUX2X1_294 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2673_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2109_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2671_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__1_));
MUX2X1 MUX2X1_295 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2675_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2112_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2671_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__2_));
MUX2X1 MUX2X1_296 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2677_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2115_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2671_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__3_));
MUX2X1 MUX2X1_297 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2679_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2118_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2671_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__4_));
MUX2X1 MUX2X1_298 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2681_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2121_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2671_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__5_));
MUX2X1 MUX2X1_299 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2683_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2124_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2671_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__6_));
MUX2X1 MUX2X1_3 ( .A(_abc_40298_new_n1153_), .B(_abc_40298_new_n1154_), .S(_abc_40298_new_n1082_), .Y(_abc_40298_new_n1155_));
MUX2X1 MUX2X1_30 ( .A(epc_q_27_), .B(REGFILE_SIM_reg_bank_reg_rb_o_27_), .S(_abc_40298_new_n1187_), .Y(_abc_40298_new_n1906_));
MUX2X1 MUX2X1_300 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2685_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2127_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2671_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__7_));
MUX2X1 MUX2X1_301 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2687_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2130_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2671_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__8_));
MUX2X1 MUX2X1_302 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2689_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2133_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2671_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__9_));
MUX2X1 MUX2X1_303 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2691_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2136_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2671_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__10_));
MUX2X1 MUX2X1_304 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2693_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2139_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2671_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__11_));
MUX2X1 MUX2X1_305 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2695_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2142_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2671_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__12_));
MUX2X1 MUX2X1_306 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2697_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2145_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2671_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__13_));
MUX2X1 MUX2X1_307 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2699_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2148_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2671_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__14_));
MUX2X1 MUX2X1_308 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2701_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2151_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2671_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__15_));
MUX2X1 MUX2X1_309 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2703_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2154_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2671_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__16_));
MUX2X1 MUX2X1_31 ( .A(_abc_40298_new_n1932_), .B(REGFILE_SIM_reg_bank_reg_rb_o_28_), .S(_abc_40298_new_n1175_), .Y(_abc_40298_new_n1933_));
MUX2X1 MUX2X1_310 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2705_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2157_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2671_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__17_));
MUX2X1 MUX2X1_311 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2707_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2160_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2671_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__18_));
MUX2X1 MUX2X1_312 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2709_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2163_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2671_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__19_));
MUX2X1 MUX2X1_313 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2711_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2166_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2671_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__20_));
MUX2X1 MUX2X1_314 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2713_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2169_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2671_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__21_));
MUX2X1 MUX2X1_315 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2715_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2172_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2671_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__22_));
MUX2X1 MUX2X1_316 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2717_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2175_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2671_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__23_));
MUX2X1 MUX2X1_317 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2719_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2178_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2671_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__24_));
MUX2X1 MUX2X1_318 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2721_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2181_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2671_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__25_));
MUX2X1 MUX2X1_319 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2723_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2184_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2671_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__26_));
MUX2X1 MUX2X1_32 ( .A(epc_q_28_), .B(REGFILE_SIM_reg_bank_reg_rb_o_28_), .S(_abc_40298_new_n1187_), .Y(_abc_40298_new_n1936_));
MUX2X1 MUX2X1_320 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2725_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2187_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2671_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__27_));
MUX2X1 MUX2X1_321 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2727_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2190_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2671_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__28_));
MUX2X1 MUX2X1_322 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2729_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2193_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2671_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__29_));
MUX2X1 MUX2X1_323 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2731_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2196_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2671_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__30_));
MUX2X1 MUX2X1_324 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2733_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2199_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2671_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__31_));
MUX2X1 MUX2X1_325 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2735_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2100_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2737_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__0_));
MUX2X1 MUX2X1_326 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2739_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2109_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2737_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__1_));
MUX2X1 MUX2X1_327 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2741_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2112_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2737_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__2_));
MUX2X1 MUX2X1_328 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2743_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2115_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2737_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__3_));
MUX2X1 MUX2X1_329 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2745_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2118_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2737_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__4_));
MUX2X1 MUX2X1_33 ( .A(epc_q_29_), .B(REGFILE_SIM_reg_bank_reg_rb_o_29_), .S(_abc_40298_new_n1187_), .Y(_abc_40298_new_n1955_));
MUX2X1 MUX2X1_330 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2747_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2121_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2737_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__5_));
MUX2X1 MUX2X1_331 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2749_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2124_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2737_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__6_));
MUX2X1 MUX2X1_332 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2751_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2127_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2737_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__7_));
MUX2X1 MUX2X1_333 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2753_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2130_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2737_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__8_));
MUX2X1 MUX2X1_334 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2755_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2133_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2737_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__9_));
MUX2X1 MUX2X1_335 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2757_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2136_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2737_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__10_));
MUX2X1 MUX2X1_336 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2759_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2139_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2737_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__11_));
MUX2X1 MUX2X1_337 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2761_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2142_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2737_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__12_));
MUX2X1 MUX2X1_338 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2763_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2145_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2737_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__13_));
MUX2X1 MUX2X1_339 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2765_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2148_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2737_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__14_));
MUX2X1 MUX2X1_34 ( .A(epc_q_30_), .B(REGFILE_SIM_reg_bank_reg_rb_o_30_), .S(_abc_40298_new_n1187_), .Y(_abc_40298_new_n1984_));
MUX2X1 MUX2X1_340 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2767_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2151_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2737_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__15_));
MUX2X1 MUX2X1_341 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2769_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2154_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2737_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__16_));
MUX2X1 MUX2X1_342 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2771_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2157_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2737_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__17_));
MUX2X1 MUX2X1_343 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2773_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2160_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2737_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__18_));
MUX2X1 MUX2X1_344 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2775_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2163_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2737_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__19_));
MUX2X1 MUX2X1_345 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2777_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2166_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2737_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__20_));
MUX2X1 MUX2X1_346 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2779_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2169_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2737_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__21_));
MUX2X1 MUX2X1_347 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2781_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2172_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2737_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__22_));
MUX2X1 MUX2X1_348 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2783_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2175_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2737_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__23_));
MUX2X1 MUX2X1_349 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2785_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2178_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2737_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__24_));
MUX2X1 MUX2X1_35 ( .A(_abc_40298_new_n1990_), .B(_abc_40298_new_n1989_), .S(_abc_40298_new_n1971_), .Y(_abc_40298_new_n1991_));
MUX2X1 MUX2X1_350 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2787_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2181_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2737_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__25_));
MUX2X1 MUX2X1_351 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2789_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2184_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2737_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__26_));
MUX2X1 MUX2X1_352 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2791_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2187_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2737_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__27_));
MUX2X1 MUX2X1_353 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2793_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2190_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2737_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__28_));
MUX2X1 MUX2X1_354 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2795_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2193_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2737_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__29_));
MUX2X1 MUX2X1_355 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2797_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2196_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2737_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__30_));
MUX2X1 MUX2X1_356 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2799_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2199_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2737_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__31_));
MUX2X1 MUX2X1_357 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2801_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2100_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2803_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__0_));
MUX2X1 MUX2X1_358 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2805_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2109_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2803_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__1_));
MUX2X1 MUX2X1_359 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2807_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2112_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2803_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__2_));
MUX2X1 MUX2X1_36 ( .A(epc_q_31_), .B(REGFILE_SIM_reg_bank_reg_rb_o_31_), .S(_abc_40298_new_n1187_), .Y(_abc_40298_new_n2007_));
MUX2X1 MUX2X1_360 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2809_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2115_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2803_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__3_));
MUX2X1 MUX2X1_361 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2811_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2118_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2803_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__4_));
MUX2X1 MUX2X1_362 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2813_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2121_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2803_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__5_));
MUX2X1 MUX2X1_363 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2815_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2124_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2803_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__6_));
MUX2X1 MUX2X1_364 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2817_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2127_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2803_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__7_));
MUX2X1 MUX2X1_365 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2819_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2130_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2803_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__8_));
MUX2X1 MUX2X1_366 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2821_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2133_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2803_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__9_));
MUX2X1 MUX2X1_367 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2823_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2136_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2803_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__10_));
MUX2X1 MUX2X1_368 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2825_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2139_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2803_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__11_));
MUX2X1 MUX2X1_369 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2827_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2142_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2803_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__12_));
MUX2X1 MUX2X1_37 ( .A(_abc_40298_new_n676_), .B(_abc_40298_new_n2516_), .S(_abc_40298_new_n669_), .Y(_0mem_offset_q_1_0__0_));
MUX2X1 MUX2X1_370 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2829_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2145_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2803_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__13_));
MUX2X1 MUX2X1_371 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2831_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2148_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2803_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__14_));
MUX2X1 MUX2X1_372 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2833_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2151_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2803_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__15_));
MUX2X1 MUX2X1_373 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2835_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2154_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2803_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__16_));
MUX2X1 MUX2X1_374 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2837_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2157_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2803_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__17_));
MUX2X1 MUX2X1_375 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2839_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2160_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2803_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__18_));
MUX2X1 MUX2X1_376 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2841_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2163_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2803_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__19_));
MUX2X1 MUX2X1_377 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2843_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2166_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2803_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__20_));
MUX2X1 MUX2X1_378 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2845_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2169_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2803_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__21_));
MUX2X1 MUX2X1_379 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2847_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2172_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2803_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__22_));
MUX2X1 MUX2X1_38 ( .A(_abc_40298_new_n672_), .B(_abc_40298_new_n2522_), .S(_abc_40298_new_n669_), .Y(_0mem_offset_q_1_0__1_));
MUX2X1 MUX2X1_380 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2849_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2175_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2803_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__23_));
MUX2X1 MUX2X1_381 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2851_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2178_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2803_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__24_));
MUX2X1 MUX2X1_382 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2853_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2181_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2803_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__25_));
MUX2X1 MUX2X1_383 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2855_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2184_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2803_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__26_));
MUX2X1 MUX2X1_384 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2857_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2187_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2803_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__27_));
MUX2X1 MUX2X1_385 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2859_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2190_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2803_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__28_));
MUX2X1 MUX2X1_386 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2861_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2193_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2803_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__29_));
MUX2X1 MUX2X1_387 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2863_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2196_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2803_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__30_));
MUX2X1 MUX2X1_388 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2865_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2199_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2803_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__31_));
MUX2X1 MUX2X1_389 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2100_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2867_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2868_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__0_));
MUX2X1 MUX2X1_39 ( .A(_abc_40298_new_n2524_), .B(_abc_40298_new_n911_), .S(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2420), .Y(_0opcode_q_31_0__0_));
MUX2X1 MUX2X1_390 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2109_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2870_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2868_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__1_));
MUX2X1 MUX2X1_391 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2112_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2872_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2868_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__2_));
MUX2X1 MUX2X1_392 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2115_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2874_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2868_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__3_));
MUX2X1 MUX2X1_393 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2118_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2876_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2868_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__4_));
MUX2X1 MUX2X1_394 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2121_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2878_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2868_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__5_));
MUX2X1 MUX2X1_395 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2124_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2880_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2868_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__6_));
MUX2X1 MUX2X1_396 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2127_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2882_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2868_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__7_));
MUX2X1 MUX2X1_397 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2130_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2884_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2868_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__8_));
MUX2X1 MUX2X1_398 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2133_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2886_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2868_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__9_));
MUX2X1 MUX2X1_399 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2136_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2888_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2868_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__10_));
MUX2X1 MUX2X1_4 ( .A(_abc_40298_new_n1155_), .B(_abc_40298_new_n1152_), .S(_abc_40298_new_n1135_), .Y(_abc_40298_new_n1156_));
MUX2X1 MUX2X1_40 ( .A(_abc_40298_new_n694_), .B(_abc_40298_new_n909_), .S(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2420), .Y(_0opcode_q_31_0__1_));
MUX2X1 MUX2X1_400 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2139_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2890_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2868_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__11_));
MUX2X1 MUX2X1_401 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2142_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2892_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2868_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__12_));
MUX2X1 MUX2X1_402 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2145_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2894_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2868_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__13_));
MUX2X1 MUX2X1_403 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2148_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2896_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2868_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__14_));
MUX2X1 MUX2X1_404 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2151_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2898_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2868_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__15_));
MUX2X1 MUX2X1_405 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2154_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2900_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2868_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__16_));
MUX2X1 MUX2X1_406 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2157_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2902_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2868_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__17_));
MUX2X1 MUX2X1_407 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2160_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2904_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2868_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__18_));
MUX2X1 MUX2X1_408 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2163_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2906_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2868_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__19_));
MUX2X1 MUX2X1_409 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2166_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2908_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2868_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__20_));
MUX2X1 MUX2X1_41 ( .A(_abc_40298_new_n707_), .B(_abc_40298_new_n898_), .S(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2420), .Y(_0opcode_q_31_0__2_));
MUX2X1 MUX2X1_410 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2169_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2910_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2868_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__21_));
MUX2X1 MUX2X1_411 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2172_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2912_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2868_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__22_));
MUX2X1 MUX2X1_412 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2175_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2914_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2868_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__23_));
MUX2X1 MUX2X1_413 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2178_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2916_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2868_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__24_));
MUX2X1 MUX2X1_414 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2181_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2918_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2868_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__25_));
MUX2X1 MUX2X1_415 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2184_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2920_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2868_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__26_));
MUX2X1 MUX2X1_416 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2187_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2922_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2868_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__27_));
MUX2X1 MUX2X1_417 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2190_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2924_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2868_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__28_));
MUX2X1 MUX2X1_418 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2193_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2926_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2868_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__29_));
MUX2X1 MUX2X1_419 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2196_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2928_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2868_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__30_));
MUX2X1 MUX2X1_42 ( .A(_abc_40298_new_n718_), .B(_abc_40298_new_n903_), .S(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2420), .Y(_0opcode_q_31_0__3_));
MUX2X1 MUX2X1_420 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2199_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2930_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2868_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__31_));
MUX2X1 MUX2X1_421 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2932_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2100_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2936_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__0_));
MUX2X1 MUX2X1_422 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2938_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2109_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2936_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__1_));
MUX2X1 MUX2X1_423 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2940_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2112_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2936_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__2_));
MUX2X1 MUX2X1_424 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2942_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2115_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2936_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__3_));
MUX2X1 MUX2X1_425 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2944_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2118_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2936_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__4_));
MUX2X1 MUX2X1_426 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2946_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2121_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2936_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__5_));
MUX2X1 MUX2X1_427 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2948_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2124_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2936_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__6_));
MUX2X1 MUX2X1_428 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2950_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2127_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2936_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__7_));
MUX2X1 MUX2X1_429 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2952_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2130_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2936_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__8_));
MUX2X1 MUX2X1_43 ( .A(_abc_40298_new_n2530_), .B(_abc_40298_new_n1315_), .S(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2420), .Y(_0opcode_q_31_0__4_));
MUX2X1 MUX2X1_430 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2954_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2133_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2936_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__9_));
MUX2X1 MUX2X1_431 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2956_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2136_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2936_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__10_));
MUX2X1 MUX2X1_432 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2958_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2139_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2936_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__11_));
MUX2X1 MUX2X1_433 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2960_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2142_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2936_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__12_));
MUX2X1 MUX2X1_434 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2962_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2145_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2936_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__13_));
MUX2X1 MUX2X1_435 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2964_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2148_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2936_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__14_));
MUX2X1 MUX2X1_436 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2966_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2151_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2936_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__15_));
MUX2X1 MUX2X1_437 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2968_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2154_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2936_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__16_));
MUX2X1 MUX2X1_438 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2970_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2157_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2936_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__17_));
MUX2X1 MUX2X1_439 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2972_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2160_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2936_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__18_));
MUX2X1 MUX2X1_44 ( .A(_abc_40298_new_n2532_), .B(_abc_40298_new_n1341_), .S(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2420), .Y(_0opcode_q_31_0__5_));
MUX2X1 MUX2X1_440 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2974_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2163_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2936_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__19_));
MUX2X1 MUX2X1_441 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2976_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2166_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2936_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__20_));
MUX2X1 MUX2X1_442 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2978_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2169_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2936_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__21_));
MUX2X1 MUX2X1_443 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2980_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2172_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2936_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__22_));
MUX2X1 MUX2X1_444 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2982_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2175_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2936_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__23_));
MUX2X1 MUX2X1_445 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2984_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2178_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2936_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__24_));
MUX2X1 MUX2X1_446 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2986_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2181_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2936_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__25_));
MUX2X1 MUX2X1_447 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2988_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2184_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2936_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__26_));
MUX2X1 MUX2X1_448 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2990_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2187_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2936_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__27_));
MUX2X1 MUX2X1_449 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2992_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2190_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2936_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__28_));
MUX2X1 MUX2X1_45 ( .A(_abc_40298_new_n747_), .B(_abc_40298_new_n917_), .S(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2420), .Y(_0opcode_q_31_0__6_));
MUX2X1 MUX2X1_450 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2994_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2193_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2936_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__29_));
MUX2X1 MUX2X1_451 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2996_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2196_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2936_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__30_));
MUX2X1 MUX2X1_452 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2998_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2199_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2936_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__31_));
MUX2X1 MUX2X1_453 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2100_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3000_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3002_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__0_));
MUX2X1 MUX2X1_454 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2109_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3004_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3002_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__1_));
MUX2X1 MUX2X1_455 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2112_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3006_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3002_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__2_));
MUX2X1 MUX2X1_456 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2115_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3008_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3002_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__3_));
MUX2X1 MUX2X1_457 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2118_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3010_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3002_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__4_));
MUX2X1 MUX2X1_458 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2121_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3012_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3002_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__5_));
MUX2X1 MUX2X1_459 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2124_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3014_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3002_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__6_));
MUX2X1 MUX2X1_46 ( .A(_abc_40298_new_n2535_), .B(_abc_40298_new_n973_), .S(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2420), .Y(_0opcode_q_31_0__7_));
MUX2X1 MUX2X1_460 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2127_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3016_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3002_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__7_));
MUX2X1 MUX2X1_461 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2130_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3018_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3002_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__8_));
MUX2X1 MUX2X1_462 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2133_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3020_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3002_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__9_));
MUX2X1 MUX2X1_463 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2136_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3022_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3002_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__10_));
MUX2X1 MUX2X1_464 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2139_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3024_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3002_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__11_));
MUX2X1 MUX2X1_465 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2142_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3026_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3002_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__12_));
MUX2X1 MUX2X1_466 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2145_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3028_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3002_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__13_));
MUX2X1 MUX2X1_467 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2148_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3030_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3002_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__14_));
MUX2X1 MUX2X1_468 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2151_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3032_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3002_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__15_));
MUX2X1 MUX2X1_469 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2154_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3034_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3002_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__16_));
MUX2X1 MUX2X1_47 ( .A(_abc_40298_new_n2537_), .B(_abc_40298_new_n1455_), .S(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2420), .Y(_0opcode_q_31_0__8_));
MUX2X1 MUX2X1_470 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2157_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3036_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3002_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__17_));
MUX2X1 MUX2X1_471 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2160_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3038_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3002_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__18_));
MUX2X1 MUX2X1_472 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2163_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3040_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3002_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__19_));
MUX2X1 MUX2X1_473 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2166_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3042_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3002_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__20_));
MUX2X1 MUX2X1_474 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2169_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3044_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3002_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__21_));
MUX2X1 MUX2X1_475 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2172_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3046_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3002_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__22_));
MUX2X1 MUX2X1_476 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2175_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3048_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3002_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__23_));
MUX2X1 MUX2X1_477 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2178_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3050_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3002_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__24_));
MUX2X1 MUX2X1_478 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2181_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3052_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3002_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__25_));
MUX2X1 MUX2X1_479 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2184_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3054_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3002_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__26_));
MUX2X1 MUX2X1_48 ( .A(_abc_40298_new_n770_), .B(_abc_40298_new_n1457_), .S(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2420), .Y(_0opcode_q_31_0__9_));
MUX2X1 MUX2X1_480 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2187_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3056_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3002_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__27_));
MUX2X1 MUX2X1_481 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2190_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3058_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3002_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__28_));
MUX2X1 MUX2X1_482 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2193_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3060_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3002_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__29_));
MUX2X1 MUX2X1_483 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2196_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3062_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3002_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__30_));
MUX2X1 MUX2X1_484 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2199_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3064_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3002_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__31_));
MUX2X1 MUX2X1_485 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2100_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3066_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3068_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__0_));
MUX2X1 MUX2X1_486 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2109_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3070_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3068_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__1_));
MUX2X1 MUX2X1_487 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2112_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3072_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3068_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__2_));
MUX2X1 MUX2X1_488 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2115_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3074_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3068_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__3_));
MUX2X1 MUX2X1_489 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2118_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3076_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3068_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__4_));
MUX2X1 MUX2X1_49 ( .A(_abc_40298_new_n776_), .B(_abc_40298_new_n2456_), .S(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2420), .Y(_0opcode_q_31_0__10_));
MUX2X1 MUX2X1_490 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2121_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3078_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3068_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__5_));
MUX2X1 MUX2X1_491 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2124_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3080_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3068_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__6_));
MUX2X1 MUX2X1_492 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2127_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3082_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3068_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__7_));
MUX2X1 MUX2X1_493 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2130_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3084_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3068_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__8_));
MUX2X1 MUX2X1_494 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2133_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3086_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3068_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__9_));
MUX2X1 MUX2X1_495 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2136_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3088_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3068_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__10_));
MUX2X1 MUX2X1_496 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2139_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3090_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3068_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__11_));
MUX2X1 MUX2X1_497 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2142_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3092_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3068_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__12_));
MUX2X1 MUX2X1_498 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2145_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3094_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3068_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__13_));
MUX2X1 MUX2X1_499 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2148_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3096_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3068_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__14_));
MUX2X1 MUX2X1_5 ( .A(epc_q_2_), .B(REGFILE_SIM_reg_bank_reg_rb_o_2_), .S(_abc_40298_new_n1187_), .Y(_abc_40298_new_n1208_));
MUX2X1 MUX2X1_50 ( .A(_abc_40298_new_n781_), .B(_abc_40298_new_n1513_), .S(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2420), .Y(_0opcode_q_31_0__11_));
MUX2X1 MUX2X1_500 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2151_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3098_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3068_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__15_));
MUX2X1 MUX2X1_501 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2154_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3100_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3068_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__16_));
MUX2X1 MUX2X1_502 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2157_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3102_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3068_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__17_));
MUX2X1 MUX2X1_503 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2160_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3104_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3068_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__18_));
MUX2X1 MUX2X1_504 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2163_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3106_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3068_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__19_));
MUX2X1 MUX2X1_505 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2166_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3108_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3068_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__20_));
MUX2X1 MUX2X1_506 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2169_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3110_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3068_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__21_));
MUX2X1 MUX2X1_507 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2172_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3112_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3068_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__22_));
MUX2X1 MUX2X1_508 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2175_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3114_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3068_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__23_));
MUX2X1 MUX2X1_509 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2178_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3116_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3068_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__24_));
MUX2X1 MUX2X1_51 ( .A(_abc_40298_new_n2542_), .B(_abc_40298_new_n2471_), .S(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2420), .Y(_0opcode_q_31_0__12_));
MUX2X1 MUX2X1_510 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2181_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3118_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3068_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__25_));
MUX2X1 MUX2X1_511 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2184_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3120_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3068_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__26_));
MUX2X1 MUX2X1_512 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2187_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3122_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3068_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__27_));
MUX2X1 MUX2X1_513 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2190_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3124_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3068_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__28_));
MUX2X1 MUX2X1_514 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2193_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3126_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3068_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__29_));
MUX2X1 MUX2X1_515 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2196_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3128_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3068_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__30_));
MUX2X1 MUX2X1_516 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2199_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3130_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3068_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__31_));
MUX2X1 MUX2X1_517 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3132_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2100_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3133_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__0_));
MUX2X1 MUX2X1_518 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3135_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2109_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3133_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__1_));
MUX2X1 MUX2X1_519 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3137_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2112_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3133_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__2_));
MUX2X1 MUX2X1_52 ( .A(_abc_40298_new_n2544_), .B(_abc_40298_new_n2479_), .S(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2420), .Y(_0opcode_q_31_0__13_));
MUX2X1 MUX2X1_520 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3139_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2115_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3133_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__3_));
MUX2X1 MUX2X1_521 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3141_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2118_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3133_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__4_));
MUX2X1 MUX2X1_522 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3143_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2121_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3133_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__5_));
MUX2X1 MUX2X1_523 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3145_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2124_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3133_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__6_));
MUX2X1 MUX2X1_524 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3147_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2127_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3133_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__7_));
MUX2X1 MUX2X1_525 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3149_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2130_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3133_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__8_));
MUX2X1 MUX2X1_526 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3151_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2133_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3133_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__9_));
MUX2X1 MUX2X1_527 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3153_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2136_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3133_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__10_));
MUX2X1 MUX2X1_528 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3155_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2139_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3133_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__11_));
MUX2X1 MUX2X1_529 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3157_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2142_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3133_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__12_));
MUX2X1 MUX2X1_53 ( .A(_abc_40298_new_n794_), .B(_abc_40298_new_n1604_), .S(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2420), .Y(_0opcode_q_31_0__14_));
MUX2X1 MUX2X1_530 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3159_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2145_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3133_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__13_));
MUX2X1 MUX2X1_531 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3161_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2148_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3133_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__14_));
MUX2X1 MUX2X1_532 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3163_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2151_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3133_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__15_));
MUX2X1 MUX2X1_533 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3165_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2154_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3133_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__16_));
MUX2X1 MUX2X1_534 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3167_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2157_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3133_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__17_));
MUX2X1 MUX2X1_535 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3169_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2160_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3133_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__18_));
MUX2X1 MUX2X1_536 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3171_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2163_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3133_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__19_));
MUX2X1 MUX2X1_537 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3173_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2166_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3133_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__20_));
MUX2X1 MUX2X1_538 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3175_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2169_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3133_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__21_));
MUX2X1 MUX2X1_539 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3177_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2172_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3133_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__22_));
MUX2X1 MUX2X1_54 ( .A(_abc_40298_new_n2547_), .B(_abc_40298_new_n1628_), .S(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2420), .Y(_0opcode_q_31_0__15_));
MUX2X1 MUX2X1_540 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3179_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2175_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3133_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__23_));
MUX2X1 MUX2X1_541 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3181_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2178_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3133_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__24_));
MUX2X1 MUX2X1_542 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3183_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2181_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3133_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__25_));
MUX2X1 MUX2X1_543 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3185_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2184_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3133_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__26_));
MUX2X1 MUX2X1_544 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3187_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2187_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3133_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__27_));
MUX2X1 MUX2X1_545 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3189_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2190_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3133_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__28_));
MUX2X1 MUX2X1_546 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3191_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2193_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3133_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__29_));
MUX2X1 MUX2X1_547 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3193_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2196_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3133_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__30_));
MUX2X1 MUX2X1_548 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3195_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2199_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3133_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__31_));
MUX2X1 MUX2X1_549 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3197_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2100_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3200_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__0_));
MUX2X1 MUX2X1_55 ( .A(_abc_40298_new_n805_), .B(_abc_40298_new_n1658_), .S(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2420), .Y(_0opcode_q_31_0__16_));
MUX2X1 MUX2X1_550 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3202_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2109_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3200_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__1_));
MUX2X1 MUX2X1_551 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3204_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2112_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3200_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__2_));
MUX2X1 MUX2X1_552 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3206_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2115_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3200_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__3_));
MUX2X1 MUX2X1_553 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3208_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2118_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3200_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__4_));
MUX2X1 MUX2X1_554 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3210_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2121_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3200_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__5_));
MUX2X1 MUX2X1_555 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3212_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2124_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3200_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__6_));
MUX2X1 MUX2X1_556 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3214_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2127_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3200_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__7_));
MUX2X1 MUX2X1_557 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3216_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2130_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3200_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__8_));
MUX2X1 MUX2X1_558 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3218_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2133_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3200_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__9_));
MUX2X1 MUX2X1_559 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3220_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2136_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3200_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__10_));
MUX2X1 MUX2X1_56 ( .A(_abc_40298_new_n810_), .B(_abc_40298_new_n1683_), .S(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2420), .Y(_0opcode_q_31_0__17_));
MUX2X1 MUX2X1_560 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3222_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2139_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3200_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__11_));
MUX2X1 MUX2X1_561 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3224_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2142_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3200_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__12_));
MUX2X1 MUX2X1_562 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3226_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2145_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3200_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__13_));
MUX2X1 MUX2X1_563 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3228_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2148_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3200_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__14_));
MUX2X1 MUX2X1_564 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3230_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2151_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3200_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__15_));
MUX2X1 MUX2X1_565 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3232_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2154_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3200_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__16_));
MUX2X1 MUX2X1_566 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3234_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2157_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3200_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__17_));
MUX2X1 MUX2X1_567 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3236_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2160_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3200_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__18_));
MUX2X1 MUX2X1_568 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3238_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2163_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3200_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__19_));
MUX2X1 MUX2X1_569 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3240_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2166_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3200_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__20_));
MUX2X1 MUX2X1_57 ( .A(_abc_40298_new_n815_), .B(_abc_40298_new_n1712_), .S(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2420), .Y(_0opcode_q_31_0__18_));
MUX2X1 MUX2X1_570 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3242_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2169_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3200_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__21_));
MUX2X1 MUX2X1_571 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3244_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2172_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3200_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__22_));
MUX2X1 MUX2X1_572 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3246_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2175_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3200_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__23_));
MUX2X1 MUX2X1_573 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3248_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2178_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3200_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__24_));
MUX2X1 MUX2X1_574 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3250_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2181_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3200_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__25_));
MUX2X1 MUX2X1_575 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3252_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2184_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3200_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__26_));
MUX2X1 MUX2X1_576 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3254_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2187_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3200_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__27_));
MUX2X1 MUX2X1_577 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3256_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2190_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3200_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__28_));
MUX2X1 MUX2X1_578 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3258_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2193_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3200_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__29_));
MUX2X1 MUX2X1_579 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3260_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2196_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3200_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__30_));
MUX2X1 MUX2X1_58 ( .A(_abc_40298_new_n820_), .B(_abc_40298_new_n1735_), .S(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2420), .Y(_0opcode_q_31_0__19_));
MUX2X1 MUX2X1_580 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3262_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2199_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3200_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__31_));
MUX2X1 MUX2X1_581 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3264_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2100_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3265_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__0_));
MUX2X1 MUX2X1_582 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3267_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2109_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3265_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__1_));
MUX2X1 MUX2X1_583 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3269_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2112_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3265_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__2_));
MUX2X1 MUX2X1_584 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3271_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2115_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3265_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__3_));
MUX2X1 MUX2X1_585 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3273_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2118_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3265_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__4_));
MUX2X1 MUX2X1_586 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3275_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2121_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3265_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__5_));
MUX2X1 MUX2X1_587 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3277_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2124_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3265_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__6_));
MUX2X1 MUX2X1_588 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3279_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2127_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3265_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__7_));
MUX2X1 MUX2X1_589 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3281_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2130_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3265_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__8_));
MUX2X1 MUX2X1_59 ( .A(_abc_40298_new_n825_), .B(_abc_40298_new_n1766_), .S(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2420), .Y(_0opcode_q_31_0__20_));
MUX2X1 MUX2X1_590 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3283_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2133_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3265_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__9_));
MUX2X1 MUX2X1_591 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3285_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2136_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3265_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__10_));
MUX2X1 MUX2X1_592 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3287_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2139_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3265_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__11_));
MUX2X1 MUX2X1_593 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3289_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2142_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3265_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__12_));
MUX2X1 MUX2X1_594 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3291_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2145_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3265_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__13_));
MUX2X1 MUX2X1_595 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3293_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2148_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3265_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__14_));
MUX2X1 MUX2X1_596 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3295_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2151_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3265_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__15_));
MUX2X1 MUX2X1_597 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3297_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2154_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3265_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__16_));
MUX2X1 MUX2X1_598 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3299_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2157_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3265_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__17_));
MUX2X1 MUX2X1_599 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3301_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2160_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3265_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__18_));
MUX2X1 MUX2X1_6 ( .A(_abc_40298_new_n1244_), .B(_abc_40298_new_n1231_), .S(_abc_40298_new_n1134_), .Y(_abc_40298_new_n1245_));
MUX2X1 MUX2X1_60 ( .A(_abc_40298_new_n830_), .B(_abc_40298_new_n949_), .S(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2420), .Y(_0opcode_q_31_0__21_));
MUX2X1 MUX2X1_600 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3303_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2163_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3265_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__19_));
MUX2X1 MUX2X1_601 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3305_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2166_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3265_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__20_));
MUX2X1 MUX2X1_602 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3307_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2169_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3265_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__21_));
MUX2X1 MUX2X1_603 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3309_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2172_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3265_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__22_));
MUX2X1 MUX2X1_604 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3311_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2175_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3265_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__23_));
MUX2X1 MUX2X1_605 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3313_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2178_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3265_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__24_));
MUX2X1 MUX2X1_606 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3315_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2181_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3265_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__25_));
MUX2X1 MUX2X1_607 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3317_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2184_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3265_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__26_));
MUX2X1 MUX2X1_608 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3319_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2187_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3265_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__27_));
MUX2X1 MUX2X1_609 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3321_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2190_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3265_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__28_));
MUX2X1 MUX2X1_61 ( .A(_abc_40298_new_n835_), .B(_abc_40298_new_n944_), .S(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2420), .Y(_0opcode_q_31_0__22_));
MUX2X1 MUX2X1_610 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3323_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2193_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3265_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__29_));
MUX2X1 MUX2X1_611 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3325_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2196_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3265_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__30_));
MUX2X1 MUX2X1_612 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3327_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2199_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3265_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__31_));
MUX2X1 MUX2X1_613 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3329_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2100_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3330_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__0_));
MUX2X1 MUX2X1_614 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3332_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2109_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3330_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__1_));
MUX2X1 MUX2X1_615 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3334_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2112_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3330_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__2_));
MUX2X1 MUX2X1_616 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3336_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2115_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3330_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__3_));
MUX2X1 MUX2X1_617 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3338_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2118_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3330_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__4_));
MUX2X1 MUX2X1_618 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3340_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2121_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3330_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__5_));
MUX2X1 MUX2X1_619 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3342_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2124_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3330_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__6_));
MUX2X1 MUX2X1_62 ( .A(_abc_40298_new_n840_), .B(_abc_40298_new_n938_), .S(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2420), .Y(_0opcode_q_31_0__23_));
MUX2X1 MUX2X1_620 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3344_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2127_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3330_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__7_));
MUX2X1 MUX2X1_621 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3346_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2130_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3330_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__8_));
MUX2X1 MUX2X1_622 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3348_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2133_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3330_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__9_));
MUX2X1 MUX2X1_623 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3350_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2136_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3330_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__10_));
MUX2X1 MUX2X1_624 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3352_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2139_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3330_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__11_));
MUX2X1 MUX2X1_625 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3354_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2142_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3330_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__12_));
MUX2X1 MUX2X1_626 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3356_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2145_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3330_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__13_));
MUX2X1 MUX2X1_627 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3358_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2148_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3330_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__14_));
MUX2X1 MUX2X1_628 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3360_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2151_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3330_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__15_));
MUX2X1 MUX2X1_629 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3362_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2154_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3330_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__16_));
MUX2X1 MUX2X1_63 ( .A(_abc_40298_new_n845_), .B(_abc_40298_new_n623_), .S(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2420), .Y(_0opcode_q_31_0__24_));
MUX2X1 MUX2X1_630 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3364_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2157_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3330_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__17_));
MUX2X1 MUX2X1_631 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3366_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2160_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3330_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__18_));
MUX2X1 MUX2X1_632 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3368_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2163_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3330_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__19_));
MUX2X1 MUX2X1_633 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3370_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2166_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3330_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__20_));
MUX2X1 MUX2X1_634 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3372_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2169_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3330_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__21_));
MUX2X1 MUX2X1_635 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3374_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2172_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3330_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__22_));
MUX2X1 MUX2X1_636 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3376_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2175_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3330_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__23_));
MUX2X1 MUX2X1_637 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3378_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2178_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3330_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__24_));
MUX2X1 MUX2X1_638 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3380_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2181_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3330_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__25_));
MUX2X1 MUX2X1_639 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3382_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2184_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3330_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__26_));
MUX2X1 MUX2X1_64 ( .A(_abc_40298_new_n850_), .B(_abc_40298_new_n624_), .S(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2420), .Y(_0opcode_q_31_0__25_));
MUX2X1 MUX2X1_640 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3384_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2187_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3330_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__27_));
MUX2X1 MUX2X1_641 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3386_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2190_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3330_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__28_));
MUX2X1 MUX2X1_642 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3388_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2193_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3330_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__29_));
MUX2X1 MUX2X1_643 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3390_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2196_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3330_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__30_));
MUX2X1 MUX2X1_644 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3392_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2199_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3330_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__31_));
MUX2X1 MUX2X1_645 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2100_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3394_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3396_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__0_));
MUX2X1 MUX2X1_646 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2109_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3398_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3396_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__1_));
MUX2X1 MUX2X1_647 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2112_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3400_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3396_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__2_));
MUX2X1 MUX2X1_648 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2115_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3402_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3396_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__3_));
MUX2X1 MUX2X1_649 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2118_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3404_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3396_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__4_));
MUX2X1 MUX2X1_65 ( .A(_abc_40298_new_n860_), .B(_abc_40298_new_n656_), .S(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2420), .Y(_0opcode_q_31_0__27_));
MUX2X1 MUX2X1_650 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2121_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3406_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3396_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__5_));
MUX2X1 MUX2X1_651 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2124_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3408_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3396_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__6_));
MUX2X1 MUX2X1_652 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2127_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3410_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3396_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__7_));
MUX2X1 MUX2X1_653 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2130_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3412_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3396_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__8_));
MUX2X1 MUX2X1_654 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2133_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3414_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3396_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__9_));
MUX2X1 MUX2X1_655 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2136_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3416_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3396_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__10_));
MUX2X1 MUX2X1_656 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2139_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3418_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3396_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__11_));
MUX2X1 MUX2X1_657 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2142_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3420_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3396_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__12_));
MUX2X1 MUX2X1_658 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2145_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3422_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3396_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__13_));
MUX2X1 MUX2X1_659 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2148_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3424_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3396_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__14_));
MUX2X1 MUX2X1_66 ( .A(_abc_40298_new_n870_), .B(_abc_40298_new_n619_), .S(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2420), .Y(_0opcode_q_31_0__29_));
MUX2X1 MUX2X1_660 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2151_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3426_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3396_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__15_));
MUX2X1 MUX2X1_661 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2154_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3428_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3396_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__16_));
MUX2X1 MUX2X1_662 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2157_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3430_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3396_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__17_));
MUX2X1 MUX2X1_663 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2160_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3432_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3396_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__18_));
MUX2X1 MUX2X1_664 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2163_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3434_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3396_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__19_));
MUX2X1 MUX2X1_665 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2166_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3436_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3396_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__20_));
MUX2X1 MUX2X1_666 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2169_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3438_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3396_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__21_));
MUX2X1 MUX2X1_667 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2172_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3440_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3396_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__22_));
MUX2X1 MUX2X1_668 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2175_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3442_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3396_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__23_));
MUX2X1 MUX2X1_669 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2178_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3444_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3396_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__24_));
MUX2X1 MUX2X1_67 ( .A(_abc_40298_new_n875_), .B(_abc_40298_new_n637_), .S(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2420), .Y(_0opcode_q_31_0__30_));
MUX2X1 MUX2X1_670 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2181_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3446_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3396_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__25_));
MUX2X1 MUX2X1_671 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2184_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3448_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3396_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__26_));
MUX2X1 MUX2X1_672 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2187_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3450_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3396_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__27_));
MUX2X1 MUX2X1_673 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2190_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3452_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3396_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__28_));
MUX2X1 MUX2X1_674 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2193_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3454_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3396_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__29_));
MUX2X1 MUX2X1_675 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2196_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3456_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3396_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__30_));
MUX2X1 MUX2X1_676 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2199_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3458_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3396_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__31_));
MUX2X1 MUX2X1_677 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3460_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2100_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3461_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__0_));
MUX2X1 MUX2X1_678 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3463_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2109_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3461_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__1_));
MUX2X1 MUX2X1_679 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3465_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2112_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3461_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__2_));
MUX2X1 MUX2X1_68 ( .A(_abc_40298_new_n880_), .B(_abc_40298_new_n638_), .S(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2420), .Y(_0opcode_q_31_0__31_));
MUX2X1 MUX2X1_680 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3467_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2115_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3461_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__3_));
MUX2X1 MUX2X1_681 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3469_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2118_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3461_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__4_));
MUX2X1 MUX2X1_682 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3471_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2121_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3461_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__5_));
MUX2X1 MUX2X1_683 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3473_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2124_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3461_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__6_));
MUX2X1 MUX2X1_684 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3475_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2127_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3461_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__7_));
MUX2X1 MUX2X1_685 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3477_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2130_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3461_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__8_));
MUX2X1 MUX2X1_686 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3479_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2133_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3461_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__9_));
MUX2X1 MUX2X1_687 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3481_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2136_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3461_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__10_));
MUX2X1 MUX2X1_688 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3483_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2139_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3461_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__11_));
MUX2X1 MUX2X1_689 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3485_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2142_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3461_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__12_));
MUX2X1 MUX2X1_69 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2099_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2100_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2106_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__0_));
MUX2X1 MUX2X1_690 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3487_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2145_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3461_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__13_));
MUX2X1 MUX2X1_691 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3489_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2148_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3461_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__14_));
MUX2X1 MUX2X1_692 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3491_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2151_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3461_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__15_));
MUX2X1 MUX2X1_693 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3493_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2154_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3461_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__16_));
MUX2X1 MUX2X1_694 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3495_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2157_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3461_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__17_));
MUX2X1 MUX2X1_695 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3497_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2160_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3461_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__18_));
MUX2X1 MUX2X1_696 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3499_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2163_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3461_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__19_));
MUX2X1 MUX2X1_697 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3501_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2166_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3461_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__20_));
MUX2X1 MUX2X1_698 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3503_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2169_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3461_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__21_));
MUX2X1 MUX2X1_699 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3505_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2172_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3461_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__22_));
MUX2X1 MUX2X1_7 ( .A(epc_q_6_), .B(REGFILE_SIM_reg_bank_reg_rb_o_6_), .S(_abc_40298_new_n1187_), .Y(_abc_40298_new_n1326_));
MUX2X1 MUX2X1_70 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2108_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2109_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2106_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__1_));
MUX2X1 MUX2X1_700 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3507_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2175_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3461_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__23_));
MUX2X1 MUX2X1_701 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3509_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2178_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3461_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__24_));
MUX2X1 MUX2X1_702 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3511_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2181_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3461_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__25_));
MUX2X1 MUX2X1_703 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3513_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2184_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3461_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__26_));
MUX2X1 MUX2X1_704 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3515_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2187_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3461_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__27_));
MUX2X1 MUX2X1_705 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3517_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2190_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3461_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__28_));
MUX2X1 MUX2X1_706 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3519_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2193_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3461_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__29_));
MUX2X1 MUX2X1_707 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3521_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2196_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3461_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__30_));
MUX2X1 MUX2X1_708 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3523_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2199_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3461_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__31_));
MUX2X1 MUX2X1_709 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3525_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2100_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3526_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__0_));
MUX2X1 MUX2X1_71 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2111_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2112_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2106_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__2_));
MUX2X1 MUX2X1_710 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3528_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2109_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3526_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__1_));
MUX2X1 MUX2X1_711 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3530_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2112_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3526_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__2_));
MUX2X1 MUX2X1_712 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3532_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2115_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3526_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__3_));
MUX2X1 MUX2X1_713 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3534_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2118_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3526_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__4_));
MUX2X1 MUX2X1_714 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3536_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2121_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3526_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__5_));
MUX2X1 MUX2X1_715 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3538_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2124_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3526_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__6_));
MUX2X1 MUX2X1_716 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3540_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2127_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3526_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__7_));
MUX2X1 MUX2X1_717 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3542_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2130_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3526_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__8_));
MUX2X1 MUX2X1_718 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3544_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2133_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3526_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__9_));
MUX2X1 MUX2X1_719 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3546_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2136_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3526_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__10_));
MUX2X1 MUX2X1_72 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2114_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2115_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2106_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__3_));
MUX2X1 MUX2X1_720 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3548_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2139_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3526_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__11_));
MUX2X1 MUX2X1_721 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3550_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2142_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3526_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__12_));
MUX2X1 MUX2X1_722 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3552_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2145_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3526_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__13_));
MUX2X1 MUX2X1_723 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3554_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2148_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3526_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__14_));
MUX2X1 MUX2X1_724 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3556_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2151_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3526_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__15_));
MUX2X1 MUX2X1_725 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3558_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2154_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3526_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__16_));
MUX2X1 MUX2X1_726 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3560_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2157_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3526_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__17_));
MUX2X1 MUX2X1_727 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3562_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2160_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3526_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__18_));
MUX2X1 MUX2X1_728 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3564_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2163_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3526_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__19_));
MUX2X1 MUX2X1_729 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3566_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2166_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3526_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__20_));
MUX2X1 MUX2X1_73 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2117_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2118_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2106_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__4_));
MUX2X1 MUX2X1_730 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3568_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2169_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3526_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__21_));
MUX2X1 MUX2X1_731 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3570_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2172_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3526_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__22_));
MUX2X1 MUX2X1_732 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3572_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2175_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3526_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__23_));
MUX2X1 MUX2X1_733 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3574_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2178_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3526_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__24_));
MUX2X1 MUX2X1_734 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3576_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2181_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3526_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__25_));
MUX2X1 MUX2X1_735 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3578_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2184_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3526_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__26_));
MUX2X1 MUX2X1_736 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3580_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2187_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3526_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__27_));
MUX2X1 MUX2X1_737 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3582_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2190_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3526_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__28_));
MUX2X1 MUX2X1_738 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3584_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2193_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3526_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__29_));
MUX2X1 MUX2X1_739 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3586_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2196_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3526_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__30_));
MUX2X1 MUX2X1_74 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2120_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2121_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2106_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__5_));
MUX2X1 MUX2X1_740 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3588_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2199_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3526_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__31_));
MUX2X1 MUX2X1_741 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2100_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3590_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3592_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__0_));
MUX2X1 MUX2X1_742 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2109_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3594_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3592_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__1_));
MUX2X1 MUX2X1_743 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2112_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3596_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3592_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__2_));
MUX2X1 MUX2X1_744 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2115_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3598_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3592_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__3_));
MUX2X1 MUX2X1_745 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2118_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3600_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3592_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__4_));
MUX2X1 MUX2X1_746 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2121_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3602_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3592_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__5_));
MUX2X1 MUX2X1_747 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2124_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3604_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3592_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__6_));
MUX2X1 MUX2X1_748 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2127_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3606_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3592_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__7_));
MUX2X1 MUX2X1_749 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2130_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3608_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3592_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__8_));
MUX2X1 MUX2X1_75 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2123_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2124_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2106_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__6_));
MUX2X1 MUX2X1_750 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2133_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3610_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3592_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__9_));
MUX2X1 MUX2X1_751 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2136_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3612_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3592_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__10_));
MUX2X1 MUX2X1_752 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2139_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3614_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3592_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__11_));
MUX2X1 MUX2X1_753 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2142_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3616_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3592_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__12_));
MUX2X1 MUX2X1_754 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2145_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3618_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3592_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__13_));
MUX2X1 MUX2X1_755 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2148_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3620_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3592_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__14_));
MUX2X1 MUX2X1_756 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2151_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3622_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3592_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__15_));
MUX2X1 MUX2X1_757 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2154_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3624_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3592_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__16_));
MUX2X1 MUX2X1_758 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2157_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3626_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3592_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__17_));
MUX2X1 MUX2X1_759 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2160_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3628_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3592_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__18_));
MUX2X1 MUX2X1_76 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2126_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2127_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2106_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__7_));
MUX2X1 MUX2X1_760 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2163_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3630_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3592_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__19_));
MUX2X1 MUX2X1_761 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2166_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3632_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3592_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__20_));
MUX2X1 MUX2X1_762 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2169_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3634_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3592_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__21_));
MUX2X1 MUX2X1_763 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2172_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3636_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3592_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__22_));
MUX2X1 MUX2X1_764 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2175_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3638_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3592_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__23_));
MUX2X1 MUX2X1_765 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2178_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3640_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3592_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__24_));
MUX2X1 MUX2X1_766 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2181_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3642_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3592_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__25_));
MUX2X1 MUX2X1_767 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2184_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3644_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3592_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__26_));
MUX2X1 MUX2X1_768 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2187_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3646_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3592_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__27_));
MUX2X1 MUX2X1_769 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2190_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3648_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3592_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__28_));
MUX2X1 MUX2X1_77 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2129_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2130_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2106_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__8_));
MUX2X1 MUX2X1_770 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2193_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3650_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3592_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__29_));
MUX2X1 MUX2X1_771 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2196_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3652_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3592_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__30_));
MUX2X1 MUX2X1_772 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2199_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3654_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3592_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__31_));
MUX2X1 MUX2X1_773 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3656_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2100_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3657_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__0_));
MUX2X1 MUX2X1_774 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3659_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2109_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3657_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__1_));
MUX2X1 MUX2X1_775 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3661_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2112_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3657_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__2_));
MUX2X1 MUX2X1_776 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3663_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2115_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3657_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__3_));
MUX2X1 MUX2X1_777 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3665_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2118_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3657_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__4_));
MUX2X1 MUX2X1_778 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3667_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2121_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3657_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__5_));
MUX2X1 MUX2X1_779 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3669_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2124_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3657_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__6_));
MUX2X1 MUX2X1_78 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2132_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2133_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2106_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__9_));
MUX2X1 MUX2X1_780 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3671_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2127_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3657_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__7_));
MUX2X1 MUX2X1_781 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3673_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2130_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3657_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__8_));
MUX2X1 MUX2X1_782 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3675_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2133_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3657_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__9_));
MUX2X1 MUX2X1_783 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3677_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2136_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3657_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__10_));
MUX2X1 MUX2X1_784 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3679_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2139_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3657_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__11_));
MUX2X1 MUX2X1_785 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3681_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2142_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3657_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__12_));
MUX2X1 MUX2X1_786 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3683_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2145_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3657_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__13_));
MUX2X1 MUX2X1_787 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3685_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2148_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3657_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__14_));
MUX2X1 MUX2X1_788 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3687_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2151_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3657_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__15_));
MUX2X1 MUX2X1_789 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3689_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2154_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3657_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__16_));
MUX2X1 MUX2X1_79 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2135_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2136_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2106_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__10_));
MUX2X1 MUX2X1_790 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3691_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2157_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3657_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__17_));
MUX2X1 MUX2X1_791 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3693_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2160_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3657_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__18_));
MUX2X1 MUX2X1_792 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3695_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2163_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3657_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__19_));
MUX2X1 MUX2X1_793 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3697_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2166_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3657_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__20_));
MUX2X1 MUX2X1_794 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3699_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2169_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3657_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__21_));
MUX2X1 MUX2X1_795 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3701_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2172_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3657_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__22_));
MUX2X1 MUX2X1_796 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3703_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2175_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3657_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__23_));
MUX2X1 MUX2X1_797 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3705_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2178_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3657_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__24_));
MUX2X1 MUX2X1_798 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3707_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2181_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3657_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__25_));
MUX2X1 MUX2X1_799 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3709_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2184_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3657_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__26_));
MUX2X1 MUX2X1_8 ( .A(epc_q_7_), .B(REGFILE_SIM_reg_bank_reg_rb_o_7_), .S(_abc_40298_new_n1187_), .Y(_abc_40298_new_n1336_));
MUX2X1 MUX2X1_80 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2138_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2139_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2106_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__11_));
MUX2X1 MUX2X1_800 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3711_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2187_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3657_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__27_));
MUX2X1 MUX2X1_801 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3713_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2190_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3657_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__28_));
MUX2X1 MUX2X1_802 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3715_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2193_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3657_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__29_));
MUX2X1 MUX2X1_803 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3717_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2196_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3657_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__30_));
MUX2X1 MUX2X1_804 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3719_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2199_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3657_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__31_));
MUX2X1 MUX2X1_805 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2100_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3721_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3722_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__0_));
MUX2X1 MUX2X1_806 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2109_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3724_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3722_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__1_));
MUX2X1 MUX2X1_807 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2112_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3726_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3722_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__2_));
MUX2X1 MUX2X1_808 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2115_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3728_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3722_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__3_));
MUX2X1 MUX2X1_809 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2118_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3730_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3722_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__4_));
MUX2X1 MUX2X1_81 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2141_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2142_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2106_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__12_));
MUX2X1 MUX2X1_810 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2121_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3732_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3722_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__5_));
MUX2X1 MUX2X1_811 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2124_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3734_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3722_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__6_));
MUX2X1 MUX2X1_812 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2127_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3736_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3722_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__7_));
MUX2X1 MUX2X1_813 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2130_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3738_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3722_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__8_));
MUX2X1 MUX2X1_814 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2133_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3740_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3722_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__9_));
MUX2X1 MUX2X1_815 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2136_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3742_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3722_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__10_));
MUX2X1 MUX2X1_816 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2139_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3744_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3722_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__11_));
MUX2X1 MUX2X1_817 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2142_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3746_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3722_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__12_));
MUX2X1 MUX2X1_818 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2145_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3748_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3722_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__13_));
MUX2X1 MUX2X1_819 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2148_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3750_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3722_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__14_));
MUX2X1 MUX2X1_82 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2144_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2145_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2106_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__13_));
MUX2X1 MUX2X1_820 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2151_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3752_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3722_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__15_));
MUX2X1 MUX2X1_821 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2154_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3754_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3722_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__16_));
MUX2X1 MUX2X1_822 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2157_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3756_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3722_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__17_));
MUX2X1 MUX2X1_823 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2160_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3758_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3722_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__18_));
MUX2X1 MUX2X1_824 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2163_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3760_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3722_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__19_));
MUX2X1 MUX2X1_825 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2166_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3762_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3722_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__20_));
MUX2X1 MUX2X1_826 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2169_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3764_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3722_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__21_));
MUX2X1 MUX2X1_827 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2172_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3766_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3722_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__22_));
MUX2X1 MUX2X1_828 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2175_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3768_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3722_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__23_));
MUX2X1 MUX2X1_829 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2178_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3770_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3722_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__24_));
MUX2X1 MUX2X1_83 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2147_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2148_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2106_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__14_));
MUX2X1 MUX2X1_830 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2181_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3772_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3722_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__25_));
MUX2X1 MUX2X1_831 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2184_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3774_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3722_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__26_));
MUX2X1 MUX2X1_832 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2187_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3776_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3722_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__27_));
MUX2X1 MUX2X1_833 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2190_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3778_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3722_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__28_));
MUX2X1 MUX2X1_834 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2193_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3780_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3722_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__29_));
MUX2X1 MUX2X1_835 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2196_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3782_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3722_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__30_));
MUX2X1 MUX2X1_836 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2199_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3784_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3722_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__31_));
MUX2X1 MUX2X1_837 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3786_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2100_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3787_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__0_));
MUX2X1 MUX2X1_838 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3789_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2109_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3787_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__1_));
MUX2X1 MUX2X1_839 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3791_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2112_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3787_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__2_));
MUX2X1 MUX2X1_84 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2150_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2151_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2106_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__15_));
MUX2X1 MUX2X1_840 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3793_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2115_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3787_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__3_));
MUX2X1 MUX2X1_841 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3795_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2118_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3787_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__4_));
MUX2X1 MUX2X1_842 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3797_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2121_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3787_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__5_));
MUX2X1 MUX2X1_843 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3799_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2124_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3787_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__6_));
MUX2X1 MUX2X1_844 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3801_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2127_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3787_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__7_));
MUX2X1 MUX2X1_845 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3803_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2130_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3787_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__8_));
MUX2X1 MUX2X1_846 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3805_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2133_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3787_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__9_));
MUX2X1 MUX2X1_847 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3807_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2136_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3787_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__10_));
MUX2X1 MUX2X1_848 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3809_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2139_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3787_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__11_));
MUX2X1 MUX2X1_849 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3811_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2142_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3787_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__12_));
MUX2X1 MUX2X1_85 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2153_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2154_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2106_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__16_));
MUX2X1 MUX2X1_850 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3813_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2145_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3787_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__13_));
MUX2X1 MUX2X1_851 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3815_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2148_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3787_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__14_));
MUX2X1 MUX2X1_852 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3817_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2151_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3787_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__15_));
MUX2X1 MUX2X1_853 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3819_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2154_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3787_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__16_));
MUX2X1 MUX2X1_854 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3821_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2157_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3787_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__17_));
MUX2X1 MUX2X1_855 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3823_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2160_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3787_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__18_));
MUX2X1 MUX2X1_856 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3825_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2163_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3787_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__19_));
MUX2X1 MUX2X1_857 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3827_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2166_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3787_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__20_));
MUX2X1 MUX2X1_858 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3829_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2169_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3787_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__21_));
MUX2X1 MUX2X1_859 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3831_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2172_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3787_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__22_));
MUX2X1 MUX2X1_86 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2156_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2157_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2106_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__17_));
MUX2X1 MUX2X1_860 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3833_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2175_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3787_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__23_));
MUX2X1 MUX2X1_861 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3835_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2178_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3787_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__24_));
MUX2X1 MUX2X1_862 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3837_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2181_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3787_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__25_));
MUX2X1 MUX2X1_863 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3839_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2184_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3787_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__26_));
MUX2X1 MUX2X1_864 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3841_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2187_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3787_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__27_));
MUX2X1 MUX2X1_865 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3843_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2190_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3787_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__28_));
MUX2X1 MUX2X1_866 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3845_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2193_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3787_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__29_));
MUX2X1 MUX2X1_867 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3847_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2196_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3787_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__30_));
MUX2X1 MUX2X1_868 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3849_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2199_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3787_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__31_));
MUX2X1 MUX2X1_869 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3851_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2100_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3852_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__0_));
MUX2X1 MUX2X1_87 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2159_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2160_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2106_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__18_));
MUX2X1 MUX2X1_870 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3854_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2109_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3852_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__1_));
MUX2X1 MUX2X1_871 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3856_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2112_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3852_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__2_));
MUX2X1 MUX2X1_872 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3858_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2115_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3852_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__3_));
MUX2X1 MUX2X1_873 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3860_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2118_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3852_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__4_));
MUX2X1 MUX2X1_874 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3862_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2121_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3852_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__5_));
MUX2X1 MUX2X1_875 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3864_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2124_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3852_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__6_));
MUX2X1 MUX2X1_876 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3866_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2127_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3852_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__7_));
MUX2X1 MUX2X1_877 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3868_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2130_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3852_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__8_));
MUX2X1 MUX2X1_878 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3870_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2133_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3852_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__9_));
MUX2X1 MUX2X1_879 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3872_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2136_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3852_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__10_));
MUX2X1 MUX2X1_88 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2162_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2163_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2106_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__19_));
MUX2X1 MUX2X1_880 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3874_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2139_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3852_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__11_));
MUX2X1 MUX2X1_881 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3876_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2142_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3852_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__12_));
MUX2X1 MUX2X1_882 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3878_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2145_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3852_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__13_));
MUX2X1 MUX2X1_883 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3880_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2148_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3852_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__14_));
MUX2X1 MUX2X1_884 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3882_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2151_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3852_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__15_));
MUX2X1 MUX2X1_885 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3884_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2154_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3852_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__16_));
MUX2X1 MUX2X1_886 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3886_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2157_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3852_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__17_));
MUX2X1 MUX2X1_887 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3888_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2160_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3852_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__18_));
MUX2X1 MUX2X1_888 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3890_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2163_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3852_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__19_));
MUX2X1 MUX2X1_889 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3892_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2166_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3852_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__20_));
MUX2X1 MUX2X1_89 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2165_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2166_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2106_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__20_));
MUX2X1 MUX2X1_890 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3894_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2169_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3852_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__21_));
MUX2X1 MUX2X1_891 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3896_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2172_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3852_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__22_));
MUX2X1 MUX2X1_892 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3898_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2175_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3852_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__23_));
MUX2X1 MUX2X1_893 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3900_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2178_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3852_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__24_));
MUX2X1 MUX2X1_894 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3902_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2181_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3852_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__25_));
MUX2X1 MUX2X1_895 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3904_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2184_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3852_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__26_));
MUX2X1 MUX2X1_896 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3906_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2187_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3852_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__27_));
MUX2X1 MUX2X1_897 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3908_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2190_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3852_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__28_));
MUX2X1 MUX2X1_898 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3910_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2193_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3852_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__29_));
MUX2X1 MUX2X1_899 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3912_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2196_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3852_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__30_));
MUX2X1 MUX2X1_9 ( .A(epc_q_8_), .B(REGFILE_SIM_reg_bank_reg_rb_o_8_), .S(_abc_40298_new_n1187_), .Y(_abc_40298_new_n1367_));
MUX2X1 MUX2X1_90 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2168_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2169_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2106_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__21_));
MUX2X1 MUX2X1_900 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3914_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2199_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3852_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__31_));
MUX2X1 MUX2X1_901 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3916_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2100_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3917_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__0_));
MUX2X1 MUX2X1_902 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3919_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2109_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3917_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__1_));
MUX2X1 MUX2X1_903 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3921_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2112_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3917_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__2_));
MUX2X1 MUX2X1_904 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3923_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2115_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3917_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__3_));
MUX2X1 MUX2X1_905 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3925_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2118_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3917_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__4_));
MUX2X1 MUX2X1_906 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3927_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2121_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3917_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__5_));
MUX2X1 MUX2X1_907 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3929_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2124_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3917_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__6_));
MUX2X1 MUX2X1_908 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3931_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2127_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3917_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__7_));
MUX2X1 MUX2X1_909 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3933_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2130_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3917_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__8_));
MUX2X1 MUX2X1_91 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2171_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2172_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2106_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__22_));
MUX2X1 MUX2X1_910 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3935_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2133_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3917_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__9_));
MUX2X1 MUX2X1_911 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3937_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2136_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3917_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__10_));
MUX2X1 MUX2X1_912 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3939_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2139_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3917_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__11_));
MUX2X1 MUX2X1_913 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3941_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2142_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3917_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__12_));
MUX2X1 MUX2X1_914 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3943_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2145_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3917_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__13_));
MUX2X1 MUX2X1_915 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3945_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2148_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3917_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__14_));
MUX2X1 MUX2X1_916 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3947_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2151_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3917_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__15_));
MUX2X1 MUX2X1_917 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3949_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2154_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3917_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__16_));
MUX2X1 MUX2X1_918 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3951_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2157_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3917_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__17_));
MUX2X1 MUX2X1_919 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3953_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2160_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3917_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__18_));
MUX2X1 MUX2X1_92 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2174_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2175_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2106_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__23_));
MUX2X1 MUX2X1_920 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3955_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2163_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3917_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__19_));
MUX2X1 MUX2X1_921 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3957_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2166_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3917_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__20_));
MUX2X1 MUX2X1_922 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3959_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2169_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3917_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__21_));
MUX2X1 MUX2X1_923 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3961_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2172_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3917_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__22_));
MUX2X1 MUX2X1_924 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3963_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2175_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3917_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__23_));
MUX2X1 MUX2X1_925 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3965_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2178_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3917_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__24_));
MUX2X1 MUX2X1_926 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3967_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2181_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3917_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__25_));
MUX2X1 MUX2X1_927 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3969_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2184_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3917_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__26_));
MUX2X1 MUX2X1_928 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3971_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2187_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3917_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__27_));
MUX2X1 MUX2X1_929 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3973_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2190_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3917_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__28_));
MUX2X1 MUX2X1_93 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2177_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2178_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2106_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__24_));
MUX2X1 MUX2X1_930 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3975_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2193_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3917_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__29_));
MUX2X1 MUX2X1_931 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3977_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2196_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3917_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__30_));
MUX2X1 MUX2X1_932 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3979_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2199_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3917_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__31_));
MUX2X1 MUX2X1_933 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2100_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3981_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3982_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__0_));
MUX2X1 MUX2X1_934 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2109_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3984_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3982_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__1_));
MUX2X1 MUX2X1_935 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2112_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3986_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3982_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__2_));
MUX2X1 MUX2X1_936 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2115_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3988_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3982_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__3_));
MUX2X1 MUX2X1_937 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2118_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3990_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3982_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__4_));
MUX2X1 MUX2X1_938 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2121_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3992_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3982_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__5_));
MUX2X1 MUX2X1_939 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2124_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3994_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3982_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__6_));
MUX2X1 MUX2X1_94 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2180_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2181_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2106_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__25_));
MUX2X1 MUX2X1_940 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2127_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3996_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3982_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__7_));
MUX2X1 MUX2X1_941 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2130_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3998_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3982_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__8_));
MUX2X1 MUX2X1_942 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2133_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4000_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3982_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__9_));
MUX2X1 MUX2X1_943 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2136_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4002_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3982_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__10_));
MUX2X1 MUX2X1_944 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2139_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4004_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3982_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__11_));
MUX2X1 MUX2X1_945 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2142_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4006_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3982_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__12_));
MUX2X1 MUX2X1_946 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2145_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4008_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3982_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__13_));
MUX2X1 MUX2X1_947 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2148_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4010_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3982_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__14_));
MUX2X1 MUX2X1_948 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2151_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4012_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3982_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__15_));
MUX2X1 MUX2X1_949 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2154_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4014_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3982_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__16_));
MUX2X1 MUX2X1_95 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2183_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2184_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2106_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__26_));
MUX2X1 MUX2X1_950 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2157_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4016_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3982_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__17_));
MUX2X1 MUX2X1_951 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2160_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4018_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3982_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__18_));
MUX2X1 MUX2X1_952 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2163_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4020_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3982_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__19_));
MUX2X1 MUX2X1_953 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2166_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4022_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3982_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__20_));
MUX2X1 MUX2X1_954 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2169_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4024_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3982_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__21_));
MUX2X1 MUX2X1_955 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2172_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4026_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3982_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__22_));
MUX2X1 MUX2X1_956 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2175_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4028_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3982_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__23_));
MUX2X1 MUX2X1_957 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2178_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4030_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3982_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__24_));
MUX2X1 MUX2X1_958 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2181_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4032_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3982_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__25_));
MUX2X1 MUX2X1_959 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2184_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4034_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3982_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__26_));
MUX2X1 MUX2X1_96 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2186_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2187_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2106_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__27_));
MUX2X1 MUX2X1_960 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2187_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4036_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3982_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__27_));
MUX2X1 MUX2X1_961 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2190_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4038_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3982_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__28_));
MUX2X1 MUX2X1_962 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2193_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4040_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3982_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__29_));
MUX2X1 MUX2X1_963 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2196_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4042_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3982_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__30_));
MUX2X1 MUX2X1_964 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2199_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4044_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n3982_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__31_));
MUX2X1 MUX2X1_965 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4046_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2100_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4047_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__0_));
MUX2X1 MUX2X1_966 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4049_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2109_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4047_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__1_));
MUX2X1 MUX2X1_967 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4051_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2112_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4047_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__2_));
MUX2X1 MUX2X1_968 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4053_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2115_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4047_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__3_));
MUX2X1 MUX2X1_969 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4055_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2118_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4047_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__4_));
MUX2X1 MUX2X1_97 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2189_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2190_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2106_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__28_));
MUX2X1 MUX2X1_970 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4057_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2121_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4047_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__5_));
MUX2X1 MUX2X1_971 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4059_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2124_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4047_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__6_));
MUX2X1 MUX2X1_972 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4061_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2127_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4047_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__7_));
MUX2X1 MUX2X1_973 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4063_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2130_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4047_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__8_));
MUX2X1 MUX2X1_974 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4065_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2133_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4047_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__9_));
MUX2X1 MUX2X1_975 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4067_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2136_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4047_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__10_));
MUX2X1 MUX2X1_976 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4069_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2139_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4047_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__11_));
MUX2X1 MUX2X1_977 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4071_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2142_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4047_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__12_));
MUX2X1 MUX2X1_978 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4073_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2145_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4047_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__13_));
MUX2X1 MUX2X1_979 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4075_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2148_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4047_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__14_));
MUX2X1 MUX2X1_98 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2192_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2193_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2106_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__29_));
MUX2X1 MUX2X1_980 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4077_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2151_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4047_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__15_));
MUX2X1 MUX2X1_981 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4079_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2154_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4047_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__16_));
MUX2X1 MUX2X1_982 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4081_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2157_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4047_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__17_));
MUX2X1 MUX2X1_983 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4083_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2160_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4047_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__18_));
MUX2X1 MUX2X1_984 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4085_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2163_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4047_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__19_));
MUX2X1 MUX2X1_985 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4087_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2166_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4047_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__20_));
MUX2X1 MUX2X1_986 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4089_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2169_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4047_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__21_));
MUX2X1 MUX2X1_987 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4091_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2172_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4047_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__22_));
MUX2X1 MUX2X1_988 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4093_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2175_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4047_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__23_));
MUX2X1 MUX2X1_989 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4095_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2178_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4047_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__24_));
MUX2X1 MUX2X1_99 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2195_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2196_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n2106_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__30_));
MUX2X1 MUX2X1_990 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4097_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2181_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4047_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__25_));
MUX2X1 MUX2X1_991 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4099_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2184_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4047_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__26_));
MUX2X1 MUX2X1_992 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4101_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2187_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4047_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__27_));
MUX2X1 MUX2X1_993 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4103_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2190_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4047_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__28_));
MUX2X1 MUX2X1_994 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4105_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2193_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4047_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__29_));
MUX2X1 MUX2X1_995 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4107_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2196_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4047_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__30_));
MUX2X1 MUX2X1_996 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4109_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2199_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4047_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__31_));
MUX2X1 MUX2X1_997 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2100_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4111_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4112_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__0_));
MUX2X1 MUX2X1_998 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2109_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4114_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4112_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__1_));
MUX2X1 MUX2X1_999 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2112_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4116_), .S(REGFILE_SIM_reg_bank__abc_34451_new_n4112_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__2_));
NAND2X1 NAND2X1_1 ( .A(_abc_40298_new_n624_), .B(_abc_40298_new_n625_), .Y(_abc_40298_new_n626_));
NAND2X1 NAND2X1_10 ( .A(\mem_dat_i[0] ), .B(_abc_40298_new_n679_), .Y(_abc_40298_new_n680_));
NAND2X1 NAND2X1_100 ( .A(_abc_40298_new_n1375_), .B(_abc_40298_new_n1403_), .Y(_abc_40298_new_n1425_));
NAND2X1 NAND2X1_101 ( .A(alu_op_r_6_), .B(pc_q_10_), .Y(_abc_40298_new_n1428_));
NAND2X1 NAND2X1_102 ( .A(_abc_40298_new_n1213_), .B(_abc_40298_new_n1439_), .Y(_abc_40298_new_n1440_));
NAND2X1 NAND2X1_103 ( .A(_abc_40298_new_n1457_), .B(_abc_40298_new_n1447_), .Y(_abc_40298_new_n1458_));
NAND2X1 NAND2X1_104 ( .A(alu_op_r_7_), .B(pc_q_11_), .Y(_abc_40298_new_n1459_));
NAND2X1 NAND2X1_105 ( .A(_abc_40298_new_n1459_), .B(_abc_40298_new_n1458_), .Y(_abc_40298_new_n1460_));
NAND2X1 NAND2X1_106 ( .A(_abc_40298_new_n1480_), .B(_abc_40298_new_n1426_), .Y(_abc_40298_new_n1481_));
NAND2X1 NAND2X1_107 ( .A(_abc_40298_new_n1483_), .B(_abc_40298_new_n1481_), .Y(_abc_40298_new_n1484_));
NAND2X1 NAND2X1_108 ( .A(int32_r_10_), .B(pc_q_12_), .Y(_abc_40298_new_n1491_));
NAND2X1 NAND2X1_109 ( .A(_abc_40298_new_n1175_), .B(_abc_40298_new_n1498_), .Y(_abc_40298_new_n1499_));
NAND2X1 NAND2X1_11 ( .A(_abc_40298_new_n644_), .B(_abc_40298_new_n684_), .Y(_abc_40298_new_n685_));
NAND2X1 NAND2X1_110 ( .A(_abc_40298_new_n1509_), .B(_abc_40298_new_n1232_), .Y(_abc_40298_new_n1525_));
NAND2X1 NAND2X1_111 ( .A(_abc_40298_new_n1533_), .B(_abc_40298_new_n1535_), .Y(_abc_40298_new_n1536_));
NAND2X1 NAND2X1_112 ( .A(epc_q_14_), .B(_abc_40298_new_n1065_), .Y(_abc_40298_new_n1539_));
NAND2X1 NAND2X1_113 ( .A(pc_q_13_), .B(REGFILE_SIM_reg_bank_rb_i_0_), .Y(_abc_40298_new_n1541_));
NAND2X1 NAND2X1_114 ( .A(pc_q_14_), .B(REGFILE_SIM_reg_bank_rb_i_1_), .Y(_abc_40298_new_n1544_));
NAND2X1 NAND2X1_115 ( .A(_abc_40298_new_n1175_), .B(_abc_40298_new_n1552_), .Y(_abc_40298_new_n1553_));
NAND2X1 NAND2X1_116 ( .A(pc_q_15_), .B(REGFILE_SIM_reg_bank_rb_i_2_), .Y(_abc_40298_new_n1571_));
NAND2X1 NAND2X1_117 ( .A(_abc_40298_new_n1175_), .B(_abc_40298_new_n1578_), .Y(_abc_40298_new_n1579_));
NAND2X1 NAND2X1_118 ( .A(_abc_40298_new_n1546_), .B(_abc_40298_new_n1573_), .Y(_abc_40298_new_n1596_));
NAND2X1 NAND2X1_119 ( .A(_abc_40298_new_n1594_), .B(_abc_40298_new_n1486_), .Y(_abc_40298_new_n1600_));
NAND2X1 NAND2X1_12 ( .A(alu_p_o_1_), .B(_abc_40298_new_n631_), .Y(_abc_40298_new_n693_));
NAND2X1 NAND2X1_120 ( .A(epc_q_17_), .B(_abc_40298_new_n1065_), .Y(_abc_40298_new_n1626_));
NAND2X1 NAND2X1_121 ( .A(_abc_40298_new_n1175_), .B(_abc_40298_new_n1635_), .Y(_abc_40298_new_n1636_));
NAND2X1 NAND2X1_122 ( .A(_abc_40298_new_n1645_), .B(_abc_40298_new_n1647_), .Y(_abc_40298_new_n1648_));
NAND2X1 NAND2X1_123 ( .A(epc_q_18_), .B(_abc_40298_new_n1065_), .Y(_abc_40298_new_n1651_));
NAND2X1 NAND2X1_124 ( .A(_abc_40298_new_n1175_), .B(_abc_40298_new_n1665_), .Y(_abc_40298_new_n1666_));
NAND2X1 NAND2X1_125 ( .A(epc_q_19_), .B(_abc_40298_new_n1065_), .Y(_abc_40298_new_n1680_));
NAND2X1 NAND2X1_126 ( .A(_abc_40298_new_n1175_), .B(_abc_40298_new_n1688_), .Y(_abc_40298_new_n1689_));
NAND2X1 NAND2X1_127 ( .A(_abc_40298_new_n1699_), .B(_abc_40298_new_n1698_), .Y(_abc_40298_new_n1700_));
NAND2X1 NAND2X1_128 ( .A(epc_q_20_), .B(_abc_40298_new_n1065_), .Y(_abc_40298_new_n1703_));
NAND2X1 NAND2X1_129 ( .A(_abc_40298_new_n1660_), .B(_abc_40298_new_n1685_), .Y(_abc_40298_new_n1704_));
NAND2X1 NAND2X1_13 ( .A(\mem_dat_i[17] ), .B(_abc_40298_new_n688_), .Y(_abc_40298_new_n696_));
NAND2X1 NAND2X1_130 ( .A(_abc_40298_new_n1175_), .B(_abc_40298_new_n1717_), .Y(_abc_40298_new_n1718_));
NAND2X1 NAND2X1_131 ( .A(_abc_40298_new_n1726_), .B(_abc_40298_new_n1699_), .Y(_abc_40298_new_n1727_));
NAND2X1 NAND2X1_132 ( .A(epc_q_21_), .B(_abc_40298_new_n1065_), .Y(_abc_40298_new_n1732_));
NAND2X1 NAND2X1_133 ( .A(_abc_40298_new_n1714_), .B(_abc_40298_new_n1740_), .Y(_abc_40298_new_n1741_));
NAND2X1 NAND2X1_134 ( .A(_abc_40298_new_n1175_), .B(_abc_40298_new_n1744_), .Y(_abc_40298_new_n1745_));
NAND2X1 NAND2X1_135 ( .A(_abc_40298_new_n1754_), .B(_abc_40298_new_n1756_), .Y(_abc_40298_new_n1757_));
NAND2X1 NAND2X1_136 ( .A(epc_q_22_), .B(_abc_40298_new_n1065_), .Y(_abc_40298_new_n1760_));
NAND2X1 NAND2X1_137 ( .A(_abc_40298_new_n1713_), .B(_abc_40298_new_n1740_), .Y(_abc_40298_new_n1762_));
NAND2X1 NAND2X1_138 ( .A(_abc_40298_new_n1175_), .B(_abc_40298_new_n1773_), .Y(_abc_40298_new_n1774_));
NAND2X1 NAND2X1_139 ( .A(epc_q_23_), .B(_abc_40298_new_n1065_), .Y(_abc_40298_new_n1788_));
NAND2X1 NAND2X1_14 ( .A(\mem_dat_i[25] ), .B(_abc_40298_new_n674_), .Y(_abc_40298_new_n698_));
NAND2X1 NAND2X1_140 ( .A(_abc_40298_new_n1175_), .B(_abc_40298_new_n1796_), .Y(_abc_40298_new_n1797_));
NAND2X1 NAND2X1_141 ( .A(_abc_40298_new_n1807_), .B(_abc_40298_new_n1806_), .Y(_abc_40298_new_n1808_));
NAND2X1 NAND2X1_142 ( .A(_abc_40298_new_n1768_), .B(_abc_40298_new_n1792_), .Y(_abc_40298_new_n1812_));
NAND2X1 NAND2X1_143 ( .A(_abc_40298_new_n1817_), .B(_abc_40298_new_n1820_), .Y(_abc_40298_new_n1821_));
NAND2X1 NAND2X1_144 ( .A(epc_q_24_), .B(_abc_40298_new_n1065_), .Y(_abc_40298_new_n1829_));
NAND2X1 NAND2X1_145 ( .A(_abc_40298_new_n1175_), .B(_abc_40298_new_n1830_), .Y(_abc_40298_new_n1831_));
NAND2X1 NAND2X1_146 ( .A(_abc_40298_new_n1232_), .B(_abc_40298_new_n1808_), .Y(_abc_40298_new_n1833_));
NAND2X1 NAND2X1_147 ( .A(_abc_40298_new_n1858_), .B(_abc_40298_new_n1856_), .Y(_abc_40298_new_n1859_));
NAND2X1 NAND2X1_148 ( .A(_abc_40298_new_n1887_), .B(_abc_40298_new_n1885_), .Y(_abc_40298_new_n1888_));
NAND2X1 NAND2X1_149 ( .A(epc_q_27_), .B(_abc_40298_new_n1065_), .Y(_abc_40298_new_n1901_));
NAND2X1 NAND2X1_15 ( .A(alu_p_o_2_), .B(_abc_40298_new_n631_), .Y(_abc_40298_new_n706_));
NAND2X1 NAND2X1_150 ( .A(_abc_40298_new_n1232_), .B(_abc_40298_new_n1892_), .Y(_abc_40298_new_n1904_));
NAND2X1 NAND2X1_151 ( .A(_abc_40298_new_n1232_), .B(_abc_40298_new_n1914_), .Y(_abc_40298_new_n1934_));
NAND2X1 NAND2X1_152 ( .A(_abc_40298_new_n1232_), .B(_abc_40298_new_n1941_), .Y(_abc_40298_new_n1953_));
NAND2X1 NAND2X1_153 ( .A(_abc_40298_new_n1953_), .B(_abc_40298_new_n1952_), .Y(_abc_40298_new_n1954_));
NAND2X1 NAND2X1_154 ( .A(pc_q_30_), .B(_abc_40298_new_n1963_), .Y(_abc_40298_new_n1964_));
NAND2X1 NAND2X1_155 ( .A(_abc_40298_new_n1970_), .B(_abc_40298_new_n1969_), .Y(_abc_40298_new_n1971_));
NAND2X1 NAND2X1_156 ( .A(_abc_40298_new_n1213_), .B(_abc_40298_new_n1980_), .Y(_abc_40298_new_n1981_));
NAND2X1 NAND2X1_157 ( .A(_abc_40298_new_n1982_), .B(_abc_40298_new_n1981_), .Y(_abc_40298_new_n1983_));
NAND2X1 NAND2X1_158 ( .A(_abc_40298_new_n2008_), .B(_abc_40298_new_n2006_), .Y(_abc_40298_new_n2009_));
NAND2X1 NAND2X1_159 ( .A(_abc_40298_new_n1179_), .B(_abc_40298_new_n2014_), .Y(_abc_40298_new_n2015_));
NAND2X1 NAND2X1_16 ( .A(\mem_dat_i[18] ), .B(_abc_40298_new_n688_), .Y(_abc_40298_new_n708_));
NAND2X1 NAND2X1_160 ( .A(_abc_40298_new_n1198_), .B(_abc_40298_new_n2014_), .Y(_abc_40298_new_n2018_));
NAND2X1 NAND2X1_161 ( .A(_abc_40298_new_n1222_), .B(_abc_40298_new_n2014_), .Y(_abc_40298_new_n2021_));
NAND2X1 NAND2X1_162 ( .A(_abc_40298_new_n1271_), .B(_abc_40298_new_n2014_), .Y(_abc_40298_new_n2028_));
NAND2X1 NAND2X1_163 ( .A(_abc_40298_new_n1325_), .B(_abc_40298_new_n2014_), .Y(_abc_40298_new_n2034_));
NAND2X1 NAND2X1_164 ( .A(REGFILE_SIM_reg_bank_wr_i), .B(_abc_40298_new_n2050_), .Y(_abc_40298_new_n2051_));
NAND2X1 NAND2X1_165 ( .A(_abc_40298_new_n1025_), .B(_abc_40298_new_n2054_), .Y(_abc_40298_new_n2055_));
NAND2X1 NAND2X1_166 ( .A(_abc_40298_new_n2014_), .B(_abc_40298_new_n1526_), .Y(_abc_40298_new_n2061_));
NAND2X1 NAND2X1_167 ( .A(_abc_40298_new_n2014_), .B(_abc_40298_new_n1555_), .Y(_abc_40298_new_n2064_));
NAND2X1 NAND2X1_168 ( .A(_abc_40298_new_n2014_), .B(_abc_40298_new_n1581_), .Y(_abc_40298_new_n2067_));
NAND2X1 NAND2X1_169 ( .A(_abc_40298_new_n2014_), .B(_abc_40298_new_n1638_), .Y(_abc_40298_new_n2073_));
NAND2X1 NAND2X1_17 ( .A(\mem_dat_i[26] ), .B(_abc_40298_new_n674_), .Y(_abc_40298_new_n710_));
NAND2X1 NAND2X1_170 ( .A(_abc_40298_new_n2014_), .B(_abc_40298_new_n1668_), .Y(_abc_40298_new_n2076_));
NAND2X1 NAND2X1_171 ( .A(_abc_40298_new_n2014_), .B(_abc_40298_new_n1691_), .Y(_abc_40298_new_n2079_));
NAND2X1 NAND2X1_172 ( .A(_abc_40298_new_n2014_), .B(_abc_40298_new_n1720_), .Y(_abc_40298_new_n2082_));
NAND2X1 NAND2X1_173 ( .A(_abc_40298_new_n2014_), .B(_abc_40298_new_n1747_), .Y(_abc_40298_new_n2085_));
NAND2X1 NAND2X1_174 ( .A(_abc_40298_new_n2014_), .B(_abc_40298_new_n1776_), .Y(_abc_40298_new_n2088_));
NAND2X1 NAND2X1_175 ( .A(_abc_40298_new_n2014_), .B(_abc_40298_new_n1799_), .Y(_abc_40298_new_n2091_));
NAND2X1 NAND2X1_176 ( .A(_abc_40298_new_n2014_), .B(_abc_40298_new_n1905_), .Y(_abc_40298_new_n2103_));
NAND2X1 NAND2X1_177 ( .A(_abc_40298_new_n2014_), .B(_abc_40298_new_n1935_), .Y(_abc_40298_new_n2106_));
NAND2X1 NAND2X1_178 ( .A(_abc_40298_new_n2014_), .B(_abc_40298_new_n1954_), .Y(_abc_40298_new_n2109_));
NAND2X1 NAND2X1_179 ( .A(_abc_40298_new_n2014_), .B(_abc_40298_new_n1983_), .Y(_abc_40298_new_n2112_));
NAND2X1 NAND2X1_18 ( .A(alu_p_o_3_), .B(_abc_40298_new_n631_), .Y(_abc_40298_new_n717_));
NAND2X1 NAND2X1_180 ( .A(_abc_40298_new_n1998_), .B(_abc_40298_new_n2005_), .Y(_abc_40298_new_n2115_));
NAND2X1 NAND2X1_181 ( .A(_abc_40298_new_n2014_), .B(_abc_40298_new_n2115_), .Y(_abc_40298_new_n2116_));
NAND2X1 NAND2X1_182 ( .A(_abc_40298_new_n904_), .B(_abc_40298_new_n912_), .Y(_abc_40298_new_n2122_));
NAND2X1 NAND2X1_183 ( .A(alu_op_r_7_), .B(_abc_40298_new_n889_), .Y(_abc_40298_new_n2124_));
NAND2X1 NAND2X1_184 ( .A(opcode_q_22_), .B(_abc_40298_new_n1013_), .Y(_abc_40298_new_n2132_));
NAND2X1 NAND2X1_185 ( .A(opcode_q_23_), .B(_abc_40298_new_n1013_), .Y(_abc_40298_new_n2134_));
NAND2X1 NAND2X1_186 ( .A(opcode_q_25_), .B(_abc_40298_new_n1013_), .Y(_abc_40298_new_n2137_));
NAND2X1 NAND2X1_187 ( .A(_abc_40298_new_n2148_), .B(_abc_40298_new_n927_), .Y(_abc_40298_new_n2149_));
NAND2X1 NAND2X1_188 ( .A(_abc_40298_new_n893_), .B(_abc_40298_new_n899_), .Y(_abc_40298_new_n2162_));
NAND2X1 NAND2X1_189 ( .A(_abc_40298_new_n893_), .B(_abc_40298_new_n901_), .Y(_abc_40298_new_n2164_));
NAND2X1 NAND2X1_19 ( .A(\mem_dat_i[19] ), .B(_abc_40298_new_n688_), .Y(_abc_40298_new_n719_));
NAND2X1 NAND2X1_190 ( .A(_abc_40298_new_n897_), .B(_abc_40298_new_n2169_), .Y(_abc_40298_new_n2170_));
NAND2X1 NAND2X1_191 ( .A(_abc_40298_new_n892_), .B(_abc_40298_new_n926_), .Y(_abc_40298_new_n2174_));
NAND2X1 NAND2X1_192 ( .A(_abc_40298_new_n1628_), .B(_abc_40298_new_n930_), .Y(_abc_40298_new_n2204_));
NAND2X1 NAND2X1_193 ( .A(_abc_40298_new_n2143_), .B(_abc_40298_new_n2285_), .Y(_abc_40298_new_n2286_));
NAND2X1 NAND2X1_194 ( .A(_abc_40298_new_n2309_), .B(_abc_40298_new_n2308_), .Y(_abc_40298_new_n2310_));
NAND2X1 NAND2X1_195 ( .A(_abc_40298_new_n2316_), .B(_abc_40298_new_n2315_), .Y(_abc_40298_new_n2317_));
NAND2X1 NAND2X1_196 ( .A(_abc_40298_new_n2329_), .B(_abc_40298_new_n2328_), .Y(_abc_40298_new_n2330_));
NAND2X1 NAND2X1_197 ( .A(_abc_40298_new_n2337_), .B(_abc_40298_new_n2336_), .Y(_abc_40298_new_n2338_));
NAND2X1 NAND2X1_198 ( .A(_abc_40298_new_n2344_), .B(_abc_40298_new_n2343_), .Y(_abc_40298_new_n2345_));
NAND2X1 NAND2X1_199 ( .A(_abc_40298_new_n1012_), .B(_abc_40298_new_n1391_), .Y(_abc_40298_new_n2355_));
NAND2X1 NAND2X1_2 ( .A(_abc_40298_new_n627_), .B(_abc_40298_new_n622_), .Y(_abc_40298_new_n628_));
NAND2X1 NAND2X1_20 ( .A(\mem_dat_i[27] ), .B(_abc_40298_new_n674_), .Y(_abc_40298_new_n721_));
NAND2X1 NAND2X1_200 ( .A(epc_q_16_), .B(_abc_40298_new_n1001_), .Y(_abc_40298_new_n2388_));
NAND2X1 NAND2X1_201 ( .A(epc_q_17_), .B(_abc_40298_new_n1001_), .Y(_abc_40298_new_n2395_));
NAND2X1 NAND2X1_202 ( .A(epc_q_18_), .B(_abc_40298_new_n1001_), .Y(_abc_40298_new_n2402_));
NAND2X1 NAND2X1_203 ( .A(epc_q_19_), .B(_abc_40298_new_n1001_), .Y(_abc_40298_new_n2409_));
NAND2X1 NAND2X1_204 ( .A(epc_q_20_), .B(_abc_40298_new_n1001_), .Y(_abc_40298_new_n2416_));
NAND2X1 NAND2X1_205 ( .A(epc_q_21_), .B(_abc_40298_new_n1001_), .Y(_abc_40298_new_n2423_));
NAND2X1 NAND2X1_206 ( .A(epc_q_22_), .B(_abc_40298_new_n1001_), .Y(_abc_40298_new_n2430_));
NAND2X1 NAND2X1_207 ( .A(epc_q_23_), .B(_abc_40298_new_n1001_), .Y(_abc_40298_new_n2437_));
NAND2X1 NAND2X1_208 ( .A(epc_q_24_), .B(_abc_40298_new_n1001_), .Y(_abc_40298_new_n2444_));
NAND2X1 NAND2X1_209 ( .A(epc_q_25_), .B(_abc_40298_new_n1001_), .Y(_abc_40298_new_n2451_));
NAND2X1 NAND2X1_21 ( .A(\mem_dat_i[20] ), .B(_abc_40298_new_n677_), .Y(_abc_40298_new_n730_));
NAND2X1 NAND2X1_210 ( .A(epc_q_26_), .B(_abc_40298_new_n1001_), .Y(_abc_40298_new_n2459_));
NAND2X1 NAND2X1_211 ( .A(epc_q_27_), .B(_abc_40298_new_n1001_), .Y(_abc_40298_new_n2466_));
NAND2X1 NAND2X1_212 ( .A(epc_q_28_), .B(_abc_40298_new_n1001_), .Y(_abc_40298_new_n2474_));
NAND2X1 NAND2X1_213 ( .A(epc_q_29_), .B(_abc_40298_new_n1001_), .Y(_abc_40298_new_n2482_));
NAND2X1 NAND2X1_214 ( .A(epc_q_30_), .B(_abc_40298_new_n1001_), .Y(_abc_40298_new_n2489_));
NAND2X1 NAND2X1_215 ( .A(epc_q_31_), .B(_abc_40298_new_n1001_), .Y(_abc_40298_new_n2496_));
NAND2X1 NAND2X1_216 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_0_), .B(alu_op_r_0_), .Y(_abc_40298_new_n2513_));
NAND2X1 NAND2X1_217 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_1_), .B(alu_op_r_1_), .Y(_abc_40298_new_n2518_));
NAND2X1 NAND2X1_218 ( .A(inst_r_0_), .B(_abc_40298_new_n641_), .Y(_abc_40298_new_n2569_));
NAND2X1 NAND2X1_219 ( .A(_abc_40298_new_n2515_), .B(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2579_));
NAND2X1 NAND2X1_22 ( .A(\mem_dat_i[4] ), .B(_abc_40298_new_n679_), .Y(_abc_40298_new_n731_));
NAND2X1 NAND2X1_220 ( .A(_abc_40298_new_n2680_), .B(_abc_40298_new_n2576_), .Y(_abc_40298_new_n2681_));
NAND2X1 NAND2X1_221 ( .A(_abc_40298_new_n2689_), .B(_abc_40298_new_n2576_), .Y(_abc_40298_new_n2690_));
NAND2X1 NAND2X1_222 ( .A(_abc_40298_new_n2698_), .B(_abc_40298_new_n2576_), .Y(_abc_40298_new_n2699_));
NAND2X1 NAND2X1_223 ( .A(_abc_40298_new_n2707_), .B(_abc_40298_new_n2576_), .Y(_abc_40298_new_n2708_));
NAND2X1 NAND2X1_224 ( .A(_abc_40298_new_n2716_), .B(_abc_40298_new_n2576_), .Y(_abc_40298_new_n2717_));
NAND2X1 NAND2X1_225 ( .A(_abc_40298_new_n2725_), .B(_abc_40298_new_n2576_), .Y(_abc_40298_new_n2726_));
NAND2X1 NAND2X1_226 ( .A(_abc_40298_new_n2734_), .B(_abc_40298_new_n2576_), .Y(_abc_40298_new_n2735_));
NAND2X1 NAND2X1_227 ( .A(_abc_40298_new_n2743_), .B(_abc_40298_new_n2576_), .Y(_abc_40298_new_n2744_));
NAND2X1 NAND2X1_228 ( .A(_abc_40298_new_n2816_), .B(_abc_40298_new_n2576_), .Y(_abc_40298_new_n2817_));
NAND2X1 NAND2X1_229 ( .A(_abc_40298_new_n2825_), .B(_abc_40298_new_n2576_), .Y(_abc_40298_new_n2826_));
NAND2X1 NAND2X1_23 ( .A(\mem_dat_i[21] ), .B(_abc_40298_new_n677_), .Y(_abc_40298_new_n739_));
NAND2X1 NAND2X1_230 ( .A(_abc_40298_new_n2834_), .B(_abc_40298_new_n2576_), .Y(_abc_40298_new_n2835_));
NAND2X1 NAND2X1_231 ( .A(_abc_40298_new_n2843_), .B(_abc_40298_new_n2576_), .Y(_abc_40298_new_n2844_));
NAND2X1 NAND2X1_232 ( .A(_abc_40298_new_n2852_), .B(_abc_40298_new_n2576_), .Y(_abc_40298_new_n2853_));
NAND2X1 NAND2X1_233 ( .A(_abc_40298_new_n2861_), .B(_abc_40298_new_n2576_), .Y(_abc_40298_new_n2862_));
NAND2X1 NAND2X1_234 ( .A(_abc_40298_new_n2870_), .B(_abc_40298_new_n2576_), .Y(_abc_40298_new_n2871_));
NAND2X1 NAND2X1_235 ( .A(_abc_40298_new_n2879_), .B(_abc_40298_new_n2576_), .Y(_abc_40298_new_n2880_));
NAND2X1 NAND2X1_236 ( .A(_abc_40298_new_n2889_), .B(_abc_40298_new_n2888_), .Y(_0mem_stb_o_0_0_));
NAND2X1 NAND2X1_237 ( .A(_abc_40298_new_n2893_), .B(_abc_40298_new_n2888_), .Y(_0mem_cyc_o_0_0_));
NAND2X1 NAND2X1_238 ( .A(\mem_addr_o[0] ), .B(_abc_40298_new_n2895_), .Y(_abc_40298_new_n2896_));
NAND2X1 NAND2X1_239 ( .A(\mem_addr_o[1] ), .B(_abc_40298_new_n2895_), .Y(_abc_40298_new_n2898_));
NAND2X1 NAND2X1_24 ( .A(\mem_dat_i[5] ), .B(_abc_40298_new_n679_), .Y(_abc_40298_new_n740_));
NAND2X1 NAND2X1_240 ( .A(\mem_addr_o[2] ), .B(_abc_40298_new_n2895_), .Y(_abc_40298_new_n2900_));
NAND2X1 NAND2X1_241 ( .A(state_q_3_), .B(pc_q_2_), .Y(_abc_40298_new_n2901_));
NAND2X1 NAND2X1_242 ( .A(_abc_40298_new_n2921_), .B(_abc_40298_new_n2923_), .Y(_abc_40298_new_n2927_));
NAND2X1 NAND2X1_243 ( .A(_abc_40298_new_n2944_), .B(_abc_40298_new_n2942_), .Y(_abc_40298_new_n2945_));
NAND2X1 NAND2X1_244 ( .A(state_q_3_), .B(pc_q_7_), .Y(_abc_40298_new_n2955_));
NAND2X1 NAND2X1_245 ( .A(\mem_addr_o[7] ), .B(_abc_40298_new_n2895_), .Y(_abc_40298_new_n2956_));
NAND2X1 NAND2X1_246 ( .A(_abc_40298_new_n2943_), .B(_abc_40298_new_n2949_), .Y(_abc_40298_new_n2958_));
NAND2X1 NAND2X1_247 ( .A(_abc_40298_new_n2962_), .B(_abc_40298_new_n2960_), .Y(_abc_40298_new_n2964_));
NAND2X1 NAND2X1_248 ( .A(_abc_40298_new_n2902_), .B(_abc_40298_new_n2964_), .Y(_abc_40298_new_n2965_));
NAND2X1 NAND2X1_249 ( .A(_abc_40298_new_n2977_), .B(_abc_40298_new_n2979_), .Y(_abc_40298_new_n2980_));
NAND2X1 NAND2X1_25 ( .A(alu_p_o_6_), .B(_abc_40298_new_n631_), .Y(_abc_40298_new_n746_));
NAND2X1 NAND2X1_250 ( .A(_abc_40298_new_n2962_), .B(_abc_40298_new_n2970_), .Y(_abc_40298_new_n2994_));
NAND2X1 NAND2X1_251 ( .A(_abc_40298_new_n2977_), .B(_abc_40298_new_n2989_), .Y(_abc_40298_new_n2995_));
NAND2X1 NAND2X1_252 ( .A(_abc_40298_new_n3004_), .B(_abc_40298_new_n3001_), .Y(_abc_40298_new_n3005_));
NAND2X1 NAND2X1_253 ( .A(_abc_40298_new_n3005_), .B(_abc_40298_new_n3006_), .Y(_abc_40298_new_n3007_));
NAND2X1 NAND2X1_254 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_12_), .B(_abc_40298_new_n3003_), .Y(_abc_40298_new_n3010_));
NAND2X1 NAND2X1_255 ( .A(_abc_40298_new_n1039_), .B(_abc_40298_new_n3012_), .Y(_abc_40298_new_n3014_));
NAND2X1 NAND2X1_256 ( .A(_abc_40298_new_n3014_), .B(_abc_40298_new_n3013_), .Y(_abc_40298_new_n3015_));
NAND2X1 NAND2X1_257 ( .A(state_q_3_), .B(pc_q_13_), .Y(_abc_40298_new_n3020_));
NAND2X1 NAND2X1_258 ( .A(\mem_addr_o[13] ), .B(_abc_40298_new_n2895_), .Y(_abc_40298_new_n3021_));
NAND2X1 NAND2X1_259 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_14_), .B(_abc_40298_new_n3025_), .Y(_abc_40298_new_n3033_));
NAND2X1 NAND2X1_26 ( .A(\mem_dat_i[22] ), .B(_abc_40298_new_n688_), .Y(_abc_40298_new_n748_));
NAND2X1 NAND2X1_260 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_15_), .B(_abc_40298_new_n3036_), .Y(_abc_40298_new_n3037_));
NAND2X1 NAND2X1_261 ( .A(_abc_40298_new_n1035_), .B(_abc_40298_new_n3039_), .Y(_abc_40298_new_n3040_));
NAND2X1 NAND2X1_262 ( .A(_abc_40298_new_n3037_), .B(_abc_40298_new_n3040_), .Y(_abc_40298_new_n3041_));
NAND2X1 NAND2X1_263 ( .A(_abc_40298_new_n3046_), .B(_abc_40298_new_n3049_), .Y(_abc_40298_new_n3050_));
NAND2X1 NAND2X1_264 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_16_), .B(_abc_40298_new_n3036_), .Y(_abc_40298_new_n3052_));
NAND2X1 NAND2X1_265 ( .A(_abc_40298_new_n2385_), .B(_abc_40298_new_n3039_), .Y(_abc_40298_new_n3053_));
NAND2X1 NAND2X1_266 ( .A(_abc_40298_new_n3052_), .B(_abc_40298_new_n3053_), .Y(_abc_40298_new_n3054_));
NAND2X1 NAND2X1_267 ( .A(_abc_40298_new_n3066_), .B(_abc_40298_new_n3069_), .Y(_abc_40298_new_n3070_));
NAND2X1 NAND2X1_268 ( .A(_abc_40298_new_n3070_), .B(_abc_40298_new_n3071_), .Y(_abc_40298_new_n3072_));
NAND2X1 NAND2X1_269 ( .A(_abc_40298_new_n3068_), .B(_abc_40298_new_n3082_), .Y(_abc_40298_new_n3083_));
NAND2X1 NAND2X1_27 ( .A(_abc_40298_new_n755_), .B(_abc_40298_new_n756_), .Y(_abc_40298_new_n757_));
NAND2X1 NAND2X1_270 ( .A(_abc_40298_new_n3067_), .B(_abc_40298_new_n3082_), .Y(_abc_40298_new_n3085_));
NAND2X1 NAND2X1_271 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_20_), .B(_abc_40298_new_n3036_), .Y(_abc_40298_new_n3090_));
NAND2X1 NAND2X1_272 ( .A(_abc_40298_new_n2413_), .B(_abc_40298_new_n3039_), .Y(_abc_40298_new_n3091_));
NAND2X1 NAND2X1_273 ( .A(_abc_40298_new_n3090_), .B(_abc_40298_new_n3091_), .Y(_abc_40298_new_n3092_));
NAND2X1 NAND2X1_274 ( .A(_abc_40298_new_n3104_), .B(_abc_40298_new_n3108_), .Y(_abc_40298_new_n3110_));
NAND2X1 NAND2X1_275 ( .A(_abc_40298_new_n2902_), .B(_abc_40298_new_n3110_), .Y(_abc_40298_new_n3111_));
NAND2X1 NAND2X1_276 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_22_), .B(_abc_40298_new_n3036_), .Y(_abc_40298_new_n3114_));
NAND2X1 NAND2X1_277 ( .A(_abc_40298_new_n3115_), .B(_abc_40298_new_n3104_), .Y(_abc_40298_new_n3122_));
NAND2X1 NAND2X1_278 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_24_), .B(_abc_40298_new_n3036_), .Y(_abc_40298_new_n3135_));
NAND2X1 NAND2X1_279 ( .A(state_q_3_), .B(pc_q_26_), .Y(_abc_40298_new_n3152_));
NAND2X1 NAND2X1_28 ( .A(_abc_40298_new_n655_), .B(_abc_40298_new_n758_), .Y(_abc_40298_new_n759_));
NAND2X1 NAND2X1_280 ( .A(\mem_addr_o[26] ), .B(_abc_40298_new_n2895_), .Y(_abc_40298_new_n3153_));
NAND2X1 NAND2X1_281 ( .A(_abc_40298_new_n3149_), .B(_abc_40298_new_n3148_), .Y(_abc_40298_new_n3155_));
NAND2X1 NAND2X1_282 ( .A(_abc_40298_new_n3149_), .B(_abc_40298_new_n3157_), .Y(_abc_40298_new_n3161_));
NAND2X1 NAND2X1_283 ( .A(_abc_40298_new_n3166_), .B(_abc_40298_new_n3165_), .Y(_abc_40298_new_n3168_));
NAND2X1 NAND2X1_284 ( .A(_abc_40298_new_n2902_), .B(_abc_40298_new_n3168_), .Y(_abc_40298_new_n3169_));
NAND2X1 NAND2X1_285 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_30_), .B(_abc_40298_new_n3036_), .Y(_abc_40298_new_n3177_));
NAND2X1 NAND2X1_286 ( .A(_abc_40298_new_n2486_), .B(_abc_40298_new_n3039_), .Y(_abc_40298_new_n3178_));
NAND2X1 NAND2X1_287 ( .A(_abc_40298_new_n3177_), .B(_abc_40298_new_n3178_), .Y(_abc_40298_new_n3179_));
NAND2X1 NAND2X1_288 ( .A(_abc_40298_new_n2470_), .B(_abc_40298_new_n2478_), .Y(_abc_40298_new_n3180_));
NAND2X1 NAND2X1_289 ( .A(_abc_40298_new_n3179_), .B(_abc_40298_new_n3183_), .Y(_abc_40298_new_n3185_));
NAND2X1 NAND2X1_29 ( .A(alu_p_o_7_), .B(_abc_40298_new_n631_), .Y(_abc_40298_new_n761_));
NAND2X1 NAND2X1_290 ( .A(REGFILE_SIM_reg_bank_rd_i_3_), .B(REGFILE_SIM_reg_bank_rd_i_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2101_));
NAND2X1 NAND2X1_291 ( .A(REGFILE_SIM_reg_bank_rd_i_0_), .B(REGFILE_SIM_reg_bank_rd_i_1_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2102_));
NAND2X1 NAND2X1_292 ( .A(REGFILE_SIM_reg_bank_rd_i_4_), .B(REGFILE_SIM_reg_bank_wr_i), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2104_));
NAND2X1 NAND2X1_293 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2105_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2103_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2106_));
NAND2X1 NAND2X1_294 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2105_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2204_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2205_));
NAND2X1 NAND2X1_295 ( .A(REGFILE_SIM_reg_bank_rd_i_0_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2202_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2270_));
NAND2X1 NAND2X1_296 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2105_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2271_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2272_));
NAND2X1 NAND2X1_297 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2337_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2105_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2338_));
NAND2X1 NAND2X1_298 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2105_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2406_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2407_));
NAND2X1 NAND2X1_299 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2105_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2472_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2473_));
NAND2X1 NAND2X1_3 ( .A(inst_r_2_), .B(_abc_40298_new_n619_), .Y(_abc_40298_new_n636_));
NAND2X1 NAND2X1_30 ( .A(_abc_40298_new_n655_), .B(_abc_40298_new_n772_), .Y(_abc_40298_new_n773_));
NAND2X1 NAND2X1_300 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2105_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2538_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2539_));
NAND2X1 NAND2X1_301 ( .A(REGFILE_SIM_reg_bank_rd_i_2_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2404_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2669_));
NAND2X1 NAND2X1_302 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2105_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2670_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2671_));
NAND2X1 NAND2X1_303 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2105_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2736_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2737_));
NAND2X1 NAND2X1_304 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2105_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2802_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2803_));
NAND2X1 NAND2X1_305 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2105_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2935_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2936_));
NAND2X1 NAND2X1_306 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3199_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2103_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3200_));
NAND2X1 NAND2X1_307 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3199_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2204_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3265_));
NAND2X1 NAND2X1_308 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3199_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2271_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3330_));
NAND2X1 NAND2X1_309 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2337_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3199_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3395_));
NAND2X1 NAND2X1_31 ( .A(_abc_40298_new_n655_), .B(_abc_40298_new_n777_), .Y(_abc_40298_new_n778_));
NAND2X1 NAND2X1_310 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3199_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2406_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3461_));
NAND2X1 NAND2X1_311 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3199_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2472_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3526_));
NAND2X1 NAND2X1_312 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3199_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2538_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3657_));
NAND2X1 NAND2X1_313 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3199_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2670_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3787_));
NAND2X1 NAND2X1_314 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3199_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2736_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3852_));
NAND2X1 NAND2X1_315 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3199_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2802_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3917_));
NAND2X1 NAND2X1_316 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3199_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2935_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4047_));
NAND2X1 NAND2X1_317 ( .A(REGFILE_SIM_reg_bank_rb_i_3_), .B(REGFILE_SIM_reg_bank_rb_i_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4178_));
NAND2X1 NAND2X1_318 ( .A(REGFILE_SIM_reg_bank_rb_i_1_), .B(REGFILE_SIM_reg_bank_rb_i_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4196_));
NAND2X1 NAND2X1_319 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4192_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4204_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4205_));
NAND2X1 NAND2X1_32 ( .A(_abc_40298_new_n655_), .B(_abc_40298_new_n782_), .Y(_abc_40298_new_n783_));
NAND2X1 NAND2X1_320 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4215_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4194_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4216_));
NAND2X1 NAND2X1_321 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4213_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4221_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4222_));
NAND2X1 NAND2X1_322 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4189_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4194_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4232_));
NAND2X1 NAND2X1_323 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4237_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4231_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4238_));
NAND2X1 NAND2X1_324 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4179_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4215_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4239_));
NAND2X1 NAND2X1_325 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4215_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4243_));
NAND2X1 NAND2X1_326 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4245_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4252_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4253_));
NAND2X1 NAND2X1_327 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4254_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4223_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_0_));
NAND2X1 NAND2X1_328 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4259_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4262_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4263_));
NAND2X1 NAND2X1_329 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4267_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4270_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4271_));
NAND2X1 NAND2X1_33 ( .A(\mem_dat_i[30] ), .B(_abc_40298_new_n674_), .Y(_abc_40298_new_n795_));
NAND2X1 NAND2X1_330 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4277_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4275_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4278_));
NAND2X1 NAND2X1_331 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4281_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4284_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4285_));
NAND2X1 NAND2X1_332 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4286_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4272_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_1_));
NAND2X1 NAND2X1_333 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4291_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4294_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4295_));
NAND2X1 NAND2X1_334 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4299_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4302_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4303_));
NAND2X1 NAND2X1_335 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4309_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4307_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4310_));
NAND2X1 NAND2X1_336 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4313_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4316_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4317_));
NAND2X1 NAND2X1_337 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4318_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4304_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_2_));
NAND2X1 NAND2X1_338 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4323_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4326_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4327_));
NAND2X1 NAND2X1_339 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4331_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4334_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4335_));
NAND2X1 NAND2X1_34 ( .A(_abc_40298_new_n655_), .B(_abc_40298_new_n796_), .Y(_abc_40298_new_n797_));
NAND2X1 NAND2X1_340 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4341_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4339_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4342_));
NAND2X1 NAND2X1_341 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4345_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4348_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4349_));
NAND2X1 NAND2X1_342 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4350_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4336_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_3_));
NAND2X1 NAND2X1_343 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4355_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4358_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4359_));
NAND2X1 NAND2X1_344 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4363_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4366_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4367_));
NAND2X1 NAND2X1_345 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4373_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4371_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4374_));
NAND2X1 NAND2X1_346 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4377_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4380_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4381_));
NAND2X1 NAND2X1_347 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4382_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4368_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_4_));
NAND2X1 NAND2X1_348 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4387_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4390_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4391_));
NAND2X1 NAND2X1_349 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4395_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4398_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4399_));
NAND2X1 NAND2X1_35 ( .A(_abc_40298_new_n889_), .B(_abc_40298_new_n890_), .Y(_abc_40298_new_n891_));
NAND2X1 NAND2X1_350 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4405_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4403_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4406_));
NAND2X1 NAND2X1_351 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4409_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4412_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4413_));
NAND2X1 NAND2X1_352 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4414_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4400_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_5_));
NAND2X1 NAND2X1_353 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4419_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4422_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4423_));
NAND2X1 NAND2X1_354 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4427_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4430_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4431_));
NAND2X1 NAND2X1_355 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4437_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4435_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4438_));
NAND2X1 NAND2X1_356 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4441_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4444_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4445_));
NAND2X1 NAND2X1_357 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4446_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4432_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_6_));
NAND2X1 NAND2X1_358 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4451_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4454_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4455_));
NAND2X1 NAND2X1_359 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4459_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4462_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4463_));
NAND2X1 NAND2X1_36 ( .A(_abc_40298_new_n893_), .B(_abc_40298_new_n892_), .Y(_abc_40298_new_n894_));
NAND2X1 NAND2X1_360 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4469_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4467_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4470_));
NAND2X1 NAND2X1_361 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4473_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4476_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4477_));
NAND2X1 NAND2X1_362 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4478_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4464_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_7_));
NAND2X1 NAND2X1_363 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4483_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4486_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4487_));
NAND2X1 NAND2X1_364 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4491_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4494_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4495_));
NAND2X1 NAND2X1_365 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4501_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4499_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4502_));
NAND2X1 NAND2X1_366 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4505_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4508_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4509_));
NAND2X1 NAND2X1_367 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4510_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4496_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_8_));
NAND2X1 NAND2X1_368 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4515_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4518_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4519_));
NAND2X1 NAND2X1_369 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4523_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4526_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4527_));
NAND2X1 NAND2X1_37 ( .A(_abc_40298_new_n620_), .B(_abc_40298_new_n639_), .Y(_abc_40298_new_n896_));
NAND2X1 NAND2X1_370 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4533_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4531_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4534_));
NAND2X1 NAND2X1_371 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4537_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4540_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4541_));
NAND2X1 NAND2X1_372 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4542_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4528_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_9_));
NAND2X1 NAND2X1_373 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4547_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4550_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4551_));
NAND2X1 NAND2X1_374 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4555_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4558_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4559_));
NAND2X1 NAND2X1_375 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4565_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4563_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4566_));
NAND2X1 NAND2X1_376 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4569_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4572_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4573_));
NAND2X1 NAND2X1_377 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4574_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4560_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_10_));
NAND2X1 NAND2X1_378 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4579_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4582_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4583_));
NAND2X1 NAND2X1_379 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4587_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4590_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4591_));
NAND2X1 NAND2X1_38 ( .A(alu_op_r_0_), .B(_abc_40298_new_n909_), .Y(_abc_40298_new_n910_));
NAND2X1 NAND2X1_380 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4597_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4595_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4598_));
NAND2X1 NAND2X1_381 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4601_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4604_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4605_));
NAND2X1 NAND2X1_382 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4606_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4592_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_11_));
NAND2X1 NAND2X1_383 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4611_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4614_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4615_));
NAND2X1 NAND2X1_384 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4619_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4622_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4623_));
NAND2X1 NAND2X1_385 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4629_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4627_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4630_));
NAND2X1 NAND2X1_386 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4633_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4636_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4637_));
NAND2X1 NAND2X1_387 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4638_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4624_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_12_));
NAND2X1 NAND2X1_388 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4643_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4646_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4647_));
NAND2X1 NAND2X1_389 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4651_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4654_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4655_));
NAND2X1 NAND2X1_39 ( .A(_abc_40298_new_n901_), .B(_abc_40298_new_n912_), .Y(_abc_40298_new_n913_));
NAND2X1 NAND2X1_390 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4661_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4659_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4662_));
NAND2X1 NAND2X1_391 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4665_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4668_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4669_));
NAND2X1 NAND2X1_392 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4670_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4656_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_13_));
NAND2X1 NAND2X1_393 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4675_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4678_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4679_));
NAND2X1 NAND2X1_394 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4683_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4686_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4687_));
NAND2X1 NAND2X1_395 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4693_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4691_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4694_));
NAND2X1 NAND2X1_396 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4697_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4700_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4701_));
NAND2X1 NAND2X1_397 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4702_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4688_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_14_));
NAND2X1 NAND2X1_398 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4707_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4710_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4711_));
NAND2X1 NAND2X1_399 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4715_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4718_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4719_));
NAND2X1 NAND2X1_4 ( .A(inst_r_1_), .B(inst_r_0_), .Y(_abc_40298_new_n646_));
NAND2X1 NAND2X1_40 ( .A(_abc_40298_new_n890_), .B(_abc_40298_new_n905_), .Y(_abc_40298_new_n920_));
NAND2X1 NAND2X1_400 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4725_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4723_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4726_));
NAND2X1 NAND2X1_401 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4729_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4732_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4733_));
NAND2X1 NAND2X1_402 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4734_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4720_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_15_));
NAND2X1 NAND2X1_403 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4739_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4742_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4743_));
NAND2X1 NAND2X1_404 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4747_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4750_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4751_));
NAND2X1 NAND2X1_405 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4757_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4755_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4758_));
NAND2X1 NAND2X1_406 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4761_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4764_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4765_));
NAND2X1 NAND2X1_407 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4766_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4752_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_16_));
NAND2X1 NAND2X1_408 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4771_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4774_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4775_));
NAND2X1 NAND2X1_409 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4779_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4782_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4783_));
NAND2X1 NAND2X1_41 ( .A(_abc_40298_new_n897_), .B(_abc_40298_new_n921_), .Y(_abc_40298_new_n922_));
NAND2X1 NAND2X1_410 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4789_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4787_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4790_));
NAND2X1 NAND2X1_411 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4793_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4796_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4797_));
NAND2X1 NAND2X1_412 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4798_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4784_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_17_));
NAND2X1 NAND2X1_413 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4803_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4806_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4807_));
NAND2X1 NAND2X1_414 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4811_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4814_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4815_));
NAND2X1 NAND2X1_415 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4821_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4819_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4822_));
NAND2X1 NAND2X1_416 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4825_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4828_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4829_));
NAND2X1 NAND2X1_417 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4830_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4816_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_18_));
NAND2X1 NAND2X1_418 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4835_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4838_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4839_));
NAND2X1 NAND2X1_419 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4843_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4846_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4847_));
NAND2X1 NAND2X1_42 ( .A(alu_op_r_1_), .B(_abc_40298_new_n911_), .Y(_abc_40298_new_n923_));
NAND2X1 NAND2X1_420 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4853_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4851_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4854_));
NAND2X1 NAND2X1_421 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4857_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4860_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4861_));
NAND2X1 NAND2X1_422 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4862_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4848_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_19_));
NAND2X1 NAND2X1_423 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4867_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4870_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4871_));
NAND2X1 NAND2X1_424 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4875_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4878_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4879_));
NAND2X1 NAND2X1_425 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4885_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4883_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4886_));
NAND2X1 NAND2X1_426 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4889_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4892_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4893_));
NAND2X1 NAND2X1_427 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4894_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4880_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_20_));
NAND2X1 NAND2X1_428 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4899_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4902_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4903_));
NAND2X1 NAND2X1_429 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4907_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4910_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4911_));
NAND2X1 NAND2X1_43 ( .A(inst_r_3_), .B(inst_r_5_), .Y(_abc_40298_new_n935_));
NAND2X1 NAND2X1_430 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4917_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4915_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4918_));
NAND2X1 NAND2X1_431 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4921_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4924_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4925_));
NAND2X1 NAND2X1_432 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4926_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4912_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_21_));
NAND2X1 NAND2X1_433 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4931_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4934_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4935_));
NAND2X1 NAND2X1_434 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4939_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4942_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4943_));
NAND2X1 NAND2X1_435 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4949_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4947_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4950_));
NAND2X1 NAND2X1_436 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4953_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4956_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4957_));
NAND2X1 NAND2X1_437 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4958_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4944_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_22_));
NAND2X1 NAND2X1_438 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4963_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4966_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4967_));
NAND2X1 NAND2X1_439 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4971_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4974_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4975_));
NAND2X1 NAND2X1_44 ( .A(inst_r_0_), .B(_abc_40298_new_n624_), .Y(_abc_40298_new_n936_));
NAND2X1 NAND2X1_440 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4981_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4979_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4982_));
NAND2X1 NAND2X1_441 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4985_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4988_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4989_));
NAND2X1 NAND2X1_442 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4990_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4976_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_23_));
NAND2X1 NAND2X1_443 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4995_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4998_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4999_));
NAND2X1 NAND2X1_444 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5003_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5006_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5007_));
NAND2X1 NAND2X1_445 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5013_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5011_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5014_));
NAND2X1 NAND2X1_446 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5017_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5020_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5021_));
NAND2X1 NAND2X1_447 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5022_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5008_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_24_));
NAND2X1 NAND2X1_448 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5027_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5030_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5031_));
NAND2X1 NAND2X1_449 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5035_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5038_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5039_));
NAND2X1 NAND2X1_45 ( .A(_abc_40298_new_n939_), .B(_abc_40298_new_n937_), .Y(_abc_40298_new_n940_));
NAND2X1 NAND2X1_450 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5045_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5043_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5046_));
NAND2X1 NAND2X1_451 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5049_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5052_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5053_));
NAND2X1 NAND2X1_452 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5054_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5040_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_25_));
NAND2X1 NAND2X1_453 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5059_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5062_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5063_));
NAND2X1 NAND2X1_454 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5067_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5070_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5071_));
NAND2X1 NAND2X1_455 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5077_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5075_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5078_));
NAND2X1 NAND2X1_456 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5081_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5084_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5085_));
NAND2X1 NAND2X1_457 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5086_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5072_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_26_));
NAND2X1 NAND2X1_458 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5091_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5094_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5095_));
NAND2X1 NAND2X1_459 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5099_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5102_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5103_));
NAND2X1 NAND2X1_46 ( .A(_abc_40298_new_n945_), .B(_abc_40298_new_n946_), .Y(_abc_40298_new_n947_));
NAND2X1 NAND2X1_460 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5109_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5107_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5110_));
NAND2X1 NAND2X1_461 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5113_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5116_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5117_));
NAND2X1 NAND2X1_462 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5118_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5104_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_27_));
NAND2X1 NAND2X1_463 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5123_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5126_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5127_));
NAND2X1 NAND2X1_464 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5131_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5134_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5135_));
NAND2X1 NAND2X1_465 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5141_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5139_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5142_));
NAND2X1 NAND2X1_466 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5145_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5148_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5149_));
NAND2X1 NAND2X1_467 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5150_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5136_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_28_));
NAND2X1 NAND2X1_468 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5155_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5158_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5159_));
NAND2X1 NAND2X1_469 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5163_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5166_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5167_));
NAND2X1 NAND2X1_47 ( .A(_abc_40298_new_n965_), .B(_abc_40298_new_n964_), .Y(_abc_40298_new_n966_));
NAND2X1 NAND2X1_470 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5173_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5171_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5174_));
NAND2X1 NAND2X1_471 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5177_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5180_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5181_));
NAND2X1 NAND2X1_472 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5182_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5168_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_29_));
NAND2X1 NAND2X1_473 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5187_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5190_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5191_));
NAND2X1 NAND2X1_474 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5195_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5198_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5199_));
NAND2X1 NAND2X1_475 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5205_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5203_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5206_));
NAND2X1 NAND2X1_476 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5209_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5212_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5213_));
NAND2X1 NAND2X1_477 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5214_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5200_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_30_));
NAND2X1 NAND2X1_478 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5219_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5222_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5223_));
NAND2X1 NAND2X1_479 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5227_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5230_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5231_));
NAND2X1 NAND2X1_48 ( .A(_abc_40298_new_n950_), .B(_abc_40298_new_n970_), .Y(_abc_40298_new_n971_));
NAND2X1 NAND2X1_480 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5237_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5235_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5238_));
NAND2X1 NAND2X1_481 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5241_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5244_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5245_));
NAND2X1 NAND2X1_482 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5246_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5232_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_31_));
NAND2X1 NAND2X1_483 ( .A(REGFILE_SIM_reg_bank_ra_i_3_), .B(REGFILE_SIM_reg_bank_ra_i_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5250_));
NAND2X1 NAND2X1_484 ( .A(REGFILE_SIM_reg_bank_ra_i_1_), .B(REGFILE_SIM_reg_bank_ra_i_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5268_));
NAND2X1 NAND2X1_485 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5264_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5276_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5277_));
NAND2X1 NAND2X1_486 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5287_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5266_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5288_));
NAND2X1 NAND2X1_487 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5285_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5293_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5294_));
NAND2X1 NAND2X1_488 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5261_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5266_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5304_));
NAND2X1 NAND2X1_489 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5309_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5303_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5310_));
NAND2X1 NAND2X1_49 ( .A(_abc_40298_new_n897_), .B(_abc_40298_new_n976_), .Y(_abc_40298_new_n977_));
NAND2X1 NAND2X1_490 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5251_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5287_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5311_));
NAND2X1 NAND2X1_491 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5287_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5315_));
NAND2X1 NAND2X1_492 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5317_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5324_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5325_));
NAND2X1 NAND2X1_493 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5326_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5295_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_0_));
NAND2X1 NAND2X1_494 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5331_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5334_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5335_));
NAND2X1 NAND2X1_495 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5339_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5342_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5343_));
NAND2X1 NAND2X1_496 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5349_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5347_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5350_));
NAND2X1 NAND2X1_497 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5353_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5356_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5357_));
NAND2X1 NAND2X1_498 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5358_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5344_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_1_));
NAND2X1 NAND2X1_499 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5363_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5366_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5367_));
NAND2X1 NAND2X1_5 ( .A(_abc_40298_new_n644_), .B(_abc_40298_new_n652_), .Y(_abc_40298_new_n653_));
NAND2X1 NAND2X1_50 ( .A(_abc_40298_new_n978_), .B(_abc_40298_new_n979_), .Y(_abc_40298_new_n980_));
NAND2X1 NAND2X1_500 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5371_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5374_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5375_));
NAND2X1 NAND2X1_501 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5381_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5379_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5382_));
NAND2X1 NAND2X1_502 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5385_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5388_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5389_));
NAND2X1 NAND2X1_503 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5390_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5376_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_2_));
NAND2X1 NAND2X1_504 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5395_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5398_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5399_));
NAND2X1 NAND2X1_505 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5403_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5406_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5407_));
NAND2X1 NAND2X1_506 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5413_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5411_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5414_));
NAND2X1 NAND2X1_507 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5417_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5420_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5421_));
NAND2X1 NAND2X1_508 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5422_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5408_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_3_));
NAND2X1 NAND2X1_509 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5427_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5430_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5431_));
NAND2X1 NAND2X1_51 ( .A(_abc_40298_new_n950_), .B(_abc_40298_new_n964_), .Y(_abc_40298_new_n988_));
NAND2X1 NAND2X1_510 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5435_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5438_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5439_));
NAND2X1 NAND2X1_511 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5445_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5443_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5446_));
NAND2X1 NAND2X1_512 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5449_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5452_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5453_));
NAND2X1 NAND2X1_513 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5454_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5440_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_4_));
NAND2X1 NAND2X1_514 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5459_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5462_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5463_));
NAND2X1 NAND2X1_515 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5467_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5470_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5471_));
NAND2X1 NAND2X1_516 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5477_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5475_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5478_));
NAND2X1 NAND2X1_517 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5481_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5484_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5485_));
NAND2X1 NAND2X1_518 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5486_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5472_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_5_));
NAND2X1 NAND2X1_519 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5491_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5494_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5495_));
NAND2X1 NAND2X1_52 ( .A(_abc_40298_new_n639_), .B(_abc_40298_new_n991_), .Y(_abc_40298_new_n992_));
NAND2X1 NAND2X1_520 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5499_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5502_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5503_));
NAND2X1 NAND2X1_521 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5509_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5507_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5510_));
NAND2X1 NAND2X1_522 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5513_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5516_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5517_));
NAND2X1 NAND2X1_523 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5518_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5504_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_6_));
NAND2X1 NAND2X1_524 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5523_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5526_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5527_));
NAND2X1 NAND2X1_525 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5531_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5534_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5535_));
NAND2X1 NAND2X1_526 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5541_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5539_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5542_));
NAND2X1 NAND2X1_527 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5545_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5548_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5549_));
NAND2X1 NAND2X1_528 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5550_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5536_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_7_));
NAND2X1 NAND2X1_529 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5555_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5558_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5559_));
NAND2X1 NAND2X1_53 ( .A(_abc_40298_new_n946_), .B(_abc_40298_new_n1006_), .Y(_abc_40298_new_n1007_));
NAND2X1 NAND2X1_530 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5563_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5566_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5567_));
NAND2X1 NAND2X1_531 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5573_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5571_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5574_));
NAND2X1 NAND2X1_532 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5577_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5580_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5581_));
NAND2X1 NAND2X1_533 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5582_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5568_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_8_));
NAND2X1 NAND2X1_534 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5587_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5590_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5591_));
NAND2X1 NAND2X1_535 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5595_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5598_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5599_));
NAND2X1 NAND2X1_536 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5605_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5603_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5606_));
NAND2X1 NAND2X1_537 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5609_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5612_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5613_));
NAND2X1 NAND2X1_538 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5614_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5600_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_9_));
NAND2X1 NAND2X1_539 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5619_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5622_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5623_));
NAND2X1 NAND2X1_54 ( .A(_abc_40298_new_n999_), .B(_abc_40298_new_n1010_), .Y(_abc_40298_new_n1011_));
NAND2X1 NAND2X1_540 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5627_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5630_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5631_));
NAND2X1 NAND2X1_541 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5637_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5635_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5638_));
NAND2X1 NAND2X1_542 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5641_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5644_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5645_));
NAND2X1 NAND2X1_543 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5646_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5632_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_10_));
NAND2X1 NAND2X1_544 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5651_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5654_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5655_));
NAND2X1 NAND2X1_545 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5659_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5662_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5663_));
NAND2X1 NAND2X1_546 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5669_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5667_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5670_));
NAND2X1 NAND2X1_547 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5673_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5676_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5677_));
NAND2X1 NAND2X1_548 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5678_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5664_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_11_));
NAND2X1 NAND2X1_549 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5683_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5686_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5687_));
NAND2X1 NAND2X1_55 ( .A(_abc_40298_new_n617_), .B(_abc_40298_new_n684_), .Y(_abc_40298_new_n1014_));
NAND2X1 NAND2X1_550 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5691_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5694_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5695_));
NAND2X1 NAND2X1_551 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5701_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5699_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5702_));
NAND2X1 NAND2X1_552 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5705_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5708_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5709_));
NAND2X1 NAND2X1_553 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5710_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5696_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_12_));
NAND2X1 NAND2X1_554 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5715_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5718_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5719_));
NAND2X1 NAND2X1_555 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5723_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5726_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5727_));
NAND2X1 NAND2X1_556 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5733_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5731_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5734_));
NAND2X1 NAND2X1_557 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5737_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5740_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5741_));
NAND2X1 NAND2X1_558 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5742_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5728_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_13_));
NAND2X1 NAND2X1_559 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5747_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5750_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5751_));
NAND2X1 NAND2X1_56 ( .A(_abc_40298_new_n945_), .B(_abc_40298_new_n964_), .Y(_abc_40298_new_n1020_));
NAND2X1 NAND2X1_560 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5755_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5758_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5759_));
NAND2X1 NAND2X1_561 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5765_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5763_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5766_));
NAND2X1 NAND2X1_562 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5769_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5772_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5773_));
NAND2X1 NAND2X1_563 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5774_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5760_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_14_));
NAND2X1 NAND2X1_564 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5779_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5782_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5783_));
NAND2X1 NAND2X1_565 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5787_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5790_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5791_));
NAND2X1 NAND2X1_566 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5797_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5795_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5798_));
NAND2X1 NAND2X1_567 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5801_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5804_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5805_));
NAND2X1 NAND2X1_568 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5806_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5792_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_15_));
NAND2X1 NAND2X1_569 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5811_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5814_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5815_));
NAND2X1 NAND2X1_57 ( .A(_abc_40298_new_n1020_), .B(_abc_40298_new_n663_), .Y(_abc_40298_new_n1021_));
NAND2X1 NAND2X1_570 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5819_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5822_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5823_));
NAND2X1 NAND2X1_571 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5829_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5827_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5830_));
NAND2X1 NAND2X1_572 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5833_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5836_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5837_));
NAND2X1 NAND2X1_573 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5838_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5824_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_16_));
NAND2X1 NAND2X1_574 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5843_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5846_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5847_));
NAND2X1 NAND2X1_575 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5851_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5854_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5855_));
NAND2X1 NAND2X1_576 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5861_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5859_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5862_));
NAND2X1 NAND2X1_577 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5865_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5868_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5869_));
NAND2X1 NAND2X1_578 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5870_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5856_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_17_));
NAND2X1 NAND2X1_579 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5875_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5878_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5879_));
NAND2X1 NAND2X1_58 ( .A(_abc_40298_new_n990_), .B(_abc_40298_new_n1022_), .Y(_abc_40298_new_n1023_));
NAND2X1 NAND2X1_580 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5883_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5886_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5887_));
NAND2X1 NAND2X1_581 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5893_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5891_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5894_));
NAND2X1 NAND2X1_582 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5897_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5900_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5901_));
NAND2X1 NAND2X1_583 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5902_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5888_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_18_));
NAND2X1 NAND2X1_584 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5907_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5910_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5911_));
NAND2X1 NAND2X1_585 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5915_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5918_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5919_));
NAND2X1 NAND2X1_586 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5925_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5923_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5926_));
NAND2X1 NAND2X1_587 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5929_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5932_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5933_));
NAND2X1 NAND2X1_588 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5934_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5920_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_19_));
NAND2X1 NAND2X1_589 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5939_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5942_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5943_));
NAND2X1 NAND2X1_59 ( .A(_abc_40298_new_n954_), .B(_abc_40298_new_n1024_), .Y(_abc_40298_new_n1025_));
NAND2X1 NAND2X1_590 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5947_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5950_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5951_));
NAND2X1 NAND2X1_591 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5957_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5955_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5958_));
NAND2X1 NAND2X1_592 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5961_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5964_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5965_));
NAND2X1 NAND2X1_593 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5966_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5952_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_20_));
NAND2X1 NAND2X1_594 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5971_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5974_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5975_));
NAND2X1 NAND2X1_595 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5979_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5982_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5983_));
NAND2X1 NAND2X1_596 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5989_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5987_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5990_));
NAND2X1 NAND2X1_597 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5993_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5996_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5997_));
NAND2X1 NAND2X1_598 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5998_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5984_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_21_));
NAND2X1 NAND2X1_599 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6003_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6006_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6007_));
NAND2X1 NAND2X1_6 ( .A(inst_r_0_), .B(_abc_40298_new_n656_), .Y(_abc_40298_new_n657_));
NAND2X1 NAND2X1_60 ( .A(_abc_40298_new_n1026_), .B(_abc_40298_new_n1025_), .Y(_abc_40298_new_n1027_));
NAND2X1 NAND2X1_600 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6011_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6014_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6015_));
NAND2X1 NAND2X1_601 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6021_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6019_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6022_));
NAND2X1 NAND2X1_602 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6025_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6028_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6029_));
NAND2X1 NAND2X1_603 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6030_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6016_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_22_));
NAND2X1 NAND2X1_604 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6035_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6038_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6039_));
NAND2X1 NAND2X1_605 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6043_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6046_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6047_));
NAND2X1 NAND2X1_606 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6053_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6051_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6054_));
NAND2X1 NAND2X1_607 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6057_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6060_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6061_));
NAND2X1 NAND2X1_608 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6062_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6048_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_23_));
NAND2X1 NAND2X1_609 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6067_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6070_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6071_));
NAND2X1 NAND2X1_61 ( .A(_abc_40298_new_n885_), .B(_abc_40298_new_n1028_), .Y(_abc_40298_new_n1029_));
NAND2X1 NAND2X1_610 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6075_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6078_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6079_));
NAND2X1 NAND2X1_611 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6085_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6083_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6086_));
NAND2X1 NAND2X1_612 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6089_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6092_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6093_));
NAND2X1 NAND2X1_613 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6094_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6080_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_24_));
NAND2X1 NAND2X1_614 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6099_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6102_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6103_));
NAND2X1 NAND2X1_615 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6107_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6110_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6111_));
NAND2X1 NAND2X1_616 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6117_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6115_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6118_));
NAND2X1 NAND2X1_617 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6121_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6124_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6125_));
NAND2X1 NAND2X1_618 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6126_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6112_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_25_));
NAND2X1 NAND2X1_619 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6131_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6134_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6135_));
NAND2X1 NAND2X1_62 ( .A(_abc_40298_new_n1033_), .B(_abc_40298_new_n1042_), .Y(_abc_40298_new_n1043_));
NAND2X1 NAND2X1_620 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6139_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6142_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6143_));
NAND2X1 NAND2X1_621 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6149_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6147_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6150_));
NAND2X1 NAND2X1_622 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6153_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6156_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6157_));
NAND2X1 NAND2X1_623 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6158_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6144_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_26_));
NAND2X1 NAND2X1_624 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6163_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6166_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6167_));
NAND2X1 NAND2X1_625 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6171_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6174_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6175_));
NAND2X1 NAND2X1_626 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6181_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6179_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6182_));
NAND2X1 NAND2X1_627 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6185_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6188_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6189_));
NAND2X1 NAND2X1_628 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6190_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6176_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_27_));
NAND2X1 NAND2X1_629 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6195_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6198_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6199_));
NAND2X1 NAND2X1_63 ( .A(_abc_40298_new_n1052_), .B(_abc_40298_new_n1053_), .Y(_abc_40298_new_n1054_));
NAND2X1 NAND2X1_630 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6203_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6206_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6207_));
NAND2X1 NAND2X1_631 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6213_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6211_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6214_));
NAND2X1 NAND2X1_632 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6217_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6220_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6221_));
NAND2X1 NAND2X1_633 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6222_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6208_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_28_));
NAND2X1 NAND2X1_634 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6227_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6230_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6231_));
NAND2X1 NAND2X1_635 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6235_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6238_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6239_));
NAND2X1 NAND2X1_636 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6245_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6243_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6246_));
NAND2X1 NAND2X1_637 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6249_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6252_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6253_));
NAND2X1 NAND2X1_638 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6254_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6240_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_29_));
NAND2X1 NAND2X1_639 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6259_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6262_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6263_));
NAND2X1 NAND2X1_64 ( .A(_abc_40298_new_n1055_), .B(_abc_40298_new_n1056_), .Y(_abc_40298_new_n1057_));
NAND2X1 NAND2X1_640 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6267_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6270_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6271_));
NAND2X1 NAND2X1_641 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6277_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6275_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6278_));
NAND2X1 NAND2X1_642 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6281_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6284_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6285_));
NAND2X1 NAND2X1_643 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6286_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6272_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_30_));
NAND2X1 NAND2X1_644 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6291_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6294_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6295_));
NAND2X1 NAND2X1_645 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6299_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6302_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6303_));
NAND2X1 NAND2X1_646 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6309_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6307_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6310_));
NAND2X1 NAND2X1_647 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6313_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6316_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6317_));
NAND2X1 NAND2X1_648 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6318_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6304_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_31_));
NAND2X1 NAND2X1_649 ( .A(alu__abc_38674_new_n163_), .B(alu__abc_38674_new_n175_), .Y(alu__abc_38674_new_n176_));
NAND2X1 NAND2X1_65 ( .A(_abc_40298_new_n1046_), .B(_abc_40298_new_n1050_), .Y(_abc_40298_new_n1075_));
NAND2X1 NAND2X1_650 ( .A(alu__abc_38674_new_n199_), .B(alu__abc_38674_new_n154_), .Y(alu__abc_38674_new_n200_));
NAND2X1 NAND2X1_651 ( .A(alu_b_i_8_), .B(alu_a_i_8_), .Y(alu__abc_38674_new_n223_));
NAND2X1 NAND2X1_652 ( .A(alu__abc_38674_new_n223_), .B(alu__abc_38674_new_n224_), .Y(alu__abc_38674_new_n225_));
NAND2X1 NAND2X1_653 ( .A(alu_b_i_9_), .B(alu_a_i_9_), .Y(alu__abc_38674_new_n226_));
NAND2X1 NAND2X1_654 ( .A(alu__abc_38674_new_n227_), .B(alu__abc_38674_new_n228_), .Y(alu__abc_38674_new_n229_));
NAND2X1 NAND2X1_655 ( .A(alu__abc_38674_new_n226_), .B(alu__abc_38674_new_n229_), .Y(alu__abc_38674_new_n230_));
NAND2X1 NAND2X1_656 ( .A(alu_b_i_10_), .B(alu_a_i_10_), .Y(alu__abc_38674_new_n231_));
NAND2X1 NAND2X1_657 ( .A(alu__abc_38674_new_n232_), .B(alu__abc_38674_new_n233_), .Y(alu__abc_38674_new_n234_));
NAND2X1 NAND2X1_658 ( .A(alu__abc_38674_new_n231_), .B(alu__abc_38674_new_n234_), .Y(alu__abc_38674_new_n235_));
NAND2X1 NAND2X1_659 ( .A(alu_b_i_11_), .B(alu_a_i_11_), .Y(alu__abc_38674_new_n237_));
NAND2X1 NAND2X1_66 ( .A(_abc_40298_new_n1079_), .B(_abc_40298_new_n1074_), .Y(_abc_40298_new_n1080_));
NAND2X1 NAND2X1_660 ( .A(alu__abc_38674_new_n237_), .B(alu__abc_38674_new_n238_), .Y(alu__abc_38674_new_n239_));
NAND2X1 NAND2X1_661 ( .A(alu_b_i_6_), .B(alu_a_i_6_), .Y(alu__abc_38674_new_n245_));
NAND2X1 NAND2X1_662 ( .A(alu__abc_38674_new_n245_), .B(alu__abc_38674_new_n246_), .Y(alu__abc_38674_new_n247_));
NAND2X1 NAND2X1_663 ( .A(alu_b_i_5_), .B(alu_a_i_5_), .Y(alu__abc_38674_new_n251_));
NAND2X1 NAND2X1_664 ( .A(alu__abc_38674_new_n251_), .B(alu__abc_38674_new_n252_), .Y(alu__abc_38674_new_n253_));
NAND2X1 NAND2X1_665 ( .A(alu_a_i_1_), .B(alu_b_i_1_), .Y(alu__abc_38674_new_n260_));
NAND2X1 NAND2X1_666 ( .A(alu_b_i_0_), .B(alu__abc_38674_new_n258_), .Y(alu__abc_38674_new_n263_));
NAND2X1 NAND2X1_667 ( .A(alu__abc_38674_new_n272_), .B(alu__abc_38674_new_n265_), .Y(alu__abc_38674_new_n273_));
NAND2X1 NAND2X1_668 ( .A(alu_a_i_2_), .B(alu__abc_38674_new_n338_), .Y(alu__abc_38674_new_n339_));
NAND2X1 NAND2X1_669 ( .A(alu_a_i_3_), .B(alu__abc_38674_new_n340_), .Y(alu__abc_38674_new_n341_));
NAND2X1 NAND2X1_67 ( .A(_abc_40298_new_n993_), .B(_abc_40298_new_n1081_), .Y(_abc_40298_new_n1082_));
NAND2X1 NAND2X1_670 ( .A(alu__abc_38674_new_n352_), .B(alu__abc_38674_new_n230_), .Y(alu__abc_38674_new_n353_));
NAND2X1 NAND2X1_671 ( .A(alu_a_i_14_), .B(alu__abc_38674_new_n201_), .Y(alu__abc_38674_new_n366_));
NAND2X1 NAND2X1_672 ( .A(alu__abc_38674_new_n385_), .B(alu__abc_38674_new_n391_), .Y(alu__abc_38674_new_n392_));
NAND2X1 NAND2X1_673 ( .A(alu__abc_38674_new_n114_), .B(alu__abc_38674_new_n321_), .Y(alu__abc_38674_new_n405_));
NAND2X1 NAND2X1_674 ( .A(alu__abc_38674_new_n125_), .B(alu__abc_38674_new_n410_), .Y(alu__abc_38674_new_n411_));
NAND2X1 NAND2X1_675 ( .A(alu__abc_38674_new_n149_), .B(alu__abc_38674_new_n306_), .Y(alu__abc_38674_new_n413_));
NAND2X1 NAND2X1_676 ( .A(alu__abc_38674_new_n417_), .B(alu__abc_38674_new_n412_), .Y(alu__abc_38674_new_n418_));
NAND2X1 NAND2X1_677 ( .A(alu_b_i_0_), .B(alu_a_i_0_), .Y(alu__abc_38674_new_n420_));
NAND2X1 NAND2X1_678 ( .A(alu__abc_38674_new_n424_), .B(alu__abc_38674_new_n422_), .Y(alu__abc_38674_new_n425_));
NAND2X1 NAND2X1_679 ( .A(alu__abc_38674_new_n428_), .B(alu__abc_38674_new_n429_), .Y(alu__abc_38674_new_n430_));
NAND2X1 NAND2X1_68 ( .A(_abc_40298_new_n1092_), .B(_abc_40298_new_n1095_), .Y(_abc_40298_new_n1101_));
NAND2X1 NAND2X1_680 ( .A(alu__abc_38674_new_n433_), .B(alu__abc_38674_new_n335_), .Y(alu__abc_38674_new_n434_));
NAND2X1 NAND2X1_681 ( .A(alu_b_i_4_), .B(alu_a_i_4_), .Y(alu__abc_38674_new_n436_));
NAND2X1 NAND2X1_682 ( .A(alu__abc_38674_new_n240_), .B(alu__abc_38674_new_n236_), .Y(alu__abc_38674_new_n443_));
NAND2X1 NAND2X1_683 ( .A(alu__abc_38674_new_n207_), .B(alu__abc_38674_new_n453_), .Y(alu__abc_38674_new_n454_));
NAND2X1 NAND2X1_684 ( .A(alu__abc_38674_new_n214_), .B(alu__abc_38674_new_n451_), .Y(alu__abc_38674_new_n456_));
NAND2X1 NAND2X1_685 ( .A(alu__abc_38674_new_n459_), .B(alu__abc_38674_new_n460_), .Y(alu__abc_38674_new_n461_));
NAND2X1 NAND2X1_686 ( .A(alu__abc_38674_new_n457_), .B(alu__abc_38674_new_n462_), .Y(alu__abc_38674_new_n463_));
NAND2X1 NAND2X1_687 ( .A(alu__abc_38674_new_n140_), .B(alu__abc_38674_new_n465_), .Y(alu__abc_38674_new_n466_));
NAND2X1 NAND2X1_688 ( .A(alu__abc_38674_new_n473_), .B(alu__abc_38674_new_n398_), .Y(alu__abc_38674_new_n479_));
NAND2X1 NAND2X1_689 ( .A(alu__abc_38674_new_n389_), .B(alu__abc_38674_new_n480_), .Y(alu__abc_38674_new_n481_));
NAND2X1 NAND2X1_69 ( .A(_abc_40298_new_n1020_), .B(_abc_40298_new_n1104_), .Y(_abc_40298_new_n1105_));
NAND2X1 NAND2X1_690 ( .A(alu__abc_38674_new_n506_), .B(alu__abc_38674_new_n505_), .Y(alu__abc_38674_new_n507_));
NAND2X1 NAND2X1_691 ( .A(alu_b_i_7_), .B(alu_a_i_7_), .Y(alu__abc_38674_new_n516_));
NAND2X1 NAND2X1_692 ( .A(alu__abc_38674_new_n516_), .B(alu__abc_38674_new_n439_), .Y(alu__abc_38674_new_n517_));
NAND2X1 NAND2X1_693 ( .A(alu__abc_38674_new_n519_), .B(alu__abc_38674_new_n345_), .Y(alu__abc_38674_new_n520_));
NAND2X1 NAND2X1_694 ( .A(alu__abc_38674_new_n436_), .B(alu__abc_38674_new_n520_), .Y(alu__abc_38674_new_n521_));
NAND2X1 NAND2X1_695 ( .A(alu__abc_38674_new_n518_), .B(alu__abc_38674_new_n522_), .Y(alu__abc_38674_new_n523_));
NAND2X1 NAND2X1_696 ( .A(alu__abc_38674_new_n207_), .B(alu__abc_38674_new_n533_), .Y(alu__abc_38674_new_n534_));
NAND2X1 NAND2X1_697 ( .A(alu__abc_38674_new_n245_), .B(alu__abc_38674_new_n542_), .Y(alu__abc_38674_new_n543_));
NAND2X1 NAND2X1_698 ( .A(alu__abc_38674_new_n522_), .B(alu__abc_38674_new_n425_), .Y(alu__abc_38674_new_n545_));
NAND2X1 NAND2X1_699 ( .A(alu__abc_38674_new_n542_), .B(alu__abc_38674_new_n546_), .Y(alu__abc_38674_new_n547_));
NAND2X1 NAND2X1_7 ( .A(_abc_40298_new_n657_), .B(_abc_40298_new_n659_), .Y(_abc_40298_new_n660_));
NAND2X1 NAND2X1_70 ( .A(_abc_40298_new_n1006_), .B(_abc_40298_new_n964_), .Y(_abc_40298_new_n1113_));
NAND2X1 NAND2X1_700 ( .A(alu__abc_38674_new_n335_), .B(alu__abc_38674_new_n425_), .Y(alu__abc_38674_new_n548_));
NAND2X1 NAND2X1_701 ( .A(alu__abc_38674_new_n551_), .B(alu__abc_38674_new_n549_), .Y(alu__abc_38674_new_n552_));
NAND2X1 NAND2X1_702 ( .A(alu__abc_38674_new_n271_), .B(alu__abc_38674_new_n553_), .Y(alu__abc_38674_new_n554_));
NAND2X1 NAND2X1_703 ( .A(alu__abc_38674_new_n554_), .B(alu__abc_38674_new_n557_), .Y(alu__abc_38674_new_n558_));
NAND2X1 NAND2X1_704 ( .A(alu__abc_38674_new_n336_), .B(alu__abc_38674_new_n559_), .Y(alu__abc_38674_new_n560_));
NAND2X1 NAND2X1_705 ( .A(alu__abc_38674_new_n260_), .B(alu__abc_38674_new_n560_), .Y(alu__abc_38674_new_n561_));
NAND2X1 NAND2X1_706 ( .A(alu__abc_38674_new_n562_), .B(alu__abc_38674_new_n258_), .Y(alu__abc_38674_new_n563_));
NAND2X1 NAND2X1_707 ( .A(alu__abc_38674_new_n268_), .B(alu__abc_38674_new_n421_), .Y(alu__abc_38674_new_n567_));
NAND2X1 NAND2X1_708 ( .A(alu__abc_38674_new_n567_), .B(alu__abc_38674_new_n568_), .Y(alu__abc_38674_new_n569_));
NAND2X1 NAND2X1_709 ( .A(alu__abc_38674_new_n575_), .B(alu__abc_38674_new_n527_), .Y(alu__abc_38674_new_n576_));
NAND2X1 NAND2X1_71 ( .A(_abc_40298_new_n992_), .B(_abc_40298_new_n1147_), .Y(_abc_40298_new_n1148_));
NAND2X1 NAND2X1_710 ( .A(alu__abc_38674_new_n214_), .B(alu__abc_38674_new_n531_), .Y(alu__abc_38674_new_n580_));
NAND2X1 NAND2X1_711 ( .A(alu__abc_38674_new_n581_), .B(alu__abc_38674_new_n583_), .Y(alu__abc_38674_new_n584_));
NAND2X1 NAND2X1_712 ( .A(alu__abc_38674_new_n236_), .B(alu__abc_38674_new_n586_), .Y(alu__abc_38674_new_n587_));
NAND2X1 NAND2X1_713 ( .A(alu__abc_38674_new_n588_), .B(alu__abc_38674_new_n591_), .Y(alu__abc_38674_new_n592_));
NAND2X1 NAND2X1_714 ( .A(alu__abc_38674_new_n595_), .B(alu__abc_38674_new_n594_), .Y(alu__abc_38674_new_n596_));
NAND2X1 NAND2X1_715 ( .A(alu__abc_38674_new_n465_), .B(alu__abc_38674_new_n464_), .Y(alu__abc_38674_new_n601_));
NAND2X1 NAND2X1_716 ( .A(alu__abc_38674_new_n508_), .B(alu__abc_38674_new_n605_), .Y(alu__abc_38674_new_n606_));
NAND2X1 NAND2X1_717 ( .A(alu__abc_38674_new_n162_), .B(alu__abc_38674_new_n612_), .Y(alu__abc_38674_new_n614_));
NAND2X1 NAND2X1_718 ( .A(alu__abc_38674_new_n190_), .B(alu__abc_38674_new_n498_), .Y(alu__abc_38674_new_n617_));
NAND2X1 NAND2X1_719 ( .A(alu__abc_38674_new_n114_), .B(alu__abc_38674_new_n495_), .Y(alu__abc_38674_new_n621_));
NAND2X1 NAND2X1_72 ( .A(_abc_40298_new_n1073_), .B(_abc_40298_new_n1159_), .Y(_abc_40298_new_n1160_));
NAND2X1 NAND2X1_720 ( .A(alu_b_i_0_), .B(alu__abc_38674_new_n356_), .Y(alu__abc_38674_new_n629_));
NAND2X1 NAND2X1_721 ( .A(alu_b_i_0_), .B(alu__abc_38674_new_n228_), .Y(alu__abc_38674_new_n631_));
NAND2X1 NAND2X1_722 ( .A(alu_b_i_0_), .B(alu__abc_38674_new_n217_), .Y(alu__abc_38674_new_n635_));
NAND2X1 NAND2X1_723 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n636_), .Y(alu__abc_38674_new_n637_));
NAND2X1 NAND2X1_724 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n638_), .Y(alu__abc_38674_new_n639_));
NAND2X1 NAND2X1_725 ( .A(alu_b_i_0_), .B(alu__abc_38674_new_n641_), .Y(alu__abc_38674_new_n642_));
NAND2X1 NAND2X1_726 ( .A(alu_b_i_0_), .B(alu__abc_38674_new_n334_), .Y(alu__abc_38674_new_n649_));
NAND2X1 NAND2X1_727 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n650_), .Y(alu__abc_38674_new_n651_));
NAND2X1 NAND2X1_728 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n662_), .Y(alu__abc_38674_new_n663_));
NAND2X1 NAND2X1_729 ( .A(alu_b_i_0_), .B(alu__abc_38674_new_n193_), .Y(alu__abc_38674_new_n665_));
NAND2X1 NAND2X1_73 ( .A(alu_c_i), .B(_abc_40298_new_n1138_), .Y(_abc_40298_new_n1167_));
NAND2X1 NAND2X1_730 ( .A(alu_b_i_0_), .B(alu__abc_38674_new_n295_), .Y(alu__abc_38674_new_n668_));
NAND2X1 NAND2X1_731 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n669_), .Y(alu__abc_38674_new_n670_));
NAND2X1 NAND2X1_732 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n671_), .Y(alu__abc_38674_new_n672_));
NAND2X1 NAND2X1_733 ( .A(alu_b_i_0_), .B(alu__abc_38674_new_n128_), .Y(alu__abc_38674_new_n676_));
NAND2X1 NAND2X1_734 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n677_), .Y(alu__abc_38674_new_n678_));
NAND2X1 NAND2X1_735 ( .A(alu_b_i_0_), .B(alu__abc_38674_new_n312_), .Y(alu__abc_38674_new_n682_));
NAND2X1 NAND2X1_736 ( .A(alu_b_i_1_), .B(alu__abc_38674_new_n683_), .Y(alu__abc_38674_new_n684_));
NAND2X1 NAND2X1_737 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n685_), .Y(alu__abc_38674_new_n686_));
NAND2X1 NAND2X1_738 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n687_), .Y(alu__abc_38674_new_n688_));
NAND2X1 NAND2X1_739 ( .A(alu__abc_38674_new_n278_), .B(alu__abc_38674_new_n657_), .Y(alu__abc_38674_new_n710_));
NAND2X1 NAND2X1_74 ( .A(REGFILE_SIM_reg_bank_wr_i), .B(_abc_40298_new_n1028_), .Y(_abc_40298_new_n1169_));
NAND2X1 NAND2X1_740 ( .A(alu_b_i_0_), .B(alu__abc_38674_new_n135_), .Y(alu__abc_38674_new_n727_));
NAND2X1 NAND2X1_741 ( .A(alu_b_i_0_), .B(alu__abc_38674_new_n202_), .Y(alu__abc_38674_new_n730_));
NAND2X1 NAND2X1_742 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n731_), .Y(alu__abc_38674_new_n732_));
NAND2X1 NAND2X1_743 ( .A(alu_b_i_0_), .B(alu__abc_38674_new_n211_), .Y(alu__abc_38674_new_n735_));
NAND2X1 NAND2X1_744 ( .A(alu_b_i_1_), .B(alu__abc_38674_new_n736_), .Y(alu__abc_38674_new_n737_));
NAND2X1 NAND2X1_745 ( .A(alu_b_i_0_), .B(alu__abc_38674_new_n178_), .Y(alu__abc_38674_new_n742_));
NAND2X1 NAND2X1_746 ( .A(alu_b_i_0_), .B(alu__abc_38674_new_n111_), .Y(alu__abc_38674_new_n745_));
NAND2X1 NAND2X1_747 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n746_), .Y(alu__abc_38674_new_n747_));
NAND2X1 NAND2X1_748 ( .A(alu_b_i_0_), .B(alu__abc_38674_new_n122_), .Y(alu__abc_38674_new_n750_));
NAND2X1 NAND2X1_749 ( .A(alu_b_i_1_), .B(alu__abc_38674_new_n751_), .Y(alu__abc_38674_new_n752_));
NAND2X1 NAND2X1_75 ( .A(_abc_40298_new_n1074_), .B(_abc_40298_new_n1184_), .Y(_abc_40298_new_n1185_));
NAND2X1 NAND2X1_750 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n754_), .Y(alu__abc_38674_new_n755_));
NAND2X1 NAND2X1_751 ( .A(alu_b_i_0_), .B(alu__abc_38674_new_n171_), .Y(alu__abc_38674_new_n757_));
NAND2X1 NAND2X1_752 ( .A(alu_b_i_0_), .B(alu__abc_38674_new_n187_), .Y(alu__abc_38674_new_n760_));
NAND2X1 NAND2X1_753 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n761_), .Y(alu__abc_38674_new_n762_));
NAND2X1 NAND2X1_754 ( .A(alu_a_i_31_), .B(alu__abc_38674_new_n657_), .Y(alu__abc_38674_new_n765_));
NAND2X1 NAND2X1_755 ( .A(alu_a_i_31_), .B(alu__abc_38674_new_n562_), .Y(alu__abc_38674_new_n766_));
NAND2X1 NAND2X1_756 ( .A(alu_b_i_0_), .B(alu__abc_38674_new_n156_), .Y(alu__abc_38674_new_n768_));
NAND2X1 NAND2X1_757 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n769_), .Y(alu__abc_38674_new_n770_));
NAND2X1 NAND2X1_758 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n771_), .Y(alu__abc_38674_new_n772_));
NAND2X1 NAND2X1_759 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n773_), .Y(alu__abc_38674_new_n774_));
NAND2X1 NAND2X1_76 ( .A(_abc_40298_new_n993_), .B(_abc_40298_new_n1186_), .Y(_abc_40298_new_n1187_));
NAND2X1 NAND2X1_760 ( .A(alu_b_i_4_), .B(alu__abc_38674_new_n775_), .Y(alu__abc_38674_new_n776_));
NAND2X1 NAND2X1_761 ( .A(alu__abc_38674_new_n741_), .B(alu__abc_38674_new_n776_), .Y(alu__abc_38674_new_n777_));
NAND2X1 NAND2X1_762 ( .A(alu__abc_38674_new_n780_), .B(alu__abc_38674_new_n701_), .Y(alu__abc_38674_new_n781_));
NAND2X1 NAND2X1_763 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n800_), .Y(alu__abc_38674_new_n801_));
NAND2X1 NAND2X1_764 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n666_), .Y(alu__abc_38674_new_n802_));
NAND2X1 NAND2X1_765 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n683_), .Y(alu__abc_38674_new_n806_));
NAND2X1 NAND2X1_766 ( .A(alu_b_i_1_), .B(alu__abc_38674_new_n669_), .Y(alu__abc_38674_new_n809_));
NAND2X1 NAND2X1_767 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n810_), .Y(alu__abc_38674_new_n811_));
NAND2X1 NAND2X1_768 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n812_), .Y(alu__abc_38674_new_n813_));
NAND2X1 NAND2X1_769 ( .A(alu_b_i_1_), .B(alu__abc_38674_new_n632_), .Y(alu__abc_38674_new_n816_));
NAND2X1 NAND2X1_77 ( .A(_abc_40298_new_n1191_), .B(_abc_40298_new_n1028_), .Y(_abc_40298_new_n1192_));
NAND2X1 NAND2X1_770 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n643_), .Y(alu__abc_38674_new_n820_));
NAND2X1 NAND2X1_771 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n821_), .Y(alu__abc_38674_new_n822_));
NAND2X1 NAND2X1_772 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n630_), .Y(alu__abc_38674_new_n826_));
NAND2X1 NAND2X1_773 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n837_), .Y(alu__abc_38674_new_n838_));
NAND2X1 NAND2X1_774 ( .A(alu__abc_38674_new_n701_), .B(alu__abc_38674_new_n841_), .Y(alu__abc_38674_new_n842_));
NAND2X1 NAND2X1_775 ( .A(alu_a_i_2_), .B(alu__abc_38674_new_n712_), .Y(alu__abc_38674_new_n843_));
NAND2X1 NAND2X1_776 ( .A(alu_b_i_1_), .B(alu__abc_38674_new_n769_), .Y(alu__abc_38674_new_n852_));
NAND2X1 NAND2X1_777 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n853_), .Y(alu__abc_38674_new_n854_));
NAND2X1 NAND2X1_778 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n856_), .Y(alu__abc_38674_new_n857_));
NAND2X1 NAND2X1_779 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n744_), .Y(alu__abc_38674_new_n858_));
NAND2X1 NAND2X1_78 ( .A(_abc_40298_new_n1203_), .B(_abc_40298_new_n1028_), .Y(_abc_40298_new_n1204_));
NAND2X1 NAND2X1_780 ( .A(alu_b_i_1_), .B(alu__abc_38674_new_n746_), .Y(alu__abc_38674_new_n861_));
NAND2X1 NAND2X1_781 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n862_), .Y(alu__abc_38674_new_n863_));
NAND2X1 NAND2X1_782 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n728_), .Y(alu__abc_38674_new_n869_));
NAND2X1 NAND2X1_783 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n736_), .Y(alu__abc_38674_new_n873_));
NAND2X1 NAND2X1_784 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n874_), .Y(alu__abc_38674_new_n875_));
NAND2X1 NAND2X1_785 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n876_), .Y(alu__abc_38674_new_n877_));
NAND2X1 NAND2X1_786 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n885_), .Y(alu__abc_38674_new_n886_));
NAND2X1 NAND2X1_787 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n887_), .Y(alu__abc_38674_new_n888_));
NAND2X1 NAND2X1_788 ( .A(alu__abc_38674_new_n558_), .B(alu__abc_38674_new_n570_), .Y(alu__abc_38674_new_n902_));
NAND2X1 NAND2X1_789 ( .A(alu__abc_38674_new_n903_), .B(alu__abc_38674_new_n902_), .Y(alu__abc_38674_new_n904_));
NAND2X1 NAND2X1_79 ( .A(_abc_40298_new_n617_), .B(_abc_40298_new_n649_), .Y(_abc_40298_new_n1209_));
NAND2X1 NAND2X1_790 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n652_), .Y(alu__abc_38674_new_n909_));
NAND2X1 NAND2X1_791 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n638_), .Y(alu__abc_38674_new_n913_));
NAND2X1 NAND2X1_792 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n671_), .Y(alu__abc_38674_new_n920_));
NAND2X1 NAND2X1_793 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n921_), .Y(alu__abc_38674_new_n922_));
NAND2X1 NAND2X1_794 ( .A(alu_b_i_1_), .B(alu__abc_38674_new_n837_), .Y(alu__abc_38674_new_n928_));
NAND2X1 NAND2X1_795 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n748_), .Y(alu__abc_38674_new_n943_));
NAND2X1 NAND2X1_796 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n944_), .Y(alu__abc_38674_new_n945_));
NAND2X1 NAND2X1_797 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n733_), .Y(alu__abc_38674_new_n948_));
NAND2X1 NAND2X1_798 ( .A(alu_b_i_0_), .B(alu__abc_38674_new_n345_), .Y(alu__abc_38674_new_n954_));
NAND2X1 NAND2X1_799 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n955_), .Y(alu__abc_38674_new_n956_));
NAND2X1 NAND2X1_8 ( .A(_abc_40298_new_n661_), .B(_abc_40298_new_n655_), .Y(_abc_40298_new_n662_));
NAND2X1 NAND2X1_80 ( .A(_abc_40298_new_n1212_), .B(_abc_40298_new_n1211_), .Y(_abc_40298_new_n1213_));
NAND2X1 NAND2X1_800 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n818_), .Y(alu__abc_38674_new_n982_));
NAND2X1 NAND2X1_801 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n824_), .Y(alu__abc_38674_new_n984_));
NAND2X1 NAND2X1_802 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n985_), .Y(alu__abc_38674_new_n986_));
NAND2X1 NAND2X1_803 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n989_), .Y(alu__abc_38674_new_n990_));
NAND2X1 NAND2X1_804 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n993_), .Y(alu__abc_38674_new_n994_));
NAND2X1 NAND2X1_805 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n996_), .Y(alu__abc_38674_new_n997_));
NAND2X1 NAND2X1_806 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n1013_), .Y(alu__abc_38674_new_n1014_));
NAND2X1 NAND2X1_807 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n862_), .Y(alu__abc_38674_new_n1015_));
NAND2X1 NAND2X1_808 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n853_), .Y(alu__abc_38674_new_n1018_));
NAND2X1 NAND2X1_809 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n1021_), .Y(alu__abc_38674_new_n1022_));
NAND2X1 NAND2X1_81 ( .A(_abc_40298_new_n1217_), .B(_abc_40298_new_n985_), .Y(_abc_40298_new_n1218_));
NAND2X1 NAND2X1_810 ( .A(alu_b_i_4_), .B(alu__abc_38674_new_n1023_), .Y(alu__abc_38674_new_n1024_));
NAND2X1 NAND2X1_811 ( .A(alu_b_i_0_), .B(alu__abc_38674_new_n330_), .Y(alu__abc_38674_new_n1027_));
NAND2X1 NAND2X1_812 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n1028_), .Y(alu__abc_38674_new_n1029_));
NAND2X1 NAND2X1_813 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n887_), .Y(alu__abc_38674_new_n1031_));
NAND2X1 NAND2X1_814 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n1032_), .Y(alu__abc_38674_new_n1033_));
NAND2X1 NAND2X1_815 ( .A(alu__abc_38674_new_n429_), .B(alu__abc_38674_new_n543_), .Y(alu__abc_38674_new_n1045_));
NAND2X1 NAND2X1_816 ( .A(alu__abc_38674_new_n1044_), .B(alu__abc_38674_new_n1045_), .Y(alu__abc_38674_new_n1046_));
NAND2X1 NAND2X1_817 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n1050_), .Y(alu__abc_38674_new_n1051_));
NAND2X1 NAND2X1_818 ( .A(alu_b_i_0_), .B(alu__abc_38674_new_n329_), .Y(alu__abc_38674_new_n1060_));
NAND2X1 NAND2X1_819 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n1061_), .Y(alu__abc_38674_new_n1062_));
NAND2X1 NAND2X1_82 ( .A(_abc_40298_new_n1213_), .B(_abc_40298_new_n1220_), .Y(_abc_40298_new_n1221_));
NAND2X1 NAND2X1_820 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n1064_), .Y(alu__abc_38674_new_n1065_));
NAND2X1 NAND2X1_821 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n958_), .Y(alu__abc_38674_new_n1085_));
NAND2X1 NAND2X1_822 ( .A(alu_b_i_0_), .B(alu__abc_38674_new_n351_), .Y(alu__abc_38674_new_n1087_));
NAND2X1 NAND2X1_823 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n1088_), .Y(alu__abc_38674_new_n1089_));
NAND2X1 NAND2X1_824 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n779_), .Y(alu__abc_38674_new_n1092_));
NAND2X1 NAND2X1_825 ( .A(alu__abc_38674_new_n353_), .B(alu__abc_38674_new_n706_), .Y(alu__abc_38674_new_n1102_));
NAND2X1 NAND2X1_826 ( .A(alu__abc_38674_new_n594_), .B(alu__abc_38674_new_n1075_), .Y(alu__abc_38674_new_n1112_));
NAND2X1 NAND2X1_827 ( .A(alu__abc_38674_new_n593_), .B(alu__abc_38674_new_n587_), .Y(alu__abc_38674_new_n1116_));
NAND2X1 NAND2X1_828 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n828_), .Y(alu__abc_38674_new_n1117_));
NAND2X1 NAND2X1_829 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n840_), .Y(alu__abc_38674_new_n1122_));
NAND2X1 NAND2X1_83 ( .A(_abc_40298_new_n1216_), .B(_abc_40298_new_n1234_), .Y(_abc_40298_new_n1236_));
NAND2X1 NAND2X1_830 ( .A(alu_b_i_1_), .B(alu__abc_38674_new_n1061_), .Y(alu__abc_38674_new_n1125_));
NAND2X1 NAND2X1_831 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n1126_), .Y(alu__abc_38674_new_n1127_));
NAND2X1 NAND2X1_832 ( .A(alu__abc_38674_new_n1143_), .B(alu__abc_38674_new_n1144_), .Y(alu__abc_38674_new_n1145_));
NAND2X1 NAND2X1_833 ( .A(alu_b_i_0_), .B(alu__abc_38674_new_n233_), .Y(alu__abc_38674_new_n1152_));
NAND2X1 NAND2X1_834 ( .A(alu_b_i_1_), .B(alu__abc_38674_new_n1088_), .Y(alu__abc_38674_new_n1155_));
NAND2X1 NAND2X1_835 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n1156_), .Y(alu__abc_38674_new_n1157_));
NAND2X1 NAND2X1_836 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n888_), .Y(alu__abc_38674_new_n1160_));
NAND2X1 NAND2X1_837 ( .A(alu__abc_38674_new_n1145_), .B(alu__abc_38674_new_n1113_), .Y(alu__abc_38674_new_n1174_));
NAND2X1 NAND2X1_838 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n1180_), .Y(alu__abc_38674_new_n1181_));
NAND2X1 NAND2X1_839 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n1182_), .Y(alu__abc_38674_new_n1183_));
NAND2X1 NAND2X1_84 ( .A(_abc_40298_new_n1175_), .B(_abc_40298_new_n1238_), .Y(_abc_40298_new_n1239_));
NAND2X1 NAND2X1_840 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n931_), .Y(alu__abc_38674_new_n1186_));
NAND2X1 NAND2X1_841 ( .A(alu__abc_38674_new_n1201_), .B(alu__abc_38674_new_n1202_), .Y(alu__abc_38674_new_n1203_));
NAND2X1 NAND2X1_842 ( .A(alu__abc_38674_new_n1203_), .B(alu__abc_38674_new_n1177_), .Y(alu__abc_38674_new_n1204_));
NAND2X1 NAND2X1_843 ( .A(alu__abc_38674_new_n1200_), .B(alu__abc_38674_new_n1204_), .Y(alu__abc_38674_new_n1205_));
NAND2X1 NAND2X1_844 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n1217_), .Y(alu__abc_38674_new_n1218_));
NAND2X1 NAND2X1_845 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n1090_), .Y(alu__abc_38674_new_n1221_));
NAND2X1 NAND2X1_846 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n959_), .Y(alu__abc_38674_new_n1224_));
NAND2X1 NAND2X1_847 ( .A(alu__abc_38674_new_n453_), .B(alu__abc_38674_new_n1234_), .Y(alu__abc_38674_new_n1235_));
NAND2X1 NAND2X1_848 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n985_), .Y(alu__abc_38674_new_n1242_));
NAND2X1 NAND2X1_849 ( .A(alu__abc_38674_new_n519_), .B(alu__abc_38674_new_n1243_), .Y(alu__abc_38674_new_n1244_));
NAND2X1 NAND2X1_85 ( .A(_abc_40298_new_n1258_), .B(_abc_40298_new_n1257_), .Y(_abc_40298_new_n1259_));
NAND2X1 NAND2X1_850 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n1248_), .Y(alu__abc_38674_new_n1249_));
NAND2X1 NAND2X1_851 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n1250_), .Y(alu__abc_38674_new_n1251_));
NAND2X1 NAND2X1_852 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n1252_), .Y(alu__abc_38674_new_n1253_));
NAND2X1 NAND2X1_853 ( .A(alu__abc_38674_new_n528_), .B(alu__abc_38674_new_n534_), .Y(alu__abc_38674_new_n1266_));
NAND2X1 NAND2X1_854 ( .A(alu__abc_38674_new_n1271_), .B(alu__abc_38674_new_n1267_), .Y(alu__abc_38674_new_n1272_));
NAND2X1 NAND2X1_855 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n1032_), .Y(alu__abc_38674_new_n1279_));
NAND2X1 NAND2X1_856 ( .A(alu_b_i_1_), .B(alu__abc_38674_new_n1217_), .Y(alu__abc_38674_new_n1281_));
NAND2X1 NAND2X1_857 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n1156_), .Y(alu__abc_38674_new_n1284_));
NAND2X1 NAND2X1_858 ( .A(alu__abc_38674_new_n701_), .B(alu__abc_38674_new_n1286_), .Y(alu__abc_38674_new_n1287_));
NAND2X1 NAND2X1_859 ( .A(alu__abc_38674_new_n205_), .B(alu__abc_38674_new_n844_), .Y(alu__abc_38674_new_n1288_));
NAND2X1 NAND2X1_86 ( .A(_abc_40298_new_n1213_), .B(_abc_40298_new_n1269_), .Y(_abc_40298_new_n1270_));
NAND2X1 NAND2X1_860 ( .A(alu__abc_38674_new_n519_), .B(alu__abc_38674_new_n689_), .Y(alu__abc_38674_new_n1307_));
NAND2X1 NAND2X1_861 ( .A(alu_b_i_0_), .B(alu__abc_38674_new_n364_), .Y(alu__abc_38674_new_n1308_));
NAND2X1 NAND2X1_862 ( .A(alu_b_i_1_), .B(alu__abc_38674_new_n1248_), .Y(alu__abc_38674_new_n1311_));
NAND2X1 NAND2X1_863 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n1313_), .Y(alu__abc_38674_new_n1314_));
NAND2X1 NAND2X1_864 ( .A(alu__abc_38674_new_n136_), .B(alu__abc_38674_new_n844_), .Y(alu__abc_38674_new_n1319_));
NAND2X1 NAND2X1_865 ( .A(alu__abc_38674_new_n510_), .B(alu__abc_38674_new_n1270_), .Y(alu__abc_38674_new_n1330_));
NAND2X1 NAND2X1_866 ( .A(alu__abc_38674_new_n706_), .B(alu__abc_38674_new_n309_), .Y(alu__abc_38674_new_n1338_));
NAND2X1 NAND2X1_867 ( .A(alu__abc_38674_new_n519_), .B(alu__abc_38674_new_n775_), .Y(alu__abc_38674_new_n1341_));
NAND2X1 NAND2X1_868 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n1220_), .Y(alu__abc_38674_new_n1342_));
NAND2X1 NAND2X1_869 ( .A(alu__abc_38674_new_n600_), .B(alu__abc_38674_new_n1331_), .Y(alu__abc_38674_new_n1359_));
NAND2X1 NAND2X1_87 ( .A(alu_op_r_3_), .B(pc_q_5_), .Y(_abc_40298_new_n1279_));
NAND2X1 NAND2X1_870 ( .A(alu__abc_38674_new_n381_), .B(alu__abc_38674_new_n1359_), .Y(alu__abc_38674_new_n1360_));
NAND2X1 NAND2X1_871 ( .A(alu_b_i_0_), .B(alu__abc_38674_new_n308_), .Y(alu__abc_38674_new_n1368_));
NAND2X1 NAND2X1_872 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n1369_), .Y(alu__abc_38674_new_n1370_));
NAND2X1 NAND2X1_873 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n1250_), .Y(alu__abc_38674_new_n1373_));
NAND2X1 NAND2X1_874 ( .A(alu__abc_38674_new_n1384_), .B(alu__abc_38674_new_n1359_), .Y(alu__abc_38674_new_n1386_));
NAND2X1 NAND2X1_875 ( .A(alu__abc_38674_new_n282_), .B(alu__abc_38674_new_n490_), .Y(alu__abc_38674_new_n1388_));
NAND2X1 NAND2X1_876 ( .A(alu_b_i_0_), .B(alu__abc_38674_new_n144_), .Y(alu__abc_38674_new_n1389_));
NAND2X1 NAND2X1_877 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n1390_), .Y(alu__abc_38674_new_n1391_));
NAND2X1 NAND2X1_878 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n1392_), .Y(alu__abc_38674_new_n1393_));
NAND2X1 NAND2X1_879 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n1394_), .Y(alu__abc_38674_new_n1395_));
NAND2X1 NAND2X1_88 ( .A(_abc_40298_new_n1287_), .B(_abc_40298_new_n1258_), .Y(_abc_40298_new_n1288_));
NAND2X1 NAND2X1_880 ( .A(alu_b_i_4_), .B(alu__abc_38674_new_n889_), .Y(alu__abc_38674_new_n1397_));
NAND2X1 NAND2X1_881 ( .A(alu__abc_38674_new_n147_), .B(alu__abc_38674_new_n844_), .Y(alu__abc_38674_new_n1407_));
NAND2X1 NAND2X1_882 ( .A(alu__abc_38674_new_n315_), .B(alu__abc_38674_new_n311_), .Y(alu__abc_38674_new_n1420_));
NAND2X1 NAND2X1_883 ( .A(alu_b_i_1_), .B(alu__abc_38674_new_n1369_), .Y(alu__abc_38674_new_n1427_));
NAND2X1 NAND2X1_884 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n1428_), .Y(alu__abc_38674_new_n1429_));
NAND2X1 NAND2X1_885 ( .A(alu__abc_38674_new_n1444_), .B(alu__abc_38674_new_n1446_), .Y(alu__abc_38674_new_n1447_));
NAND2X1 NAND2X1_886 ( .A(alu__abc_38674_new_n519_), .B(alu__abc_38674_new_n946_), .Y(alu__abc_38674_new_n1452_));
NAND2X1 NAND2X1_887 ( .A(alu_b_i_1_), .B(alu__abc_38674_new_n1390_), .Y(alu__abc_38674_new_n1455_));
NAND2X1 NAND2X1_888 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n1475_), .Y(alu__abc_38674_new_n1476_));
NAND2X1 NAND2X1_889 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n1477_), .Y(alu__abc_38674_new_n1478_));
NAND2X1 NAND2X1_89 ( .A(_abc_40298_new_n1288_), .B(_abc_40298_new_n1289_), .Y(_abc_40298_new_n1290_));
NAND2X1 NAND2X1_890 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n1479_), .Y(alu__abc_38674_new_n1480_));
NAND2X1 NAND2X1_891 ( .A(alu_b_i_4_), .B(alu__abc_38674_new_n999_), .Y(alu__abc_38674_new_n1482_));
NAND2X1 NAND2X1_892 ( .A(alu__abc_38674_new_n519_), .B(alu__abc_38674_new_n991_), .Y(alu__abc_38674_new_n1484_));
NAND2X1 NAND2X1_893 ( .A(alu__abc_38674_new_n112_), .B(alu__abc_38674_new_n844_), .Y(alu__abc_38674_new_n1491_));
NAND2X1 NAND2X1_894 ( .A(alu__abc_38674_new_n282_), .B(alu__abc_38674_new_n623_), .Y(alu__abc_38674_new_n1497_));
NAND2X1 NAND2X1_895 ( .A(alu__abc_38674_new_n1500_), .B(alu__abc_38674_new_n1499_), .Y(alu__abc_38674_new_n1501_));
NAND2X1 NAND2X1_896 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n1507_), .Y(alu__abc_38674_new_n1508_));
NAND2X1 NAND2X1_897 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n1509_), .Y(alu__abc_38674_new_n1510_));
NAND2X1 NAND2X1_898 ( .A(alu__abc_38674_new_n327_), .B(alu__abc_38674_new_n370_), .Y(alu__abc_38674_new_n1528_));
NAND2X1 NAND2X1_899 ( .A(alu__abc_38674_new_n519_), .B(alu__abc_38674_new_n1054_), .Y(alu__abc_38674_new_n1532_));
NAND2X1 NAND2X1_9 ( .A(\mem_dat_i[16] ), .B(_abc_40298_new_n677_), .Y(_abc_40298_new_n678_));
NAND2X1 NAND2X1_90 ( .A(_abc_40298_new_n1290_), .B(_abc_40298_new_n1232_), .Y(_abc_40298_new_n1291_));
NAND2X1 NAND2X1_900 ( .A(alu_b_i_0_), .B(alu__abc_38674_new_n117_), .Y(alu__abc_38674_new_n1533_));
NAND2X1 NAND2X1_901 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n1428_), .Y(alu__abc_38674_new_n1536_));
NAND2X1 NAND2X1_902 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n1315_), .Y(alu__abc_38674_new_n1538_));
NAND2X1 NAND2X1_903 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n1456_), .Y(alu__abc_38674_new_n1550_));
NAND2X1 NAND2X1_904 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n1552_), .Y(alu__abc_38674_new_n1553_));
NAND2X1 NAND2X1_905 ( .A(alu__abc_38674_new_n519_), .B(alu__abc_38674_new_n1119_), .Y(alu__abc_38674_new_n1583_));
NAND2X1 NAND2X1_906 ( .A(alu_b_i_1_), .B(alu__abc_38674_new_n1534_), .Y(alu__abc_38674_new_n1587_));
NAND2X1 NAND2X1_907 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n1588_), .Y(alu__abc_38674_new_n1589_));
NAND2X1 NAND2X1_908 ( .A(alu__abc_38674_new_n1317_), .B(alu__abc_38674_new_n1129_), .Y(alu__abc_38674_new_n1594_));
NAND2X1 NAND2X1_909 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n1608_), .Y(alu__abc_38674_new_n1609_));
NAND2X1 NAND2X1_91 ( .A(_abc_40298_new_n1295_), .B(_abc_40298_new_n1168_), .Y(_abc_40298_new_n1296_));
NAND2X1 NAND2X1_910 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n1509_), .Y(alu__abc_38674_new_n1611_));
NAND2X1 NAND2X1_911 ( .A(alu__abc_38674_new_n1614_), .B(alu__abc_38674_new_n1618_), .Y(alu__abc_38674_new_n1619_));
NAND2X1 NAND2X1_912 ( .A(alu__abc_38674_new_n381_), .B(alu__abc_38674_new_n1626_), .Y(alu__abc_38674_new_n1627_));
NAND2X1 NAND2X1_913 ( .A(alu__abc_38674_new_n282_), .B(alu__abc_38674_new_n484_), .Y(alu__abc_38674_new_n1628_));
NAND2X1 NAND2X1_914 ( .A(alu__abc_38674_new_n389_), .B(alu__abc_38674_new_n372_), .Y(alu__abc_38674_new_n1630_));
NAND2X1 NAND2X1_915 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n1430_), .Y(alu__abc_38674_new_n1633_));
NAND2X1 NAND2X1_916 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n1656_), .Y(alu__abc_38674_new_n1657_));
NAND2X1 NAND2X1_917 ( .A(alu__abc_38674_new_n519_), .B(alu__abc_38674_new_n1215_), .Y(alu__abc_38674_new_n1663_));
NAND2X1 NAND2X1_918 ( .A(alu__abc_38674_new_n282_), .B(alu__abc_38674_new_n616_), .Y(alu__abc_38674_new_n1678_));
NAND2X1 NAND2X1_919 ( .A(alu_b_i_1_), .B(alu__abc_38674_new_n1634_), .Y(alu__abc_38674_new_n1681_));
NAND2X1 NAND2X1_92 ( .A(_abc_40298_new_n1261_), .B(_abc_40298_new_n1310_), .Y(_abc_40298_new_n1311_));
NAND2X1 NAND2X1_920 ( .A(alu__abc_38674_new_n1693_), .B(alu__abc_38674_new_n1674_), .Y(alu_p_o_30_));
NAND2X1 NAND2X1_921 ( .A(alu__abc_38674_new_n1701_), .B(alu__abc_38674_new_n1702_), .Y(alu__abc_38674_new_n1703_));
NAND2X1 NAND2X1_922 ( .A(alu__abc_38674_new_n519_), .B(alu__abc_38674_new_n1277_), .Y(alu__abc_38674_new_n1704_));
NAND2X1 NAND2X1_923 ( .A(alu__abc_38674_new_n160_), .B(alu__abc_38674_new_n844_), .Y(alu__abc_38674_new_n1712_));
NAND2X1 NAND2X1_93 ( .A(_abc_40298_new_n1312_), .B(_abc_40298_new_n1311_), .Y(_abc_40298_new_n1313_));
NAND2X1 NAND2X1_94 ( .A(_abc_40298_new_n1175_), .B(_abc_40298_new_n1353_), .Y(_abc_40298_new_n1354_));
NAND2X1 NAND2X1_95 ( .A(_abc_40298_new_n1364_), .B(_abc_40298_new_n1363_), .Y(_abc_40298_new_n1365_));
NAND2X1 NAND2X1_96 ( .A(_abc_40298_new_n1175_), .B(_abc_40298_new_n1380_), .Y(_abc_40298_new_n1381_));
NAND2X1 NAND2X1_97 ( .A(_abc_40298_new_n1365_), .B(_abc_40298_new_n1232_), .Y(_abc_40298_new_n1383_));
NAND2X1 NAND2X1_98 ( .A(_abc_40298_new_n1415_), .B(_abc_40298_new_n1417_), .Y(_abc_40298_new_n1418_));
NAND2X1 NAND2X1_99 ( .A(_abc_40298_new_n1376_), .B(_abc_40298_new_n1403_), .Y(_abc_40298_new_n1423_));
NAND3X1 NAND3X1_1 ( .A(_abc_40298_new_n619_), .B(_abc_40298_new_n644_), .C(_abc_40298_new_n660_), .Y(_abc_40298_new_n661_));
NAND3X1 NAND3X1_10 ( .A(_abc_40298_new_n942_), .B(_abc_40298_new_n952_), .C(_abc_40298_new_n928_), .Y(_abc_40298_new_n953_));
NAND3X1 NAND3X1_100 ( .A(REGFILE_SIM_reg_bank_rb_i_4_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4200_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4225_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4226_));
NAND3X1 NAND3X1_101 ( .A(REGFILE_SIM_reg_bank_rb_i_4_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4197_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4179_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4228_));
NAND3X1 NAND3X1_102 ( .A(REGFILE_SIM_reg_bank_rb_i_4_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4225_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4179_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4229_));
NAND3X1 NAND3X1_103 ( .A(REGFILE_SIM_reg_bank_rb_i_4_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4225_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4194_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4234_));
NAND3X1 NAND3X1_104 ( .A(REGFILE_SIM_reg_bank_rb_i_4_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4200_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4197_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4235_));
NAND3X1 NAND3X1_105 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4179_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4177_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4240_));
NAND3X1 NAND3X1_106 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4177_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4242_));
NAND3X1 NAND3X1_107 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4200_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4189_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4246_));
NAND3X1 NAND3X1_108 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4200_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4197_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4247_));
NAND3X1 NAND3X1_109 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4197_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4194_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4249_));
NAND3X1 NAND3X1_11 ( .A(_abc_40298_new_n623_), .B(_abc_40298_new_n938_), .C(_abc_40298_new_n937_), .Y(_abc_40298_new_n963_));
NAND3X1 NAND3X1_110 ( .A(REGFILE_SIM_reg_bank_rb_i_4_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4179_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4189_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4250_));
NAND3X1 NAND3X1_111 ( .A(REGFILE_SIM_reg_bank_reg_r24_1_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4184_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4256_));
NAND3X1 NAND3X1_112 ( .A(REGFILE_SIM_reg_bank_reg_r15_1_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4209_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4265_));
NAND3X1 NAND3X1_113 ( .A(REGFILE_SIM_reg_bank_reg_r24_2_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4184_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4288_));
NAND3X1 NAND3X1_114 ( .A(REGFILE_SIM_reg_bank_reg_r15_2_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4209_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4297_));
NAND3X1 NAND3X1_115 ( .A(REGFILE_SIM_reg_bank_reg_r24_3_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4184_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4320_));
NAND3X1 NAND3X1_116 ( .A(REGFILE_SIM_reg_bank_reg_r15_3_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4209_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4329_));
NAND3X1 NAND3X1_117 ( .A(REGFILE_SIM_reg_bank_reg_r24_4_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4184_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4352_));
NAND3X1 NAND3X1_118 ( .A(REGFILE_SIM_reg_bank_reg_r15_4_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4209_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4361_));
NAND3X1 NAND3X1_119 ( .A(REGFILE_SIM_reg_bank_reg_r24_5_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4184_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4384_));
NAND3X1 NAND3X1_12 ( .A(_abc_40298_new_n966_), .B(_abc_40298_new_n971_), .C(_abc_40298_new_n962_), .Y(_abc_40298_new_n972_));
NAND3X1 NAND3X1_120 ( .A(REGFILE_SIM_reg_bank_reg_r15_5_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4209_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4393_));
NAND3X1 NAND3X1_121 ( .A(REGFILE_SIM_reg_bank_reg_r24_6_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4184_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4416_));
NAND3X1 NAND3X1_122 ( .A(REGFILE_SIM_reg_bank_reg_r15_6_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4209_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4425_));
NAND3X1 NAND3X1_123 ( .A(REGFILE_SIM_reg_bank_reg_r24_7_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4184_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4448_));
NAND3X1 NAND3X1_124 ( .A(REGFILE_SIM_reg_bank_reg_r15_7_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4209_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4457_));
NAND3X1 NAND3X1_125 ( .A(REGFILE_SIM_reg_bank_reg_r24_8_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4184_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4480_));
NAND3X1 NAND3X1_126 ( .A(REGFILE_SIM_reg_bank_reg_r15_8_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4209_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4489_));
NAND3X1 NAND3X1_127 ( .A(REGFILE_SIM_reg_bank_reg_r24_9_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4184_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4512_));
NAND3X1 NAND3X1_128 ( .A(REGFILE_SIM_reg_bank_reg_r15_9_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4209_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4521_));
NAND3X1 NAND3X1_129 ( .A(REGFILE_SIM_reg_bank_reg_r24_10_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4184_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4544_));
NAND3X1 NAND3X1_13 ( .A(_abc_40298_new_n977_), .B(_abc_40298_new_n985_), .C(_abc_40298_new_n982_), .Y(_abc_40298_new_n986_));
NAND3X1 NAND3X1_130 ( .A(REGFILE_SIM_reg_bank_reg_r15_10_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4209_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4553_));
NAND3X1 NAND3X1_131 ( .A(REGFILE_SIM_reg_bank_reg_r24_11_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4184_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4576_));
NAND3X1 NAND3X1_132 ( .A(REGFILE_SIM_reg_bank_reg_r15_11_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4209_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4585_));
NAND3X1 NAND3X1_133 ( .A(REGFILE_SIM_reg_bank_reg_r24_12_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4184_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4608_));
NAND3X1 NAND3X1_134 ( .A(REGFILE_SIM_reg_bank_reg_r15_12_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4209_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4617_));
NAND3X1 NAND3X1_135 ( .A(REGFILE_SIM_reg_bank_reg_r24_13_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4184_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4640_));
NAND3X1 NAND3X1_136 ( .A(REGFILE_SIM_reg_bank_reg_r15_13_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4209_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4649_));
NAND3X1 NAND3X1_137 ( .A(REGFILE_SIM_reg_bank_reg_r24_14_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4184_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4672_));
NAND3X1 NAND3X1_138 ( .A(REGFILE_SIM_reg_bank_reg_r15_14_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4209_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4681_));
NAND3X1 NAND3X1_139 ( .A(REGFILE_SIM_reg_bank_reg_r24_15_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4184_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4704_));
NAND3X1 NAND3X1_14 ( .A(_abc_40298_new_n1014_), .B(_abc_40298_new_n1013_), .C(_abc_40298_new_n1016_), .Y(_abc_40298_new_n1017_));
NAND3X1 NAND3X1_140 ( .A(REGFILE_SIM_reg_bank_reg_r15_15_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4209_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4713_));
NAND3X1 NAND3X1_141 ( .A(REGFILE_SIM_reg_bank_reg_r24_16_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4184_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4736_));
NAND3X1 NAND3X1_142 ( .A(REGFILE_SIM_reg_bank_reg_r15_16_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4209_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4745_));
NAND3X1 NAND3X1_143 ( .A(REGFILE_SIM_reg_bank_reg_r24_17_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4184_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4768_));
NAND3X1 NAND3X1_144 ( .A(REGFILE_SIM_reg_bank_reg_r15_17_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4209_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4777_));
NAND3X1 NAND3X1_145 ( .A(REGFILE_SIM_reg_bank_reg_r24_18_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4184_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4800_));
NAND3X1 NAND3X1_146 ( .A(REGFILE_SIM_reg_bank_reg_r15_18_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4209_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4809_));
NAND3X1 NAND3X1_147 ( .A(REGFILE_SIM_reg_bank_reg_r24_19_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4184_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4832_));
NAND3X1 NAND3X1_148 ( .A(REGFILE_SIM_reg_bank_reg_r15_19_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4209_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4841_));
NAND3X1 NAND3X1_149 ( .A(REGFILE_SIM_reg_bank_reg_r24_20_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4184_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4864_));
NAND3X1 NAND3X1_15 ( .A(_abc_40298_new_n997_), .B(_abc_40298_new_n1005_), .C(_abc_40298_new_n1018_), .Y(_abc_40298_new_n1019_));
NAND3X1 NAND3X1_150 ( .A(REGFILE_SIM_reg_bank_reg_r15_20_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4209_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4873_));
NAND3X1 NAND3X1_151 ( .A(REGFILE_SIM_reg_bank_reg_r24_21_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4184_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4896_));
NAND3X1 NAND3X1_152 ( .A(REGFILE_SIM_reg_bank_reg_r15_21_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4209_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4905_));
NAND3X1 NAND3X1_153 ( .A(REGFILE_SIM_reg_bank_reg_r24_22_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4184_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4928_));
NAND3X1 NAND3X1_154 ( .A(REGFILE_SIM_reg_bank_reg_r15_22_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4209_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4937_));
NAND3X1 NAND3X1_155 ( .A(REGFILE_SIM_reg_bank_reg_r24_23_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4184_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4960_));
NAND3X1 NAND3X1_156 ( .A(REGFILE_SIM_reg_bank_reg_r15_23_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4209_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4969_));
NAND3X1 NAND3X1_157 ( .A(REGFILE_SIM_reg_bank_reg_r24_24_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4184_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4992_));
NAND3X1 NAND3X1_158 ( .A(REGFILE_SIM_reg_bank_reg_r15_24_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4209_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5001_));
NAND3X1 NAND3X1_159 ( .A(REGFILE_SIM_reg_bank_reg_r24_25_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4184_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5024_));
NAND3X1 NAND3X1_16 ( .A(_abc_40298_new_n1034_), .B(_abc_40298_new_n1035_), .C(_abc_40298_new_n1036_), .Y(_abc_40298_new_n1037_));
NAND3X1 NAND3X1_160 ( .A(REGFILE_SIM_reg_bank_reg_r15_25_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4209_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5033_));
NAND3X1 NAND3X1_161 ( .A(REGFILE_SIM_reg_bank_reg_r24_26_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4184_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5056_));
NAND3X1 NAND3X1_162 ( .A(REGFILE_SIM_reg_bank_reg_r15_26_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4209_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5065_));
NAND3X1 NAND3X1_163 ( .A(REGFILE_SIM_reg_bank_reg_r24_27_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4184_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5088_));
NAND3X1 NAND3X1_164 ( .A(REGFILE_SIM_reg_bank_reg_r15_27_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4209_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5097_));
NAND3X1 NAND3X1_165 ( .A(REGFILE_SIM_reg_bank_reg_r24_28_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4184_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5120_));
NAND3X1 NAND3X1_166 ( .A(REGFILE_SIM_reg_bank_reg_r15_28_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4209_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5129_));
NAND3X1 NAND3X1_167 ( .A(REGFILE_SIM_reg_bank_reg_r24_29_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4184_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5152_));
NAND3X1 NAND3X1_168 ( .A(REGFILE_SIM_reg_bank_reg_r15_29_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4209_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5161_));
NAND3X1 NAND3X1_169 ( .A(REGFILE_SIM_reg_bank_reg_r24_30_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4184_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5184_));
NAND3X1 NAND3X1_17 ( .A(_abc_40298_new_n1038_), .B(_abc_40298_new_n1039_), .C(_abc_40298_new_n1040_), .Y(_abc_40298_new_n1041_));
NAND3X1 NAND3X1_170 ( .A(REGFILE_SIM_reg_bank_reg_r15_30_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4209_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5193_));
NAND3X1 NAND3X1_171 ( .A(REGFILE_SIM_reg_bank_reg_r24_31_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4184_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5216_));
NAND3X1 NAND3X1_172 ( .A(REGFILE_SIM_reg_bank_reg_r15_31_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4209_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5225_));
NAND3X1 NAND3X1_173 ( .A(REGFILE_SIM_reg_bank_ra_i_4_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5251_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5249_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5252_));
NAND3X1 NAND3X1_174 ( .A(REGFILE_SIM_reg_bank_reg_r24_0_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5256_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5257_));
NAND3X1 NAND3X1_175 ( .A(REGFILE_SIM_reg_bank_ra_i_4_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5249_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5259_));
NAND3X1 NAND3X1_176 ( .A(REGFILE_SIM_reg_bank_ra_i_4_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5261_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5262_));
NAND3X1 NAND3X1_177 ( .A(REGFILE_SIM_reg_bank_ra_i_4_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5249_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5266_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5267_));
NAND3X1 NAND3X1_178 ( .A(REGFILE_SIM_reg_bank_ra_i_4_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5269_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5266_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5270_));
NAND3X1 NAND3X1_179 ( .A(REGFILE_SIM_reg_bank_ra_i_4_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5272_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5249_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5273_));
NAND3X1 NAND3X1_18 ( .A(_abc_40298_new_n1047_), .B(_abc_40298_new_n1051_), .C(_abc_40298_new_n1058_), .Y(_abc_40298_new_n1059_));
NAND3X1 NAND3X1_180 ( .A(REGFILE_SIM_reg_bank_ra_i_4_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5272_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5261_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5274_));
NAND3X1 NAND3X1_181 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5261_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5278_));
NAND3X1 NAND3X1_182 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5269_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5279_));
NAND3X1 NAND3X1_183 ( .A(REGFILE_SIM_reg_bank_reg_r15_0_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5281_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5282_));
NAND3X1 NAND3X1_184 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5251_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5261_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5283_));
NAND3X1 NAND3X1_185 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5272_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5249_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5286_));
NAND3X1 NAND3X1_186 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5261_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5266_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5290_));
NAND3X1 NAND3X1_187 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5249_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5266_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5291_));
NAND3X1 NAND3X1_188 ( .A(REGFILE_SIM_reg_bank_ra_i_4_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5269_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5296_));
NAND3X1 NAND3X1_189 ( .A(REGFILE_SIM_reg_bank_ra_i_4_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5272_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5297_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5298_));
NAND3X1 NAND3X1_19 ( .A(_abc_40298_new_n1044_), .B(_abc_40298_new_n1048_), .C(_abc_40298_new_n1052_), .Y(_abc_40298_new_n1077_));
NAND3X1 NAND3X1_190 ( .A(REGFILE_SIM_reg_bank_ra_i_4_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5269_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5251_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5300_));
NAND3X1 NAND3X1_191 ( .A(REGFILE_SIM_reg_bank_ra_i_4_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5297_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5251_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5301_));
NAND3X1 NAND3X1_192 ( .A(REGFILE_SIM_reg_bank_ra_i_4_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5297_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5266_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5306_));
NAND3X1 NAND3X1_193 ( .A(REGFILE_SIM_reg_bank_ra_i_4_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5272_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5269_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5307_));
NAND3X1 NAND3X1_194 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5251_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5249_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5312_));
NAND3X1 NAND3X1_195 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5249_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5314_));
NAND3X1 NAND3X1_196 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5272_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5261_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5318_));
NAND3X1 NAND3X1_197 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5272_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5269_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5319_));
NAND3X1 NAND3X1_198 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5269_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5266_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5321_));
NAND3X1 NAND3X1_199 ( .A(REGFILE_SIM_reg_bank_ra_i_4_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5251_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5261_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5322_));
NAND3X1 NAND3X1_2 ( .A(_abc_40298_new_n678_), .B(_abc_40298_new_n680_), .C(_abc_40298_new_n675_), .Y(_abc_40298_new_n681_));
NAND3X1 NAND3X1_20 ( .A(_abc_40298_new_n1095_), .B(_abc_40298_new_n934_), .C(_abc_40298_new_n970_), .Y(_abc_40298_new_n1096_));
NAND3X1 NAND3X1_200 ( .A(REGFILE_SIM_reg_bank_reg_r24_1_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5256_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5328_));
NAND3X1 NAND3X1_201 ( .A(REGFILE_SIM_reg_bank_reg_r15_1_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5281_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5337_));
NAND3X1 NAND3X1_202 ( .A(REGFILE_SIM_reg_bank_reg_r24_2_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5256_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5360_));
NAND3X1 NAND3X1_203 ( .A(REGFILE_SIM_reg_bank_reg_r15_2_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5281_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5369_));
NAND3X1 NAND3X1_204 ( .A(REGFILE_SIM_reg_bank_reg_r24_3_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5256_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5392_));
NAND3X1 NAND3X1_205 ( .A(REGFILE_SIM_reg_bank_reg_r15_3_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5281_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5401_));
NAND3X1 NAND3X1_206 ( .A(REGFILE_SIM_reg_bank_reg_r24_4_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5256_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5424_));
NAND3X1 NAND3X1_207 ( .A(REGFILE_SIM_reg_bank_reg_r15_4_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5281_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5433_));
NAND3X1 NAND3X1_208 ( .A(REGFILE_SIM_reg_bank_reg_r24_5_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5256_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5456_));
NAND3X1 NAND3X1_209 ( .A(REGFILE_SIM_reg_bank_reg_r15_5_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5281_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5465_));
NAND3X1 NAND3X1_21 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1152_), .C(_abc_40298_new_n1170_), .Y(_abc_40298_new_n1171_));
NAND3X1 NAND3X1_210 ( .A(REGFILE_SIM_reg_bank_reg_r24_6_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5256_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5488_));
NAND3X1 NAND3X1_211 ( .A(REGFILE_SIM_reg_bank_reg_r15_6_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5281_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5497_));
NAND3X1 NAND3X1_212 ( .A(REGFILE_SIM_reg_bank_reg_r24_7_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5256_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5520_));
NAND3X1 NAND3X1_213 ( .A(REGFILE_SIM_reg_bank_reg_r15_7_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5281_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5529_));
NAND3X1 NAND3X1_214 ( .A(REGFILE_SIM_reg_bank_reg_r24_8_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5256_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5552_));
NAND3X1 NAND3X1_215 ( .A(REGFILE_SIM_reg_bank_reg_r15_8_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5281_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5561_));
NAND3X1 NAND3X1_216 ( .A(REGFILE_SIM_reg_bank_reg_r24_9_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5256_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5584_));
NAND3X1 NAND3X1_217 ( .A(REGFILE_SIM_reg_bank_reg_r15_9_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5281_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5593_));
NAND3X1 NAND3X1_218 ( .A(REGFILE_SIM_reg_bank_reg_r24_10_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5256_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5616_));
NAND3X1 NAND3X1_219 ( .A(REGFILE_SIM_reg_bank_reg_r15_10_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5281_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5625_));
NAND3X1 NAND3X1_22 ( .A(_abc_40298_new_n1045_), .B(_abc_40298_new_n1048_), .C(_abc_40298_new_n1182_), .Y(_abc_40298_new_n1183_));
NAND3X1 NAND3X1_220 ( .A(REGFILE_SIM_reg_bank_reg_r24_11_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5256_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5648_));
NAND3X1 NAND3X1_221 ( .A(REGFILE_SIM_reg_bank_reg_r15_11_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5281_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5657_));
NAND3X1 NAND3X1_222 ( .A(REGFILE_SIM_reg_bank_reg_r24_12_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5256_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5680_));
NAND3X1 NAND3X1_223 ( .A(REGFILE_SIM_reg_bank_reg_r15_12_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5281_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5689_));
NAND3X1 NAND3X1_224 ( .A(REGFILE_SIM_reg_bank_reg_r24_13_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5256_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5712_));
NAND3X1 NAND3X1_225 ( .A(REGFILE_SIM_reg_bank_reg_r15_13_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5281_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5721_));
NAND3X1 NAND3X1_226 ( .A(REGFILE_SIM_reg_bank_reg_r24_14_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5256_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5744_));
NAND3X1 NAND3X1_227 ( .A(REGFILE_SIM_reg_bank_reg_r15_14_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5281_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5753_));
NAND3X1 NAND3X1_228 ( .A(REGFILE_SIM_reg_bank_reg_r24_15_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5256_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5776_));
NAND3X1 NAND3X1_229 ( .A(REGFILE_SIM_reg_bank_reg_r15_15_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5281_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5785_));
NAND3X1 NAND3X1_23 ( .A(sr_q_9_), .B(_abc_40298_new_n617_), .C(_abc_40298_new_n652_), .Y(_abc_40298_new_n1212_));
NAND3X1 NAND3X1_230 ( .A(REGFILE_SIM_reg_bank_reg_r24_16_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5256_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5808_));
NAND3X1 NAND3X1_231 ( .A(REGFILE_SIM_reg_bank_reg_r15_16_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5281_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5817_));
NAND3X1 NAND3X1_232 ( .A(REGFILE_SIM_reg_bank_reg_r24_17_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5256_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5840_));
NAND3X1 NAND3X1_233 ( .A(REGFILE_SIM_reg_bank_reg_r15_17_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5281_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5849_));
NAND3X1 NAND3X1_234 ( .A(REGFILE_SIM_reg_bank_reg_r24_18_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5256_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5872_));
NAND3X1 NAND3X1_235 ( .A(REGFILE_SIM_reg_bank_reg_r15_18_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5281_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5881_));
NAND3X1 NAND3X1_236 ( .A(REGFILE_SIM_reg_bank_reg_r24_19_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5256_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5904_));
NAND3X1 NAND3X1_237 ( .A(REGFILE_SIM_reg_bank_reg_r15_19_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5281_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5913_));
NAND3X1 NAND3X1_238 ( .A(REGFILE_SIM_reg_bank_reg_r24_20_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5256_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5936_));
NAND3X1 NAND3X1_239 ( .A(REGFILE_SIM_reg_bank_reg_r15_20_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5281_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5945_));
NAND3X1 NAND3X1_24 ( .A(_abc_40298_new_n1235_), .B(_abc_40298_new_n1236_), .C(_abc_40298_new_n985_), .Y(_abc_40298_new_n1237_));
NAND3X1 NAND3X1_240 ( .A(REGFILE_SIM_reg_bank_reg_r24_21_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5256_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5968_));
NAND3X1 NAND3X1_241 ( .A(REGFILE_SIM_reg_bank_reg_r15_21_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5281_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5977_));
NAND3X1 NAND3X1_242 ( .A(REGFILE_SIM_reg_bank_reg_r24_22_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5256_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6000_));
NAND3X1 NAND3X1_243 ( .A(REGFILE_SIM_reg_bank_reg_r15_22_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5281_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6009_));
NAND3X1 NAND3X1_244 ( .A(REGFILE_SIM_reg_bank_reg_r24_23_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5256_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6032_));
NAND3X1 NAND3X1_245 ( .A(REGFILE_SIM_reg_bank_reg_r15_23_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5281_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6041_));
NAND3X1 NAND3X1_246 ( .A(REGFILE_SIM_reg_bank_reg_r24_24_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5256_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6064_));
NAND3X1 NAND3X1_247 ( .A(REGFILE_SIM_reg_bank_reg_r15_24_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5281_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6073_));
NAND3X1 NAND3X1_248 ( .A(REGFILE_SIM_reg_bank_reg_r24_25_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5256_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6096_));
NAND3X1 NAND3X1_249 ( .A(REGFILE_SIM_reg_bank_reg_r15_25_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5281_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6105_));
NAND3X1 NAND3X1_25 ( .A(pc_q_2_), .B(pc_q_3_), .C(pc_q_4_), .Y(_abc_40298_new_n1258_));
NAND3X1 NAND3X1_250 ( .A(REGFILE_SIM_reg_bank_reg_r24_26_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5256_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6128_));
NAND3X1 NAND3X1_251 ( .A(REGFILE_SIM_reg_bank_reg_r15_26_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5281_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6137_));
NAND3X1 NAND3X1_252 ( .A(REGFILE_SIM_reg_bank_reg_r24_27_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5256_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6160_));
NAND3X1 NAND3X1_253 ( .A(REGFILE_SIM_reg_bank_reg_r15_27_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5281_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6169_));
NAND3X1 NAND3X1_254 ( .A(REGFILE_SIM_reg_bank_reg_r24_28_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5256_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6192_));
NAND3X1 NAND3X1_255 ( .A(REGFILE_SIM_reg_bank_reg_r15_28_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5281_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6201_));
NAND3X1 NAND3X1_256 ( .A(REGFILE_SIM_reg_bank_reg_r24_29_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5256_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6224_));
NAND3X1 NAND3X1_257 ( .A(REGFILE_SIM_reg_bank_reg_r15_29_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5281_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6233_));
NAND3X1 NAND3X1_258 ( .A(REGFILE_SIM_reg_bank_reg_r24_30_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5256_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6256_));
NAND3X1 NAND3X1_259 ( .A(REGFILE_SIM_reg_bank_reg_r15_30_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5281_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6265_));
NAND3X1 NAND3X1_26 ( .A(pc_q_4_), .B(pc_q_5_), .C(_abc_40298_new_n1242_), .Y(_abc_40298_new_n1289_));
NAND3X1 NAND3X1_260 ( .A(REGFILE_SIM_reg_bank_reg_r24_31_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5254_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5256_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6288_));
NAND3X1 NAND3X1_261 ( .A(REGFILE_SIM_reg_bank_reg_r15_31_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5281_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6297_));
NAND3X1 NAND3X1_262 ( .A(alu__abc_38674_new_n225_), .B(alu__abc_38674_new_n230_), .C(alu__abc_38674_new_n241_), .Y(alu__abc_38674_new_n242_));
NAND3X1 NAND3X1_263 ( .A(alu__abc_38674_new_n257_), .B(alu__abc_38674_new_n274_), .C(alu__abc_38674_new_n244_), .Y(alu__abc_38674_new_n275_));
NAND3X1 NAND3X1_264 ( .A(alu__abc_38674_new_n134_), .B(alu_a_i_16_), .C(alu__abc_38674_new_n141_), .Y(alu__abc_38674_new_n309_));
NAND3X1 NAND3X1_265 ( .A(alu__abc_38674_new_n307_), .B(alu__abc_38674_new_n150_), .C(alu__abc_38674_new_n310_), .Y(alu__abc_38674_new_n311_));
NAND3X1 NAND3X1_266 ( .A(alu__abc_38674_new_n232_), .B(alu_a_i_10_), .C(alu__abc_38674_new_n239_), .Y(alu__abc_38674_new_n357_));
NAND3X1 NAND3X1_267 ( .A(alu__abc_38674_new_n268_), .B(alu__abc_38674_new_n271_), .C(alu__abc_38674_new_n421_), .Y(alu__abc_38674_new_n422_));
NAND3X1 NAND3X1_268 ( .A(alu__abc_38674_new_n412_), .B(alu__abc_38674_new_n467_), .C(alu__abc_38674_new_n464_), .Y(alu__abc_38674_new_n468_));
NAND3X1 NAND3X1_269 ( .A(alu__abc_38674_new_n418_), .B(alu__abc_38674_new_n419_), .C(alu__abc_38674_new_n468_), .Y(alu__abc_38674_new_n469_));
NAND3X1 NAND3X1_27 ( .A(pc_q_7_), .B(pc_q_8_), .C(_abc_40298_new_n1304_), .Y(_abc_40298_new_n1364_));
NAND3X1 NAND3X1_270 ( .A(alu__abc_38674_new_n385_), .B(alu__abc_38674_new_n391_), .C(alu__abc_38674_new_n398_), .Y(alu__abc_38674_new_n476_));
NAND3X1 NAND3X1_271 ( .A(alu__abc_38674_new_n490_), .B(alu__abc_38674_new_n497_), .C(alu__abc_38674_new_n499_), .Y(alu__abc_38674_new_n500_));
NAND3X1 NAND3X1_272 ( .A(alu__abc_38674_new_n229_), .B(alu__abc_38674_new_n444_), .C(alu__abc_38674_new_n459_), .Y(alu__abc_38674_new_n514_));
NAND3X1 NAND3X1_273 ( .A(alu__abc_38674_new_n512_), .B(alu__abc_38674_new_n208_), .C(alu__abc_38674_new_n527_), .Y(alu__abc_38674_new_n528_));
NAND3X1 NAND3X1_274 ( .A(alu__abc_38674_new_n247_), .B(alu__abc_38674_new_n438_), .C(alu__abc_38674_new_n545_), .Y(alu__abc_38674_new_n546_));
NAND3X1 NAND3X1_275 ( .A(alu__abc_38674_new_n253_), .B(alu__abc_38674_new_n436_), .C(alu__abc_38674_new_n548_), .Y(alu__abc_38674_new_n549_));
NAND3X1 NAND3X1_276 ( .A(alu_c_i), .B(alu__abc_38674_new_n420_), .C(alu__abc_38674_new_n563_), .Y(alu__abc_38674_new_n564_));
NAND3X1 NAND3X1_277 ( .A(alu__abc_38674_new_n558_), .B(alu__abc_38674_new_n570_), .C(alu__abc_38674_new_n571_), .Y(alu__abc_38674_new_n572_));
NAND3X1 NAND3X1_278 ( .A(alu__abc_38674_new_n540_), .B(alu__abc_38674_new_n544_), .C(alu__abc_38674_new_n573_), .Y(alu__abc_38674_new_n574_));
NAND3X1 NAND3X1_279 ( .A(alu__abc_38674_new_n578_), .B(alu__abc_38674_new_n579_), .C(alu__abc_38674_new_n580_), .Y(alu__abc_38674_new_n581_));
NAND3X1 NAND3X1_28 ( .A(pc_q_8_), .B(pc_q_9_), .C(_abc_40298_new_n1333_), .Y(_abc_40298_new_n1448_));
NAND3X1 NAND3X1_280 ( .A(alu__abc_38674_new_n231_), .B(alu__abc_38674_new_n239_), .C(alu__abc_38674_new_n587_), .Y(alu__abc_38674_new_n588_));
NAND3X1 NAND3X1_281 ( .A(alu__abc_38674_new_n235_), .B(alu__abc_38674_new_n445_), .C(alu__abc_38674_new_n589_), .Y(alu__abc_38674_new_n593_));
NAND3X1 NAND3X1_282 ( .A(alu__abc_38674_new_n535_), .B(alu__abc_38674_new_n577_), .C(alu__abc_38674_new_n597_), .Y(alu__abc_38674_new_n598_));
NAND3X1 NAND3X1_283 ( .A(alu__abc_38674_new_n599_), .B(alu__abc_38674_new_n600_), .C(alu__abc_38674_new_n603_), .Y(alu__abc_38674_new_n604_));
NAND3X1 NAND3X1_284 ( .A(alu__abc_38674_new_n483_), .B(alu__abc_38674_new_n484_), .C(alu__abc_38674_new_n608_), .Y(alu__abc_38674_new_n609_));
NAND3X1 NAND3X1_285 ( .A(alu__abc_38674_new_n615_), .B(alu__abc_38674_new_n616_), .C(alu__abc_38674_new_n625_), .Y(alu__abc_38674_new_n626_));
NAND3X1 NAND3X1_286 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n563_), .C(alu__abc_38674_new_n645_), .Y(alu__abc_38674_new_n646_));
NAND3X1 NAND3X1_287 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n338_), .C(alu__abc_38674_new_n696_), .Y(alu__abc_38674_new_n697_));
NAND3X1 NAND3X1_288 ( .A(alu__abc_38674_new_n694_), .B(alu__abc_38674_new_n715_), .C(alu__abc_38674_new_n691_), .Y(alu_p_o_0_));
NAND3X1 NAND3X1_289 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n559_), .C(alu__abc_38674_new_n778_), .Y(alu__abc_38674_new_n779_));
NAND3X1 NAND3X1_29 ( .A(pc_q_11_), .B(pc_q_12_), .C(_abc_40298_new_n1416_), .Y(_abc_40298_new_n1475_));
NAND3X1 NAND3X1_290 ( .A(alu__abc_38674_new_n781_), .B(alu__abc_38674_new_n794_), .C(alu__abc_38674_new_n792_), .Y(alu__abc_38674_new_n795_));
NAND3X1 NAND3X1_291 ( .A(alu__abc_38674_new_n836_), .B(alu__abc_38674_new_n847_), .C(alu__abc_38674_new_n842_), .Y(alu__abc_38674_new_n848_));
NAND3X1 NAND3X1_292 ( .A(alu__abc_38674_new_n880_), .B(alu__abc_38674_new_n882_), .C(alu__abc_38674_new_n900_), .Y(alu_p_o_3_));
NAND3X1 NAND3X1_293 ( .A(alu__abc_38674_new_n381_), .B(alu__abc_38674_new_n572_), .C(alu__abc_38674_new_n904_), .Y(alu__abc_38674_new_n905_));
NAND3X1 NAND3X1_294 ( .A(alu__abc_38674_new_n905_), .B(alu__abc_38674_new_n907_), .C(alu__abc_38674_new_n939_), .Y(alu_p_o_4_));
NAND3X1 NAND3X1_295 ( .A(alu__abc_38674_new_n706_), .B(alu__abc_38674_new_n973_), .C(alu__abc_38674_new_n347_), .Y(alu__abc_38674_new_n974_));
NAND3X1 NAND3X1_296 ( .A(alu__abc_38674_new_n971_), .B(alu__abc_38674_new_n974_), .C(alu__abc_38674_new_n966_), .Y(alu_p_o_5_));
NAND3X1 NAND3X1_297 ( .A(alu__abc_38674_new_n978_), .B(alu__abc_38674_new_n981_), .C(alu__abc_38674_new_n1005_), .Y(alu_p_o_6_));
NAND3X1 NAND3X1_298 ( .A(alu__abc_38674_new_n1012_), .B(alu__abc_38674_new_n1039_), .C(alu__abc_38674_new_n1010_), .Y(alu_p_o_7_));
NAND3X1 NAND3X1_299 ( .A(alu__abc_38674_new_n245_), .B(alu__abc_38674_new_n517_), .C(alu__abc_38674_new_n542_), .Y(alu__abc_38674_new_n1044_));
NAND3X1 NAND3X1_3 ( .A(_abc_40298_new_n730_), .B(_abc_40298_new_n731_), .C(_abc_40298_new_n729_), .Y(_abc_40298_new_n732_));
NAND3X1 NAND3X1_30 ( .A(pc_q_12_), .B(pc_q_13_), .C(_abc_40298_new_n1449_), .Y(_abc_40298_new_n1562_));
NAND3X1 NAND3X1_300 ( .A(alu__abc_38674_new_n979_), .B(alu__abc_38674_new_n968_), .C(alu__abc_38674_new_n967_), .Y(alu__abc_38674_new_n1047_));
NAND3X1 NAND3X1_301 ( .A(alu__abc_38674_new_n381_), .B(alu__abc_38674_new_n574_), .C(alu__abc_38674_new_n1048_), .Y(alu__abc_38674_new_n1049_));
NAND3X1 NAND3X1_302 ( .A(alu__abc_38674_new_n1068_), .B(alu__abc_38674_new_n1071_), .C(alu__abc_38674_new_n1056_), .Y(alu__abc_38674_new_n1072_));
NAND3X1 NAND3X1_303 ( .A(alu__abc_38674_new_n1042_), .B(alu__abc_38674_new_n1049_), .C(alu__abc_38674_new_n1073_), .Y(alu_p_o_8_));
NAND3X1 NAND3X1_304 ( .A(alu__abc_38674_new_n1115_), .B(alu__abc_38674_new_n1135_), .C(alu__abc_38674_new_n1111_), .Y(alu_p_o_10_));
NAND3X1 NAND3X1_305 ( .A(alu__abc_38674_new_n231_), .B(alu__abc_38674_new_n240_), .C(alu__abc_38674_new_n587_), .Y(alu__abc_38674_new_n1143_));
NAND3X1 NAND3X1_306 ( .A(alu__abc_38674_new_n1142_), .B(alu__abc_38674_new_n1169_), .C(alu__abc_38674_new_n1140_), .Y(alu_p_o_11_));
NAND3X1 NAND3X1_307 ( .A(alu__abc_38674_new_n1173_), .B(alu__abc_38674_new_n1198_), .C(alu__abc_38674_new_n1179_), .Y(alu_p_o_12_));
NAND3X1 NAND3X1_308 ( .A(alu__abc_38674_new_n578_), .B(alu__abc_38674_new_n451_), .C(alu__abc_38674_new_n580_), .Y(alu__abc_38674_new_n1201_));
NAND3X1 NAND3X1_309 ( .A(alu__abc_38674_new_n451_), .B(alu__abc_38674_new_n1209_), .C(alu__abc_38674_new_n1207_), .Y(alu__abc_38674_new_n1210_));
NAND3X1 NAND3X1_31 ( .A(_abc_40298_new_n1544_), .B(_abc_40298_new_n1574_), .C(_abc_40298_new_n1547_), .Y(_abc_40298_new_n1575_));
NAND3X1 NAND3X1_310 ( .A(alu__abc_38674_new_n362_), .B(alu__abc_38674_new_n706_), .C(alu__abc_38674_new_n1210_), .Y(alu__abc_38674_new_n1211_));
NAND3X1 NAND3X1_311 ( .A(alu__abc_38674_new_n706_), .B(alu__abc_38674_new_n1236_), .C(alu__abc_38674_new_n1235_), .Y(alu__abc_38674_new_n1237_));
NAND3X1 NAND3X1_312 ( .A(alu__abc_38674_new_n1237_), .B(alu__abc_38674_new_n1261_), .C(alu__abc_38674_new_n1239_), .Y(alu_p_o_14_));
NAND3X1 NAND3X1_313 ( .A(alu__abc_38674_new_n1145_), .B(alu__abc_38674_new_n1240_), .C(alu__abc_38674_new_n1268_), .Y(alu__abc_38674_new_n1269_));
NAND3X1 NAND3X1_314 ( .A(alu__abc_38674_new_n1288_), .B(alu__abc_38674_new_n1290_), .C(alu__abc_38674_new_n1287_), .Y(alu__abc_38674_new_n1291_));
NAND3X1 NAND3X1_315 ( .A(alu__abc_38674_new_n1292_), .B(alu__abc_38674_new_n1265_), .C(alu__abc_38674_new_n1272_), .Y(alu_p_o_15_));
NAND3X1 NAND3X1_316 ( .A(alu__abc_38674_new_n537_), .B(alu__abc_38674_new_n1240_), .C(alu__abc_38674_new_n1076_), .Y(alu__abc_38674_new_n1294_));
NAND3X1 NAND3X1_317 ( .A(alu__abc_38674_new_n1295_), .B(alu__abc_38674_new_n1203_), .C(alu__abc_38674_new_n1145_), .Y(alu__abc_38674_new_n1296_));
NAND3X1 NAND3X1_318 ( .A(alu__abc_38674_new_n1303_), .B(alu__abc_38674_new_n1325_), .C(alu__abc_38674_new_n1300_), .Y(alu_p_o_16_));
NAND3X1 NAND3X1_319 ( .A(alu__abc_38674_new_n1340_), .B(alu__abc_38674_new_n1356_), .C(alu__abc_38674_new_n1333_), .Y(alu_p_o_17_));
NAND3X1 NAND3X1_32 ( .A(_abc_40298_new_n985_), .B(_abc_40298_new_n1575_), .C(_abc_40298_new_n1576_), .Y(_abc_40298_new_n1577_));
NAND3X1 NAND3X1_320 ( .A(alu__abc_38674_new_n1365_), .B(alu__abc_38674_new_n1382_), .C(alu__abc_38674_new_n1362_), .Y(alu_p_o_18_));
NAND3X1 NAND3X1_321 ( .A(alu__abc_38674_new_n381_), .B(alu__abc_38674_new_n1386_), .C(alu__abc_38674_new_n1385_), .Y(alu__abc_38674_new_n1387_));
NAND3X1 NAND3X1_322 ( .A(alu__abc_38674_new_n1388_), .B(alu__abc_38674_new_n1400_), .C(alu__abc_38674_new_n1387_), .Y(alu__abc_38674_new_n1401_));
NAND3X1 NAND3X1_323 ( .A(alu__abc_38674_new_n1406_), .B(alu__abc_38674_new_n1407_), .C(alu__abc_38674_new_n1405_), .Y(alu__abc_38674_new_n1408_));
NAND3X1 NAND3X1_324 ( .A(alu__abc_38674_new_n510_), .B(alu__abc_38674_new_n577_), .C(alu__abc_38674_new_n1415_), .Y(alu__abc_38674_new_n1416_));
NAND3X1 NAND3X1_325 ( .A(alu__abc_38674_new_n1424_), .B(alu__abc_38674_new_n1440_), .C(alu__abc_38674_new_n1419_), .Y(alu_p_o_20_));
NAND3X1 NAND3X1_326 ( .A(alu__abc_38674_new_n510_), .B(alu__abc_38674_new_n1442_), .C(alu__abc_38674_new_n1297_), .Y(alu__abc_38674_new_n1443_));
NAND3X1 NAND3X1_327 ( .A(alu__abc_38674_new_n490_), .B(alu__abc_38674_new_n497_), .C(alu__abc_38674_new_n605_), .Y(alu__abc_38674_new_n1472_));
NAND3X1 NAND3X1_328 ( .A(alu__abc_38674_new_n1491_), .B(alu__abc_38674_new_n1493_), .C(alu__abc_38674_new_n1490_), .Y(alu__abc_38674_new_n1494_));
NAND3X1 NAND3X1_329 ( .A(alu__abc_38674_new_n497_), .B(alu__abc_38674_new_n623_), .C(alu__abc_38674_new_n1417_), .Y(alu__abc_38674_new_n1500_));
NAND3X1 NAND3X1_33 ( .A(pc_q_15_), .B(pc_q_16_), .C(_abc_40298_new_n1534_), .Y(_abc_40298_new_n1589_));
NAND3X1 NAND3X1_330 ( .A(alu__abc_38674_new_n1531_), .B(alu__abc_38674_new_n1545_), .C(alu__abc_38674_new_n1527_), .Y(alu_p_o_24_));
NAND3X1 NAND3X1_331 ( .A(alu__abc_38674_new_n297_), .B(alu__abc_38674_new_n706_), .C(alu__abc_38674_new_n1561_), .Y(alu__abc_38674_new_n1562_));
NAND3X1 NAND3X1_332 ( .A(alu__abc_38674_new_n1557_), .B(alu__abc_38674_new_n1570_), .C(alu__abc_38674_new_n1549_), .Y(alu_p_o_25_));
NAND3X1 NAND3X1_333 ( .A(alu__abc_38674_new_n508_), .B(alu__abc_38674_new_n623_), .C(alu__abc_38674_new_n1574_), .Y(alu__abc_38674_new_n1575_));
NAND3X1 NAND3X1_334 ( .A(alu__abc_38674_new_n1593_), .B(alu__abc_38674_new_n1597_), .C(alu__abc_38674_new_n1594_), .Y(alu__abc_38674_new_n1598_));
NAND3X1 NAND3X1_335 ( .A(alu__abc_38674_new_n1582_), .B(alu__abc_38674_new_n1599_), .C(alu__abc_38674_new_n1578_), .Y(alu_p_o_26_));
NAND3X1 NAND3X1_336 ( .A(alu__abc_38674_new_n503_), .B(alu__abc_38674_new_n499_), .C(alu__abc_38674_new_n1525_), .Y(alu__abc_38674_new_n1602_));
NAND3X1 NAND3X1_337 ( .A(alu__abc_38674_new_n1629_), .B(alu__abc_38674_new_n706_), .C(alu__abc_38674_new_n1630_), .Y(alu__abc_38674_new_n1631_));
NAND3X1 NAND3X1_338 ( .A(alu__abc_38674_new_n1628_), .B(alu__abc_38674_new_n1645_), .C(alu__abc_38674_new_n1631_), .Y(alu__abc_38674_new_n1646_));
NAND3X1 NAND3X1_339 ( .A(alu__abc_38674_new_n484_), .B(alu__abc_38674_new_n619_), .C(alu__abc_38674_new_n1576_), .Y(alu__abc_38674_new_n1650_));
NAND3X1 NAND3X1_34 ( .A(pc_q_16_), .B(pc_q_17_), .C(_abc_40298_new_n1564_), .Y(_abc_40298_new_n1622_));
NAND3X1 NAND3X1_340 ( .A(alu__abc_38674_new_n1662_), .B(alu__abc_38674_new_n1667_), .C(alu__abc_38674_new_n1654_), .Y(alu__abc_38674_new_n1668_));
NAND3X1 NAND3X1_341 ( .A(alu__abc_38674_new_n616_), .B(alu__abc_38674_new_n483_), .C(alu__abc_38674_new_n1625_), .Y(alu__abc_38674_new_n1673_));
NAND3X1 NAND3X1_342 ( .A(alu__abc_38674_new_n381_), .B(alu__abc_38674_new_n1672_), .C(alu__abc_38674_new_n1673_), .Y(alu__abc_38674_new_n1674_));
NAND3X1 NAND3X1_343 ( .A(alu__abc_38674_new_n1678_), .B(alu__abc_38674_new_n1691_), .C(alu__abc_38674_new_n1677_), .Y(alu__abc_38674_new_n1692_));
NAND3X1 NAND3X1_344 ( .A(alu__abc_38674_new_n619_), .B(alu__abc_38674_new_n499_), .C(alu__abc_38674_new_n1547_), .Y(alu__abc_38674_new_n1695_));
NAND3X1 NAND3X1_345 ( .A(alu__abc_38674_new_n162_), .B(alu__abc_38674_new_n1700_), .C(alu__abc_38674_new_n377_), .Y(alu__abc_38674_new_n1701_));
NAND3X1 NAND3X1_346 ( .A(alu__abc_38674_new_n1725_), .B(alu__abc_38674_new_n1729_), .C(alu__abc_38674_new_n1724_), .Y(alu__abc_38674_new_n1730_));
NAND3X1 NAND3X1_35 ( .A(pc_q_19_), .B(pc_q_20_), .C(_abc_40298_new_n1646_), .Y(_abc_40298_new_n1699_));
NAND3X1 NAND3X1_36 ( .A(pc_q_20_), .B(pc_q_21_), .C(_abc_40298_new_n1676_), .Y(_abc_40298_new_n1728_));
NAND3X1 NAND3X1_37 ( .A(pc_q_23_), .B(pc_q_24_), .C(_abc_40298_new_n1755_), .Y(_abc_40298_new_n1807_));
NAND3X1 NAND3X1_38 ( .A(pc_q_27_), .B(pc_q_28_), .C(_abc_40298_new_n1864_), .Y(_abc_40298_new_n1913_));
NAND3X1 NAND3X1_39 ( .A(_abc_40298_new_n1213_), .B(_abc_40298_new_n1951_), .C(_abc_40298_new_n1949_), .Y(_abc_40298_new_n1952_));
NAND3X1 NAND3X1_4 ( .A(_abc_40298_new_n739_), .B(_abc_40298_new_n740_), .C(_abc_40298_new_n738_), .Y(_abc_40298_new_n741_));
NAND3X1 NAND3X1_40 ( .A(_abc_40298_new_n1232_), .B(_abc_40298_new_n1962_), .C(_abc_40298_new_n1964_), .Y(_abc_40298_new_n1982_));
NAND3X1 NAND3X1_41 ( .A(_abc_40298_new_n1213_), .B(_abc_40298_new_n1997_), .C(_abc_40298_new_n1995_), .Y(_abc_40298_new_n1998_));
NAND3X1 NAND3X1_42 ( .A(pc_q_24_), .B(pc_q_25_), .C(_abc_40298_new_n1784_), .Y(_abc_40298_new_n2000_));
NAND3X1 NAND3X1_43 ( .A(pc_q_28_), .B(pc_q_29_), .C(_abc_40298_new_n2001_), .Y(_abc_40298_new_n2002_));
NAND3X1 NAND3X1_44 ( .A(pc_q_30_), .B(pc_q_31_), .C(_abc_40298_new_n1963_), .Y(_abc_40298_new_n2004_));
NAND3X1 NAND3X1_45 ( .A(_abc_40298_new_n1232_), .B(_abc_40298_new_n2004_), .C(_abc_40298_new_n2003_), .Y(_abc_40298_new_n2005_));
NAND3X1 NAND3X1_46 ( .A(_abc_40298_new_n1134_), .B(_abc_40298_new_n1998_), .C(_abc_40298_new_n2005_), .Y(_abc_40298_new_n2006_));
NAND3X1 NAND3X1_47 ( .A(_abc_40298_new_n977_), .B(_abc_40298_new_n982_), .C(_abc_40298_new_n928_), .Y(_abc_40298_new_n2119_));
NAND3X1 NAND3X1_48 ( .A(_abc_40298_new_n1080_), .B(_abc_40298_new_n1185_), .C(_abc_40298_new_n1061_), .Y(_abc_40298_new_n2121_));
NAND3X1 NAND3X1_49 ( .A(_abc_40298_new_n2125_), .B(_abc_40298_new_n2123_), .C(_abc_40298_new_n897_), .Y(_abc_40298_new_n2126_));
NAND3X1 NAND3X1_5 ( .A(_abc_40298_new_n897_), .B(_abc_40298_new_n899_), .C(_abc_40298_new_n895_), .Y(_abc_40298_new_n900_));
NAND3X1 NAND3X1_50 ( .A(_abc_40298_new_n2126_), .B(_abc_40298_new_n962_), .C(_abc_40298_new_n2127_), .Y(_abc_40298_new_n2128_));
NAND3X1 NAND3X1_51 ( .A(_abc_40298_new_n2143_), .B(_abc_40298_new_n2144_), .C(_abc_40298_new_n2141_), .Y(_abc_40298_new_n2145_));
NAND3X1 NAND3X1_52 ( .A(_abc_40298_new_n892_), .B(_abc_40298_new_n924_), .C(_abc_40298_new_n897_), .Y(_abc_40298_new_n2173_));
NAND3X1 NAND3X1_53 ( .A(_abc_40298_new_n2355_), .B(_abc_40298_new_n2356_), .C(_abc_40298_new_n2354_), .Y(alu_input_a_r_9_));
NAND3X1 NAND3X1_54 ( .A(epc_q_13_), .B(_abc_40298_new_n1001_), .C(_abc_40298_new_n1186_), .Y(_abc_40298_new_n2373_));
NAND3X1 NAND3X1_55 ( .A(epc_q_14_), .B(_abc_40298_new_n1001_), .C(_abc_40298_new_n1186_), .Y(_abc_40298_new_n2377_));
NAND3X1 NAND3X1_56 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_16_), .B(_abc_40298_new_n1014_), .C(_abc_40298_new_n2286_), .Y(_abc_40298_new_n2386_));
NAND3X1 NAND3X1_57 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_17_), .B(_abc_40298_new_n1014_), .C(_abc_40298_new_n2286_), .Y(_abc_40298_new_n2393_));
NAND3X1 NAND3X1_58 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_18_), .B(_abc_40298_new_n1014_), .C(_abc_40298_new_n2286_), .Y(_abc_40298_new_n2400_));
NAND3X1 NAND3X1_59 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_19_), .B(_abc_40298_new_n1014_), .C(_abc_40298_new_n2286_), .Y(_abc_40298_new_n2407_));
NAND3X1 NAND3X1_6 ( .A(_abc_40298_new_n897_), .B(_abc_40298_new_n901_), .C(_abc_40298_new_n895_), .Y(_abc_40298_new_n902_));
NAND3X1 NAND3X1_60 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_20_), .B(_abc_40298_new_n1014_), .C(_abc_40298_new_n2286_), .Y(_abc_40298_new_n2414_));
NAND3X1 NAND3X1_61 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_21_), .B(_abc_40298_new_n1014_), .C(_abc_40298_new_n2286_), .Y(_abc_40298_new_n2421_));
NAND3X1 NAND3X1_62 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_22_), .B(_abc_40298_new_n1014_), .C(_abc_40298_new_n2286_), .Y(_abc_40298_new_n2428_));
NAND3X1 NAND3X1_63 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_23_), .B(_abc_40298_new_n1014_), .C(_abc_40298_new_n2286_), .Y(_abc_40298_new_n2435_));
NAND3X1 NAND3X1_64 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_24_), .B(_abc_40298_new_n1014_), .C(_abc_40298_new_n2286_), .Y(_abc_40298_new_n2442_));
NAND3X1 NAND3X1_65 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_25_), .B(_abc_40298_new_n1014_), .C(_abc_40298_new_n2286_), .Y(_abc_40298_new_n2449_));
NAND3X1 NAND3X1_66 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_26_), .B(_abc_40298_new_n1014_), .C(_abc_40298_new_n2286_), .Y(_abc_40298_new_n2457_));
NAND3X1 NAND3X1_67 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_27_), .B(_abc_40298_new_n1014_), .C(_abc_40298_new_n2286_), .Y(_abc_40298_new_n2464_));
NAND3X1 NAND3X1_68 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_28_), .B(_abc_40298_new_n1014_), .C(_abc_40298_new_n2286_), .Y(_abc_40298_new_n2472_));
NAND3X1 NAND3X1_69 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_29_), .B(_abc_40298_new_n1014_), .C(_abc_40298_new_n2286_), .Y(_abc_40298_new_n2480_));
NAND3X1 NAND3X1_7 ( .A(_abc_40298_new_n900_), .B(_abc_40298_new_n902_), .C(_abc_40298_new_n915_), .Y(_abc_40298_new_n916_));
NAND3X1 NAND3X1_70 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_30_), .B(_abc_40298_new_n1014_), .C(_abc_40298_new_n2286_), .Y(_abc_40298_new_n2487_));
NAND3X1 NAND3X1_71 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_31_), .B(_abc_40298_new_n1014_), .C(_abc_40298_new_n2286_), .Y(_abc_40298_new_n2494_));
NAND3X1 NAND3X1_72 ( .A(_abc_40298_new_n2501_), .B(_abc_40298_new_n2502_), .C(_abc_40298_new_n2503_), .Y(alu_func_r_0_));
NAND3X1 NAND3X1_73 ( .A(_abc_40298_new_n2506_), .B(_abc_40298_new_n2507_), .C(_abc_40298_new_n2505_), .Y(alu_func_r_1_));
NAND3X1 NAND3X1_74 ( .A(_abc_40298_new_n982_), .B(_abc_40298_new_n2173_), .C(_abc_40298_new_n2171_), .Y(alu_func_r_2_));
NAND3X1 NAND3X1_75 ( .A(_abc_40298_new_n900_), .B(_abc_40298_new_n2510_), .C(_abc_40298_new_n2511_), .Y(alu_func_r_3_));
NAND3X1 NAND3X1_76 ( .A(_abc_40298_new_n2906_), .B(_abc_40298_new_n2908_), .C(_abc_40298_new_n2902_), .Y(_abc_40298_new_n2909_));
NAND3X1 NAND3X1_77 ( .A(_abc_40298_new_n2901_), .B(_abc_40298_new_n2909_), .C(_abc_40298_new_n2900_), .Y(_0mem_addr_o_31_0__2_));
NAND3X1 NAND3X1_78 ( .A(_abc_40298_new_n2955_), .B(_abc_40298_new_n2956_), .C(_abc_40298_new_n2954_), .Y(_0mem_addr_o_31_0__7_));
NAND3X1 NAND3X1_79 ( .A(_abc_40298_new_n3010_), .B(_abc_40298_new_n3015_), .C(_abc_40298_new_n3006_), .Y(_abc_40298_new_n3016_));
NAND3X1 NAND3X1_8 ( .A(inst_r_2_), .B(inst_r_3_), .C(_abc_40298_new_n644_), .Y(_abc_40298_new_n929_));
NAND3X1 NAND3X1_80 ( .A(_abc_40298_new_n3013_), .B(_abc_40298_new_n3014_), .C(_abc_40298_new_n3017_), .Y(_abc_40298_new_n3018_));
NAND3X1 NAND3X1_81 ( .A(_abc_40298_new_n2902_), .B(_abc_40298_new_n3018_), .C(_abc_40298_new_n3016_), .Y(_abc_40298_new_n3019_));
NAND3X1 NAND3X1_82 ( .A(_abc_40298_new_n3020_), .B(_abc_40298_new_n3021_), .C(_abc_40298_new_n3019_), .Y(_0mem_addr_o_31_0__13_));
NAND3X1 NAND3X1_83 ( .A(_abc_40298_new_n3152_), .B(_abc_40298_new_n3153_), .C(_abc_40298_new_n3151_), .Y(_0mem_addr_o_31_0__26_));
NAND3X1 NAND3X1_84 ( .A(REGFILE_SIM_reg_bank_rb_i_4_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4179_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4177_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4180_));
NAND3X1 NAND3X1_85 ( .A(REGFILE_SIM_reg_bank_reg_r24_0_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4184_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4185_));
NAND3X1 NAND3X1_86 ( .A(REGFILE_SIM_reg_bank_rb_i_4_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4177_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4187_));
NAND3X1 NAND3X1_87 ( .A(REGFILE_SIM_reg_bank_rb_i_4_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4189_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4190_));
NAND3X1 NAND3X1_88 ( .A(REGFILE_SIM_reg_bank_rb_i_4_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4177_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4194_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4195_));
NAND3X1 NAND3X1_89 ( .A(REGFILE_SIM_reg_bank_rb_i_4_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4197_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4194_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4198_));
NAND3X1 NAND3X1_9 ( .A(_abc_40298_new_n934_), .B(_abc_40298_new_n941_), .C(_abc_40298_new_n933_), .Y(_abc_40298_new_n942_));
NAND3X1 NAND3X1_90 ( .A(REGFILE_SIM_reg_bank_rb_i_4_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4200_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4177_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4201_));
NAND3X1 NAND3X1_91 ( .A(REGFILE_SIM_reg_bank_rb_i_4_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4200_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4189_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4202_));
NAND3X1 NAND3X1_92 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4189_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4206_));
NAND3X1 NAND3X1_93 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4197_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4207_));
NAND3X1 NAND3X1_94 ( .A(REGFILE_SIM_reg_bank_reg_r15_0_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4209_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4210_));
NAND3X1 NAND3X1_95 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4179_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4189_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4211_));
NAND3X1 NAND3X1_96 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4200_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4177_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4214_));
NAND3X1 NAND3X1_97 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4189_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4194_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4218_));
NAND3X1 NAND3X1_98 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4177_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4194_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4219_));
NAND3X1 NAND3X1_99 ( .A(REGFILE_SIM_reg_bank_rb_i_4_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4197_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4182_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4224_));
NOR2X1 NOR2X1_1 ( .A(inst_r_4_), .B(inst_r_5_), .Y(_abc_40298_new_n617_));
NOR2X1 NOR2X1_10 ( .A(_abc_40298_new_n646_), .B(_abc_40298_new_n648_), .Y(_abc_40298_new_n649_));
NOR2X1 NOR2X1_100 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_3_), .B(alu_op_r_3_), .Y(_abc_40298_new_n1055_));
NOR2X1 NOR2X1_1000 ( .A(alu_b_i_23_), .B(alu_a_i_23_), .Y(alu__abc_38674_new_n119_));
NOR2X1 NOR2X1_1001 ( .A(alu__abc_38674_new_n121_), .B(alu__abc_38674_new_n122_), .Y(alu__abc_38674_new_n123_));
NOR2X1 NOR2X1_1002 ( .A(alu_b_i_20_), .B(alu_a_i_20_), .Y(alu__abc_38674_new_n124_));
NOR2X1 NOR2X1_1003 ( .A(alu__abc_38674_new_n124_), .B(alu__abc_38674_new_n123_), .Y(alu__abc_38674_new_n125_));
NOR2X1 NOR2X1_1004 ( .A(alu__abc_38674_new_n127_), .B(alu__abc_38674_new_n128_), .Y(alu__abc_38674_new_n129_));
NOR2X1 NOR2X1_1005 ( .A(alu_b_i_21_), .B(alu_a_i_21_), .Y(alu__abc_38674_new_n130_));
NOR2X1 NOR2X1_1006 ( .A(alu__abc_38674_new_n120_), .B(alu__abc_38674_new_n131_), .Y(alu__abc_38674_new_n132_));
NOR2X1 NOR2X1_1007 ( .A(alu__abc_38674_new_n134_), .B(alu__abc_38674_new_n135_), .Y(alu__abc_38674_new_n136_));
NOR2X1 NOR2X1_1008 ( .A(alu_b_i_16_), .B(alu_a_i_16_), .Y(alu__abc_38674_new_n137_));
NOR2X1 NOR2X1_1009 ( .A(alu_b_i_17_), .B(alu_a_i_17_), .Y(alu__abc_38674_new_n139_));
NOR2X1 NOR2X1_101 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_2_), .B(alu_op_r_2_), .Y(_abc_40298_new_n1056_));
NOR2X1 NOR2X1_1010 ( .A(alu__abc_38674_new_n139_), .B(alu__abc_38674_new_n138_), .Y(alu__abc_38674_new_n140_));
NOR2X1 NOR2X1_1011 ( .A(alu__abc_38674_new_n143_), .B(alu__abc_38674_new_n144_), .Y(alu__abc_38674_new_n145_));
NOR2X1 NOR2X1_1012 ( .A(alu_b_i_18_), .B(alu_a_i_18_), .Y(alu__abc_38674_new_n146_));
NOR2X1 NOR2X1_1013 ( .A(alu_b_i_19_), .B(alu_a_i_19_), .Y(alu__abc_38674_new_n148_));
NOR2X1 NOR2X1_1014 ( .A(alu__abc_38674_new_n148_), .B(alu__abc_38674_new_n147_), .Y(alu__abc_38674_new_n149_));
NOR2X1 NOR2X1_1015 ( .A(alu__abc_38674_new_n142_), .B(alu__abc_38674_new_n151_), .Y(alu__abc_38674_new_n152_));
NOR2X1 NOR2X1_1016 ( .A(alu__abc_38674_new_n153_), .B(alu__abc_38674_new_n133_), .Y(alu__abc_38674_new_n154_));
NOR2X1 NOR2X1_1017 ( .A(alu__abc_38674_new_n155_), .B(alu__abc_38674_new_n156_), .Y(alu__abc_38674_new_n157_));
NOR2X1 NOR2X1_1018 ( .A(alu_b_i_30_), .B(alu_a_i_30_), .Y(alu__abc_38674_new_n158_));
NOR2X1 NOR2X1_1019 ( .A(alu__abc_38674_new_n158_), .B(alu__abc_38674_new_n157_), .Y(alu__abc_38674_new_n159_));
NOR2X1 NOR2X1_102 ( .A(_abc_40298_new_n1054_), .B(_abc_40298_new_n1057_), .Y(_abc_40298_new_n1058_));
NOR2X1 NOR2X1_1020 ( .A(alu_b_i_31_), .B(alu_a_i_31_), .Y(alu__abc_38674_new_n161_));
NOR2X1 NOR2X1_1021 ( .A(alu__abc_38674_new_n161_), .B(alu__abc_38674_new_n160_), .Y(alu__abc_38674_new_n162_));
NOR2X1 NOR2X1_1022 ( .A(alu__abc_38674_new_n162_), .B(alu__abc_38674_new_n159_), .Y(alu__abc_38674_new_n163_));
NOR2X1 NOR2X1_1023 ( .A(alu__abc_38674_new_n164_), .B(alu__abc_38674_new_n165_), .Y(alu__abc_38674_new_n166_));
NOR2X1 NOR2X1_1024 ( .A(alu_b_i_29_), .B(alu_a_i_29_), .Y(alu__abc_38674_new_n167_));
NOR2X1 NOR2X1_1025 ( .A(alu__abc_38674_new_n167_), .B(alu__abc_38674_new_n166_), .Y(alu__abc_38674_new_n168_));
NOR2X1 NOR2X1_1026 ( .A(alu__abc_38674_new_n170_), .B(alu__abc_38674_new_n171_), .Y(alu__abc_38674_new_n172_));
NOR2X1 NOR2X1_1027 ( .A(alu_b_i_28_), .B(alu_a_i_28_), .Y(alu__abc_38674_new_n173_));
NOR2X1 NOR2X1_1028 ( .A(alu__abc_38674_new_n177_), .B(alu__abc_38674_new_n178_), .Y(alu__abc_38674_new_n179_));
NOR2X1 NOR2X1_1029 ( .A(alu_b_i_24_), .B(alu_a_i_24_), .Y(alu__abc_38674_new_n180_));
NOR2X1 NOR2X1_103 ( .A(_abc_40298_new_n1043_), .B(_abc_40298_new_n1059_), .Y(_abc_40298_new_n1060_));
NOR2X1 NOR2X1_1030 ( .A(alu_b_i_25_), .B(alu_a_i_25_), .Y(alu__abc_38674_new_n182_));
NOR2X1 NOR2X1_1031 ( .A(alu__abc_38674_new_n182_), .B(alu__abc_38674_new_n181_), .Y(alu__abc_38674_new_n183_));
NOR2X1 NOR2X1_1032 ( .A(alu__abc_38674_new_n186_), .B(alu__abc_38674_new_n187_), .Y(alu__abc_38674_new_n188_));
NOR2X1 NOR2X1_1033 ( .A(alu_b_i_26_), .B(alu_a_i_26_), .Y(alu__abc_38674_new_n189_));
NOR2X1 NOR2X1_1034 ( .A(alu__abc_38674_new_n189_), .B(alu__abc_38674_new_n188_), .Y(alu__abc_38674_new_n190_));
NOR2X1 NOR2X1_1035 ( .A(alu__abc_38674_new_n192_), .B(alu__abc_38674_new_n193_), .Y(alu__abc_38674_new_n194_));
NOR2X1 NOR2X1_1036 ( .A(alu_b_i_27_), .B(alu_a_i_27_), .Y(alu__abc_38674_new_n195_));
NOR2X1 NOR2X1_1037 ( .A(alu__abc_38674_new_n185_), .B(alu__abc_38674_new_n196_), .Y(alu__abc_38674_new_n197_));
NOR2X1 NOR2X1_1038 ( .A(alu__abc_38674_new_n176_), .B(alu__abc_38674_new_n198_), .Y(alu__abc_38674_new_n199_));
NOR2X1 NOR2X1_1039 ( .A(alu__abc_38674_new_n201_), .B(alu__abc_38674_new_n202_), .Y(alu__abc_38674_new_n203_));
NOR2X1 NOR2X1_104 ( .A(_abc_40298_new_n657_), .B(_abc_40298_new_n983_), .Y(_abc_40298_new_n1065_));
NOR2X1 NOR2X1_1040 ( .A(alu_b_i_14_), .B(alu_a_i_14_), .Y(alu__abc_38674_new_n204_));
NOR2X1 NOR2X1_1041 ( .A(alu_b_i_15_), .B(alu_a_i_15_), .Y(alu__abc_38674_new_n206_));
NOR2X1 NOR2X1_1042 ( .A(alu__abc_38674_new_n206_), .B(alu__abc_38674_new_n205_), .Y(alu__abc_38674_new_n207_));
NOR2X1 NOR2X1_1043 ( .A(alu__abc_38674_new_n210_), .B(alu__abc_38674_new_n211_), .Y(alu__abc_38674_new_n212_));
NOR2X1 NOR2X1_1044 ( .A(alu_b_i_12_), .B(alu_a_i_12_), .Y(alu__abc_38674_new_n213_));
NOR2X1 NOR2X1_1045 ( .A(alu__abc_38674_new_n213_), .B(alu__abc_38674_new_n212_), .Y(alu__abc_38674_new_n214_));
NOR2X1 NOR2X1_1046 ( .A(alu__abc_38674_new_n216_), .B(alu__abc_38674_new_n217_), .Y(alu__abc_38674_new_n218_));
NOR2X1 NOR2X1_1047 ( .A(alu_b_i_13_), .B(alu_a_i_13_), .Y(alu__abc_38674_new_n219_));
NOR2X1 NOR2X1_1048 ( .A(alu__abc_38674_new_n209_), .B(alu__abc_38674_new_n220_), .Y(alu__abc_38674_new_n221_));
NOR2X1 NOR2X1_1049 ( .A(alu__abc_38674_new_n240_), .B(alu__abc_38674_new_n236_), .Y(alu__abc_38674_new_n241_));
NOR2X1 NOR2X1_105 ( .A(_abc_40298_new_n1057_), .B(_abc_40298_new_n1075_), .Y(_abc_40298_new_n1076_));
NOR2X1 NOR2X1_1050 ( .A(alu_b_i_7_), .B(alu_a_i_7_), .Y(alu__abc_38674_new_n249_));
NOR2X1 NOR2X1_1051 ( .A(alu_b_i_4_), .B(alu_a_i_4_), .Y(alu__abc_38674_new_n255_));
NOR2X1 NOR2X1_1052 ( .A(alu__abc_38674_new_n250_), .B(alu__abc_38674_new_n256_), .Y(alu__abc_38674_new_n257_));
NOR2X1 NOR2X1_1053 ( .A(alu_b_i_0_), .B(alu__abc_38674_new_n258_), .Y(alu__abc_38674_new_n259_));
NOR2X1 NOR2X1_1054 ( .A(alu_a_i_1_), .B(alu_b_i_1_), .Y(alu__abc_38674_new_n262_));
NOR2X1 NOR2X1_1055 ( .A(alu_a_i_2_), .B(alu_b_i_2_), .Y(alu__abc_38674_new_n267_));
NOR2X1 NOR2X1_1056 ( .A(alu__abc_38674_new_n267_), .B(alu__abc_38674_new_n266_), .Y(alu__abc_38674_new_n268_));
NOR2X1 NOR2X1_1057 ( .A(alu_a_i_3_), .B(alu_b_i_3_), .Y(alu__abc_38674_new_n270_));
NOR2X1 NOR2X1_1058 ( .A(alu__abc_38674_new_n270_), .B(alu__abc_38674_new_n269_), .Y(alu__abc_38674_new_n271_));
NOR2X1 NOR2X1_1059 ( .A(alu__abc_38674_new_n268_), .B(alu__abc_38674_new_n271_), .Y(alu__abc_38674_new_n272_));
NOR2X1 NOR2X1_106 ( .A(_abc_40298_new_n1053_), .B(_abc_40298_new_n1077_), .Y(_abc_40298_new_n1078_));
NOR2X1 NOR2X1_1060 ( .A(alu__abc_38674_new_n259_), .B(alu__abc_38674_new_n273_), .Y(alu__abc_38674_new_n274_));
NOR2X1 NOR2X1_1061 ( .A(alu__abc_38674_new_n200_), .B(alu__abc_38674_new_n275_), .Y(alu_equal_o));
NOR2X1 NOR2X1_1062 ( .A(alu_op_i_3_), .B(alu__abc_38674_new_n277_), .Y(alu__abc_38674_new_n278_));
NOR2X1 NOR2X1_1063 ( .A(alu_op_i_1_), .B(alu_op_i_0_), .Y(alu__abc_38674_new_n280_));
NOR2X1 NOR2X1_1064 ( .A(alu__abc_38674_new_n281_), .B(alu__abc_38674_new_n279_), .Y(alu__abc_38674_new_n282_));
NOR2X1 NOR2X1_1065 ( .A(alu_op_i_1_), .B(alu__abc_38674_new_n284_), .Y(alu__abc_38674_new_n285_));
NOR2X1 NOR2X1_1066 ( .A(alu_op_i_0_), .B(alu__abc_38674_new_n288_), .Y(alu__abc_38674_new_n289_));
NOR2X1 NOR2X1_1067 ( .A(alu__abc_38674_new_n290_), .B(alu__abc_38674_new_n292_), .Y(alu_flag_update_o));
NOR2X1 NOR2X1_1068 ( .A(alu_b_i_24_), .B(alu__abc_38674_new_n178_), .Y(alu__abc_38674_new_n296_));
NOR2X1 NOR2X1_1069 ( .A(alu__abc_38674_new_n299_), .B(alu__abc_38674_new_n196_), .Y(alu__abc_38674_new_n300_));
NOR2X1 NOR2X1_107 ( .A(_abc_40298_new_n940_), .B(_abc_40298_new_n1090_), .Y(_abc_40298_new_n1091_));
NOR2X1 NOR2X1_1070 ( .A(alu_b_i_26_), .B(alu__abc_38674_new_n187_), .Y(alu__abc_38674_new_n301_));
NOR2X1 NOR2X1_1071 ( .A(alu__abc_38674_new_n303_), .B(alu__abc_38674_new_n300_), .Y(alu__abc_38674_new_n304_));
NOR2X1 NOR2X1_1072 ( .A(alu__abc_38674_new_n146_), .B(alu__abc_38674_new_n145_), .Y(alu__abc_38674_new_n306_));
NOR2X1 NOR2X1_1073 ( .A(alu_b_i_19_), .B(alu__abc_38674_new_n312_), .Y(alu__abc_38674_new_n313_));
NOR2X1 NOR2X1_1074 ( .A(alu_b_i_18_), .B(alu__abc_38674_new_n144_), .Y(alu__abc_38674_new_n314_));
NOR2X1 NOR2X1_1075 ( .A(alu_b_i_20_), .B(alu__abc_38674_new_n122_), .Y(alu__abc_38674_new_n317_));
NOR2X1 NOR2X1_1076 ( .A(alu__abc_38674_new_n119_), .B(alu__abc_38674_new_n118_), .Y(alu__abc_38674_new_n321_));
NOR2X1 NOR2X1_1077 ( .A(alu_b_i_23_), .B(alu__abc_38674_new_n117_), .Y(alu__abc_38674_new_n323_));
NOR2X1 NOR2X1_1078 ( .A(alu_b_i_22_), .B(alu__abc_38674_new_n111_), .Y(alu__abc_38674_new_n324_));
NOR2X1 NOR2X1_1079 ( .A(alu__abc_38674_new_n326_), .B(alu__abc_38674_new_n316_), .Y(alu__abc_38674_new_n327_));
NOR2X1 NOR2X1_108 ( .A(_abc_40298_new_n1101_), .B(_abc_40298_new_n971_), .Y(_abc_40298_new_n1102_));
NOR2X1 NOR2X1_1080 ( .A(alu_b_i_6_), .B(alu__abc_38674_new_n330_), .Y(alu__abc_38674_new_n331_));
NOR2X1 NOR2X1_1081 ( .A(alu__abc_38674_new_n255_), .B(alu__abc_38674_new_n254_), .Y(alu__abc_38674_new_n335_));
NOR2X1 NOR2X1_1082 ( .A(alu__abc_38674_new_n335_), .B(alu__abc_38674_new_n343_), .Y(alu__abc_38674_new_n344_));
NOR2X1 NOR2X1_1083 ( .A(alu_b_i_4_), .B(alu__abc_38674_new_n345_), .Y(alu__abc_38674_new_n346_));
NOR2X1 NOR2X1_1084 ( .A(alu__abc_38674_new_n243_), .B(alu__abc_38674_new_n349_), .Y(alu__abc_38674_new_n350_));
NOR2X1 NOR2X1_1085 ( .A(alu_b_i_8_), .B(alu__abc_38674_new_n351_), .Y(alu__abc_38674_new_n352_));
NOR2X1 NOR2X1_1086 ( .A(alu__abc_38674_new_n358_), .B(alu__abc_38674_new_n355_), .Y(alu__abc_38674_new_n359_));
NOR2X1 NOR2X1_1087 ( .A(alu_b_i_12_), .B(alu__abc_38674_new_n211_), .Y(alu__abc_38674_new_n361_));
NOR2X1 NOR2X1_1088 ( .A(alu__abc_38674_new_n305_), .B(alu__abc_38674_new_n371_), .Y(alu__abc_38674_new_n372_));
NOR2X1 NOR2X1_1089 ( .A(alu_b_i_29_), .B(alu__abc_38674_new_n165_), .Y(alu__abc_38674_new_n373_));
NOR2X1 NOR2X1_109 ( .A(alu_greater_than_o), .B(_abc_40298_new_n1020_), .Y(_abc_40298_new_n1108_));
NOR2X1 NOR2X1_1090 ( .A(alu_b_i_28_), .B(alu__abc_38674_new_n171_), .Y(alu__abc_38674_new_n374_));
NOR2X1 NOR2X1_1091 ( .A(alu__abc_38674_new_n279_), .B(alu__abc_38674_new_n286_), .Y(alu__abc_38674_new_n381_));
NOR2X1 NOR2X1_1092 ( .A(alu__abc_38674_new_n384_), .B(alu__abc_38674_new_n383_), .Y(alu__abc_38674_new_n385_));
NOR2X1 NOR2X1_1093 ( .A(alu__abc_38674_new_n173_), .B(alu__abc_38674_new_n172_), .Y(alu__abc_38674_new_n389_));
NOR2X1 NOR2X1_1094 ( .A(alu__abc_38674_new_n169_), .B(alu__abc_38674_new_n390_), .Y(alu__abc_38674_new_n391_));
NOR2X1 NOR2X1_1095 ( .A(alu__abc_38674_new_n195_), .B(alu__abc_38674_new_n194_), .Y(alu__abc_38674_new_n395_));
NOR2X1 NOR2X1_1096 ( .A(alu__abc_38674_new_n191_), .B(alu__abc_38674_new_n396_), .Y(alu__abc_38674_new_n398_));
NOR2X1 NOR2X1_1097 ( .A(alu__abc_38674_new_n130_), .B(alu__abc_38674_new_n129_), .Y(alu__abc_38674_new_n410_));
NOR2X1 NOR2X1_1098 ( .A(alu__abc_38674_new_n405_), .B(alu__abc_38674_new_n411_), .Y(alu__abc_38674_new_n412_));
NOR2X1 NOR2X1_1099 ( .A(alu_b_i_6_), .B(alu_a_i_6_), .Y(alu__abc_38674_new_n427_));
NOR2X1 NOR2X1_11 ( .A(_abc_40298_new_n636_), .B(_abc_40298_new_n651_), .Y(_abc_40298_new_n652_));
NOR2X1 NOR2X1_110 ( .A(_abc_40298_new_n1107_), .B(_abc_40298_new_n1108_), .Y(_abc_40298_new_n1109_));
NOR2X1 NOR2X1_1100 ( .A(alu__abc_38674_new_n427_), .B(alu__abc_38674_new_n426_), .Y(alu__abc_38674_new_n428_));
NOR2X1 NOR2X1_1101 ( .A(alu__abc_38674_new_n249_), .B(alu__abc_38674_new_n248_), .Y(alu__abc_38674_new_n429_));
NOR2X1 NOR2X1_1102 ( .A(alu_b_i_5_), .B(alu_a_i_5_), .Y(alu__abc_38674_new_n432_));
NOR2X1 NOR2X1_1103 ( .A(alu__abc_38674_new_n432_), .B(alu__abc_38674_new_n431_), .Y(alu__abc_38674_new_n433_));
NOR2X1 NOR2X1_1104 ( .A(alu__abc_38674_new_n430_), .B(alu__abc_38674_new_n434_), .Y(alu__abc_38674_new_n435_));
NOR2X1 NOR2X1_1105 ( .A(alu__abc_38674_new_n219_), .B(alu__abc_38674_new_n218_), .Y(alu__abc_38674_new_n451_));
NOR2X1 NOR2X1_1106 ( .A(alu__abc_38674_new_n204_), .B(alu__abc_38674_new_n203_), .Y(alu__abc_38674_new_n453_));
NOR2X1 NOR2X1_1107 ( .A(alu__abc_38674_new_n454_), .B(alu__abc_38674_new_n456_), .Y(alu__abc_38674_new_n457_));
NOR2X1 NOR2X1_1108 ( .A(alu__abc_38674_new_n239_), .B(alu__abc_38674_new_n235_), .Y(alu__abc_38674_new_n459_));
NOR2X1 NOR2X1_1109 ( .A(alu__abc_38674_new_n225_), .B(alu__abc_38674_new_n230_), .Y(alu__abc_38674_new_n460_));
NOR2X1 NOR2X1_111 ( .A(alu_equal_o), .B(alu_greater_than_o), .Y(_abc_40298_new_n1114_));
NOR2X1 NOR2X1_1110 ( .A(alu__abc_38674_new_n137_), .B(alu__abc_38674_new_n136_), .Y(alu__abc_38674_new_n465_));
NOR2X1 NOR2X1_1111 ( .A(alu__abc_38674_new_n413_), .B(alu__abc_38674_new_n466_), .Y(alu__abc_38674_new_n467_));
NOR2X1 NOR2X1_1112 ( .A(alu__abc_38674_new_n180_), .B(alu__abc_38674_new_n179_), .Y(alu__abc_38674_new_n471_));
NOR2X1 NOR2X1_1113 ( .A(alu__abc_38674_new_n184_), .B(alu__abc_38674_new_n472_), .Y(alu__abc_38674_new_n473_));
NOR2X1 NOR2X1_1114 ( .A(alu__abc_38674_new_n493_), .B(alu__abc_38674_new_n496_), .Y(alu__abc_38674_new_n497_));
NOR2X1 NOR2X1_1115 ( .A(alu__abc_38674_new_n247_), .B(alu__abc_38674_new_n517_), .Y(alu__abc_38674_new_n518_));
NOR2X1 NOR2X1_1116 ( .A(alu__abc_38674_new_n253_), .B(alu__abc_38674_new_n521_), .Y(alu__abc_38674_new_n522_));
NOR2X1 NOR2X1_1117 ( .A(alu__abc_38674_new_n561_), .B(alu__abc_38674_new_n564_), .Y(alu__abc_38674_new_n565_));
NOR2X1 NOR2X1_1118 ( .A(alu__abc_38674_new_n566_), .B(alu__abc_38674_new_n569_), .Y(alu__abc_38674_new_n570_));
NOR2X1 NOR2X1_1119 ( .A(alu__abc_38674_new_n500_), .B(alu__abc_38674_new_n607_), .Y(alu__abc_38674_new_n608_));
NOR2X1 NOR2X1_112 ( .A(_abc_40298_new_n1134_), .B(_abc_40298_new_n1071_), .Y(_abc_40298_new_n1135_));
NOR2X1 NOR2X1_1120 ( .A(alu__abc_38674_new_n624_), .B(alu__abc_38674_new_n620_), .Y(alu__abc_38674_new_n625_));
NOR2X1 NOR2X1_1121 ( .A(alu_a_i_1_), .B(alu__abc_38674_new_n562_), .Y(alu__abc_38674_new_n644_));
NOR2X1 NOR2X1_1122 ( .A(alu_op_i_3_), .B(alu_op_i_2_), .Y(alu__abc_38674_new_n656_));
NOR2X1 NOR2X1_1123 ( .A(alu__abc_38674_new_n288_), .B(alu__abc_38674_new_n284_), .Y(alu__abc_38674_new_n657_));
NOR2X1 NOR2X1_1124 ( .A(alu_a_i_30_), .B(alu_b_i_0_), .Y(alu__abc_38674_new_n659_));
NOR2X1 NOR2X1_1125 ( .A(alu_b_i_1_), .B(alu__abc_38674_new_n695_), .Y(alu__abc_38674_new_n696_));
NOR2X1 NOR2X1_1126 ( .A(alu__abc_38674_new_n698_), .B(alu__abc_38674_new_n286_), .Y(alu__abc_38674_new_n699_));
NOR2X1 NOR2X1_1127 ( .A(alu_b_i_4_), .B(alu__abc_38674_new_n700_), .Y(alu__abc_38674_new_n701_));
NOR2X1 NOR2X1_1128 ( .A(alu__abc_38674_new_n281_), .B(alu__abc_38674_new_n292_), .Y(alu__abc_38674_new_n703_));
NOR2X1 NOR2X1_1129 ( .A(alu__abc_38674_new_n286_), .B(alu__abc_38674_new_n292_), .Y(alu__abc_38674_new_n705_));
NOR2X1 NOR2X1_113 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_10_), .B(_abc_40298_new_n1061_), .Y(_abc_40298_new_n1150_));
NOR2X1 NOR2X1_1130 ( .A(alu__abc_38674_new_n279_), .B(alu__abc_38674_new_n290_), .Y(alu__abc_38674_new_n706_));
NOR2X1 NOR2X1_1131 ( .A(alu__abc_38674_new_n714_), .B(alu__abc_38674_new_n709_), .Y(alu__abc_38674_new_n715_));
NOR2X1 NOR2X1_1132 ( .A(alu_a_i_2_), .B(alu__abc_38674_new_n562_), .Y(alu__abc_38674_new_n718_));
NOR2X1 NOR2X1_1133 ( .A(alu_a_i_1_), .B(alu_b_i_0_), .Y(alu__abc_38674_new_n719_));
NOR2X1 NOR2X1_1134 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n725_), .Y(alu__abc_38674_new_n726_));
NOR2X1 NOR2X1_1135 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n739_), .Y(alu__abc_38674_new_n740_));
NOR2X1 NOR2X1_1136 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n779_), .Y(alu__abc_38674_new_n780_));
NOR2X1 NOR2X1_1137 ( .A(alu__abc_38674_new_n265_), .B(alu__abc_38674_new_n782_), .Y(alu__abc_38674_new_n783_));
NOR2X1 NOR2X1_1138 ( .A(alu__abc_38674_new_n785_), .B(alu__abc_38674_new_n791_), .Y(alu__abc_38674_new_n792_));
NOR2X1 NOR2X1_1139 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n839_), .Y(alu__abc_38674_new_n840_));
NOR2X1 NOR2X1_114 ( .A(_abc_40298_new_n1069_), .B(_abc_40298_new_n1029_), .Y(_abc_40298_new_n1159_));
NOR2X1 NOR2X1_1140 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n888_), .Y(alu__abc_38674_new_n889_));
NOR2X1 NOR2X1_1141 ( .A(alu__abc_38674_new_n270_), .B(alu__abc_38674_new_n787_), .Y(alu__abc_38674_new_n894_));
NOR2X1 NOR2X1_1142 ( .A(alu__abc_38674_new_n893_), .B(alu__abc_38674_new_n899_), .Y(alu__abc_38674_new_n900_));
NOR2X1 NOR2X1_1143 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n910_), .Y(alu__abc_38674_new_n911_));
NOR2X1 NOR2X1_1144 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n914_), .Y(alu__abc_38674_new_n915_));
NOR2X1 NOR2X1_1145 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n931_), .Y(alu__abc_38674_new_n932_));
NOR2X1 NOR2X1_1146 ( .A(alu__abc_38674_new_n345_), .B(alu__abc_38674_new_n713_), .Y(alu__abc_38674_new_n933_));
NOR2X1 NOR2X1_1147 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n959_), .Y(alu__abc_38674_new_n960_));
NOR2X1 NOR2X1_1148 ( .A(alu__abc_38674_new_n903_), .B(alu__abc_38674_new_n902_), .Y(alu__abc_38674_new_n968_));
NOR2X1 NOR2X1_1149 ( .A(alu__abc_38674_new_n552_), .B(alu__abc_38674_new_n572_), .Y(alu__abc_38674_new_n969_));
NOR2X1 NOR2X1_115 ( .A(_abc_40298_new_n1073_), .B(_abc_40298_new_n1069_), .Y(_abc_40298_new_n1173_));
NOR2X1 NOR2X1_1150 ( .A(alu__abc_38674_new_n382_), .B(alu__abc_38674_new_n969_), .Y(alu__abc_38674_new_n970_));
NOR2X1 NOR2X1_1151 ( .A(alu__abc_38674_new_n346_), .B(alu__abc_38674_new_n253_), .Y(alu__abc_38674_new_n972_));
NOR2X1 NOR2X1_1152 ( .A(alu__abc_38674_new_n382_), .B(alu__abc_38674_new_n573_), .Y(alu__abc_38674_new_n980_));
NOR2X1 NOR2X1_1153 ( .A(alu__abc_38674_new_n538_), .B(alu__abc_38674_new_n574_), .Y(alu__abc_38674_new_n1075_));
NOR2X1 NOR2X1_1154 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n739_), .Y(alu__abc_38674_new_n1081_));
NOR2X1 NOR2X1_1155 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n756_), .Y(alu__abc_38674_new_n1082_));
NOR2X1 NOR2X1_1156 ( .A(alu__abc_38674_new_n1094_), .B(alu__abc_38674_new_n1078_), .Y(alu__abc_38674_new_n1095_));
NOR2X1 NOR2X1_1157 ( .A(alu__abc_38674_new_n539_), .B(alu__abc_38674_new_n349_), .Y(alu__abc_38674_new_n1100_));
NOR2X1 NOR2X1_1158 ( .A(alu__abc_38674_new_n1102_), .B(alu__abc_38674_new_n1101_), .Y(alu__abc_38674_new_n1103_));
NOR2X1 NOR2X1_1159 ( .A(alu__abc_38674_new_n1097_), .B(alu__abc_38674_new_n1105_), .Y(alu__abc_38674_new_n1106_));
NOR2X1 NOR2X1_116 ( .A(_abc_40298_new_n1183_), .B(_abc_40298_new_n1181_), .Y(_abc_40298_new_n1184_));
NOR2X1 NOR2X1_1160 ( .A(alu__abc_38674_new_n354_), .B(alu__abc_38674_new_n1101_), .Y(alu__abc_38674_new_n1109_));
NOR2X1 NOR2X1_1161 ( .A(alu__abc_38674_new_n382_), .B(alu__abc_38674_new_n1113_), .Y(alu__abc_38674_new_n1114_));
NOR2X1 NOR2X1_1162 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n876_), .Y(alu__abc_38674_new_n1146_));
NOR2X1 NOR2X1_1163 ( .A(alu__abc_38674_new_n1176_), .B(alu__abc_38674_new_n1174_), .Y(alu__abc_38674_new_n1177_));
NOR2X1 NOR2X1_1164 ( .A(alu__abc_38674_new_n382_), .B(alu__abc_38674_new_n1177_), .Y(alu__abc_38674_new_n1178_));
NOR2X1 NOR2X1_1165 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n914_), .Y(alu__abc_38674_new_n1193_));
NOR2X1 NOR2X1_1166 ( .A(alu__abc_38674_new_n451_), .B(alu__abc_38674_new_n1207_), .Y(alu__abc_38674_new_n1208_));
NOR2X1 NOR2X1_1167 ( .A(alu__abc_38674_new_n363_), .B(alu__abc_38674_new_n1208_), .Y(alu__abc_38674_new_n1234_));
NOR2X1 NOR2X1_1168 ( .A(alu__abc_38674_new_n1176_), .B(alu__abc_38674_new_n584_), .Y(alu__abc_38674_new_n1268_));
NOR2X1 NOR2X1_1169 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n1016_), .Y(alu__abc_38674_new_n1273_));
NOR2X1 NOR2X1_117 ( .A(next_pc_r_0_), .B(_abc_40298_new_n1138_), .Y(_abc_40298_new_n1193_));
NOR2X1 NOR2X1_1170 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n1019_), .Y(alu__abc_38674_new_n1274_));
NOR2X1 NOR2X1_1171 ( .A(alu__abc_38674_new_n1116_), .B(alu__abc_38674_new_n1176_), .Y(alu__abc_38674_new_n1295_));
NOR2X1 NOR2X1_1172 ( .A(alu__abc_38674_new_n369_), .B(alu__abc_38674_new_n350_), .Y(alu__abc_38674_new_n1301_));
NOR2X1 NOR2X1_1173 ( .A(alu__abc_38674_new_n698_), .B(alu__abc_38674_new_n765_), .Y(alu__abc_38674_new_n1304_));
NOR2X1 NOR2X1_1174 ( .A(alu__abc_38674_new_n519_), .B(alu__abc_38674_new_n700_), .Y(alu__abc_38674_new_n1317_));
NOR2X1 NOR2X1_1175 ( .A(alu__abc_38674_new_n283_), .B(alu__abc_38674_new_n1327_), .Y(alu__abc_38674_new_n1329_));
NOR2X1 NOR2X1_1176 ( .A(alu__abc_38674_new_n1327_), .B(alu__abc_38674_new_n1330_), .Y(alu__abc_38674_new_n1331_));
NOR2X1 NOR2X1_1177 ( .A(alu__abc_38674_new_n382_), .B(alu__abc_38674_new_n1331_), .Y(alu__abc_38674_new_n1332_));
NOR2X1 NOR2X1_1178 ( .A(alu__abc_38674_new_n465_), .B(alu__abc_38674_new_n1301_), .Y(alu__abc_38674_new_n1334_));
NOR2X1 NOR2X1_1179 ( .A(alu__abc_38674_new_n1338_), .B(alu__abc_38674_new_n1337_), .Y(alu__abc_38674_new_n1339_));
NOR2X1 NOR2X1_118 ( .A(next_pc_r_1_), .B(_abc_40298_new_n1138_), .Y(_abc_40298_new_n1205_));
NOR2X1 NOR2X1_1180 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n1345_), .Y(alu__abc_38674_new_n1346_));
NOR2X1 NOR2X1_1181 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n1091_), .Y(alu__abc_38674_new_n1347_));
NOR2X1 NOR2X1_1182 ( .A(alu__abc_38674_new_n310_), .B(alu__abc_38674_new_n1337_), .Y(alu__abc_38674_new_n1363_));
NOR2X1 NOR2X1_1183 ( .A(alu__abc_38674_new_n146_), .B(alu__abc_38674_new_n787_), .Y(alu__abc_38674_new_n1367_));
NOR2X1 NOR2X1_1184 ( .A(alu__abc_38674_new_n1401_), .B(alu__abc_38674_new_n1408_), .Y(alu__abc_38674_new_n1409_));
NOR2X1 NOR2X1_1185 ( .A(alu__abc_38674_new_n153_), .B(alu__abc_38674_new_n1301_), .Y(alu__abc_38674_new_n1421_));
NOR2X1 NOR2X1_1186 ( .A(alu__abc_38674_new_n1420_), .B(alu__abc_38674_new_n1421_), .Y(alu__abc_38674_new_n1422_));
NOR2X1 NOR2X1_1187 ( .A(alu__abc_38674_new_n1439_), .B(alu__abc_38674_new_n1436_), .Y(alu__abc_38674_new_n1440_));
NOR2X1 NOR2X1_1188 ( .A(alu__abc_38674_new_n283_), .B(alu__abc_38674_new_n493_), .Y(alu__abc_38674_new_n1451_));
NOR2X1 NOR2X1_1189 ( .A(alu__abc_38674_new_n283_), .B(alu__abc_38674_new_n496_), .Y(alu__abc_38674_new_n1471_));
NOR2X1 NOR2X1_119 ( .A(alu_op_r_0_), .B(pc_q_2_), .Y(_abc_40298_new_n1214_));
NOR2X1 NOR2X1_1190 ( .A(alu__abc_38674_new_n782_), .B(alu__abc_38674_new_n1488_), .Y(alu__abc_38674_new_n1489_));
NOR2X1 NOR2X1_1191 ( .A(alu__abc_38674_new_n1486_), .B(alu__abc_38674_new_n1494_), .Y(alu__abc_38674_new_n1495_));
NOR2X1 NOR2X1_1192 ( .A(alu__abc_38674_new_n324_), .B(alu__abc_38674_new_n1488_), .Y(alu__abc_38674_new_n1503_));
NOR2X1 NOR2X1_1193 ( .A(alu__abc_38674_new_n382_), .B(alu__abc_38674_new_n1547_), .Y(alu__abc_38674_new_n1548_));
NOR2X1 NOR2X1_1194 ( .A(alu__abc_38674_new_n296_), .B(alu__abc_38674_new_n184_), .Y(alu__abc_38674_new_n1560_));
NOR2X1 NOR2X1_1195 ( .A(alu__abc_38674_new_n499_), .B(alu__abc_38674_new_n1547_), .Y(alu__abc_38674_new_n1572_));
NOR2X1 NOR2X1_1196 ( .A(alu__abc_38674_new_n1576_), .B(alu__abc_38674_new_n1572_), .Y(alu__abc_38674_new_n1577_));
NOR2X1 NOR2X1_1197 ( .A(alu__abc_38674_new_n782_), .B(alu__abc_38674_new_n1580_), .Y(alu__abc_38674_new_n1581_));
NOR2X1 NOR2X1_1198 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n1590_), .Y(alu__abc_38674_new_n1591_));
NOR2X1 NOR2X1_1199 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n1374_), .Y(alu__abc_38674_new_n1592_));
NOR2X1 NOR2X1_12 ( .A(inst_r_0_), .B(_abc_40298_new_n656_), .Y(_abc_40298_new_n658_));
NOR2X1 NOR2X1_120 ( .A(_abc_40298_new_n911_), .B(_abc_40298_new_n1215_), .Y(_abc_40298_new_n1216_));
NOR2X1 NOR2X1_1200 ( .A(alu__abc_38674_new_n619_), .B(alu__abc_38674_new_n1576_), .Y(alu__abc_38674_new_n1601_));
NOR2X1 NOR2X1_1201 ( .A(alu__abc_38674_new_n301_), .B(alu__abc_38674_new_n1580_), .Y(alu__abc_38674_new_n1604_));
NOR2X1 NOR2X1_1202 ( .A(alu_b_i_1_), .B(alu__abc_38674_new_n1634_), .Y(alu__abc_38674_new_n1635_));
NOR2X1 NOR2X1_1203 ( .A(alu__abc_38674_new_n782_), .B(alu__abc_38674_new_n1675_), .Y(alu__abc_38674_new_n1676_));
NOR2X1 NOR2X1_1204 ( .A(alu_b_i_30_), .B(alu__abc_38674_new_n156_), .Y(alu__abc_38674_new_n1699_));
NOR2X1 NOR2X1_1205 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n1707_), .Y(alu__abc_38674_new_n1708_));
NOR2X1 NOR2X1_1206 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n1610_), .Y(alu__abc_38674_new_n1709_));
NOR2X1 NOR2X1_1207 ( .A(alu_equal_o), .B(alu_less_than_signed_o), .Y(alu_greater_than_signed_o));
NOR2X1 NOR2X1_1208 ( .A(alu__abc_38674_new_n200_), .B(alu__abc_38674_new_n1301_), .Y(alu__abc_38674_new_n1723_));
NOR2X1 NOR2X1_1209 ( .A(alu__abc_38674_new_n1730_), .B(alu__abc_38674_new_n1723_), .Y(alu_less_than_o));
NOR2X1 NOR2X1_121 ( .A(_abc_40298_new_n1214_), .B(_abc_40298_new_n1216_), .Y(_abc_40298_new_n1217_));
NOR2X1 NOR2X1_1210 ( .A(alu_equal_o), .B(alu_less_than_o), .Y(alu_greater_than_o));
NOR2X1 NOR2X1_122 ( .A(pc_q_2_), .B(pc_q_3_), .Y(_abc_40298_new_n1241_));
NOR2X1 NOR2X1_123 ( .A(_abc_40298_new_n1241_), .B(_abc_40298_new_n1242_), .Y(_abc_40298_new_n1246_));
NOR2X1 NOR2X1_124 ( .A(alu_op_r_2_), .B(pc_q_4_), .Y(_abc_40298_new_n1262_));
NOR2X1 NOR2X1_125 ( .A(_abc_40298_new_n898_), .B(_abc_40298_new_n1256_), .Y(_abc_40298_new_n1263_));
NOR2X1 NOR2X1_126 ( .A(_abc_40298_new_n1262_), .B(_abc_40298_new_n1263_), .Y(_abc_40298_new_n1264_));
NOR2X1 NOR2X1_127 ( .A(_abc_40298_new_n1265_), .B(_abc_40298_new_n984_), .Y(_abc_40298_new_n1266_));
NOR2X1 NOR2X1_128 ( .A(alu_op_r_3_), .B(pc_q_5_), .Y(_abc_40298_new_n1278_));
NOR2X1 NOR2X1_129 ( .A(_abc_40298_new_n1278_), .B(_abc_40298_new_n1280_), .Y(_abc_40298_new_n1281_));
NOR2X1 NOR2X1_13 ( .A(_abc_40298_new_n643_), .B(_abc_40298_new_n662_), .Y(_abc_40298_new_n663_));
NOR2X1 NOR2X1_130 ( .A(_abc_40298_new_n1263_), .B(_abc_40298_new_n1265_), .Y(_abc_40298_new_n1282_));
NOR2X1 NOR2X1_131 ( .A(int32_r_4_), .B(pc_q_6_), .Y(_abc_40298_new_n1314_));
NOR2X1 NOR2X1_132 ( .A(_abc_40298_new_n1315_), .B(_abc_40298_new_n1302_), .Y(_abc_40298_new_n1316_));
NOR2X1 NOR2X1_133 ( .A(pc_q_7_), .B(_abc_40298_new_n1304_), .Y(_abc_40298_new_n1331_));
NOR2X1 NOR2X1_134 ( .A(_abc_40298_new_n1331_), .B(_abc_40298_new_n1333_), .Y(_abc_40298_new_n1334_));
NOR2X1 NOR2X1_135 ( .A(_abc_40298_new_n1336_), .B(_abc_40298_new_n1134_), .Y(_abc_40298_new_n1337_));
NOR2X1 NOR2X1_136 ( .A(int32_r_5_), .B(pc_q_7_), .Y(_abc_40298_new_n1340_));
NOR2X1 NOR2X1_137 ( .A(_abc_40298_new_n1341_), .B(_abc_40298_new_n1332_), .Y(_abc_40298_new_n1342_));
NOR2X1 NOR2X1_138 ( .A(_abc_40298_new_n1340_), .B(_abc_40298_new_n1342_), .Y(_abc_40298_new_n1343_));
NOR2X1 NOR2X1_139 ( .A(_abc_40298_new_n1343_), .B(_abc_40298_new_n1346_), .Y(_abc_40298_new_n1347_));
NOR2X1 NOR2X1_14 ( .A(mem_offset_q_0_), .B(_abc_40298_new_n672_), .Y(_abc_40298_new_n673_));
NOR2X1 NOR2X1_140 ( .A(_abc_40298_new_n1317_), .B(_abc_40298_new_n1348_), .Y(_abc_40298_new_n1349_));
NOR2X1 NOR2X1_141 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1357_), .Y(_abc_40298_new_n1358_));
NOR2X1 NOR2X1_142 ( .A(alu_op_r_4_), .B(pc_q_8_), .Y(_abc_40298_new_n1374_));
NOR2X1 NOR2X1_143 ( .A(_abc_40298_new_n917_), .B(_abc_40298_new_n1362_), .Y(_abc_40298_new_n1375_));
NOR2X1 NOR2X1_144 ( .A(_abc_40298_new_n1374_), .B(_abc_40298_new_n1375_), .Y(_abc_40298_new_n1376_));
NOR2X1 NOR2X1_145 ( .A(_abc_40298_new_n984_), .B(_abc_40298_new_n1377_), .Y(_abc_40298_new_n1378_));
NOR2X1 NOR2X1_146 ( .A(_abc_40298_new_n1389_), .B(_abc_40298_new_n1388_), .Y(_0epc_q_31_0__8_));
NOR2X1 NOR2X1_147 ( .A(_abc_40298_new_n1393_), .B(_abc_40298_new_n1134_), .Y(_abc_40298_new_n1394_));
NOR2X1 NOR2X1_148 ( .A(alu_op_r_5_), .B(pc_q_9_), .Y(_abc_40298_new_n1398_));
NOR2X1 NOR2X1_149 ( .A(_abc_40298_new_n973_), .B(_abc_40298_new_n1399_), .Y(_abc_40298_new_n1400_));
NOR2X1 NOR2X1_15 ( .A(mem_offset_q_1_), .B(mem_offset_q_0_), .Y(_abc_40298_new_n674_));
NOR2X1 NOR2X1_150 ( .A(_abc_40298_new_n1375_), .B(_abc_40298_new_n1377_), .Y(_abc_40298_new_n1401_));
NOR2X1 NOR2X1_151 ( .A(_abc_40298_new_n1398_), .B(_abc_40298_new_n1400_), .Y(_abc_40298_new_n1403_));
NOR2X1 NOR2X1_152 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1409_), .Y(_abc_40298_new_n1410_));
NOR2X1 NOR2X1_153 ( .A(_abc_40298_new_n1421_), .B(_abc_40298_new_n1134_), .Y(_abc_40298_new_n1422_));
NOR2X1 NOR2X1_154 ( .A(_abc_40298_new_n1423_), .B(_abc_40298_new_n1372_), .Y(_abc_40298_new_n1424_));
NOR2X1 NOR2X1_155 ( .A(alu_op_r_6_), .B(pc_q_10_), .Y(_abc_40298_new_n1427_));
NOR2X1 NOR2X1_156 ( .A(_abc_40298_new_n1427_), .B(_abc_40298_new_n1429_), .Y(_abc_40298_new_n1430_));
NOR2X1 NOR2X1_157 ( .A(_abc_40298_new_n1426_), .B(_abc_40298_new_n1424_), .Y(_abc_40298_new_n1433_));
NOR2X1 NOR2X1_158 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1441_), .Y(_abc_40298_new_n1442_));
NOR2X1 NOR2X1_159 ( .A(pc_q_11_), .B(_abc_40298_new_n1416_), .Y(_abc_40298_new_n1446_));
NOR2X1 NOR2X1_16 ( .A(mem_offset_q_1_), .B(_abc_40298_new_n676_), .Y(_abc_40298_new_n677_));
NOR2X1 NOR2X1_160 ( .A(_abc_40298_new_n1446_), .B(_abc_40298_new_n1449_), .Y(_abc_40298_new_n1450_));
NOR2X1 NOR2X1_161 ( .A(_abc_40298_new_n1452_), .B(_abc_40298_new_n1134_), .Y(_abc_40298_new_n1453_));
NOR2X1 NOR2X1_162 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1468_), .Y(_abc_40298_new_n1469_));
NOR2X1 NOR2X1_163 ( .A(_abc_40298_new_n1460_), .B(_abc_40298_new_n1434_), .Y(_abc_40298_new_n1480_));
NOR2X1 NOR2X1_164 ( .A(_abc_40298_new_n1423_), .B(_abc_40298_new_n1485_), .Y(_abc_40298_new_n1486_));
NOR2X1 NOR2X1_165 ( .A(_abc_40298_new_n1487_), .B(_abc_40298_new_n1372_), .Y(_abc_40298_new_n1488_));
NOR2X1 NOR2X1_166 ( .A(int32_r_10_), .B(pc_q_12_), .Y(_abc_40298_new_n1490_));
NOR2X1 NOR2X1_167 ( .A(_abc_40298_new_n1490_), .B(_abc_40298_new_n1492_), .Y(_abc_40298_new_n1493_));
NOR2X1 NOR2X1_168 ( .A(_abc_40298_new_n984_), .B(_abc_40298_new_n1495_), .Y(_abc_40298_new_n1496_));
NOR2X1 NOR2X1_169 ( .A(pc_q_13_), .B(REGFILE_SIM_reg_bank_rb_i_0_), .Y(_abc_40298_new_n1511_));
NOR2X1 NOR2X1_17 ( .A(_abc_40298_new_n672_), .B(_abc_40298_new_n676_), .Y(_abc_40298_new_n679_));
NOR2X1 NOR2X1_170 ( .A(_abc_40298_new_n1512_), .B(_abc_40298_new_n1513_), .Y(_abc_40298_new_n1514_));
NOR2X1 NOR2X1_171 ( .A(_abc_40298_new_n1511_), .B(_abc_40298_new_n1514_), .Y(_abc_40298_new_n1515_));
NOR2X1 NOR2X1_172 ( .A(_abc_40298_new_n1492_), .B(_abc_40298_new_n1515_), .Y(_abc_40298_new_n1518_));
NOR2X1 NOR2X1_173 ( .A(_abc_40298_new_n1176_), .B(_abc_40298_new_n1522_), .Y(_abc_40298_new_n1523_));
NOR2X1 NOR2X1_174 ( .A(pc_q_14_), .B(REGFILE_SIM_reg_bank_rb_i_1_), .Y(_abc_40298_new_n1543_));
NOR2X1 NOR2X1_175 ( .A(_abc_40298_new_n1543_), .B(_abc_40298_new_n1545_), .Y(_abc_40298_new_n1546_));
NOR2X1 NOR2X1_176 ( .A(pc_q_15_), .B(REGFILE_SIM_reg_bank_rb_i_2_), .Y(_abc_40298_new_n1570_));
NOR2X1 NOR2X1_177 ( .A(_abc_40298_new_n1570_), .B(_abc_40298_new_n1572_), .Y(_abc_40298_new_n1573_));
NOR2X1 NOR2X1_178 ( .A(_abc_40298_new_n1600_), .B(_abc_40298_new_n1372_), .Y(_abc_40298_new_n1601_));
NOR2X1 NOR2X1_179 ( .A(_abc_40298_new_n1601_), .B(_abc_40298_new_n1599_), .Y(_abc_40298_new_n1602_));
NOR2X1 NOR2X1_18 ( .A(_abc_40298_new_n636_), .B(_abc_40298_new_n657_), .Y(_abc_40298_new_n682_));
NOR2X1 NOR2X1_180 ( .A(pc_q_16_), .B(REGFILE_SIM_reg_bank_rb_i_3_), .Y(_abc_40298_new_n1603_));
NOR2X1 NOR2X1_181 ( .A(_abc_40298_new_n1587_), .B(_abc_40298_new_n1604_), .Y(_abc_40298_new_n1605_));
NOR2X1 NOR2X1_182 ( .A(_abc_40298_new_n1603_), .B(_abc_40298_new_n1605_), .Y(_abc_40298_new_n1606_));
NOR2X1 NOR2X1_183 ( .A(pc_q_17_), .B(REGFILE_SIM_reg_bank_rb_i_4_), .Y(_abc_40298_new_n1627_));
NOR2X1 NOR2X1_184 ( .A(_abc_40298_new_n1620_), .B(_abc_40298_new_n1628_), .Y(_abc_40298_new_n1629_));
NOR2X1 NOR2X1_185 ( .A(_abc_40298_new_n1627_), .B(_abc_40298_new_n1629_), .Y(_abc_40298_new_n1630_));
NOR2X1 NOR2X1_186 ( .A(_abc_40298_new_n1607_), .B(_abc_40298_new_n1602_), .Y(_abc_40298_new_n1632_));
NOR2X1 NOR2X1_187 ( .A(_abc_40298_new_n1605_), .B(_abc_40298_new_n1632_), .Y(_abc_40298_new_n1633_));
NOR2X1 NOR2X1_188 ( .A(_abc_40298_new_n1607_), .B(_abc_40298_new_n1631_), .Y(_abc_40298_new_n1653_));
NOR2X1 NOR2X1_189 ( .A(pc_q_18_), .B(REGFILE_SIM_reg_bank_ra_i_0_), .Y(_abc_40298_new_n1657_));
NOR2X1 NOR2X1_19 ( .A(_abc_40298_new_n636_), .B(_abc_40298_new_n659_), .Y(_abc_40298_new_n684_));
NOR2X1 NOR2X1_190 ( .A(_abc_40298_new_n1644_), .B(_abc_40298_new_n1658_), .Y(_abc_40298_new_n1659_));
NOR2X1 NOR2X1_191 ( .A(_abc_40298_new_n1657_), .B(_abc_40298_new_n1659_), .Y(_abc_40298_new_n1660_));
NOR2X1 NOR2X1_192 ( .A(_abc_40298_new_n1661_), .B(_abc_40298_new_n1656_), .Y(_abc_40298_new_n1662_));
NOR2X1 NOR2X1_193 ( .A(pc_q_19_), .B(_abc_40298_new_n1646_), .Y(_abc_40298_new_n1674_));
NOR2X1 NOR2X1_194 ( .A(_abc_40298_new_n1674_), .B(_abc_40298_new_n1676_), .Y(_abc_40298_new_n1677_));
NOR2X1 NOR2X1_195 ( .A(pc_q_19_), .B(REGFILE_SIM_reg_bank_ra_i_1_), .Y(_abc_40298_new_n1682_));
NOR2X1 NOR2X1_196 ( .A(_abc_40298_new_n1675_), .B(_abc_40298_new_n1683_), .Y(_abc_40298_new_n1684_));
NOR2X1 NOR2X1_197 ( .A(_abc_40298_new_n1682_), .B(_abc_40298_new_n1684_), .Y(_abc_40298_new_n1685_));
NOR2X1 NOR2X1_198 ( .A(pc_q_20_), .B(REGFILE_SIM_reg_bank_ra_i_2_), .Y(_abc_40298_new_n1711_));
NOR2X1 NOR2X1_199 ( .A(_abc_40298_new_n1697_), .B(_abc_40298_new_n1712_), .Y(_abc_40298_new_n1713_));
NOR2X1 NOR2X1_2 ( .A(inst_r_2_), .B(_abc_40298_new_n619_), .Y(_abc_40298_new_n620_));
NOR2X1 NOR2X1_20 ( .A(_abc_40298_new_n755_), .B(_abc_40298_new_n685_), .Y(_abc_40298_new_n804_));
NOR2X1 NOR2X1_200 ( .A(_abc_40298_new_n1711_), .B(_abc_40298_new_n1713_), .Y(_abc_40298_new_n1714_));
NOR2X1 NOR2X1_201 ( .A(pc_q_21_), .B(REGFILE_SIM_reg_bank_ra_i_3_), .Y(_abc_40298_new_n1734_));
NOR2X1 NOR2X1_202 ( .A(_abc_40298_new_n1726_), .B(_abc_40298_new_n1735_), .Y(_abc_40298_new_n1736_));
NOR2X1 NOR2X1_203 ( .A(_abc_40298_new_n1737_), .B(_abc_40298_new_n1715_), .Y(_abc_40298_new_n1738_));
NOR2X1 NOR2X1_204 ( .A(_abc_40298_new_n1734_), .B(_abc_40298_new_n1736_), .Y(_abc_40298_new_n1740_));
NOR2X1 NOR2X1_205 ( .A(pc_q_22_), .B(REGFILE_SIM_reg_bank_ra_i_4_), .Y(_abc_40298_new_n1765_));
NOR2X1 NOR2X1_206 ( .A(_abc_40298_new_n1753_), .B(_abc_40298_new_n1766_), .Y(_abc_40298_new_n1767_));
NOR2X1 NOR2X1_207 ( .A(_abc_40298_new_n1765_), .B(_abc_40298_new_n1767_), .Y(_abc_40298_new_n1768_));
NOR2X1 NOR2X1_208 ( .A(_abc_40298_new_n1769_), .B(_abc_40298_new_n1764_), .Y(_abc_40298_new_n1770_));
NOR2X1 NOR2X1_209 ( .A(pc_q_23_), .B(_abc_40298_new_n1755_), .Y(_abc_40298_new_n1782_));
NOR2X1 NOR2X1_21 ( .A(_abc_40298_new_n805_), .B(_abc_40298_new_n686_), .Y(_abc_40298_new_n806_));
NOR2X1 NOR2X1_210 ( .A(_abc_40298_new_n1782_), .B(_abc_40298_new_n1784_), .Y(_abc_40298_new_n1785_));
NOR2X1 NOR2X1_211 ( .A(_abc_40298_new_n1767_), .B(_abc_40298_new_n1770_), .Y(_abc_40298_new_n1789_));
NOR2X1 NOR2X1_212 ( .A(opcode_q_21_), .B(pc_q_23_), .Y(_abc_40298_new_n1790_));
NOR2X1 NOR2X1_213 ( .A(_abc_40298_new_n949_), .B(_abc_40298_new_n1783_), .Y(_abc_40298_new_n1791_));
NOR2X1 NOR2X1_214 ( .A(_abc_40298_new_n1790_), .B(_abc_40298_new_n1791_), .Y(_abc_40298_new_n1792_));
NOR2X1 NOR2X1_215 ( .A(_abc_40298_new_n1741_), .B(_abc_40298_new_n1812_), .Y(_abc_40298_new_n1813_));
NOR2X1 NOR2X1_216 ( .A(_abc_40298_new_n1818_), .B(_abc_40298_new_n1709_), .Y(_abc_40298_new_n1819_));
NOR2X1 NOR2X1_217 ( .A(opcode_q_22_), .B(pc_q_24_), .Y(_abc_40298_new_n1822_));
NOR2X1 NOR2X1_218 ( .A(_abc_40298_new_n944_), .B(_abc_40298_new_n1805_), .Y(_abc_40298_new_n1823_));
NOR2X1 NOR2X1_219 ( .A(_abc_40298_new_n1822_), .B(_abc_40298_new_n1823_), .Y(_abc_40298_new_n1824_));
NOR2X1 NOR2X1_22 ( .A(_abc_40298_new_n810_), .B(_abc_40298_new_n686_), .Y(_abc_40298_new_n811_));
NOR2X1 NOR2X1_220 ( .A(_abc_40298_new_n1824_), .B(_abc_40298_new_n1821_), .Y(_abc_40298_new_n1825_));
NOR2X1 NOR2X1_221 ( .A(opcode_q_23_), .B(pc_q_25_), .Y(_abc_40298_new_n1843_));
NOR2X1 NOR2X1_222 ( .A(_abc_40298_new_n938_), .B(_abc_40298_new_n1844_), .Y(_abc_40298_new_n1845_));
NOR2X1 NOR2X1_223 ( .A(_abc_40298_new_n1843_), .B(_abc_40298_new_n1845_), .Y(_abc_40298_new_n1846_));
NOR2X1 NOR2X1_224 ( .A(_abc_40298_new_n1176_), .B(_abc_40298_new_n1850_), .Y(_abc_40298_new_n1851_));
NOR2X1 NOR2X1_225 ( .A(_abc_40298_new_n1827_), .B(_abc_40298_new_n1869_), .Y(_abc_40298_new_n1870_));
NOR2X1 NOR2X1_226 ( .A(_abc_40298_new_n1847_), .B(_abc_40298_new_n1869_), .Y(_abc_40298_new_n1871_));
NOR2X1 NOR2X1_227 ( .A(_abc_40298_new_n1845_), .B(_abc_40298_new_n1871_), .Y(_abc_40298_new_n1872_));
NOR2X1 NOR2X1_228 ( .A(opcode_q_24_), .B(pc_q_26_), .Y(_abc_40298_new_n1875_));
NOR2X1 NOR2X1_229 ( .A(_abc_40298_new_n623_), .B(_abc_40298_new_n1862_), .Y(_abc_40298_new_n1876_));
NOR2X1 NOR2X1_23 ( .A(_abc_40298_new_n815_), .B(_abc_40298_new_n686_), .Y(_abc_40298_new_n816_));
NOR2X1 NOR2X1_230 ( .A(_abc_40298_new_n1875_), .B(_abc_40298_new_n1876_), .Y(_abc_40298_new_n1877_));
NOR2X1 NOR2X1_231 ( .A(opcode_q_25_), .B(pc_q_27_), .Y(_abc_40298_new_n1894_));
NOR2X1 NOR2X1_232 ( .A(_abc_40298_new_n624_), .B(_abc_40298_new_n1895_), .Y(_abc_40298_new_n1896_));
NOR2X1 NOR2X1_233 ( .A(_abc_40298_new_n1894_), .B(_abc_40298_new_n1896_), .Y(_abc_40298_new_n1897_));
NOR2X1 NOR2X1_234 ( .A(_abc_40298_new_n1917_), .B(_abc_40298_new_n1878_), .Y(_abc_40298_new_n1918_));
NOR2X1 NOR2X1_235 ( .A(opcode_q_25_), .B(pc_q_28_), .Y(_abc_40298_new_n1926_));
NOR2X1 NOR2X1_236 ( .A(_abc_40298_new_n624_), .B(_abc_40298_new_n1911_), .Y(_abc_40298_new_n1927_));
NOR2X1 NOR2X1_237 ( .A(_abc_40298_new_n1926_), .B(_abc_40298_new_n1927_), .Y(_abc_40298_new_n1928_));
NOR2X1 NOR2X1_238 ( .A(_abc_40298_new_n1928_), .B(_abc_40298_new_n1925_), .Y(_abc_40298_new_n1929_));
NOR2X1 NOR2X1_239 ( .A(_abc_40298_new_n1927_), .B(_abc_40298_new_n1930_), .Y(_abc_40298_new_n1943_));
NOR2X1 NOR2X1_24 ( .A(_abc_40298_new_n820_), .B(_abc_40298_new_n686_), .Y(_abc_40298_new_n821_));
NOR2X1 NOR2X1_240 ( .A(_abc_40298_new_n1960_), .B(_abc_40298_new_n1913_), .Y(_abc_40298_new_n1963_));
NOR2X1 NOR2X1_241 ( .A(pc_q_30_), .B(_abc_40298_new_n624_), .Y(_abc_40298_new_n1972_));
NOR2X1 NOR2X1_242 ( .A(opcode_q_25_), .B(_abc_40298_new_n1961_), .Y(_abc_40298_new_n1973_));
NOR2X1 NOR2X1_243 ( .A(_abc_40298_new_n1972_), .B(_abc_40298_new_n1973_), .Y(_abc_40298_new_n1974_));
NOR2X1 NOR2X1_244 ( .A(_abc_40298_new_n1134_), .B(_abc_40298_new_n1027_), .Y(_abc_40298_new_n2014_));
NOR2X1 NOR2X1_245 ( .A(_abc_40298_new_n1166_), .B(_abc_40298_new_n2026_), .Y(_0pc_q_31_0__3_));
NOR2X1 NOR2X1_246 ( .A(_abc_40298_new_n1166_), .B(_abc_40298_new_n2032_), .Y(_0pc_q_31_0__5_));
NOR2X1 NOR2X1_247 ( .A(_abc_40298_new_n1166_), .B(_abc_40298_new_n2038_), .Y(_0pc_q_31_0__7_));
NOR2X1 NOR2X1_248 ( .A(_abc_40298_new_n1166_), .B(_abc_40298_new_n2052_), .Y(_0pc_q_31_0__10_));
NOR2X1 NOR2X1_249 ( .A(_abc_40298_new_n1166_), .B(_abc_40298_new_n2059_), .Y(_0pc_q_31_0__12_));
NOR2X1 NOR2X1_25 ( .A(_abc_40298_new_n825_), .B(_abc_40298_new_n686_), .Y(_abc_40298_new_n826_));
NOR2X1 NOR2X1_250 ( .A(_abc_40298_new_n1166_), .B(_abc_40298_new_n2071_), .Y(_0pc_q_31_0__16_));
NOR2X1 NOR2X1_251 ( .A(_abc_40298_new_n1166_), .B(_abc_40298_new_n2095_), .Y(_0pc_q_31_0__24_));
NOR2X1 NOR2X1_252 ( .A(_abc_40298_new_n1166_), .B(_abc_40298_new_n2098_), .Y(_0pc_q_31_0__25_));
NOR2X1 NOR2X1_253 ( .A(_abc_40298_new_n1166_), .B(_abc_40298_new_n2101_), .Y(_0pc_q_31_0__26_));
NOR2X1 NOR2X1_254 ( .A(_abc_40298_new_n916_), .B(_abc_40298_new_n2119_), .Y(_abc_40298_new_n2120_));
NOR2X1 NOR2X1_255 ( .A(_abc_40298_new_n1455_), .B(_abc_40298_new_n2124_), .Y(_abc_40298_new_n2125_));
NOR2X1 NOR2X1_256 ( .A(_abc_40298_new_n662_), .B(_abc_40298_new_n1017_), .Y(_abc_40298_new_n2127_));
NOR2X1 NOR2X1_257 ( .A(_abc_40298_new_n2132_), .B(_abc_40298_new_n2130_), .Y(_0ex_rd_q_4_0__1_));
NOR2X1 NOR2X1_258 ( .A(_abc_40298_new_n2134_), .B(_abc_40298_new_n2130_), .Y(_0ex_rd_q_4_0__2_));
NOR2X1 NOR2X1_259 ( .A(_abc_40298_new_n2137_), .B(_abc_40298_new_n2130_), .Y(_0ex_rd_q_4_0__4_));
NOR2X1 NOR2X1_26 ( .A(_abc_40298_new_n830_), .B(_abc_40298_new_n686_), .Y(_abc_40298_new_n831_));
NOR2X1 NOR2X1_260 ( .A(alu_op_r_4_), .B(_abc_40298_new_n956_), .Y(_abc_40298_new_n2142_));
NOR2X1 NOR2X1_261 ( .A(_abc_40298_new_n959_), .B(_abc_40298_new_n2145_), .Y(_abc_40298_new_n2146_));
NOR2X1 NOR2X1_262 ( .A(_abc_40298_new_n2149_), .B(_abc_40298_new_n916_), .Y(_abc_40298_new_n2150_));
NOR2X1 NOR2X1_263 ( .A(_abc_40298_new_n891_), .B(_abc_40298_new_n2164_), .Y(_abc_40298_new_n2165_));
NOR2X1 NOR2X1_264 ( .A(_abc_40298_new_n910_), .B(_abc_40298_new_n908_), .Y(_abc_40298_new_n2166_));
NOR2X1 NOR2X1_265 ( .A(_abc_40298_new_n891_), .B(_abc_40298_new_n913_), .Y(_abc_40298_new_n2169_));
NOR2X1 NOR2X1_266 ( .A(_abc_40298_new_n2175_), .B(_abc_40298_new_n2172_), .Y(_abc_40298_new_n2176_));
NOR2X1 NOR2X1_267 ( .A(REGFILE_SIM_reg_bank_rb_i_4_), .B(_abc_40298_new_n980_), .Y(_abc_40298_new_n2202_));
NOR2X1 NOR2X1_268 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_16_), .B(_abc_40298_new_n2147_), .Y(_abc_40298_new_n2206_));
NOR2X1 NOR2X1_269 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_17_), .B(_abc_40298_new_n2147_), .Y(_abc_40298_new_n2211_));
NOR2X1 NOR2X1_27 ( .A(_abc_40298_new_n835_), .B(_abc_40298_new_n686_), .Y(_abc_40298_new_n836_));
NOR2X1 NOR2X1_270 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_18_), .B(_abc_40298_new_n2147_), .Y(_abc_40298_new_n2216_));
NOR2X1 NOR2X1_271 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_19_), .B(_abc_40298_new_n2147_), .Y(_abc_40298_new_n2221_));
NOR2X1 NOR2X1_272 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_20_), .B(_abc_40298_new_n2147_), .Y(_abc_40298_new_n2226_));
NOR2X1 NOR2X1_273 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_21_), .B(_abc_40298_new_n2147_), .Y(_abc_40298_new_n2231_));
NOR2X1 NOR2X1_274 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_22_), .B(_abc_40298_new_n2147_), .Y(_abc_40298_new_n2236_));
NOR2X1 NOR2X1_275 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_23_), .B(_abc_40298_new_n2147_), .Y(_abc_40298_new_n2241_));
NOR2X1 NOR2X1_276 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_24_), .B(_abc_40298_new_n2147_), .Y(_abc_40298_new_n2246_));
NOR2X1 NOR2X1_277 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_25_), .B(_abc_40298_new_n2147_), .Y(_abc_40298_new_n2250_));
NOR2X1 NOR2X1_278 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_26_), .B(_abc_40298_new_n2147_), .Y(_abc_40298_new_n2254_));
NOR2X1 NOR2X1_279 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_27_), .B(_abc_40298_new_n2147_), .Y(_abc_40298_new_n2258_));
NOR2X1 NOR2X1_28 ( .A(_abc_40298_new_n840_), .B(_abc_40298_new_n686_), .Y(_abc_40298_new_n841_));
NOR2X1 NOR2X1_280 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_28_), .B(_abc_40298_new_n2147_), .Y(_abc_40298_new_n2263_));
NOR2X1 NOR2X1_281 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_29_), .B(_abc_40298_new_n2147_), .Y(_abc_40298_new_n2268_));
NOR2X1 NOR2X1_282 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_30_), .B(_abc_40298_new_n2147_), .Y(_abc_40298_new_n2272_));
NOR2X1 NOR2X1_283 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_31_), .B(_abc_40298_new_n2147_), .Y(_abc_40298_new_n2276_));
NOR2X1 NOR2X1_284 ( .A(_abc_40298_new_n2283_), .B(_abc_40298_new_n2284_), .Y(_abc_40298_new_n2285_));
NOR2X1 NOR2X1_285 ( .A(_abc_40298_new_n1188_), .B(_abc_40298_new_n1002_), .Y(_abc_40298_new_n2287_));
NOR2X1 NOR2X1_286 ( .A(_abc_40298_new_n1200_), .B(_abc_40298_new_n1002_), .Y(_abc_40298_new_n2294_));
NOR2X1 NOR2X1_287 ( .A(_abc_40298_new_n657_), .B(_abc_40298_new_n958_), .Y(_abc_40298_new_n2500_));
NOR2X1 NOR2X1_288 ( .A(_abc_40298_new_n2500_), .B(_abc_40298_new_n2283_), .Y(_abc_40298_new_n2507_));
NOR2X1 NOR2X1_289 ( .A(_abc_40298_new_n1046_), .B(_abc_40298_new_n2514_), .Y(_abc_40298_new_n2515_));
NOR2X1 NOR2X1_29 ( .A(_abc_40298_new_n845_), .B(_abc_40298_new_n686_), .Y(_abc_40298_new_n846_));
NOR2X1 NOR2X1_290 ( .A(_abc_40298_new_n1050_), .B(_abc_40298_new_n2519_), .Y(_abc_40298_new_n2520_));
NOR2X1 NOR2X1_291 ( .A(_abc_40298_new_n630_), .B(_abc_40298_new_n666_), .Y(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2420));
NOR2X1 NOR2X1_292 ( .A(inst_r_0_), .B(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2420), .Y(_abc_40298_new_n2559_));
NOR2X1 NOR2X1_293 ( .A(inst_r_2_), .B(_abc_27663_auto_fsm_map_cc_118_implement_pattern_cache_2420), .Y(_abc_40298_new_n2562_));
NOR2X1 NOR2X1_294 ( .A(_abc_40298_new_n646_), .B(_abc_40298_new_n2568_), .Y(_abc_40298_new_n2571_));
NOR2X1 NOR2X1_295 ( .A(_abc_40298_new_n635_), .B(_abc_40298_new_n662_), .Y(_abc_40298_new_n2576_));
NOR2X1 NOR2X1_296 ( .A(_abc_40298_new_n659_), .B(_abc_40298_new_n2568_), .Y(_abc_40298_new_n2578_));
NOR2X1 NOR2X1_297 ( .A(_abc_40298_new_n2580_), .B(_abc_40298_new_n2579_), .Y(_abc_40298_new_n2581_));
NOR2X1 NOR2X1_298 ( .A(_abc_40298_new_n2581_), .B(_abc_40298_new_n2577_), .Y(_abc_40298_new_n2582_));
NOR2X1 NOR2X1_299 ( .A(_abc_40298_new_n2520_), .B(_abc_40298_new_n2579_), .Y(_abc_40298_new_n2597_));
NOR2X1 NOR2X1_3 ( .A(_abc_40298_new_n618_), .B(_abc_40298_new_n621_), .Y(_abc_40298_new_n622_));
NOR2X1 NOR2X1_30 ( .A(_abc_40298_new_n850_), .B(_abc_40298_new_n686_), .Y(_abc_40298_new_n851_));
NOR2X1 NOR2X1_300 ( .A(_abc_40298_new_n2597_), .B(_abc_40298_new_n2577_), .Y(_abc_40298_new_n2598_));
NOR2X1 NOR2X1_301 ( .A(_abc_40298_new_n640_), .B(_abc_40298_new_n683_), .Y(_abc_40298_new_n2611_));
NOR2X1 NOR2X1_302 ( .A(state_q_5_), .B(state_q_3_), .Y(_abc_40298_new_n2883_));
NOR2X1 NOR2X1_303 ( .A(state_q_5_), .B(_abc_40298_new_n630_), .Y(_abc_40298_new_n2891_));
NOR2X1 NOR2X1_304 ( .A(_abc_40298_new_n2299_), .B(_abc_40298_new_n898_), .Y(_abc_40298_new_n2904_));
NOR2X1 NOR2X1_305 ( .A(_abc_40298_new_n1056_), .B(_abc_40298_new_n2904_), .Y(_abc_40298_new_n2905_));
NOR2X1 NOR2X1_306 ( .A(_abc_40298_new_n2904_), .B(_abc_40298_new_n2907_), .Y(_abc_40298_new_n2911_));
NOR2X1 NOR2X1_307 ( .A(_abc_40298_new_n2307_), .B(_abc_40298_new_n903_), .Y(_abc_40298_new_n2912_));
NOR2X1 NOR2X1_308 ( .A(_abc_40298_new_n1055_), .B(_abc_40298_new_n2912_), .Y(_abc_40298_new_n2914_));
NOR2X1 NOR2X1_309 ( .A(_abc_40298_new_n2314_), .B(_abc_40298_new_n1315_), .Y(_abc_40298_new_n2920_));
NOR2X1 NOR2X1_31 ( .A(_abc_40298_new_n855_), .B(_abc_40298_new_n686_), .Y(_abc_40298_new_n856_));
NOR2X1 NOR2X1_310 ( .A(_abc_40298_new_n1048_), .B(_abc_40298_new_n2920_), .Y(_abc_40298_new_n2921_));
NOR2X1 NOR2X1_311 ( .A(_abc_40298_new_n2321_), .B(_abc_40298_new_n1341_), .Y(_abc_40298_new_n2929_));
NOR2X1 NOR2X1_312 ( .A(_abc_40298_new_n1044_), .B(_abc_40298_new_n2929_), .Y(_abc_40298_new_n2930_));
NOR2X1 NOR2X1_313 ( .A(_abc_40298_new_n2930_), .B(_abc_40298_new_n2928_), .Y(_abc_40298_new_n2931_));
NOR2X1 NOR2X1_314 ( .A(_abc_40298_new_n2934_), .B(_abc_40298_new_n2931_), .Y(_abc_40298_new_n2935_));
NOR2X1 NOR2X1_315 ( .A(_abc_40298_new_n663_), .B(_abc_40298_new_n2935_), .Y(_abc_40298_new_n2936_));
NOR2X1 NOR2X1_316 ( .A(_abc_40298_new_n2929_), .B(_abc_40298_new_n2934_), .Y(_abc_40298_new_n2940_));
NOR2X1 NOR2X1_317 ( .A(_abc_40298_new_n2327_), .B(_abc_40298_new_n917_), .Y(_abc_40298_new_n2941_));
NOR2X1 NOR2X1_318 ( .A(_abc_40298_new_n1053_), .B(_abc_40298_new_n2941_), .Y(_abc_40298_new_n2943_));
NOR2X1 NOR2X1_319 ( .A(_abc_40298_new_n2334_), .B(_abc_40298_new_n973_), .Y(_abc_40298_new_n2948_));
NOR2X1 NOR2X1_32 ( .A(_abc_40298_new_n860_), .B(_abc_40298_new_n686_), .Y(_abc_40298_new_n861_));
NOR2X1 NOR2X1_320 ( .A(_abc_40298_new_n1052_), .B(_abc_40298_new_n2948_), .Y(_abc_40298_new_n2949_));
NOR2X1 NOR2X1_321 ( .A(_abc_40298_new_n2342_), .B(_abc_40298_new_n1455_), .Y(_abc_40298_new_n2961_));
NOR2X1 NOR2X1_322 ( .A(_abc_40298_new_n1031_), .B(_abc_40298_new_n2961_), .Y(_abc_40298_new_n2962_));
NOR2X1 NOR2X1_323 ( .A(_abc_40298_new_n2962_), .B(_abc_40298_new_n2960_), .Y(_abc_40298_new_n2963_));
NOR2X1 NOR2X1_324 ( .A(_abc_40298_new_n2352_), .B(_abc_40298_new_n1457_), .Y(_abc_40298_new_n2969_));
NOR2X1 NOR2X1_325 ( .A(_abc_40298_new_n1032_), .B(_abc_40298_new_n2969_), .Y(_abc_40298_new_n2970_));
NOR2X1 NOR2X1_326 ( .A(_abc_40298_new_n663_), .B(_abc_40298_new_n2971_), .Y(_abc_40298_new_n2972_));
NOR2X1 NOR2X1_327 ( .A(_abc_40298_new_n2358_), .B(_abc_40298_new_n2456_), .Y(_abc_40298_new_n2976_));
NOR2X1 NOR2X1_328 ( .A(_abc_40298_new_n1040_), .B(_abc_40298_new_n2976_), .Y(_abc_40298_new_n2977_));
NOR2X1 NOR2X1_329 ( .A(_abc_40298_new_n2969_), .B(_abc_40298_new_n2968_), .Y(_abc_40298_new_n2978_));
NOR2X1 NOR2X1_33 ( .A(_abc_40298_new_n865_), .B(_abc_40298_new_n686_), .Y(_abc_40298_new_n866_));
NOR2X1 NOR2X1_330 ( .A(_abc_40298_new_n1032_), .B(_abc_40298_new_n2978_), .Y(_abc_40298_new_n2979_));
NOR2X1 NOR2X1_331 ( .A(_abc_40298_new_n2994_), .B(_abc_40298_new_n2995_), .Y(_abc_40298_new_n2996_));
NOR2X1 NOR2X1_332 ( .A(_abc_40298_new_n1038_), .B(_abc_40298_new_n2988_), .Y(_abc_40298_new_n2998_));
NOR2X1 NOR2X1_333 ( .A(_abc_40298_new_n663_), .B(_abc_40298_new_n3027_), .Y(_abc_40298_new_n3028_));
NOR2X1 NOR2X1_334 ( .A(_abc_40298_new_n3041_), .B(_abc_40298_new_n3026_), .Y(_abc_40298_new_n3046_));
NOR2X1 NOR2X1_335 ( .A(_abc_40298_new_n3004_), .B(_abc_40298_new_n3015_), .Y(_abc_40298_new_n3049_));
NOR2X1 NOR2X1_336 ( .A(_abc_40298_new_n3055_), .B(_abc_40298_new_n3051_), .Y(_abc_40298_new_n3056_));
NOR2X1 NOR2X1_337 ( .A(_abc_40298_new_n3054_), .B(_abc_40298_new_n3062_), .Y(_abc_40298_new_n3068_));
NOR2X1 NOR2X1_338 ( .A(_abc_40298_new_n3066_), .B(_abc_40298_new_n3076_), .Y(_abc_40298_new_n3082_));
NOR2X1 NOR2X1_339 ( .A(_abc_40298_new_n3083_), .B(_abc_40298_new_n3057_), .Y(_abc_40298_new_n3084_));
NOR2X1 NOR2X1_34 ( .A(_abc_40298_new_n870_), .B(_abc_40298_new_n686_), .Y(_abc_40298_new_n871_));
NOR2X1 NOR2X1_340 ( .A(_abc_40298_new_n3088_), .B(_abc_40298_new_n3084_), .Y(_abc_40298_new_n3089_));
NOR2X1 NOR2X1_341 ( .A(_abc_40298_new_n3092_), .B(_abc_40298_new_n3098_), .Y(_abc_40298_new_n3106_));
NOR2X1 NOR2X1_342 ( .A(_abc_40298_new_n3104_), .B(_abc_40298_new_n3108_), .Y(_abc_40298_new_n3109_));
NOR2X1 NOR2X1_343 ( .A(_abc_40298_new_n3083_), .B(_abc_40298_new_n3125_), .Y(_abc_40298_new_n3127_));
NOR2X1 NOR2X1_344 ( .A(_abc_40298_new_n3139_), .B(_abc_40298_new_n3140_), .Y(_abc_40298_new_n3141_));
NOR2X1 NOR2X1_345 ( .A(_abc_40298_new_n3130_), .B(_abc_40298_new_n3138_), .Y(_abc_40298_new_n3145_));
NOR2X1 NOR2X1_346 ( .A(_abc_40298_new_n3166_), .B(_abc_40298_new_n3165_), .Y(_abc_40298_new_n3167_));
NOR2X1 NOR2X1_347 ( .A(_abc_40298_new_n3173_), .B(_abc_40298_new_n3181_), .Y(_abc_40298_new_n3182_));
NOR2X1 NOR2X1_348 ( .A(_abc_40298_new_n3198_), .B(_abc_40298_new_n1170_), .Y(_0nmi_q_0_0_));
NOR2X1 NOR2X1_349 ( .A(_abc_40298_new_n1166_), .B(_abc_40298_new_n3200_), .Y(_0fault_o_0_0_));
NOR2X1 NOR2X1_35 ( .A(_abc_40298_new_n875_), .B(_abc_40298_new_n686_), .Y(_abc_40298_new_n876_));
NOR2X1 NOR2X1_350 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2101_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2102_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2103_));
NOR2X1 NOR2X1_351 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2101_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2203_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2204_));
NOR2X1 NOR2X1_352 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2101_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2270_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2271_));
NOR2X1 NOR2X1_353 ( .A(REGFILE_SIM_reg_bank_rd_i_0_), .B(REGFILE_SIM_reg_bank_rd_i_1_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2337_));
NOR2X1 NOR2X1_354 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2102_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2405_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2406_));
NOR2X1 NOR2X1_355 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2203_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2405_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2472_));
NOR2X1 NOR2X1_356 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2270_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2405_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2538_));
NOR2X1 NOR2X1_357 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2405_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2338_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2603_));
NOR2X1 NOR2X1_358 ( .A(REGFILE_SIM_reg_bank_reg_r24_0_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2604_));
NOR2X1 NOR2X1_359 ( .A(REGFILE_SIM_reg_bank_reg_r24_1_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2606_));
NOR2X1 NOR2X1_36 ( .A(_abc_40298_new_n880_), .B(_abc_40298_new_n686_), .Y(_abc_40298_new_n881_));
NOR2X1 NOR2X1_360 ( .A(REGFILE_SIM_reg_bank_reg_r24_2_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2608_));
NOR2X1 NOR2X1_361 ( .A(REGFILE_SIM_reg_bank_reg_r24_3_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2610_));
NOR2X1 NOR2X1_362 ( .A(REGFILE_SIM_reg_bank_reg_r24_4_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2612_));
NOR2X1 NOR2X1_363 ( .A(REGFILE_SIM_reg_bank_reg_r24_5_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2614_));
NOR2X1 NOR2X1_364 ( .A(REGFILE_SIM_reg_bank_reg_r24_6_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2616_));
NOR2X1 NOR2X1_365 ( .A(REGFILE_SIM_reg_bank_reg_r24_7_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2618_));
NOR2X1 NOR2X1_366 ( .A(REGFILE_SIM_reg_bank_reg_r24_8_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2620_));
NOR2X1 NOR2X1_367 ( .A(REGFILE_SIM_reg_bank_reg_r24_9_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2622_));
NOR2X1 NOR2X1_368 ( .A(REGFILE_SIM_reg_bank_reg_r24_10_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2624_));
NOR2X1 NOR2X1_369 ( .A(REGFILE_SIM_reg_bank_reg_r24_11_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2626_));
NOR2X1 NOR2X1_37 ( .A(nmi_q), .B(nmi_i), .Y(_abc_40298_new_n885_));
NOR2X1 NOR2X1_370 ( .A(REGFILE_SIM_reg_bank_reg_r24_12_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2628_));
NOR2X1 NOR2X1_371 ( .A(REGFILE_SIM_reg_bank_reg_r24_13_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2630_));
NOR2X1 NOR2X1_372 ( .A(REGFILE_SIM_reg_bank_reg_r24_14_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2632_));
NOR2X1 NOR2X1_373 ( .A(REGFILE_SIM_reg_bank_reg_r24_15_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2634_));
NOR2X1 NOR2X1_374 ( .A(REGFILE_SIM_reg_bank_reg_r24_16_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2636_));
NOR2X1 NOR2X1_375 ( .A(REGFILE_SIM_reg_bank_reg_r24_17_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2638_));
NOR2X1 NOR2X1_376 ( .A(REGFILE_SIM_reg_bank_reg_r24_18_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2640_));
NOR2X1 NOR2X1_377 ( .A(REGFILE_SIM_reg_bank_reg_r24_19_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2642_));
NOR2X1 NOR2X1_378 ( .A(REGFILE_SIM_reg_bank_reg_r24_20_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2644_));
NOR2X1 NOR2X1_379 ( .A(REGFILE_SIM_reg_bank_reg_r24_21_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2646_));
NOR2X1 NOR2X1_38 ( .A(opcode_q_24_), .B(_abc_40298_new_n626_), .Y(_abc_40298_new_n886_));
NOR2X1 NOR2X1_380 ( .A(REGFILE_SIM_reg_bank_reg_r24_22_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2648_));
NOR2X1 NOR2X1_381 ( .A(REGFILE_SIM_reg_bank_reg_r24_23_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2650_));
NOR2X1 NOR2X1_382 ( .A(REGFILE_SIM_reg_bank_reg_r24_24_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2652_));
NOR2X1 NOR2X1_383 ( .A(REGFILE_SIM_reg_bank_reg_r24_25_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2654_));
NOR2X1 NOR2X1_384 ( .A(REGFILE_SIM_reg_bank_reg_r24_26_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2656_));
NOR2X1 NOR2X1_385 ( .A(REGFILE_SIM_reg_bank_reg_r24_27_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2658_));
NOR2X1 NOR2X1_386 ( .A(REGFILE_SIM_reg_bank_reg_r24_28_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2660_));
NOR2X1 NOR2X1_387 ( .A(REGFILE_SIM_reg_bank_reg_r24_29_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2662_));
NOR2X1 NOR2X1_388 ( .A(REGFILE_SIM_reg_bank_reg_r24_30_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2664_));
NOR2X1 NOR2X1_389 ( .A(REGFILE_SIM_reg_bank_reg_r24_31_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2603_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2666_));
NOR2X1 NOR2X1_39 ( .A(alu_op_r_4_), .B(alu_op_r_5_), .Y(_abc_40298_new_n889_));
NOR2X1 NOR2X1_390 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2102_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2669_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2670_));
NOR2X1 NOR2X1_391 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2669_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2203_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2736_));
NOR2X1 NOR2X1_392 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2270_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2669_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2802_));
NOR2X1 NOR2X1_393 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2669_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2338_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2868_));
NOR2X1 NOR2X1_394 ( .A(REGFILE_SIM_reg_bank_rd_i_3_), .B(REGFILE_SIM_reg_bank_rd_i_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2933_));
NOR2X1 NOR2X1_395 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2102_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2934_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2935_));
NOR2X1 NOR2X1_396 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2104_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3001_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3002_));
NOR2X1 NOR2X1_397 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2104_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3067_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3068_));
NOR2X1 NOR2X1_398 ( .A(REGFILE_SIM_reg_bank_rd_i_4_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3198_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3199_));
NOR2X1 NOR2X1_399 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2101_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3395_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3396_));
NOR2X1 NOR2X1_4 ( .A(inst_r_1_), .B(inst_r_0_), .Y(_abc_40298_new_n625_));
NOR2X1 NOR2X1_40 ( .A(alu_op_r_6_), .B(alu_op_r_7_), .Y(_abc_40298_new_n890_));
NOR2X1 NOR2X1_400 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3591_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3067_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3592_));
NOR2X1 NOR2X1_401 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2405_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3395_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3722_));
NOR2X1 NOR2X1_402 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2669_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3395_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3982_));
NOR2X1 NOR2X1_403 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3591_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n3001_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4112_));
NOR2X1 NOR2X1_404 ( .A(REGFILE_SIM_reg_bank_rb_i_1_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4176_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4177_));
NOR2X1 NOR2X1_405 ( .A(REGFILE_SIM_reg_bank_rb_i_2_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4181_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4182_));
NOR2X1 NOR2X1_406 ( .A(REGFILE_SIM_reg_bank_rb_i_0_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4188_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4189_));
NOR2X1 NOR2X1_407 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4186_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4191_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4192_));
NOR2X1 NOR2X1_408 ( .A(REGFILE_SIM_reg_bank_rb_i_3_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4193_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4194_));
NOR2X1 NOR2X1_409 ( .A(REGFILE_SIM_reg_bank_rb_i_3_), .B(REGFILE_SIM_reg_bank_rb_i_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4200_));
NOR2X1 NOR2X1_41 ( .A(alu_op_r_0_), .B(alu_op_r_1_), .Y(_abc_40298_new_n893_));
NOR2X1 NOR2X1_410 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4203_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4199_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4204_));
NOR2X1 NOR2X1_411 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4196_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4178_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4209_));
NOR2X1 NOR2X1_412 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4212_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4208_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4213_));
NOR2X1 NOR2X1_413 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4217_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4220_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4221_));
NOR2X1 NOR2X1_414 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4222_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4205_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4223_));
NOR2X1 NOR2X1_415 ( .A(REGFILE_SIM_reg_bank_rb_i_1_), .B(REGFILE_SIM_reg_bank_rb_i_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4225_));
NOR2X1 NOR2X1_416 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4230_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4227_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4231_));
NOR2X1 NOR2X1_417 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4232_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4233_));
NOR2X1 NOR2X1_418 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4241_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4244_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4245_));
NOR2X1 NOR2X1_419 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4248_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4251_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4252_));
NOR2X1 NOR2X1_42 ( .A(_abc_40298_new_n651_), .B(_abc_40298_new_n896_), .Y(_abc_40298_new_n897_));
NOR2X1 NOR2X1_420 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4238_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4253_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4254_));
NOR2X1 NOR2X1_421 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4257_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4258_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4259_));
NOR2X1 NOR2X1_422 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4261_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4260_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4262_));
NOR2X1 NOR2X1_423 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4266_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4264_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4267_));
NOR2X1 NOR2X1_424 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4268_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4269_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4270_));
NOR2X1 NOR2X1_425 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4271_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4263_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4272_));
NOR2X1 NOR2X1_426 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4274_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4273_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4275_));
NOR2X1 NOR2X1_427 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4279_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4280_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4281_));
NOR2X1 NOR2X1_428 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4282_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4283_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4284_));
NOR2X1 NOR2X1_429 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4278_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4285_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4286_));
NOR2X1 NOR2X1_43 ( .A(alu_op_r_3_), .B(_abc_40298_new_n898_), .Y(_abc_40298_new_n899_));
NOR2X1 NOR2X1_430 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4289_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4290_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4291_));
NOR2X1 NOR2X1_431 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4293_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4292_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4294_));
NOR2X1 NOR2X1_432 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4298_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4296_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4299_));
NOR2X1 NOR2X1_433 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4300_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4301_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4302_));
NOR2X1 NOR2X1_434 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4303_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4295_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4304_));
NOR2X1 NOR2X1_435 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4306_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4305_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4307_));
NOR2X1 NOR2X1_436 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4311_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4312_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4313_));
NOR2X1 NOR2X1_437 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4314_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4315_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4316_));
NOR2X1 NOR2X1_438 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4310_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4317_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4318_));
NOR2X1 NOR2X1_439 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4321_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4322_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4323_));
NOR2X1 NOR2X1_44 ( .A(alu_op_r_2_), .B(alu_op_r_3_), .Y(_abc_40298_new_n901_));
NOR2X1 NOR2X1_440 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4325_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4324_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4326_));
NOR2X1 NOR2X1_441 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4330_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4328_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4331_));
NOR2X1 NOR2X1_442 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4332_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4333_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4334_));
NOR2X1 NOR2X1_443 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4335_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4327_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4336_));
NOR2X1 NOR2X1_444 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4338_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4337_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4339_));
NOR2X1 NOR2X1_445 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4343_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4344_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4345_));
NOR2X1 NOR2X1_446 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4346_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4347_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4348_));
NOR2X1 NOR2X1_447 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4342_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4349_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4350_));
NOR2X1 NOR2X1_448 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4353_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4354_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4355_));
NOR2X1 NOR2X1_449 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4357_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4356_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4358_));
NOR2X1 NOR2X1_45 ( .A(alu_op_r_2_), .B(_abc_40298_new_n903_), .Y(_abc_40298_new_n904_));
NOR2X1 NOR2X1_450 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4362_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4360_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4363_));
NOR2X1 NOR2X1_451 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4364_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4365_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4366_));
NOR2X1 NOR2X1_452 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4367_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4359_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4368_));
NOR2X1 NOR2X1_453 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4370_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4369_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4371_));
NOR2X1 NOR2X1_454 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4375_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4376_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4377_));
NOR2X1 NOR2X1_455 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4378_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4379_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4380_));
NOR2X1 NOR2X1_456 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4374_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4381_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4382_));
NOR2X1 NOR2X1_457 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4385_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4386_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4387_));
NOR2X1 NOR2X1_458 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4389_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4388_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4390_));
NOR2X1 NOR2X1_459 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4394_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4392_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4395_));
NOR2X1 NOR2X1_46 ( .A(_abc_40298_new_n891_), .B(_abc_40298_new_n906_), .Y(_abc_40298_new_n907_));
NOR2X1 NOR2X1_460 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4396_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4397_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4398_));
NOR2X1 NOR2X1_461 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4399_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4391_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4400_));
NOR2X1 NOR2X1_462 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4402_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4401_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4403_));
NOR2X1 NOR2X1_463 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4407_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4408_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4409_));
NOR2X1 NOR2X1_464 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4410_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4411_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4412_));
NOR2X1 NOR2X1_465 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4406_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4413_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4414_));
NOR2X1 NOR2X1_466 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4417_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4418_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4419_));
NOR2X1 NOR2X1_467 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4421_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4420_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4422_));
NOR2X1 NOR2X1_468 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4426_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4424_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4427_));
NOR2X1 NOR2X1_469 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4428_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4429_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4430_));
NOR2X1 NOR2X1_47 ( .A(_abc_40298_new_n911_), .B(_abc_40298_new_n909_), .Y(_abc_40298_new_n912_));
NOR2X1 NOR2X1_470 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4431_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4423_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4432_));
NOR2X1 NOR2X1_471 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4434_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4433_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4435_));
NOR2X1 NOR2X1_472 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4439_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4440_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4441_));
NOR2X1 NOR2X1_473 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4442_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4443_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4444_));
NOR2X1 NOR2X1_474 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4438_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4445_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4446_));
NOR2X1 NOR2X1_475 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4449_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4450_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4451_));
NOR2X1 NOR2X1_476 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4453_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4452_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4454_));
NOR2X1 NOR2X1_477 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4458_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4456_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4459_));
NOR2X1 NOR2X1_478 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4460_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4461_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4462_));
NOR2X1 NOR2X1_479 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4463_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4455_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4464_));
NOR2X1 NOR2X1_48 ( .A(alu_op_r_5_), .B(_abc_40298_new_n917_), .Y(_abc_40298_new_n918_));
NOR2X1 NOR2X1_480 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4466_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4465_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4467_));
NOR2X1 NOR2X1_481 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4471_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4472_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4473_));
NOR2X1 NOR2X1_482 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4474_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4475_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4476_));
NOR2X1 NOR2X1_483 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4470_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4477_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4478_));
NOR2X1 NOR2X1_484 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4481_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4482_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4483_));
NOR2X1 NOR2X1_485 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4485_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4484_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4486_));
NOR2X1 NOR2X1_486 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4490_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4488_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4491_));
NOR2X1 NOR2X1_487 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4492_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4493_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4494_));
NOR2X1 NOR2X1_488 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4495_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4487_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4496_));
NOR2X1 NOR2X1_489 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4498_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4497_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4499_));
NOR2X1 NOR2X1_49 ( .A(_abc_40298_new_n919_), .B(_abc_40298_new_n920_), .Y(_abc_40298_new_n921_));
NOR2X1 NOR2X1_490 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4503_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4504_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4505_));
NOR2X1 NOR2X1_491 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4506_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4507_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4508_));
NOR2X1 NOR2X1_492 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4502_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4509_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4510_));
NOR2X1 NOR2X1_493 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4513_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4514_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4515_));
NOR2X1 NOR2X1_494 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4517_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4516_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4518_));
NOR2X1 NOR2X1_495 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4522_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4520_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4523_));
NOR2X1 NOR2X1_496 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4524_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4525_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4526_));
NOR2X1 NOR2X1_497 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4527_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4519_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4528_));
NOR2X1 NOR2X1_498 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4530_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4529_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4531_));
NOR2X1 NOR2X1_499 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4535_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4536_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4537_));
NOR2X1 NOR2X1_5 ( .A(_abc_40298_new_n623_), .B(_abc_40298_new_n626_), .Y(_abc_40298_new_n627_));
NOR2X1 NOR2X1_50 ( .A(_abc_40298_new_n923_), .B(_abc_40298_new_n908_), .Y(_abc_40298_new_n924_));
NOR2X1 NOR2X1_500 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4538_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4539_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4540_));
NOR2X1 NOR2X1_501 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4534_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4541_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4542_));
NOR2X1 NOR2X1_502 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4545_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4546_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4547_));
NOR2X1 NOR2X1_503 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4549_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4548_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4550_));
NOR2X1 NOR2X1_504 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4554_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4552_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4555_));
NOR2X1 NOR2X1_505 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4556_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4557_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4558_));
NOR2X1 NOR2X1_506 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4559_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4551_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4560_));
NOR2X1 NOR2X1_507 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4562_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4561_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4563_));
NOR2X1 NOR2X1_508 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4567_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4568_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4569_));
NOR2X1 NOR2X1_509 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4570_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4571_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4572_));
NOR2X1 NOR2X1_51 ( .A(_abc_40298_new_n910_), .B(_abc_40298_new_n925_), .Y(_abc_40298_new_n926_));
NOR2X1 NOR2X1_510 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4566_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4573_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4574_));
NOR2X1 NOR2X1_511 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4577_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4578_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4579_));
NOR2X1 NOR2X1_512 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4581_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4580_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4582_));
NOR2X1 NOR2X1_513 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4586_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4584_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4587_));
NOR2X1 NOR2X1_514 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4588_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4589_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4590_));
NOR2X1 NOR2X1_515 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4591_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4583_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4592_));
NOR2X1 NOR2X1_516 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4594_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4593_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4595_));
NOR2X1 NOR2X1_517 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4599_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4600_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4601_));
NOR2X1 NOR2X1_518 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4602_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4603_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4604_));
NOR2X1 NOR2X1_519 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4598_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4605_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4606_));
NOR2X1 NOR2X1_52 ( .A(_abc_40298_new_n646_), .B(_abc_40298_new_n929_), .Y(_abc_40298_new_n930_));
NOR2X1 NOR2X1_520 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4609_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4610_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4611_));
NOR2X1 NOR2X1_521 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4613_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4612_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4614_));
NOR2X1 NOR2X1_522 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4618_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4616_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4619_));
NOR2X1 NOR2X1_523 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4620_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4621_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4622_));
NOR2X1 NOR2X1_524 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4623_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4615_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4624_));
NOR2X1 NOR2X1_525 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4626_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4625_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4627_));
NOR2X1 NOR2X1_526 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4631_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4632_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4633_));
NOR2X1 NOR2X1_527 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4634_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4635_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4636_));
NOR2X1 NOR2X1_528 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4630_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4637_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4638_));
NOR2X1 NOR2X1_529 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4641_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4642_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4643_));
NOR2X1 NOR2X1_53 ( .A(_abc_40298_new_n657_), .B(_abc_40298_new_n896_), .Y(_abc_40298_new_n931_));
NOR2X1 NOR2X1_530 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4645_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4644_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4646_));
NOR2X1 NOR2X1_531 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4650_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4648_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4651_));
NOR2X1 NOR2X1_532 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4652_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4653_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4654_));
NOR2X1 NOR2X1_533 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4655_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4647_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4656_));
NOR2X1 NOR2X1_534 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4658_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4657_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4659_));
NOR2X1 NOR2X1_535 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4663_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4664_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4665_));
NOR2X1 NOR2X1_536 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4666_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4667_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4668_));
NOR2X1 NOR2X1_537 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4662_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4669_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4670_));
NOR2X1 NOR2X1_538 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4673_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4674_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4675_));
NOR2X1 NOR2X1_539 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4677_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4676_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4678_));
NOR2X1 NOR2X1_54 ( .A(_abc_40298_new_n931_), .B(_abc_40298_new_n930_), .Y(_abc_40298_new_n932_));
NOR2X1 NOR2X1_540 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4682_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4680_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4683_));
NOR2X1 NOR2X1_541 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4684_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4685_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4686_));
NOR2X1 NOR2X1_542 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4687_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4679_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4688_));
NOR2X1 NOR2X1_543 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4690_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4689_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4691_));
NOR2X1 NOR2X1_544 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4695_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4696_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4697_));
NOR2X1 NOR2X1_545 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4698_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4699_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4700_));
NOR2X1 NOR2X1_546 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4694_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4701_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4702_));
NOR2X1 NOR2X1_547 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4705_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4706_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4707_));
NOR2X1 NOR2X1_548 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4709_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4708_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4710_));
NOR2X1 NOR2X1_549 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4714_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4712_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4715_));
NOR2X1 NOR2X1_55 ( .A(opcode_q_22_), .B(opcode_q_21_), .Y(_abc_40298_new_n934_));
NOR2X1 NOR2X1_550 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4716_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4717_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4718_));
NOR2X1 NOR2X1_551 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4719_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4711_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4720_));
NOR2X1 NOR2X1_552 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4722_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4721_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4723_));
NOR2X1 NOR2X1_553 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4727_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4728_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4729_));
NOR2X1 NOR2X1_554 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4730_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4731_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4732_));
NOR2X1 NOR2X1_555 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4726_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4733_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4734_));
NOR2X1 NOR2X1_556 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4737_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4738_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4739_));
NOR2X1 NOR2X1_557 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4741_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4740_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4742_));
NOR2X1 NOR2X1_558 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4746_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4744_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4747_));
NOR2X1 NOR2X1_559 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4748_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4749_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4750_));
NOR2X1 NOR2X1_56 ( .A(_abc_40298_new_n935_), .B(_abc_40298_new_n936_), .Y(_abc_40298_new_n937_));
NOR2X1 NOR2X1_560 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4751_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4743_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4752_));
NOR2X1 NOR2X1_561 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4754_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4753_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4755_));
NOR2X1 NOR2X1_562 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4759_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4760_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4761_));
NOR2X1 NOR2X1_563 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4762_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4763_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4764_));
NOR2X1 NOR2X1_564 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4758_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4765_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4766_));
NOR2X1 NOR2X1_565 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4769_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4770_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4771_));
NOR2X1 NOR2X1_566 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4773_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4772_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4774_));
NOR2X1 NOR2X1_567 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4778_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4776_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4779_));
NOR2X1 NOR2X1_568 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4780_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4781_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4782_));
NOR2X1 NOR2X1_569 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4783_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4775_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4784_));
NOR2X1 NOR2X1_57 ( .A(_abc_40298_new_n623_), .B(_abc_40298_new_n938_), .Y(_abc_40298_new_n939_));
NOR2X1 NOR2X1_570 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4786_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4785_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4787_));
NOR2X1 NOR2X1_571 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4791_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4792_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4793_));
NOR2X1 NOR2X1_572 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4794_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4795_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4796_));
NOR2X1 NOR2X1_573 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4790_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4797_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4798_));
NOR2X1 NOR2X1_574 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4801_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4802_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4803_));
NOR2X1 NOR2X1_575 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4805_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4804_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4806_));
NOR2X1 NOR2X1_576 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4810_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4808_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4811_));
NOR2X1 NOR2X1_577 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4812_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4813_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4814_));
NOR2X1 NOR2X1_578 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4815_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4807_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4816_));
NOR2X1 NOR2X1_579 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4818_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4817_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4819_));
NOR2X1 NOR2X1_58 ( .A(opcode_q_21_), .B(_abc_40298_new_n944_), .Y(_abc_40298_new_n945_));
NOR2X1 NOR2X1_580 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4823_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4824_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4825_));
NOR2X1 NOR2X1_581 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4826_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4827_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4828_));
NOR2X1 NOR2X1_582 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4822_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4829_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4830_));
NOR2X1 NOR2X1_583 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4833_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4834_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4835_));
NOR2X1 NOR2X1_584 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4837_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4836_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4838_));
NOR2X1 NOR2X1_585 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4842_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4840_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4843_));
NOR2X1 NOR2X1_586 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4844_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4845_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4846_));
NOR2X1 NOR2X1_587 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4847_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4839_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4848_));
NOR2X1 NOR2X1_588 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4850_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4849_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4851_));
NOR2X1 NOR2X1_589 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4855_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4856_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4857_));
NOR2X1 NOR2X1_59 ( .A(opcode_q_23_), .B(_abc_40298_new_n623_), .Y(_abc_40298_new_n946_));
NOR2X1 NOR2X1_590 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4858_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4859_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4860_));
NOR2X1 NOR2X1_591 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4854_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4861_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4862_));
NOR2X1 NOR2X1_592 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4865_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4866_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4867_));
NOR2X1 NOR2X1_593 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4869_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4868_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4870_));
NOR2X1 NOR2X1_594 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4874_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4872_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4875_));
NOR2X1 NOR2X1_595 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4876_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4877_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4878_));
NOR2X1 NOR2X1_596 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4879_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4871_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4880_));
NOR2X1 NOR2X1_597 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4882_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4881_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4883_));
NOR2X1 NOR2X1_598 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4887_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4888_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4889_));
NOR2X1 NOR2X1_599 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4890_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4891_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4892_));
NOR2X1 NOR2X1_6 ( .A(_abc_40298_new_n637_), .B(_abc_40298_new_n638_), .Y(_abc_40298_new_n639_));
NOR2X1 NOR2X1_60 ( .A(_abc_40298_new_n947_), .B(_abc_40298_new_n943_), .Y(_abc_40298_new_n948_));
NOR2X1 NOR2X1_600 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4886_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4893_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4894_));
NOR2X1 NOR2X1_601 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4897_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4898_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4899_));
NOR2X1 NOR2X1_602 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4901_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4900_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4902_));
NOR2X1 NOR2X1_603 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4906_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4904_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4907_));
NOR2X1 NOR2X1_604 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4908_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4909_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4910_));
NOR2X1 NOR2X1_605 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4911_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4903_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4912_));
NOR2X1 NOR2X1_606 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4914_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4913_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4915_));
NOR2X1 NOR2X1_607 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4919_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4920_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4921_));
NOR2X1 NOR2X1_608 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4922_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4923_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4924_));
NOR2X1 NOR2X1_609 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4918_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4925_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4926_));
NOR2X1 NOR2X1_61 ( .A(opcode_q_22_), .B(_abc_40298_new_n949_), .Y(_abc_40298_new_n950_));
NOR2X1 NOR2X1_610 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4929_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4930_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4931_));
NOR2X1 NOR2X1_611 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4933_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4932_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4934_));
NOR2X1 NOR2X1_612 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4938_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4936_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4939_));
NOR2X1 NOR2X1_613 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4940_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4941_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4942_));
NOR2X1 NOR2X1_614 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4943_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4935_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4944_));
NOR2X1 NOR2X1_615 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4946_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4945_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4947_));
NOR2X1 NOR2X1_616 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4951_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4952_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4953_));
NOR2X1 NOR2X1_617 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4954_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4955_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4956_));
NOR2X1 NOR2X1_618 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4950_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4957_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4958_));
NOR2X1 NOR2X1_619 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4961_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4962_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4963_));
NOR2X1 NOR2X1_62 ( .A(_abc_40298_new_n916_), .B(_abc_40298_new_n953_), .Y(_abc_40298_new_n954_));
NOR2X1 NOR2X1_620 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4965_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4964_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4966_));
NOR2X1 NOR2X1_621 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4970_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4968_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4971_));
NOR2X1 NOR2X1_622 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4972_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4973_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4974_));
NOR2X1 NOR2X1_623 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4975_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4967_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4976_));
NOR2X1 NOR2X1_624 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4978_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4977_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4979_));
NOR2X1 NOR2X1_625 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4983_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4984_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4985_));
NOR2X1 NOR2X1_626 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4986_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4987_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4988_));
NOR2X1 NOR2X1_627 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4982_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4989_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4990_));
NOR2X1 NOR2X1_628 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4993_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4994_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4995_));
NOR2X1 NOR2X1_629 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4997_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4996_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4998_));
NOR2X1 NOR2X1_63 ( .A(_abc_40298_new_n659_), .B(_abc_40298_new_n929_), .Y(_abc_40298_new_n955_));
NOR2X1 NOR2X1_630 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5002_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5000_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5003_));
NOR2X1 NOR2X1_631 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5004_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5005_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5006_));
NOR2X1 NOR2X1_632 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5007_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4999_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5008_));
NOR2X1 NOR2X1_633 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5010_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5009_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5011_));
NOR2X1 NOR2X1_634 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5015_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5016_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5017_));
NOR2X1 NOR2X1_635 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5018_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5019_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5020_));
NOR2X1 NOR2X1_636 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5014_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5021_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5022_));
NOR2X1 NOR2X1_637 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5025_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5026_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5027_));
NOR2X1 NOR2X1_638 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5029_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5028_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5030_));
NOR2X1 NOR2X1_639 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5034_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5032_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5035_));
NOR2X1 NOR2X1_64 ( .A(_abc_40298_new_n621_), .B(_abc_40298_new_n645_), .Y(_abc_40298_new_n957_));
NOR2X1 NOR2X1_640 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5036_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5037_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5038_));
NOR2X1 NOR2X1_641 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5039_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5031_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5040_));
NOR2X1 NOR2X1_642 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5042_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5041_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5043_));
NOR2X1 NOR2X1_643 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5047_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5048_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5049_));
NOR2X1 NOR2X1_644 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5050_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5051_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5052_));
NOR2X1 NOR2X1_645 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5046_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5053_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5054_));
NOR2X1 NOR2X1_646 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5057_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5058_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5059_));
NOR2X1 NOR2X1_647 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5061_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5060_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5062_));
NOR2X1 NOR2X1_648 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5066_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5064_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5067_));
NOR2X1 NOR2X1_649 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5068_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5069_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5070_));
NOR2X1 NOR2X1_65 ( .A(_abc_40298_new_n646_), .B(_abc_40298_new_n958_), .Y(_abc_40298_new_n959_));
NOR2X1 NOR2X1_650 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5071_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5063_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5072_));
NOR2X1 NOR2X1_651 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5074_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5073_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5075_));
NOR2X1 NOR2X1_652 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5079_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5080_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5081_));
NOR2X1 NOR2X1_653 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5082_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5083_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5084_));
NOR2X1 NOR2X1_654 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5078_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5085_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5086_));
NOR2X1 NOR2X1_655 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5089_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5090_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5091_));
NOR2X1 NOR2X1_656 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5093_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5092_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5094_));
NOR2X1 NOR2X1_657 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5098_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5096_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5099_));
NOR2X1 NOR2X1_658 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5100_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5101_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5102_));
NOR2X1 NOR2X1_659 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5103_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5095_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5104_));
NOR2X1 NOR2X1_66 ( .A(_abc_40298_new_n963_), .B(_abc_40298_new_n932_), .Y(_abc_40298_new_n964_));
NOR2X1 NOR2X1_660 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5106_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5105_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5107_));
NOR2X1 NOR2X1_661 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5111_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5112_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5113_));
NOR2X1 NOR2X1_662 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5114_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5115_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5116_));
NOR2X1 NOR2X1_663 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5110_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5117_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5118_));
NOR2X1 NOR2X1_664 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5121_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5122_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5123_));
NOR2X1 NOR2X1_665 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5125_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5124_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5126_));
NOR2X1 NOR2X1_666 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5130_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5128_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5131_));
NOR2X1 NOR2X1_667 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5132_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5133_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5134_));
NOR2X1 NOR2X1_668 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5135_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5127_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5136_));
NOR2X1 NOR2X1_669 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5138_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5137_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5139_));
NOR2X1 NOR2X1_67 ( .A(_abc_40298_new_n945_), .B(_abc_40298_new_n950_), .Y(_abc_40298_new_n965_));
NOR2X1 NOR2X1_670 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5143_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5144_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5145_));
NOR2X1 NOR2X1_671 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5146_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5147_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5148_));
NOR2X1 NOR2X1_672 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5142_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5149_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5150_));
NOR2X1 NOR2X1_673 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5153_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5154_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5155_));
NOR2X1 NOR2X1_674 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5157_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5156_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5158_));
NOR2X1 NOR2X1_675 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5162_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5160_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5163_));
NOR2X1 NOR2X1_676 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5164_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5165_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5166_));
NOR2X1 NOR2X1_677 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5167_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5159_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5168_));
NOR2X1 NOR2X1_678 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5170_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5169_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5171_));
NOR2X1 NOR2X1_679 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5175_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5176_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5177_));
NOR2X1 NOR2X1_68 ( .A(opcode_q_24_), .B(_abc_40298_new_n938_), .Y(_abc_40298_new_n967_));
NOR2X1 NOR2X1_680 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5178_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5179_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5180_));
NOR2X1 NOR2X1_681 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5174_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5181_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5182_));
NOR2X1 NOR2X1_682 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5185_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5186_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5187_));
NOR2X1 NOR2X1_683 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5189_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5188_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5190_));
NOR2X1 NOR2X1_684 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5194_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5192_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5195_));
NOR2X1 NOR2X1_685 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5196_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5197_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5198_));
NOR2X1 NOR2X1_686 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5199_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5191_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5200_));
NOR2X1 NOR2X1_687 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5202_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5201_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5203_));
NOR2X1 NOR2X1_688 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5207_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5208_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5209_));
NOR2X1 NOR2X1_689 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5210_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5211_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5212_));
NOR2X1 NOR2X1_69 ( .A(alu_op_r_4_), .B(_abc_40298_new_n973_), .Y(_abc_40298_new_n974_));
NOR2X1 NOR2X1_690 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5206_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5213_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5214_));
NOR2X1 NOR2X1_691 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5217_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5218_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5219_));
NOR2X1 NOR2X1_692 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5221_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5220_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5222_));
NOR2X1 NOR2X1_693 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5226_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5224_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5227_));
NOR2X1 NOR2X1_694 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5228_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5229_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5230_));
NOR2X1 NOR2X1_695 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5231_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5223_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5232_));
NOR2X1 NOR2X1_696 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5234_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5233_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5235_));
NOR2X1 NOR2X1_697 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5239_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5240_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5241_));
NOR2X1 NOR2X1_698 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5242_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5243_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5244_));
NOR2X1 NOR2X1_699 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5238_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5245_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5246_));
NOR2X1 NOR2X1_7 ( .A(_abc_40298_new_n636_), .B(_abc_40298_new_n640_), .Y(_abc_40298_new_n641_));
NOR2X1 NOR2X1_70 ( .A(_abc_40298_new_n975_), .B(_abc_40298_new_n920_), .Y(_abc_40298_new_n976_));
NOR2X1 NOR2X1_700 ( .A(REGFILE_SIM_reg_bank_ra_i_1_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5248_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5249_));
NOR2X1 NOR2X1_701 ( .A(REGFILE_SIM_reg_bank_ra_i_2_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5253_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5254_));
NOR2X1 NOR2X1_702 ( .A(REGFILE_SIM_reg_bank_ra_i_0_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5260_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5261_));
NOR2X1 NOR2X1_703 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5258_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5263_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5264_));
NOR2X1 NOR2X1_704 ( .A(REGFILE_SIM_reg_bank_ra_i_3_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5265_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5266_));
NOR2X1 NOR2X1_705 ( .A(REGFILE_SIM_reg_bank_ra_i_3_), .B(REGFILE_SIM_reg_bank_ra_i_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5272_));
NOR2X1 NOR2X1_706 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5275_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5271_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5276_));
NOR2X1 NOR2X1_707 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5268_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5250_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5281_));
NOR2X1 NOR2X1_708 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5284_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5280_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5285_));
NOR2X1 NOR2X1_709 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5289_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5292_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5293_));
NOR2X1 NOR2X1_71 ( .A(_abc_40298_new_n636_), .B(_abc_40298_new_n645_), .Y(_abc_40298_new_n979_));
NOR2X1 NOR2X1_710 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5294_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5277_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5295_));
NOR2X1 NOR2X1_711 ( .A(REGFILE_SIM_reg_bank_ra_i_1_), .B(REGFILE_SIM_reg_bank_ra_i_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5297_));
NOR2X1 NOR2X1_712 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5302_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5299_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5303_));
NOR2X1 NOR2X1_713 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5304_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5305_));
NOR2X1 NOR2X1_714 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5313_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5316_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5317_));
NOR2X1 NOR2X1_715 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5320_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5323_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5324_));
NOR2X1 NOR2X1_716 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5310_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5325_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5326_));
NOR2X1 NOR2X1_717 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5329_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5330_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5331_));
NOR2X1 NOR2X1_718 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5333_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5332_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5334_));
NOR2X1 NOR2X1_719 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5338_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5336_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5339_));
NOR2X1 NOR2X1_72 ( .A(_abc_40298_new_n986_), .B(_abc_40298_new_n989_), .Y(_abc_40298_new_n990_));
NOR2X1 NOR2X1_720 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5340_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5341_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5342_));
NOR2X1 NOR2X1_721 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5343_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5335_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5344_));
NOR2X1 NOR2X1_722 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5346_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5345_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5347_));
NOR2X1 NOR2X1_723 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5351_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5352_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5353_));
NOR2X1 NOR2X1_724 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5354_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5355_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5356_));
NOR2X1 NOR2X1_725 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5350_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5357_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5358_));
NOR2X1 NOR2X1_726 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5361_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5362_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5363_));
NOR2X1 NOR2X1_727 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5365_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5364_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5366_));
NOR2X1 NOR2X1_728 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5370_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5368_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5371_));
NOR2X1 NOR2X1_729 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5372_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5373_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5374_));
NOR2X1 NOR2X1_73 ( .A(_abc_40298_new_n651_), .B(_abc_40298_new_n648_), .Y(_abc_40298_new_n991_));
NOR2X1 NOR2X1_730 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5375_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5367_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5376_));
NOR2X1 NOR2X1_731 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5378_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5377_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5379_));
NOR2X1 NOR2X1_732 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5383_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5384_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5385_));
NOR2X1 NOR2X1_733 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5386_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5387_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5388_));
NOR2X1 NOR2X1_734 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5382_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5389_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5390_));
NOR2X1 NOR2X1_735 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5393_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5394_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5395_));
NOR2X1 NOR2X1_736 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5397_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5396_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5398_));
NOR2X1 NOR2X1_737 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5402_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5400_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5403_));
NOR2X1 NOR2X1_738 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5404_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5405_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5406_));
NOR2X1 NOR2X1_739 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5407_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5399_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5408_));
NOR2X1 NOR2X1_74 ( .A(_abc_40298_new_n618_), .B(_abc_40298_new_n648_), .Y(_abc_40298_new_n994_));
NOR2X1 NOR2X1_740 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5410_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5409_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5411_));
NOR2X1 NOR2X1_741 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5415_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5416_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5417_));
NOR2X1 NOR2X1_742 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5418_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5419_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5420_));
NOR2X1 NOR2X1_743 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5414_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5421_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5422_));
NOR2X1 NOR2X1_744 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5425_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5426_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5427_));
NOR2X1 NOR2X1_745 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5429_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5428_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5430_));
NOR2X1 NOR2X1_746 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5434_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5432_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5435_));
NOR2X1 NOR2X1_747 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5436_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5437_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5438_));
NOR2X1 NOR2X1_748 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5439_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5431_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5440_));
NOR2X1 NOR2X1_749 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5442_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5441_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5443_));
NOR2X1 NOR2X1_75 ( .A(_abc_40298_new_n660_), .B(_abc_40298_new_n995_), .Y(_abc_40298_new_n996_));
NOR2X1 NOR2X1_750 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5447_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5448_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5449_));
NOR2X1 NOR2X1_751 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5450_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5451_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5452_));
NOR2X1 NOR2X1_752 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5446_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5453_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5454_));
NOR2X1 NOR2X1_753 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5457_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5458_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5459_));
NOR2X1 NOR2X1_754 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5461_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5460_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5462_));
NOR2X1 NOR2X1_755 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5466_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5464_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5467_));
NOR2X1 NOR2X1_756 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5468_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5469_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5470_));
NOR2X1 NOR2X1_757 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5471_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5463_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5472_));
NOR2X1 NOR2X1_758 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5474_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5473_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5475_));
NOR2X1 NOR2X1_759 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5479_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5480_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5481_));
NOR2X1 NOR2X1_76 ( .A(_abc_40298_new_n993_), .B(_abc_40298_new_n996_), .Y(_abc_40298_new_n997_));
NOR2X1 NOR2X1_760 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5482_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5483_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5484_));
NOR2X1 NOR2X1_761 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5478_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5485_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5486_));
NOR2X1 NOR2X1_762 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5489_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5490_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5491_));
NOR2X1 NOR2X1_763 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5493_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5492_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5494_));
NOR2X1 NOR2X1_764 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5498_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5496_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5499_));
NOR2X1 NOR2X1_765 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5500_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5501_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5502_));
NOR2X1 NOR2X1_766 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5503_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5495_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5504_));
NOR2X1 NOR2X1_767 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5506_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5505_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5507_));
NOR2X1 NOR2X1_768 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5511_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5512_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5513_));
NOR2X1 NOR2X1_769 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5514_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5515_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5516_));
NOR2X1 NOR2X1_77 ( .A(_abc_40298_new_n657_), .B(_abc_40298_new_n648_), .Y(_abc_40298_new_n998_));
NOR2X1 NOR2X1_770 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5510_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5517_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5518_));
NOR2X1 NOR2X1_771 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5521_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5522_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5523_));
NOR2X1 NOR2X1_772 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5525_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5524_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5526_));
NOR2X1 NOR2X1_773 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5530_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5528_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5531_));
NOR2X1 NOR2X1_774 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5532_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5533_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5534_));
NOR2X1 NOR2X1_775 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5535_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5527_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5536_));
NOR2X1 NOR2X1_776 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5538_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5537_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5539_));
NOR2X1 NOR2X1_777 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5543_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5544_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5545_));
NOR2X1 NOR2X1_778 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5546_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5547_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5548_));
NOR2X1 NOR2X1_779 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5542_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5549_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5550_));
NOR2X1 NOR2X1_78 ( .A(inst_r_5_), .B(_abc_40298_new_n637_), .Y(_abc_40298_new_n999_));
NOR2X1 NOR2X1_780 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5553_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5554_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5555_));
NOR2X1 NOR2X1_781 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5557_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5556_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5558_));
NOR2X1 NOR2X1_782 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5562_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5560_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5563_));
NOR2X1 NOR2X1_783 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5564_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5565_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5566_));
NOR2X1 NOR2X1_784 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5567_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5559_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5568_));
NOR2X1 NOR2X1_785 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5570_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5569_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5571_));
NOR2X1 NOR2X1_786 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5575_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5576_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5577_));
NOR2X1 NOR2X1_787 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5578_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5579_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5580_));
NOR2X1 NOR2X1_788 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5574_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5581_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5582_));
NOR2X1 NOR2X1_789 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5585_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5586_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5587_));
NOR2X1 NOR2X1_79 ( .A(_abc_40298_new_n657_), .B(_abc_40298_new_n929_), .Y(_abc_40298_new_n1001_));
NOR2X1 NOR2X1_790 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5589_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5588_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5590_));
NOR2X1 NOR2X1_791 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5594_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5592_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5595_));
NOR2X1 NOR2X1_792 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5596_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5597_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5598_));
NOR2X1 NOR2X1_793 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5599_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5591_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5600_));
NOR2X1 NOR2X1_794 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5602_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5601_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5603_));
NOR2X1 NOR2X1_795 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5607_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5608_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5609_));
NOR2X1 NOR2X1_796 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5610_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5611_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5612_));
NOR2X1 NOR2X1_797 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5606_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5613_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5614_));
NOR2X1 NOR2X1_798 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5617_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5618_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5619_));
NOR2X1 NOR2X1_799 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5621_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5620_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5622_));
NOR2X1 NOR2X1_8 ( .A(inst_r_4_), .B(_abc_40298_new_n638_), .Y(_abc_40298_new_n644_));
NOR2X1 NOR2X1_80 ( .A(_abc_40298_new_n1000_), .B(_abc_40298_new_n1004_), .Y(_abc_40298_new_n1005_));
NOR2X1 NOR2X1_800 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5626_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5624_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5627_));
NOR2X1 NOR2X1_801 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5628_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5629_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5630_));
NOR2X1 NOR2X1_802 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5631_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5623_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5632_));
NOR2X1 NOR2X1_803 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5634_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5633_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5635_));
NOR2X1 NOR2X1_804 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5639_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5640_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5641_));
NOR2X1 NOR2X1_805 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5642_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5643_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5644_));
NOR2X1 NOR2X1_806 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5638_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5645_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5646_));
NOR2X1 NOR2X1_807 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5649_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5650_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5651_));
NOR2X1 NOR2X1_808 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5653_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5652_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5654_));
NOR2X1 NOR2X1_809 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5658_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5656_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5659_));
NOR2X1 NOR2X1_81 ( .A(_abc_40298_new_n944_), .B(_abc_40298_new_n949_), .Y(_abc_40298_new_n1006_));
NOR2X1 NOR2X1_810 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5660_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5661_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5662_));
NOR2X1 NOR2X1_811 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5663_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5655_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5664_));
NOR2X1 NOR2X1_812 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5666_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5665_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5667_));
NOR2X1 NOR2X1_813 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5671_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5672_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5673_));
NOR2X1 NOR2X1_814 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5674_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5675_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5676_));
NOR2X1 NOR2X1_815 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5670_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5677_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5678_));
NOR2X1 NOR2X1_816 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5681_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5682_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5683_));
NOR2X1 NOR2X1_817 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5685_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5684_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5686_));
NOR2X1 NOR2X1_818 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5690_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5688_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5691_));
NOR2X1 NOR2X1_819 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5692_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5693_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5694_));
NOR2X1 NOR2X1_82 ( .A(_abc_40298_new_n1007_), .B(_abc_40298_new_n943_), .Y(_abc_40298_new_n1008_));
NOR2X1 NOR2X1_820 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5695_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5687_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5696_));
NOR2X1 NOR2X1_821 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5698_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5697_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5699_));
NOR2X1 NOR2X1_822 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5703_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5704_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5705_));
NOR2X1 NOR2X1_823 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5706_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5707_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5708_));
NOR2X1 NOR2X1_824 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5702_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5709_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5710_));
NOR2X1 NOR2X1_825 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5713_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5714_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5715_));
NOR2X1 NOR2X1_826 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5717_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5716_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5718_));
NOR2X1 NOR2X1_827 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5722_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5720_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5723_));
NOR2X1 NOR2X1_828 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5724_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5725_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5726_));
NOR2X1 NOR2X1_829 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5727_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5719_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5728_));
NOR2X1 NOR2X1_83 ( .A(_abc_40298_new_n648_), .B(_abc_40298_new_n659_), .Y(_abc_40298_new_n1010_));
NOR2X1 NOR2X1_830 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5730_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5729_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5731_));
NOR2X1 NOR2X1_831 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5735_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5736_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5737_));
NOR2X1 NOR2X1_832 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5738_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5739_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5740_));
NOR2X1 NOR2X1_833 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5734_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5741_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5742_));
NOR2X1 NOR2X1_834 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5745_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5746_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5747_));
NOR2X1 NOR2X1_835 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5749_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5748_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5750_));
NOR2X1 NOR2X1_836 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5754_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5752_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5755_));
NOR2X1 NOR2X1_837 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5756_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5757_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5758_));
NOR2X1 NOR2X1_838 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5759_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5751_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5760_));
NOR2X1 NOR2X1_839 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5762_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5761_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5763_));
NOR2X1 NOR2X1_84 ( .A(_abc_40298_new_n659_), .B(_abc_40298_new_n958_), .Y(_abc_40298_new_n1015_));
NOR2X1 NOR2X1_840 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5767_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5768_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5769_));
NOR2X1 NOR2X1_841 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5770_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5771_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5772_));
NOR2X1 NOR2X1_842 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5766_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5773_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5774_));
NOR2X1 NOR2X1_843 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5777_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5778_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5779_));
NOR2X1 NOR2X1_844 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5781_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5780_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5782_));
NOR2X1 NOR2X1_845 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5786_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5784_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5787_));
NOR2X1 NOR2X1_846 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5788_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5789_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5790_));
NOR2X1 NOR2X1_847 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5791_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5783_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5792_));
NOR2X1 NOR2X1_848 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5794_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5793_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5795_));
NOR2X1 NOR2X1_849 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5799_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5800_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5801_));
NOR2X1 NOR2X1_85 ( .A(_abc_40298_new_n1021_), .B(_abc_40298_new_n1019_), .Y(_abc_40298_new_n1022_));
NOR2X1 NOR2X1_850 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5802_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5803_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5804_));
NOR2X1 NOR2X1_851 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5798_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5805_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5806_));
NOR2X1 NOR2X1_852 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5809_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5810_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5811_));
NOR2X1 NOR2X1_853 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5813_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5812_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5814_));
NOR2X1 NOR2X1_854 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5818_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5816_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5819_));
NOR2X1 NOR2X1_855 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5820_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5821_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5822_));
NOR2X1 NOR2X1_856 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5823_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5815_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5824_));
NOR2X1 NOR2X1_857 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5826_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5825_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5827_));
NOR2X1 NOR2X1_858 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5831_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5832_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5833_));
NOR2X1 NOR2X1_859 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5834_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5835_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5836_));
NOR2X1 NOR2X1_86 ( .A(_abc_40298_new_n972_), .B(_abc_40298_new_n1023_), .Y(_abc_40298_new_n1024_));
NOR2X1 NOR2X1_860 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5830_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5837_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5838_));
NOR2X1 NOR2X1_861 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5841_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5842_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5843_));
NOR2X1 NOR2X1_862 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5845_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5844_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5846_));
NOR2X1 NOR2X1_863 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5850_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5848_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5851_));
NOR2X1 NOR2X1_864 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5852_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5853_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5854_));
NOR2X1 NOR2X1_865 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5855_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5847_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5856_));
NOR2X1 NOR2X1_866 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5858_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5857_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5859_));
NOR2X1 NOR2X1_867 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5863_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5864_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5865_));
NOR2X1 NOR2X1_868 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5866_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5867_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5868_));
NOR2X1 NOR2X1_869 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5862_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5869_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5870_));
NOR2X1 NOR2X1_87 ( .A(next_pc_r_1_), .B(next_pc_r_0_), .Y(_abc_40298_new_n1026_));
NOR2X1 NOR2X1_870 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5873_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5874_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5875_));
NOR2X1 NOR2X1_871 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5877_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5876_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5878_));
NOR2X1 NOR2X1_872 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5882_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5880_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5883_));
NOR2X1 NOR2X1_873 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5884_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5885_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5886_));
NOR2X1 NOR2X1_874 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5887_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5879_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5888_));
NOR2X1 NOR2X1_875 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5890_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5889_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5891_));
NOR2X1 NOR2X1_876 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5895_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5896_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5897_));
NOR2X1 NOR2X1_877 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5898_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5899_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5900_));
NOR2X1 NOR2X1_878 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5894_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5901_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5902_));
NOR2X1 NOR2X1_879 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5905_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5906_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5907_));
NOR2X1 NOR2X1_88 ( .A(_abc_40298_new_n888_), .B(_abc_40298_new_n1027_), .Y(_abc_40298_new_n1028_));
NOR2X1 NOR2X1_880 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5909_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5908_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5910_));
NOR2X1 NOR2X1_881 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5914_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5912_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5915_));
NOR2X1 NOR2X1_882 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5916_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5917_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5918_));
NOR2X1 NOR2X1_883 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5919_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5911_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5920_));
NOR2X1 NOR2X1_884 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5922_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5921_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5923_));
NOR2X1 NOR2X1_885 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5927_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5928_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5929_));
NOR2X1 NOR2X1_886 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5930_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5931_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5932_));
NOR2X1 NOR2X1_887 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5926_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5933_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5934_));
NOR2X1 NOR2X1_888 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5937_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5938_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5939_));
NOR2X1 NOR2X1_889 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5941_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5940_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5942_));
NOR2X1 NOR2X1_89 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_8_), .B(alu_op_r_6_), .Y(_abc_40298_new_n1031_));
NOR2X1 NOR2X1_890 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5946_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5944_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5947_));
NOR2X1 NOR2X1_891 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5948_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5949_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5950_));
NOR2X1 NOR2X1_892 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5951_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5943_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5952_));
NOR2X1 NOR2X1_893 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5954_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5953_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5955_));
NOR2X1 NOR2X1_894 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5959_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5960_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5961_));
NOR2X1 NOR2X1_895 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5962_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5963_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5964_));
NOR2X1 NOR2X1_896 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5958_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5965_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5966_));
NOR2X1 NOR2X1_897 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5969_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5970_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5971_));
NOR2X1 NOR2X1_898 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5973_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5972_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5974_));
NOR2X1 NOR2X1_899 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5978_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5976_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5979_));
NOR2X1 NOR2X1_9 ( .A(inst_r_2_), .B(inst_r_3_), .Y(_abc_40298_new_n647_));
NOR2X1 NOR2X1_90 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_9_), .B(alu_op_r_7_), .Y(_abc_40298_new_n1032_));
NOR2X1 NOR2X1_900 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5980_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5981_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5982_));
NOR2X1 NOR2X1_901 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5983_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5975_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5984_));
NOR2X1 NOR2X1_902 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5986_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5985_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5987_));
NOR2X1 NOR2X1_903 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5991_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5992_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5993_));
NOR2X1 NOR2X1_904 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5994_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5995_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5996_));
NOR2X1 NOR2X1_905 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n5990_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5997_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5998_));
NOR2X1 NOR2X1_906 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6001_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6002_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6003_));
NOR2X1 NOR2X1_907 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6005_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6004_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6006_));
NOR2X1 NOR2X1_908 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6010_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6008_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6011_));
NOR2X1 NOR2X1_909 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6012_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6013_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6014_));
NOR2X1 NOR2X1_91 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_10_), .B(int32_r_10_), .Y(_abc_40298_new_n1040_));
NOR2X1 NOR2X1_910 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6015_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6007_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6016_));
NOR2X1 NOR2X1_911 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6018_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6017_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6019_));
NOR2X1 NOR2X1_912 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6023_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6024_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6025_));
NOR2X1 NOR2X1_913 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6026_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6027_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6028_));
NOR2X1 NOR2X1_914 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6022_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6029_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6030_));
NOR2X1 NOR2X1_915 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6033_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6034_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6035_));
NOR2X1 NOR2X1_916 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6037_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6036_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6038_));
NOR2X1 NOR2X1_917 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6042_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6040_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6043_));
NOR2X1 NOR2X1_918 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6044_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6045_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6046_));
NOR2X1 NOR2X1_919 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6047_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6039_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6048_));
NOR2X1 NOR2X1_92 ( .A(_abc_40298_new_n1037_), .B(_abc_40298_new_n1041_), .Y(_abc_40298_new_n1042_));
NOR2X1 NOR2X1_920 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6050_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6049_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6051_));
NOR2X1 NOR2X1_921 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6055_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6056_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6057_));
NOR2X1 NOR2X1_922 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6058_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6059_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6060_));
NOR2X1 NOR2X1_923 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6054_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6061_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6062_));
NOR2X1 NOR2X1_924 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6065_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6066_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6067_));
NOR2X1 NOR2X1_925 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6069_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6068_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6070_));
NOR2X1 NOR2X1_926 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6074_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6072_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6075_));
NOR2X1 NOR2X1_927 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6076_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6077_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6078_));
NOR2X1 NOR2X1_928 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6079_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6071_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6080_));
NOR2X1 NOR2X1_929 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6082_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6081_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6083_));
NOR2X1 NOR2X1_93 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_5_), .B(int32_r_5_), .Y(_abc_40298_new_n1044_));
NOR2X1 NOR2X1_930 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6087_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6088_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6089_));
NOR2X1 NOR2X1_931 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6090_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6091_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6092_));
NOR2X1 NOR2X1_932 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6086_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6093_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6094_));
NOR2X1 NOR2X1_933 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6097_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6098_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6099_));
NOR2X1 NOR2X1_934 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6101_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6100_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6102_));
NOR2X1 NOR2X1_935 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6106_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6104_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6107_));
NOR2X1 NOR2X1_936 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6108_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6109_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6110_));
NOR2X1 NOR2X1_937 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6111_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6103_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6112_));
NOR2X1 NOR2X1_938 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6114_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6113_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6115_));
NOR2X1 NOR2X1_939 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6119_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6120_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6121_));
NOR2X1 NOR2X1_94 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_0_), .B(alu_op_r_0_), .Y(_abc_40298_new_n1046_));
NOR2X1 NOR2X1_940 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6122_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6123_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6124_));
NOR2X1 NOR2X1_941 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6118_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6125_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6126_));
NOR2X1 NOR2X1_942 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6129_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6130_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6131_));
NOR2X1 NOR2X1_943 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6133_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6132_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6134_));
NOR2X1 NOR2X1_944 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6138_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6136_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6139_));
NOR2X1 NOR2X1_945 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6140_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6141_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6142_));
NOR2X1 NOR2X1_946 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6143_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6135_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6144_));
NOR2X1 NOR2X1_947 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6146_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6145_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6147_));
NOR2X1 NOR2X1_948 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6151_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6152_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6153_));
NOR2X1 NOR2X1_949 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6154_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6155_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6156_));
NOR2X1 NOR2X1_95 ( .A(_abc_40298_new_n1046_), .B(_abc_40298_new_n1045_), .Y(_abc_40298_new_n1047_));
NOR2X1 NOR2X1_950 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6150_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6157_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6158_));
NOR2X1 NOR2X1_951 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6161_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6162_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6163_));
NOR2X1 NOR2X1_952 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6165_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6164_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6166_));
NOR2X1 NOR2X1_953 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6170_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6168_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6171_));
NOR2X1 NOR2X1_954 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6172_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6173_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6174_));
NOR2X1 NOR2X1_955 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6175_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6167_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6176_));
NOR2X1 NOR2X1_956 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6178_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6177_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6179_));
NOR2X1 NOR2X1_957 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6183_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6184_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6185_));
NOR2X1 NOR2X1_958 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6186_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6187_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6188_));
NOR2X1 NOR2X1_959 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6182_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6189_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6190_));
NOR2X1 NOR2X1_96 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_4_), .B(int32_r_4_), .Y(_abc_40298_new_n1048_));
NOR2X1 NOR2X1_960 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6193_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6194_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6195_));
NOR2X1 NOR2X1_961 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6197_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6196_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6198_));
NOR2X1 NOR2X1_962 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6202_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6200_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6203_));
NOR2X1 NOR2X1_963 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6204_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6205_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6206_));
NOR2X1 NOR2X1_964 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6207_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6199_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6208_));
NOR2X1 NOR2X1_965 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6210_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6209_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6211_));
NOR2X1 NOR2X1_966 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6215_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6216_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6217_));
NOR2X1 NOR2X1_967 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6218_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6219_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6220_));
NOR2X1 NOR2X1_968 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6214_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6221_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6222_));
NOR2X1 NOR2X1_969 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6225_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6226_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6227_));
NOR2X1 NOR2X1_97 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_1_), .B(alu_op_r_1_), .Y(_abc_40298_new_n1050_));
NOR2X1 NOR2X1_970 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6229_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6228_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6230_));
NOR2X1 NOR2X1_971 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6234_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6232_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6235_));
NOR2X1 NOR2X1_972 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6236_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6237_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6238_));
NOR2X1 NOR2X1_973 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6239_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6231_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6240_));
NOR2X1 NOR2X1_974 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6242_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6241_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6243_));
NOR2X1 NOR2X1_975 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6247_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6248_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6249_));
NOR2X1 NOR2X1_976 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6250_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6251_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6252_));
NOR2X1 NOR2X1_977 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6246_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6253_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6254_));
NOR2X1 NOR2X1_978 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6257_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6258_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6259_));
NOR2X1 NOR2X1_979 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6261_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6260_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6262_));
NOR2X1 NOR2X1_98 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_7_), .B(alu_op_r_5_), .Y(_abc_40298_new_n1052_));
NOR2X1 NOR2X1_980 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6266_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6264_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6267_));
NOR2X1 NOR2X1_981 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6268_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6269_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6270_));
NOR2X1 NOR2X1_982 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6271_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6263_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6272_));
NOR2X1 NOR2X1_983 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6274_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6273_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6275_));
NOR2X1 NOR2X1_984 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6279_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6280_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6281_));
NOR2X1 NOR2X1_985 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6282_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6283_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6284_));
NOR2X1 NOR2X1_986 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6278_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6285_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6286_));
NOR2X1 NOR2X1_987 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6289_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6290_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6291_));
NOR2X1 NOR2X1_988 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6293_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6292_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6294_));
NOR2X1 NOR2X1_989 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6298_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6296_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6299_));
NOR2X1 NOR2X1_99 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_6_), .B(alu_op_r_4_), .Y(_abc_40298_new_n1053_));
NOR2X1 NOR2X1_990 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6300_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6301_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6302_));
NOR2X1 NOR2X1_991 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6303_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6295_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6304_));
NOR2X1 NOR2X1_992 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6306_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6305_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6307_));
NOR2X1 NOR2X1_993 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6311_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6312_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6313_));
NOR2X1 NOR2X1_994 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6314_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6315_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6316_));
NOR2X1 NOR2X1_995 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n6310_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n6317_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6318_));
NOR2X1 NOR2X1_996 ( .A(alu__abc_38674_new_n110_), .B(alu__abc_38674_new_n111_), .Y(alu__abc_38674_new_n112_));
NOR2X1 NOR2X1_997 ( .A(alu_b_i_22_), .B(alu_a_i_22_), .Y(alu__abc_38674_new_n113_));
NOR2X1 NOR2X1_998 ( .A(alu__abc_38674_new_n113_), .B(alu__abc_38674_new_n112_), .Y(alu__abc_38674_new_n114_));
NOR2X1 NOR2X1_999 ( .A(alu__abc_38674_new_n116_), .B(alu__abc_38674_new_n117_), .Y(alu__abc_38674_new_n118_));
NOR3X1 NOR3X1_1 ( .A(_abc_40298_new_n1091_), .B(_abc_40298_new_n1102_), .C(_abc_40298_new_n1100_), .Y(_abc_40298_new_n1103_));
NOR3X1 NOR3X1_10 ( .A(_abc_40298_new_n1726_), .B(_abc_40298_new_n1753_), .C(_abc_40298_new_n1699_), .Y(_abc_40298_new_n1755_));
NOR3X1 NOR3X1_11 ( .A(_abc_40298_new_n1753_), .B(_abc_40298_new_n1783_), .C(_abc_40298_new_n1728_), .Y(_abc_40298_new_n1784_));
NOR3X1 NOR3X1_12 ( .A(_abc_40298_new_n1844_), .B(_abc_40298_new_n1862_), .C(_abc_40298_new_n1807_), .Y(_abc_40298_new_n1864_));
NOR3X1 NOR3X1_13 ( .A(_abc_40298_new_n1862_), .B(_abc_40298_new_n1895_), .C(_abc_40298_new_n2000_), .Y(_abc_40298_new_n2001_));
NOR3X1 NOR3X1_14 ( .A(REGFILE_SIM_reg_bank_rb_i_1_), .B(REGFILE_SIM_reg_bank_rb_i_0_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4183_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4184_));
NOR3X1 NOR3X1_15 ( .A(REGFILE_SIM_reg_bank_rb_i_1_), .B(REGFILE_SIM_reg_bank_rb_i_0_), .C(REGFILE_SIM_reg_bank_rb_i_4_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4215_));
NOR3X1 NOR3X1_16 ( .A(REGFILE_SIM_reg_bank_ra_i_1_), .B(REGFILE_SIM_reg_bank_ra_i_0_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5255_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5256_));
NOR3X1 NOR3X1_17 ( .A(REGFILE_SIM_reg_bank_ra_i_1_), .B(REGFILE_SIM_reg_bank_ra_i_0_), .C(REGFILE_SIM_reg_bank_ra_i_4_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5287_));
NOR3X1 NOR3X1_18 ( .A(alu__abc_38674_new_n547_), .B(alu__abc_38674_new_n552_), .C(alu__abc_38674_new_n572_), .Y(alu__abc_38674_new_n573_));
NOR3X1 NOR3X1_19 ( .A(alu__abc_38674_new_n538_), .B(alu__abc_38674_new_n574_), .C(alu__abc_38674_new_n576_), .Y(alu__abc_38674_new_n577_));
NOR3X1 NOR3X1_2 ( .A(_abc_40298_new_n1287_), .B(_abc_40298_new_n1302_), .C(_abc_40298_new_n1258_), .Y(_abc_40298_new_n1304_));
NOR3X1 NOR3X1_20 ( .A(alu__abc_38674_new_n596_), .B(alu__abc_38674_new_n584_), .C(alu__abc_38674_new_n592_), .Y(alu__abc_38674_new_n597_));
NOR3X1 NOR3X1_21 ( .A(alu__abc_38674_new_n511_), .B(alu__abc_38674_new_n604_), .C(alu__abc_38674_new_n598_), .Y(alu__abc_38674_new_n605_));
NOR3X1 NOR3X1_22 ( .A(alu__abc_38674_new_n1043_), .B(alu__abc_38674_new_n1046_), .C(alu__abc_38674_new_n1047_), .Y(alu__abc_38674_new_n1076_));
NOR3X1 NOR3X1_23 ( .A(alu__abc_38674_new_n1266_), .B(alu__abc_38674_new_n1112_), .C(alu__abc_38674_new_n1269_), .Y(alu__abc_38674_new_n1270_));
NOR3X1 NOR3X1_24 ( .A(alu__abc_38674_new_n1266_), .B(alu__abc_38674_new_n1296_), .C(alu__abc_38674_new_n1294_), .Y(alu__abc_38674_new_n1297_));
NOR3X1 NOR3X1_25 ( .A(alu__abc_38674_new_n1366_), .B(alu__abc_38674_new_n1367_), .C(alu__abc_38674_new_n1381_), .Y(alu__abc_38674_new_n1382_));
NOR3X1 NOR3X1_26 ( .A(alu__abc_38674_new_n1384_), .B(alu__abc_38674_new_n604_), .C(alu__abc_38674_new_n1416_), .Y(alu__abc_38674_new_n1417_));
NOR3X1 NOR3X1_27 ( .A(alu__abc_38674_new_n1358_), .B(alu__abc_38674_new_n1412_), .C(alu__abc_38674_new_n1327_), .Y(alu__abc_38674_new_n1442_));
NOR3X1 NOR3X1_28 ( .A(alu__abc_38674_new_n507_), .B(alu__abc_38674_new_n624_), .C(alu__abc_38674_new_n1472_), .Y(alu__abc_38674_new_n1525_));
NOR3X1 NOR3X1_29 ( .A(alu__abc_38674_new_n507_), .B(alu__abc_38674_new_n504_), .C(alu__abc_38674_new_n1500_), .Y(alu__abc_38674_new_n1547_));
NOR3X1 NOR3X1_3 ( .A(_abc_40298_new_n1302_), .B(_abc_40298_new_n1332_), .C(_abc_40298_new_n1289_), .Y(_abc_40298_new_n1333_));
NOR3X1 NOR3X1_30 ( .A(alu__abc_38674_new_n1384_), .B(alu__abc_38674_new_n1498_), .C(alu__abc_38674_new_n1443_), .Y(alu__abc_38674_new_n1574_));
NOR3X1 NOR3X1_31 ( .A(alu__abc_38674_new_n504_), .B(alu__abc_38674_new_n1573_), .C(alu__abc_38674_new_n1575_), .Y(alu__abc_38674_new_n1576_));
NOR3X1 NOR3X1_32 ( .A(alu__abc_38674_new_n1624_), .B(alu__abc_38674_new_n620_), .C(alu__abc_38674_new_n1602_), .Y(alu__abc_38674_new_n1625_));
NOR3X1 NOR3X1_33 ( .A(alu__abc_38674_new_n1649_), .B(alu__abc_38674_new_n1624_), .C(alu__abc_38674_new_n1695_), .Y(alu__abc_38674_new_n1696_));
NOR3X1 NOR3X1_4 ( .A(_abc_40298_new_n1399_), .B(_abc_40298_new_n1414_), .C(_abc_40298_new_n1364_), .Y(_abc_40298_new_n1416_));
NOR3X1 NOR3X1_5 ( .A(_abc_40298_new_n1414_), .B(_abc_40298_new_n1447_), .C(_abc_40298_new_n1448_), .Y(_abc_40298_new_n1449_));
NOR3X1 NOR3X1_6 ( .A(_abc_40298_new_n1512_), .B(_abc_40298_new_n1532_), .C(_abc_40298_new_n1475_), .Y(_abc_40298_new_n1534_));
NOR3X1 NOR3X1_7 ( .A(_abc_40298_new_n1532_), .B(_abc_40298_new_n1561_), .C(_abc_40298_new_n1562_), .Y(_abc_40298_new_n1564_));
NOR3X1 NOR3X1_8 ( .A(_abc_40298_new_n1620_), .B(_abc_40298_new_n1644_), .C(_abc_40298_new_n1589_), .Y(_abc_40298_new_n1646_));
NOR3X1 NOR3X1_9 ( .A(_abc_40298_new_n1644_), .B(_abc_40298_new_n1675_), .C(_abc_40298_new_n1622_), .Y(_abc_40298_new_n1676_));
OAI21X1 OAI21X1_1 ( .A(state_q_0_), .B(state_q_4_), .C(enable_i), .Y(_abc_40298_new_n632_));
OAI21X1 OAI21X1_10 ( .A(_abc_40298_new_n655_), .B(_abc_40298_new_n681_), .C(_abc_40298_new_n690_), .Y(_abc_40298_new_n691_));
OAI21X1 OAI21X1_100 ( .A(_abc_40298_new_n1176_), .B(_abc_40298_new_n1174_), .C(_abc_40298_new_n1178_), .Y(_abc_40298_new_n1179_));
OAI21X1 OAI21X1_1000 ( .A(alu_a_i_13_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n730_), .Y(alu__abc_38674_new_n731_));
OAI21X1 OAI21X1_1001 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n729_), .C(alu__abc_38674_new_n732_), .Y(alu__abc_38674_new_n733_));
OAI21X1 OAI21X1_1002 ( .A(alu_a_i_11_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n735_), .Y(alu__abc_38674_new_n736_));
OAI21X1 OAI21X1_1003 ( .A(alu_b_i_1_), .B(alu__abc_38674_new_n734_), .C(alu__abc_38674_new_n737_), .Y(alu__abc_38674_new_n738_));
OAI21X1 OAI21X1_1004 ( .A(alu__abc_38674_new_n726_), .B(alu__abc_38674_new_n740_), .C(alu__abc_38674_new_n519_), .Y(alu__abc_38674_new_n741_));
OAI21X1 OAI21X1_1005 ( .A(alu_a_i_23_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n742_), .Y(alu__abc_38674_new_n743_));
OAI21X1 OAI21X1_1006 ( .A(alu_a_i_21_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n745_), .Y(alu__abc_38674_new_n746_));
OAI21X1 OAI21X1_1007 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n744_), .C(alu__abc_38674_new_n747_), .Y(alu__abc_38674_new_n748_));
OAI21X1 OAI21X1_1008 ( .A(alu_a_i_19_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n750_), .Y(alu__abc_38674_new_n751_));
OAI21X1 OAI21X1_1009 ( .A(alu_b_i_1_), .B(alu__abc_38674_new_n749_), .C(alu__abc_38674_new_n752_), .Y(alu__abc_38674_new_n753_));
OAI21X1 OAI21X1_101 ( .A(_abc_40298_new_n1070_), .B(_abc_40298_new_n1173_), .C(_abc_40298_new_n1179_), .Y(_abc_40298_new_n1180_));
OAI21X1 OAI21X1_1010 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n748_), .C(alu__abc_38674_new_n755_), .Y(alu__abc_38674_new_n756_));
OAI21X1 OAI21X1_1011 ( .A(alu_a_i_27_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n757_), .Y(alu__abc_38674_new_n758_));
OAI21X1 OAI21X1_1012 ( .A(alu_a_i_25_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n760_), .Y(alu__abc_38674_new_n761_));
OAI21X1 OAI21X1_1013 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n759_), .C(alu__abc_38674_new_n762_), .Y(alu__abc_38674_new_n763_));
OAI21X1 OAI21X1_1014 ( .A(alu__abc_38674_new_n698_), .B(alu__abc_38674_new_n765_), .C(alu__abc_38674_new_n766_), .Y(alu__abc_38674_new_n767_));
OAI21X1 OAI21X1_1015 ( .A(alu_a_i_29_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n768_), .Y(alu__abc_38674_new_n769_));
OAI21X1 OAI21X1_1016 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n767_), .C(alu__abc_38674_new_n770_), .Y(alu__abc_38674_new_n771_));
OAI21X1 OAI21X1_1017 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n764_), .C(alu__abc_38674_new_n772_), .Y(alu__abc_38674_new_n773_));
OAI21X1 OAI21X1_1018 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n756_), .C(alu__abc_38674_new_n774_), .Y(alu__abc_38674_new_n775_));
OAI21X1 OAI21X1_1019 ( .A(alu_b_i_0_), .B(alu__abc_38674_new_n336_), .C(alu__abc_38674_new_n420_), .Y(alu__abc_38674_new_n778_));
OAI21X1 OAI21X1_102 ( .A(_abc_40298_new_n992_), .B(_abc_40298_new_n1185_), .C(_abc_40298_new_n1188_), .Y(_abc_40298_new_n1189_));
OAI21X1 OAI21X1_1020 ( .A(alu__abc_38674_new_n561_), .B(alu__abc_38674_new_n263_), .C(alu__abc_38674_new_n783_), .Y(alu__abc_38674_new_n784_));
OAI21X1 OAI21X1_1021 ( .A(alu__abc_38674_new_n260_), .B(alu__abc_38674_new_n710_), .C(alu__abc_38674_new_n784_), .Y(alu__abc_38674_new_n785_));
OAI21X1 OAI21X1_1022 ( .A(alu__abc_38674_new_n261_), .B(alu__abc_38674_new_n788_), .C(alu__abc_38674_new_n787_), .Y(alu__abc_38674_new_n789_));
OAI21X1 OAI21X1_1023 ( .A(alu_a_i_1_), .B(alu_b_i_1_), .C(alu__abc_38674_new_n789_), .Y(alu__abc_38674_new_n790_));
OAI21X1 OAI21X1_1024 ( .A(alu__abc_38674_new_n283_), .B(alu__abc_38674_new_n786_), .C(alu__abc_38674_new_n790_), .Y(alu__abc_38674_new_n791_));
OAI21X1 OAI21X1_1025 ( .A(alu__abc_38674_new_n564_), .B(alu__abc_38674_new_n786_), .C(alu__abc_38674_new_n793_), .Y(alu__abc_38674_new_n794_));
OAI21X1 OAI21X1_1026 ( .A(alu__abc_38674_new_n658_), .B(alu__abc_38674_new_n777_), .C(alu__abc_38674_new_n796_), .Y(alu_p_o_1_));
OAI21X1 OAI21X1_1027 ( .A(alu__abc_38674_new_n698_), .B(alu__abc_38674_new_n765_), .C(alu_b_i_1_), .Y(alu__abc_38674_new_n798_));
OAI21X1 OAI21X1_1028 ( .A(alu_b_i_1_), .B(alu__abc_38674_new_n660_), .C(alu__abc_38674_new_n798_), .Y(alu__abc_38674_new_n799_));
OAI21X1 OAI21X1_1029 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n662_), .C(alu__abc_38674_new_n802_), .Y(alu__abc_38674_new_n803_));
OAI21X1 OAI21X1_103 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_0_), .B(_abc_40298_new_n1187_), .C(_abc_40298_new_n1189_), .Y(_abc_40298_new_n1190_));
OAI21X1 OAI21X1_1030 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n803_), .C(alu__abc_38674_new_n801_), .Y(alu__abc_38674_new_n804_));
OAI21X1 OAI21X1_1031 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n805_), .C(alu__abc_38674_new_n806_), .Y(alu__abc_38674_new_n807_));
OAI21X1 OAI21X1_1032 ( .A(alu_b_i_1_), .B(alu__abc_38674_new_n675_), .C(alu__abc_38674_new_n809_), .Y(alu__abc_38674_new_n810_));
OAI21X1 OAI21X1_1033 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n808_), .C(alu__abc_38674_new_n811_), .Y(alu__abc_38674_new_n812_));
OAI21X1 OAI21X1_1034 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n804_), .C(alu__abc_38674_new_n813_), .Y(alu__abc_38674_new_n814_));
OAI21X1 OAI21X1_1035 ( .A(alu_b_i_1_), .B(alu__abc_38674_new_n648_), .C(alu__abc_38674_new_n816_), .Y(alu__abc_38674_new_n817_));
OAI21X1 OAI21X1_1036 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n819_), .C(alu__abc_38674_new_n820_), .Y(alu__abc_38674_new_n821_));
OAI21X1 OAI21X1_1037 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n818_), .C(alu__abc_38674_new_n822_), .Y(alu__abc_38674_new_n823_));
OAI21X1 OAI21X1_1038 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n825_), .C(alu__abc_38674_new_n826_), .Y(alu__abc_38674_new_n827_));
OAI21X1 OAI21X1_1039 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n823_), .C(alu__abc_38674_new_n829_), .Y(alu__abc_38674_new_n830_));
OAI21X1 OAI21X1_104 ( .A(_abc_40298_new_n1134_), .B(_abc_40298_new_n1190_), .C(_abc_40298_new_n1180_), .Y(_abc_40298_new_n1191_));
OAI21X1 OAI21X1_1040 ( .A(alu__abc_38674_new_n519_), .B(alu__abc_38674_new_n815_), .C(alu__abc_38674_new_n830_), .Y(alu__abc_38674_new_n831_));
OAI21X1 OAI21X1_1041 ( .A(alu__abc_38674_new_n382_), .B(alu__abc_38674_new_n566_), .C(alu__abc_38674_new_n569_), .Y(alu__abc_38674_new_n832_));
OAI21X1 OAI21X1_1042 ( .A(alu__abc_38674_new_n382_), .B(alu__abc_38674_new_n570_), .C(alu__abc_38674_new_n283_), .Y(alu__abc_38674_new_n833_));
OAI21X1 OAI21X1_1043 ( .A(alu__abc_38674_new_n834_), .B(alu__abc_38674_new_n337_), .C(alu__abc_38674_new_n835_), .Y(alu__abc_38674_new_n836_));
OAI21X1 OAI21X1_1044 ( .A(alu_a_i_2_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n645_), .Y(alu__abc_38674_new_n837_));
OAI21X1 OAI21X1_1045 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n259_), .C(alu__abc_38674_new_n838_), .Y(alu__abc_38674_new_n839_));
OAI21X1 OAI21X1_1046 ( .A(alu__abc_38674_new_n658_), .B(alu__abc_38674_new_n831_), .C(alu__abc_38674_new_n849_), .Y(alu_p_o_2_));
OAI21X1 OAI21X1_1047 ( .A(alu_b_i_1_), .B(alu__abc_38674_new_n759_), .C(alu__abc_38674_new_n852_), .Y(alu__abc_38674_new_n853_));
OAI21X1 OAI21X1_1048 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n851_), .C(alu__abc_38674_new_n854_), .Y(alu__abc_38674_new_n855_));
OAI21X1 OAI21X1_1049 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n761_), .C(alu__abc_38674_new_n858_), .Y(alu__abc_38674_new_n859_));
OAI21X1 OAI21X1_105 ( .A(epc_q_0_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n1194_));
OAI21X1 OAI21X1_1050 ( .A(alu_b_i_1_), .B(alu__abc_38674_new_n860_), .C(alu__abc_38674_new_n861_), .Y(alu__abc_38674_new_n862_));
OAI21X1 OAI21X1_1051 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n859_), .C(alu__abc_38674_new_n863_), .Y(alu__abc_38674_new_n864_));
OAI21X1 OAI21X1_1052 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n864_), .C(alu__abc_38674_new_n857_), .Y(alu__abc_38674_new_n865_));
OAI21X1 OAI21X1_1053 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n749_), .C(alu__abc_38674_new_n869_), .Y(alu__abc_38674_new_n870_));
OAI21X1 OAI21X1_1054 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n872_), .C(alu__abc_38674_new_n873_), .Y(alu__abc_38674_new_n874_));
OAI21X1 OAI21X1_1055 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n871_), .C(alu__abc_38674_new_n875_), .Y(alu__abc_38674_new_n876_));
OAI21X1 OAI21X1_1056 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n868_), .C(alu__abc_38674_new_n877_), .Y(alu__abc_38674_new_n878_));
OAI21X1 OAI21X1_1057 ( .A(alu__abc_38674_new_n519_), .B(alu__abc_38674_new_n865_), .C(alu__abc_38674_new_n879_), .Y(alu__abc_38674_new_n880_));
OAI21X1 OAI21X1_1058 ( .A(alu__abc_38674_new_n558_), .B(alu__abc_38674_new_n570_), .C(alu__abc_38674_new_n881_), .Y(alu__abc_38674_new_n882_));
OAI21X1 OAI21X1_1059 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n884_), .C(alu__abc_38674_new_n886_), .Y(alu__abc_38674_new_n887_));
OAI21X1 OAI21X1_106 ( .A(_abc_40298_new_n1000_), .B(_abc_40298_new_n1177_), .C(REGFILE_SIM_reg_bank_reg_rb_o_1_), .Y(_abc_40298_new_n1197_));
OAI21X1 OAI21X1_1060 ( .A(alu__abc_38674_new_n641_), .B(alu__abc_38674_new_n713_), .C(alu__abc_38674_new_n890_), .Y(alu__abc_38674_new_n891_));
OAI21X1 OAI21X1_1061 ( .A(alu__abc_38674_new_n283_), .B(alu__abc_38674_new_n883_), .C(alu__abc_38674_new_n892_), .Y(alu__abc_38674_new_n893_));
OAI21X1 OAI21X1_1062 ( .A(alu__abc_38674_new_n268_), .B(alu__abc_38674_new_n895_), .C(alu__abc_38674_new_n339_), .Y(alu__abc_38674_new_n896_));
OAI21X1 OAI21X1_1063 ( .A(alu__abc_38674_new_n555_), .B(alu__abc_38674_new_n896_), .C(alu__abc_38674_new_n706_), .Y(alu__abc_38674_new_n897_));
OAI21X1 OAI21X1_1064 ( .A(alu__abc_38674_new_n335_), .B(alu__abc_38674_new_n343_), .C(alu__abc_38674_new_n906_), .Y(alu__abc_38674_new_n907_));
OAI21X1 OAI21X1_1065 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n633_), .C(alu__abc_38674_new_n909_), .Y(alu__abc_38674_new_n910_));
OAI21X1 OAI21X1_1066 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n912_), .C(alu__abc_38674_new_n913_), .Y(alu__abc_38674_new_n914_));
OAI21X1 OAI21X1_1067 ( .A(alu__abc_38674_new_n911_), .B(alu__abc_38674_new_n915_), .C(alu__abc_38674_new_n519_), .Y(alu__abc_38674_new_n916_));
OAI21X1 OAI21X1_1068 ( .A(alu__abc_38674_new_n698_), .B(alu__abc_38674_new_n765_), .C(alu_b_i_2_), .Y(alu__abc_38674_new_n917_));
OAI21X1 OAI21X1_1069 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n664_), .C(alu__abc_38674_new_n917_), .Y(alu__abc_38674_new_n918_));
OAI21X1 OAI21X1_107 ( .A(_abc_40298_new_n1176_), .B(_abc_40298_new_n1196_), .C(_abc_40298_new_n1197_), .Y(_abc_40298_new_n1198_));
OAI21X1 OAI21X1_1070 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n680_), .C(alu__abc_38674_new_n920_), .Y(alu__abc_38674_new_n921_));
OAI21X1 OAI21X1_1071 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n919_), .C(alu__abc_38674_new_n922_), .Y(alu__abc_38674_new_n923_));
OAI21X1 OAI21X1_1072 ( .A(alu__abc_38674_new_n519_), .B(alu__abc_38674_new_n923_), .C(alu__abc_38674_new_n916_), .Y(alu__abc_38674_new_n924_));
OAI21X1 OAI21X1_1073 ( .A(alu_b_i_1_), .B(alu__abc_38674_new_n695_), .C(alu_b_i_2_), .Y(alu__abc_38674_new_n925_));
OAI21X1 OAI21X1_1074 ( .A(alu_a_i_4_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n642_), .Y(alu__abc_38674_new_n926_));
OAI21X1 OAI21X1_1075 ( .A(alu_b_i_1_), .B(alu__abc_38674_new_n927_), .C(alu__abc_38674_new_n928_), .Y(alu__abc_38674_new_n929_));
OAI21X1 OAI21X1_1076 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n930_), .C(alu__abc_38674_new_n925_), .Y(alu__abc_38674_new_n931_));
OAI21X1 OAI21X1_1077 ( .A(alu__abc_38674_new_n436_), .B(alu__abc_38674_new_n710_), .C(alu__abc_38674_new_n934_), .Y(alu__abc_38674_new_n935_));
OAI21X1 OAI21X1_1078 ( .A(alu__abc_38674_new_n283_), .B(alu__abc_38674_new_n903_), .C(alu__abc_38674_new_n937_), .Y(alu__abc_38674_new_n938_));
OAI21X1 OAI21X1_1079 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n764_), .C(alu__abc_38674_new_n943_), .Y(alu__abc_38674_new_n944_));
OAI21X1 OAI21X1_108 ( .A(_abc_40298_new_n1070_), .B(_abc_40298_new_n1173_), .C(_abc_40298_new_n1198_), .Y(_abc_40298_new_n1199_));
OAI21X1 OAI21X1_1080 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n942_), .C(alu__abc_38674_new_n945_), .Y(alu__abc_38674_new_n946_));
OAI21X1 OAI21X1_1081 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n754_), .C(alu__abc_38674_new_n948_), .Y(alu__abc_38674_new_n949_));
OAI21X1 OAI21X1_1082 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n949_), .C(alu__abc_38674_new_n519_), .Y(alu__abc_38674_new_n950_));
OAI21X1 OAI21X1_1083 ( .A(alu_b_i_1_), .B(alu__abc_38674_new_n884_), .C(alu_b_i_2_), .Y(alu__abc_38674_new_n953_));
OAI21X1 OAI21X1_1084 ( .A(alu_a_i_5_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n954_), .Y(alu__abc_38674_new_n955_));
OAI21X1 OAI21X1_1085 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n885_), .C(alu__abc_38674_new_n956_), .Y(alu__abc_38674_new_n957_));
OAI21X1 OAI21X1_1086 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n958_), .C(alu__abc_38674_new_n953_), .Y(alu__abc_38674_new_n959_));
OAI21X1 OAI21X1_1087 ( .A(alu__abc_38674_new_n431_), .B(alu__abc_38674_new_n788_), .C(alu__abc_38674_new_n787_), .Y(alu__abc_38674_new_n961_));
OAI21X1 OAI21X1_1088 ( .A(alu__abc_38674_new_n334_), .B(alu__abc_38674_new_n713_), .C(alu__abc_38674_new_n962_), .Y(alu__abc_38674_new_n963_));
OAI21X1 OAI21X1_1089 ( .A(alu__abc_38674_new_n283_), .B(alu__abc_38674_new_n552_), .C(alu__abc_38674_new_n964_), .Y(alu__abc_38674_new_n965_));
OAI21X1 OAI21X1_109 ( .A(_abc_40298_new_n992_), .B(_abc_40298_new_n1185_), .C(_abc_40298_new_n1200_), .Y(_abc_40298_new_n1201_));
OAI21X1 OAI21X1_1090 ( .A(alu__abc_38674_new_n967_), .B(alu__abc_38674_new_n968_), .C(alu__abc_38674_new_n970_), .Y(alu__abc_38674_new_n971_));
OAI21X1 OAI21X1_1091 ( .A(alu__abc_38674_new_n335_), .B(alu__abc_38674_new_n343_), .C(alu__abc_38674_new_n972_), .Y(alu__abc_38674_new_n973_));
OAI21X1 OAI21X1_1092 ( .A(alu__abc_38674_new_n428_), .B(alu__abc_38674_new_n976_), .C(alu__abc_38674_new_n977_), .Y(alu__abc_38674_new_n978_));
OAI21X1 OAI21X1_1093 ( .A(alu__abc_38674_new_n979_), .B(alu__abc_38674_new_n969_), .C(alu__abc_38674_new_n980_), .Y(alu__abc_38674_new_n981_));
OAI21X1 OAI21X1_1094 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n827_), .C(alu__abc_38674_new_n982_), .Y(alu__abc_38674_new_n983_));
OAI21X1 OAI21X1_1095 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n808_), .C(alu__abc_38674_new_n984_), .Y(alu__abc_38674_new_n985_));
OAI21X1 OAI21X1_1096 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n983_), .C(alu__abc_38674_new_n986_), .Y(alu__abc_38674_new_n987_));
OAI21X1 OAI21X1_1097 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n800_), .C(alu__abc_38674_new_n917_), .Y(alu__abc_38674_new_n989_));
OAI21X1 OAI21X1_1098 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n988_), .C(alu__abc_38674_new_n990_), .Y(alu__abc_38674_new_n991_));
OAI21X1 OAI21X1_1099 ( .A(alu_a_i_6_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n649_), .Y(alu__abc_38674_new_n993_));
OAI21X1 OAI21X1_11 ( .A(state_q_1_), .B(_abc_40298_new_n671_), .C(_abc_40298_new_n691_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_0_));
OAI21X1 OAI21X1_110 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_1_), .B(_abc_40298_new_n1187_), .C(_abc_40298_new_n1201_), .Y(_abc_40298_new_n1202_));
OAI21X1 OAI21X1_1100 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n927_), .C(alu__abc_38674_new_n994_), .Y(alu__abc_38674_new_n995_));
OAI21X1 OAI21X1_1101 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n839_), .C(alu__abc_38674_new_n997_), .Y(alu__abc_38674_new_n998_));
OAI21X1 OAI21X1_1102 ( .A(alu__abc_38674_new_n330_), .B(alu__abc_38674_new_n713_), .C(alu__abc_38674_new_n1001_), .Y(alu__abc_38674_new_n1002_));
OAI21X1 OAI21X1_1103 ( .A(alu__abc_38674_new_n283_), .B(alu__abc_38674_new_n547_), .C(alu__abc_38674_new_n1003_), .Y(alu__abc_38674_new_n1004_));
OAI21X1 OAI21X1_1104 ( .A(alu__abc_38674_new_n426_), .B(alu__abc_38674_new_n427_), .C(alu__abc_38674_new_n348_), .Y(alu__abc_38674_new_n1007_));
OAI21X1 OAI21X1_1105 ( .A(alu_b_i_6_), .B(alu__abc_38674_new_n330_), .C(alu__abc_38674_new_n1007_), .Y(alu__abc_38674_new_n1008_));
OAI21X1 OAI21X1_1106 ( .A(alu__abc_38674_new_n517_), .B(alu__abc_38674_new_n1008_), .C(alu__abc_38674_new_n1009_), .Y(alu__abc_38674_new_n1010_));
OAI21X1 OAI21X1_1107 ( .A(alu__abc_38674_new_n544_), .B(alu__abc_38674_new_n573_), .C(alu__abc_38674_new_n1011_), .Y(alu__abc_38674_new_n1012_));
OAI21X1 OAI21X1_1108 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n871_), .C(alu__abc_38674_new_n1015_), .Y(alu__abc_38674_new_n1016_));
OAI21X1 OAI21X1_1109 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n1016_), .C(alu__abc_38674_new_n1014_), .Y(alu__abc_38674_new_n1017_));
OAI21X1 OAI21X1_111 ( .A(_abc_40298_new_n1134_), .B(_abc_40298_new_n1202_), .C(_abc_40298_new_n1199_), .Y(_abc_40298_new_n1203_));
OAI21X1 OAI21X1_1110 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n859_), .C(alu__abc_38674_new_n1018_), .Y(alu__abc_38674_new_n1019_));
OAI21X1 OAI21X1_1111 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n851_), .C(alu__abc_38674_new_n917_), .Y(alu__abc_38674_new_n1021_));
OAI21X1 OAI21X1_1112 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n1020_), .C(alu__abc_38674_new_n1022_), .Y(alu__abc_38674_new_n1023_));
OAI21X1 OAI21X1_1113 ( .A(alu_b_i_4_), .B(alu__abc_38674_new_n1017_), .C(alu__abc_38674_new_n1024_), .Y(alu__abc_38674_new_n1025_));
OAI21X1 OAI21X1_1114 ( .A(alu_a_i_7_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n1027_), .Y(alu__abc_38674_new_n1028_));
OAI21X1 OAI21X1_1115 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n1026_), .C(alu__abc_38674_new_n1029_), .Y(alu__abc_38674_new_n1030_));
OAI21X1 OAI21X1_1116 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n1030_), .C(alu__abc_38674_new_n1031_), .Y(alu__abc_38674_new_n1032_));
OAI21X1 OAI21X1_1117 ( .A(alu__abc_38674_new_n702_), .B(alu__abc_38674_new_n1033_), .C(alu__abc_38674_new_n1035_), .Y(alu__abc_38674_new_n1036_));
OAI21X1 OAI21X1_1118 ( .A(alu__abc_38674_new_n658_), .B(alu__abc_38674_new_n1025_), .C(alu__abc_38674_new_n1037_), .Y(alu__abc_38674_new_n1038_));
OAI21X1 OAI21X1_1119 ( .A(alu__abc_38674_new_n539_), .B(alu__abc_38674_new_n349_), .C(alu__abc_38674_new_n1041_), .Y(alu__abc_38674_new_n1042_));
OAI21X1 OAI21X1_112 ( .A(epc_q_1_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n1206_));
OAI21X1 OAI21X1_1120 ( .A(alu__abc_38674_new_n1046_), .B(alu__abc_38674_new_n1047_), .C(alu__abc_38674_new_n1043_), .Y(alu__abc_38674_new_n1048_));
OAI21X1 OAI21X1_1121 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n640_), .C(alu__abc_38674_new_n1051_), .Y(alu__abc_38674_new_n1052_));
OAI21X1 OAI21X1_1122 ( .A(alu__abc_38674_new_n698_), .B(alu__abc_38674_new_n765_), .C(alu_b_i_3_), .Y(alu__abc_38674_new_n1053_));
OAI21X1 OAI21X1_1123 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n674_), .C(alu__abc_38674_new_n1053_), .Y(alu__abc_38674_new_n1054_));
OAI21X1 OAI21X1_1124 ( .A(alu_b_i_4_), .B(alu__abc_38674_new_n1052_), .C(alu__abc_38674_new_n1055_), .Y(alu__abc_38674_new_n1056_));
OAI21X1 OAI21X1_1125 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n1057_), .C(alu_b_i_3_), .Y(alu__abc_38674_new_n1058_));
OAI21X1 OAI21X1_1126 ( .A(alu_a_i_8_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n1060_), .Y(alu__abc_38674_new_n1061_));
OAI21X1 OAI21X1_1127 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n1059_), .C(alu__abc_38674_new_n1062_), .Y(alu__abc_38674_new_n1063_));
OAI21X1 OAI21X1_1128 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n929_), .C(alu__abc_38674_new_n1065_), .Y(alu__abc_38674_new_n1066_));
OAI21X1 OAI21X1_1129 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n1066_), .C(alu__abc_38674_new_n1058_), .Y(alu__abc_38674_new_n1067_));
OAI21X1 OAI21X1_113 ( .A(_abc_40298_new_n658_), .B(_abc_40298_new_n995_), .C(_abc_40298_new_n1175_), .Y(_abc_40298_new_n1210_));
OAI21X1 OAI21X1_1130 ( .A(alu__abc_38674_new_n223_), .B(alu__abc_38674_new_n710_), .C(alu__abc_38674_new_n1069_), .Y(alu__abc_38674_new_n1070_));
OAI21X1 OAI21X1_1131 ( .A(alu__abc_38674_new_n537_), .B(alu__abc_38674_new_n1076_), .C(alu__abc_38674_new_n381_), .Y(alu__abc_38674_new_n1077_));
OAI21X1 OAI21X1_1132 ( .A(alu__abc_38674_new_n1081_), .B(alu__abc_38674_new_n1082_), .C(alu__abc_38674_new_n519_), .Y(alu__abc_38674_new_n1083_));
OAI21X1 OAI21X1_1133 ( .A(alu__abc_38674_new_n519_), .B(alu__abc_38674_new_n1080_), .C(alu__abc_38674_new_n1083_), .Y(alu__abc_38674_new_n1084_));
OAI21X1 OAI21X1_1134 ( .A(alu_a_i_9_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n1087_), .Y(alu__abc_38674_new_n1088_));
OAI21X1 OAI21X1_1135 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n1086_), .C(alu__abc_38674_new_n1089_), .Y(alu__abc_38674_new_n1090_));
OAI21X1 OAI21X1_1136 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n1090_), .C(alu__abc_38674_new_n1085_), .Y(alu__abc_38674_new_n1091_));
OAI21X1 OAI21X1_1137 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n1091_), .C(alu__abc_38674_new_n1092_), .Y(alu__abc_38674_new_n1093_));
OAI21X1 OAI21X1_1138 ( .A(alu_b_i_9_), .B(alu_a_i_9_), .C(alu__abc_38674_new_n703_), .Y(alu__abc_38674_new_n1096_));
OAI21X1 OAI21X1_1139 ( .A(alu__abc_38674_new_n230_), .B(alu__abc_38674_new_n788_), .C(alu__abc_38674_new_n1096_), .Y(alu__abc_38674_new_n1097_));
OAI21X1 OAI21X1_114 ( .A(pc_q_2_), .B(_abc_40298_new_n1213_), .C(_abc_40298_new_n1221_), .Y(_abc_40298_new_n1222_));
OAI21X1 OAI21X1_1140 ( .A(alu__abc_38674_new_n539_), .B(alu__abc_38674_new_n349_), .C(alu__abc_38674_new_n1098_), .Y(alu__abc_38674_new_n1099_));
OAI21X1 OAI21X1_1141 ( .A(alu__abc_38674_new_n230_), .B(alu__abc_38674_new_n1099_), .C(alu__abc_38674_new_n1103_), .Y(alu__abc_38674_new_n1104_));
OAI21X1 OAI21X1_1142 ( .A(alu__abc_38674_new_n226_), .B(alu__abc_38674_new_n710_), .C(alu__abc_38674_new_n1104_), .Y(alu__abc_38674_new_n1105_));
OAI21X1 OAI21X1_1143 ( .A(alu__abc_38674_new_n228_), .B(alu__abc_38674_new_n713_), .C(alu__abc_38674_new_n1107_), .Y(alu_p_o_9_));
OAI21X1 OAI21X1_1144 ( .A(alu__abc_38674_new_n236_), .B(alu__abc_38674_new_n1109_), .C(alu__abc_38674_new_n1110_), .Y(alu__abc_38674_new_n1111_));
OAI21X1 OAI21X1_1145 ( .A(alu__abc_38674_new_n594_), .B(alu__abc_38674_new_n1075_), .C(alu__abc_38674_new_n1114_), .Y(alu__abc_38674_new_n1115_));
OAI21X1 OAI21X1_1146 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n812_), .C(alu__abc_38674_new_n1117_), .Y(alu__abc_38674_new_n1118_));
OAI21X1 OAI21X1_1147 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n804_), .C(alu__abc_38674_new_n1053_), .Y(alu__abc_38674_new_n1119_));
OAI21X1 OAI21X1_1148 ( .A(alu_b_i_4_), .B(alu__abc_38674_new_n1118_), .C(alu__abc_38674_new_n1120_), .Y(alu__abc_38674_new_n1121_));
OAI21X1 OAI21X1_1149 ( .A(alu_a_i_10_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n631_), .Y(alu__abc_38674_new_n1123_));
OAI21X1 OAI21X1_115 ( .A(_abc_40298_new_n1070_), .B(_abc_40298_new_n1173_), .C(_abc_40298_new_n1222_), .Y(_abc_40298_new_n1223_));
OAI21X1 OAI21X1_1150 ( .A(alu_b_i_1_), .B(alu__abc_38674_new_n1124_), .C(alu__abc_38674_new_n1125_), .Y(alu__abc_38674_new_n1126_));
OAI21X1 OAI21X1_1151 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n996_), .C(alu__abc_38674_new_n1127_), .Y(alu__abc_38674_new_n1128_));
OAI21X1 OAI21X1_1152 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n1128_), .C(alu__abc_38674_new_n1122_), .Y(alu__abc_38674_new_n1129_));
OAI21X1 OAI21X1_1153 ( .A(alu__abc_38674_new_n233_), .B(alu__abc_38674_new_n713_), .C(alu__abc_38674_new_n1130_), .Y(alu__abc_38674_new_n1131_));
OAI21X1 OAI21X1_1154 ( .A(alu__abc_38674_new_n283_), .B(alu__abc_38674_new_n1116_), .C(alu__abc_38674_new_n1133_), .Y(alu__abc_38674_new_n1134_));
OAI21X1 OAI21X1_1155 ( .A(alu__abc_38674_new_n354_), .B(alu__abc_38674_new_n1101_), .C(alu__abc_38674_new_n235_), .Y(alu__abc_38674_new_n1137_));
OAI21X1 OAI21X1_1156 ( .A(alu_b_i_10_), .B(alu__abc_38674_new_n233_), .C(alu__abc_38674_new_n1137_), .Y(alu__abc_38674_new_n1138_));
OAI21X1 OAI21X1_1157 ( .A(alu__abc_38674_new_n239_), .B(alu__abc_38674_new_n1138_), .C(alu__abc_38674_new_n1139_), .Y(alu__abc_38674_new_n1140_));
OAI21X1 OAI21X1_1158 ( .A(alu__abc_38674_new_n1112_), .B(alu__abc_38674_new_n592_), .C(alu__abc_38674_new_n1141_), .Y(alu__abc_38674_new_n1142_));
OAI21X1 OAI21X1_1159 ( .A(alu__abc_38674_new_n446_), .B(alu__abc_38674_new_n590_), .C(alu__abc_38674_new_n239_), .Y(alu__abc_38674_new_n1144_));
OAI21X1 OAI21X1_116 ( .A(_abc_40298_new_n1134_), .B(_abc_40298_new_n1208_), .C(_abc_40298_new_n1223_), .Y(_abc_40298_new_n1224_));
OAI21X1 OAI21X1_1160 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n856_), .C(alu__abc_38674_new_n1053_), .Y(alu__abc_38674_new_n1147_));
OAI21X1 OAI21X1_1161 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n864_), .C(alu__abc_38674_new_n519_), .Y(alu__abc_38674_new_n1149_));
OAI21X1 OAI21X1_1162 ( .A(alu_a_i_11_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n1152_), .Y(alu__abc_38674_new_n1153_));
OAI21X1 OAI21X1_1163 ( .A(alu_b_i_1_), .B(alu__abc_38674_new_n1154_), .C(alu__abc_38674_new_n1155_), .Y(alu__abc_38674_new_n1156_));
OAI21X1 OAI21X1_1164 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n1151_), .C(alu__abc_38674_new_n1157_), .Y(alu__abc_38674_new_n1158_));
OAI21X1 OAI21X1_1165 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n1159_), .C(alu__abc_38674_new_n1160_), .Y(alu__abc_38674_new_n1161_));
OAI21X1 OAI21X1_1166 ( .A(alu_b_i_11_), .B(alu_a_i_11_), .C(alu__abc_38674_new_n703_), .Y(alu__abc_38674_new_n1163_));
OAI21X1 OAI21X1_1167 ( .A(alu__abc_38674_new_n237_), .B(alu__abc_38674_new_n710_), .C(alu__abc_38674_new_n1163_), .Y(alu__abc_38674_new_n1164_));
OAI21X1 OAI21X1_1168 ( .A(alu__abc_38674_new_n356_), .B(alu__abc_38674_new_n713_), .C(alu__abc_38674_new_n1165_), .Y(alu__abc_38674_new_n1166_));
OAI21X1 OAI21X1_1169 ( .A(alu__abc_38674_new_n658_), .B(alu__abc_38674_new_n1150_), .C(alu__abc_38674_new_n1167_), .Y(alu__abc_38674_new_n1168_));
OAI21X1 OAI21X1_117 ( .A(_abc_40298_new_n888_), .B(_abc_40298_new_n1027_), .C(pc_q_2_), .Y(_abc_40298_new_n1225_));
OAI21X1 OAI21X1_1170 ( .A(alu__abc_38674_new_n242_), .B(alu__abc_38674_new_n349_), .C(alu__abc_38674_new_n359_), .Y(alu__abc_38674_new_n1171_));
OAI21X1 OAI21X1_1171 ( .A(alu__abc_38674_new_n215_), .B(alu__abc_38674_new_n1171_), .C(alu__abc_38674_new_n1172_), .Y(alu__abc_38674_new_n1173_));
OAI21X1 OAI21X1_1172 ( .A(alu__abc_38674_new_n595_), .B(alu__abc_38674_new_n1175_), .C(alu__abc_38674_new_n1178_), .Y(alu__abc_38674_new_n1179_));
OAI21X1 OAI21X1_1173 ( .A(alu_a_i_12_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n629_), .Y(alu__abc_38674_new_n1180_));
OAI21X1 OAI21X1_1174 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n1124_), .C(alu__abc_38674_new_n1181_), .Y(alu__abc_38674_new_n1182_));
OAI21X1 OAI21X1_1175 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n1064_), .C(alu__abc_38674_new_n1183_), .Y(alu__abc_38674_new_n1184_));
OAI21X1 OAI21X1_1176 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n1185_), .C(alu__abc_38674_new_n1186_), .Y(alu__abc_38674_new_n1187_));
OAI21X1 OAI21X1_1177 ( .A(alu__abc_38674_new_n702_), .B(alu__abc_38674_new_n1187_), .C(alu__abc_38674_new_n1189_), .Y(alu__abc_38674_new_n1190_));
OAI21X1 OAI21X1_1178 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n919_), .C(alu__abc_38674_new_n1053_), .Y(alu__abc_38674_new_n1191_));
OAI21X1 OAI21X1_1179 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n921_), .C(alu__abc_38674_new_n519_), .Y(alu__abc_38674_new_n1194_));
OAI21X1 OAI21X1_118 ( .A(_abc_40298_new_n1224_), .B(_abc_40298_new_n1071_), .C(_abc_40298_new_n1225_), .Y(_abc_40298_new_n1226_));
OAI21X1 OAI21X1_1180 ( .A(alu__abc_38674_new_n1176_), .B(alu__abc_38674_new_n1174_), .C(alu__abc_38674_new_n584_), .Y(alu__abc_38674_new_n1200_));
OAI21X1 OAI21X1_1181 ( .A(alu__abc_38674_new_n212_), .B(alu__abc_38674_new_n582_), .C(alu__abc_38674_new_n579_), .Y(alu__abc_38674_new_n1202_));
OAI21X1 OAI21X1_1182 ( .A(alu__abc_38674_new_n212_), .B(alu__abc_38674_new_n213_), .C(alu__abc_38674_new_n1171_), .Y(alu__abc_38674_new_n1207_));
OAI21X1 OAI21X1_1183 ( .A(alu__abc_38674_new_n1212_), .B(alu__abc_38674_new_n1213_), .C(alu__abc_38674_new_n519_), .Y(alu__abc_38674_new_n1214_));
OAI21X1 OAI21X1_1184 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n942_), .C(alu__abc_38674_new_n1053_), .Y(alu__abc_38674_new_n1215_));
OAI21X1 OAI21X1_1185 ( .A(alu_a_i_13_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n735_), .Y(alu__abc_38674_new_n1217_));
OAI21X1 OAI21X1_1186 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n1154_), .C(alu__abc_38674_new_n1218_), .Y(alu__abc_38674_new_n1219_));
OAI21X1 OAI21X1_1187 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n1220_), .C(alu__abc_38674_new_n1221_), .Y(alu__abc_38674_new_n1222_));
OAI21X1 OAI21X1_1188 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n1223_), .C(alu__abc_38674_new_n1224_), .Y(alu__abc_38674_new_n1225_));
OAI21X1 OAI21X1_1189 ( .A(alu__abc_38674_new_n219_), .B(alu__abc_38674_new_n787_), .C(alu__abc_38674_new_n1227_), .Y(alu__abc_38674_new_n1228_));
OAI21X1 OAI21X1_119 ( .A(epc_q_2_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n1227_));
OAI21X1 OAI21X1_1190 ( .A(alu__abc_38674_new_n702_), .B(alu__abc_38674_new_n1225_), .C(alu__abc_38674_new_n1229_), .Y(alu__abc_38674_new_n1230_));
OAI21X1 OAI21X1_1191 ( .A(alu__abc_38674_new_n1208_), .B(alu__abc_38674_new_n1211_), .C(alu__abc_38674_new_n1231_), .Y(alu__abc_38674_new_n1232_));
OAI21X1 OAI21X1_1192 ( .A(alu__abc_38674_new_n363_), .B(alu__abc_38674_new_n1208_), .C(alu__abc_38674_new_n529_), .Y(alu__abc_38674_new_n1236_));
OAI21X1 OAI21X1_1193 ( .A(alu__abc_38674_new_n576_), .B(alu__abc_38674_new_n1204_), .C(alu__abc_38674_new_n1238_), .Y(alu__abc_38674_new_n1239_));
OAI21X1 OAI21X1_1194 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n988_), .C(alu__abc_38674_new_n1242_), .Y(alu__abc_38674_new_n1243_));
OAI21X1 OAI21X1_1195 ( .A(alu__abc_38674_new_n519_), .B(alu__abc_38674_new_n1241_), .C(alu__abc_38674_new_n1244_), .Y(alu__abc_38674_new_n1245_));
OAI21X1 OAI21X1_1196 ( .A(alu_a_i_14_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n635_), .Y(alu__abc_38674_new_n1248_));
OAI21X1 OAI21X1_1197 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n1247_), .C(alu__abc_38674_new_n1249_), .Y(alu__abc_38674_new_n1250_));
OAI21X1 OAI21X1_1198 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n1246_), .C(alu__abc_38674_new_n1251_), .Y(alu__abc_38674_new_n1252_));
OAI21X1 OAI21X1_1199 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n998_), .C(alu__abc_38674_new_n1253_), .Y(alu__abc_38674_new_n1254_));
OAI21X1 OAI21X1_12 ( .A(_abc_40298_new_n694_), .B(_abc_40298_new_n695_), .C(_abc_40298_new_n696_), .Y(_abc_40298_new_n697_));
OAI21X1 OAI21X1_120 ( .A(_abc_40298_new_n992_), .B(_abc_40298_new_n1185_), .C(_abc_40298_new_n1229_), .Y(_abc_40298_new_n1230_));
OAI21X1 OAI21X1_1200 ( .A(alu__abc_38674_new_n202_), .B(alu__abc_38674_new_n713_), .C(alu__abc_38674_new_n1257_), .Y(alu__abc_38674_new_n1258_));
OAI21X1 OAI21X1_1201 ( .A(alu__abc_38674_new_n658_), .B(alu__abc_38674_new_n1245_), .C(alu__abc_38674_new_n1259_), .Y(alu__abc_38674_new_n1260_));
OAI21X1 OAI21X1_1202 ( .A(alu_b_i_14_), .B(alu__abc_38674_new_n202_), .C(alu__abc_38674_new_n1236_), .Y(alu__abc_38674_new_n1263_));
OAI21X1 OAI21X1_1203 ( .A(alu__abc_38674_new_n208_), .B(alu__abc_38674_new_n1263_), .C(alu__abc_38674_new_n1264_), .Y(alu__abc_38674_new_n1265_));
OAI21X1 OAI21X1_1204 ( .A(alu__abc_38674_new_n576_), .B(alu__abc_38674_new_n1204_), .C(alu__abc_38674_new_n1266_), .Y(alu__abc_38674_new_n1267_));
OAI21X1 OAI21X1_1205 ( .A(alu__abc_38674_new_n1273_), .B(alu__abc_38674_new_n1274_), .C(alu__abc_38674_new_n519_), .Y(alu__abc_38674_new_n1275_));
OAI21X1 OAI21X1_1206 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n1276_), .C(alu__abc_38674_new_n1053_), .Y(alu__abc_38674_new_n1277_));
OAI21X1 OAI21X1_1207 ( .A(alu__abc_38674_new_n519_), .B(alu__abc_38674_new_n1277_), .C(alu__abc_38674_new_n1275_), .Y(alu__abc_38674_new_n1278_));
OAI21X1 OAI21X1_1208 ( .A(alu_b_i_1_), .B(alu__abc_38674_new_n1280_), .C(alu__abc_38674_new_n1281_), .Y(alu__abc_38674_new_n1282_));
OAI21X1 OAI21X1_1209 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n1283_), .C(alu__abc_38674_new_n1284_), .Y(alu__abc_38674_new_n1285_));
OAI21X1 OAI21X1_121 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_3_), .B(_abc_40298_new_n1187_), .C(_abc_40298_new_n1230_), .Y(_abc_40298_new_n1231_));
OAI21X1 OAI21X1_1210 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n1285_), .C(alu__abc_38674_new_n1279_), .Y(alu__abc_38674_new_n1286_));
OAI21X1 OAI21X1_1211 ( .A(alu__abc_38674_new_n511_), .B(alu__abc_38674_new_n598_), .C(alu__abc_38674_new_n381_), .Y(alu__abc_38674_new_n1298_));
OAI21X1 OAI21X1_1212 ( .A(alu__abc_38674_new_n283_), .B(alu__abc_38674_new_n511_), .C(alu__abc_38674_new_n1298_), .Y(alu__abc_38674_new_n1299_));
OAI21X1 OAI21X1_1213 ( .A(alu__abc_38674_new_n510_), .B(alu__abc_38674_new_n1297_), .C(alu__abc_38674_new_n1299_), .Y(alu__abc_38674_new_n1300_));
OAI21X1 OAI21X1_1214 ( .A(alu__abc_38674_new_n465_), .B(alu__abc_38674_new_n1301_), .C(alu__abc_38674_new_n1302_), .Y(alu__abc_38674_new_n1303_));
OAI21X1 OAI21X1_1215 ( .A(alu__abc_38674_new_n519_), .B(alu__abc_38674_new_n1304_), .C(alu__abc_38674_new_n908_), .Y(alu__abc_38674_new_n1305_));
OAI21X1 OAI21X1_1216 ( .A(alu_a_i_16_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n1308_), .Y(alu__abc_38674_new_n1309_));
OAI21X1 OAI21X1_1217 ( .A(alu_b_i_1_), .B(alu__abc_38674_new_n1310_), .C(alu__abc_38674_new_n1311_), .Y(alu__abc_38674_new_n1312_));
OAI21X1 OAI21X1_1218 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n1182_), .C(alu__abc_38674_new_n1314_), .Y(alu__abc_38674_new_n1315_));
OAI21X1 OAI21X1_1219 ( .A(alu__abc_38674_new_n137_), .B(alu__abc_38674_new_n787_), .C(alu__abc_38674_new_n1319_), .Y(alu__abc_38674_new_n1320_));
OAI21X1 OAI21X1_122 ( .A(_abc_40298_new_n1229_), .B(_abc_40298_new_n1066_), .C(_abc_40298_new_n1237_), .Y(_abc_40298_new_n1238_));
OAI21X1 OAI21X1_1220 ( .A(alu__abc_38674_new_n697_), .B(alu__abc_38674_new_n1318_), .C(alu__abc_38674_new_n1321_), .Y(alu__abc_38674_new_n1322_));
OAI21X1 OAI21X1_1221 ( .A(alu__abc_38674_new_n702_), .B(alu__abc_38674_new_n1316_), .C(alu__abc_38674_new_n1323_), .Y(alu__abc_38674_new_n1324_));
OAI21X1 OAI21X1_1222 ( .A(alu__abc_38674_new_n511_), .B(alu__abc_38674_new_n598_), .C(alu__abc_38674_new_n1327_), .Y(alu__abc_38674_new_n1328_));
OAI21X1 OAI21X1_1223 ( .A(alu__abc_38674_new_n1329_), .B(alu__abc_38674_new_n1332_), .C(alu__abc_38674_new_n1328_), .Y(alu__abc_38674_new_n1333_));
OAI21X1 OAI21X1_1224 ( .A(alu_b_i_16_), .B(alu__abc_38674_new_n135_), .C(alu__abc_38674_new_n140_), .Y(alu__abc_38674_new_n1335_));
OAI21X1 OAI21X1_1225 ( .A(alu__abc_38674_new_n138_), .B(alu__abc_38674_new_n139_), .C(alu__abc_38674_new_n1334_), .Y(alu__abc_38674_new_n1336_));
OAI21X1 OAI21X1_1226 ( .A(alu__abc_38674_new_n1334_), .B(alu__abc_38674_new_n1335_), .C(alu__abc_38674_new_n1339_), .Y(alu__abc_38674_new_n1340_));
OAI21X1 OAI21X1_1227 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n1344_), .C(alu__abc_38674_new_n1342_), .Y(alu__abc_38674_new_n1345_));
OAI21X1 OAI21X1_1228 ( .A(alu__abc_38674_new_n1347_), .B(alu__abc_38674_new_n1346_), .C(alu__abc_38674_new_n519_), .Y(alu__abc_38674_new_n1348_));
OAI21X1 OAI21X1_1229 ( .A(alu__abc_38674_new_n519_), .B(alu__abc_38674_new_n780_), .C(alu__abc_38674_new_n1348_), .Y(alu__abc_38674_new_n1349_));
OAI21X1 OAI21X1_123 ( .A(_abc_40298_new_n1233_), .B(_abc_40298_new_n1175_), .C(_abc_40298_new_n1239_), .Y(_abc_40298_new_n1240_));
OAI21X1 OAI21X1_1230 ( .A(alu__abc_38674_new_n1350_), .B(alu__abc_38674_new_n710_), .C(alu__abc_38674_new_n1352_), .Y(alu__abc_38674_new_n1353_));
OAI21X1 OAI21X1_1231 ( .A(alu__abc_38674_new_n700_), .B(alu__abc_38674_new_n1349_), .C(alu__abc_38674_new_n1354_), .Y(alu__abc_38674_new_n1355_));
OAI21X1 OAI21X1_1232 ( .A(alu__abc_38674_new_n283_), .B(alu__abc_38674_new_n1358_), .C(alu__abc_38674_new_n1360_), .Y(alu__abc_38674_new_n1361_));
OAI21X1 OAI21X1_1233 ( .A(alu__abc_38674_new_n600_), .B(alu__abc_38674_new_n1331_), .C(alu__abc_38674_new_n1361_), .Y(alu__abc_38674_new_n1362_));
OAI21X1 OAI21X1_1234 ( .A(alu__abc_38674_new_n306_), .B(alu__abc_38674_new_n1363_), .C(alu__abc_38674_new_n1364_), .Y(alu__abc_38674_new_n1365_));
OAI21X1 OAI21X1_1235 ( .A(alu_a_i_18_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n1368_), .Y(alu__abc_38674_new_n1369_));
OAI21X1 OAI21X1_1236 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n1310_), .C(alu__abc_38674_new_n1370_), .Y(alu__abc_38674_new_n1371_));
OAI21X1 OAI21X1_1237 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n1372_), .C(alu__abc_38674_new_n1373_), .Y(alu__abc_38674_new_n1374_));
OAI21X1 OAI21X1_1238 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n1374_), .C(alu__abc_38674_new_n1376_), .Y(alu__abc_38674_new_n1377_));
OAI21X1 OAI21X1_1239 ( .A(alu__abc_38674_new_n519_), .B(alu__abc_38674_new_n841_), .C(alu__abc_38674_new_n1377_), .Y(alu__abc_38674_new_n1378_));
OAI21X1 OAI21X1_124 ( .A(_abc_40298_new_n1241_), .B(_abc_40298_new_n1242_), .C(_abc_40298_new_n1232_), .Y(_abc_40298_new_n1243_));
OAI21X1 OAI21X1_1240 ( .A(alu__abc_38674_new_n700_), .B(alu__abc_38674_new_n1378_), .C(alu__abc_38674_new_n1380_), .Y(alu__abc_38674_new_n1381_));
OAI21X1 OAI21X1_1241 ( .A(alu_a_i_19_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n1389_), .Y(alu__abc_38674_new_n1390_));
OAI21X1 OAI21X1_1242 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n1343_), .C(alu__abc_38674_new_n1391_), .Y(alu__abc_38674_new_n1392_));
OAI21X1 OAI21X1_1243 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n1283_), .C(alu__abc_38674_new_n1393_), .Y(alu__abc_38674_new_n1394_));
OAI21X1 OAI21X1_1244 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n1159_), .C(alu__abc_38674_new_n1395_), .Y(alu__abc_38674_new_n1396_));
OAI21X1 OAI21X1_1245 ( .A(alu_b_i_4_), .B(alu__abc_38674_new_n1396_), .C(alu__abc_38674_new_n1397_), .Y(alu__abc_38674_new_n1398_));
OAI21X1 OAI21X1_1246 ( .A(alu__abc_38674_new_n310_), .B(alu__abc_38674_new_n1337_), .C(alu__abc_38674_new_n307_), .Y(alu__abc_38674_new_n1402_));
OAI21X1 OAI21X1_1247 ( .A(alu_b_i_18_), .B(alu__abc_38674_new_n144_), .C(alu__abc_38674_new_n1402_), .Y(alu__abc_38674_new_n1403_));
OAI21X1 OAI21X1_1248 ( .A(alu__abc_38674_new_n150_), .B(alu__abc_38674_new_n1403_), .C(alu__abc_38674_new_n1404_), .Y(alu__abc_38674_new_n1405_));
OAI21X1 OAI21X1_1249 ( .A(alu__abc_38674_new_n312_), .B(alu__abc_38674_new_n713_), .C(alu__abc_38674_new_n1409_), .Y(alu_p_o_19_));
OAI21X1 OAI21X1_125 ( .A(_abc_40298_new_n1232_), .B(_abc_40298_new_n1240_), .C(_abc_40298_new_n1243_), .Y(_abc_40298_new_n1244_));
OAI21X1 OAI21X1_1250 ( .A(alu__abc_38674_new_n205_), .B(alu__abc_38674_new_n206_), .C(alu__abc_38674_new_n533_), .Y(alu__abc_38674_new_n1414_));
OAI21X1 OAI21X1_1251 ( .A(alu__abc_38674_new_n599_), .B(alu__abc_38674_new_n1411_), .C(alu__abc_38674_new_n1418_), .Y(alu__abc_38674_new_n1419_));
OAI21X1 OAI21X1_1252 ( .A(alu__abc_38674_new_n125_), .B(alu__abc_38674_new_n1422_), .C(alu__abc_38674_new_n1423_), .Y(alu__abc_38674_new_n1424_));
OAI21X1 OAI21X1_1253 ( .A(alu_a_i_20_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n682_), .Y(alu__abc_38674_new_n1425_));
OAI21X1 OAI21X1_1254 ( .A(alu_b_i_1_), .B(alu__abc_38674_new_n1426_), .C(alu__abc_38674_new_n1427_), .Y(alu__abc_38674_new_n1428_));
OAI21X1 OAI21X1_1255 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n1313_), .C(alu__abc_38674_new_n1429_), .Y(alu__abc_38674_new_n1430_));
OAI21X1 OAI21X1_1256 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n1430_), .C(alu__abc_38674_new_n1431_), .Y(alu__abc_38674_new_n1432_));
OAI21X1 OAI21X1_1257 ( .A(alu__abc_38674_new_n519_), .B(alu__abc_38674_new_n932_), .C(alu__abc_38674_new_n1432_), .Y(alu__abc_38674_new_n1433_));
OAI21X1 OAI21X1_1258 ( .A(alu__abc_38674_new_n700_), .B(alu__abc_38674_new_n1433_), .C(alu__abc_38674_new_n1435_), .Y(alu__abc_38674_new_n1436_));
OAI21X1 OAI21X1_1259 ( .A(alu_b_i_4_), .B(alu__abc_38674_new_n1437_), .C(alu__abc_38674_new_n1306_), .Y(alu__abc_38674_new_n1438_));
OAI21X1 OAI21X1_126 ( .A(_abc_40298_new_n888_), .B(_abc_40298_new_n1027_), .C(_abc_40298_new_n1247_), .Y(_abc_40298_new_n1248_));
OAI21X1 OAI21X1_1260 ( .A(alu__abc_38674_new_n407_), .B(alu__abc_38674_new_n710_), .C(alu__abc_38674_new_n1438_), .Y(alu__abc_38674_new_n1439_));
OAI21X1 OAI21X1_1261 ( .A(alu__abc_38674_new_n1384_), .B(alu__abc_38674_new_n1443_), .C(alu__abc_38674_new_n493_), .Y(alu__abc_38674_new_n1444_));
OAI21X1 OAI21X1_1262 ( .A(alu__abc_38674_new_n1420_), .B(alu__abc_38674_new_n1421_), .C(alu__abc_38674_new_n126_), .Y(alu__abc_38674_new_n1448_));
OAI21X1 OAI21X1_1263 ( .A(alu_b_i_20_), .B(alu__abc_38674_new_n122_), .C(alu__abc_38674_new_n1448_), .Y(alu__abc_38674_new_n1449_));
OAI21X1 OAI21X1_1264 ( .A(alu_a_i_21_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n750_), .Y(alu__abc_38674_new_n1453_));
OAI21X1 OAI21X1_1265 ( .A(alu_b_i_1_), .B(alu__abc_38674_new_n1454_), .C(alu__abc_38674_new_n1455_), .Y(alu__abc_38674_new_n1456_));
OAI21X1 OAI21X1_1266 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n1222_), .C(alu__abc_38674_new_n519_), .Y(alu__abc_38674_new_n1458_));
OAI21X1 OAI21X1_1267 ( .A(alu__abc_38674_new_n519_), .B(alu__abc_38674_new_n960_), .C(alu__abc_38674_new_n699_), .Y(alu__abc_38674_new_n1460_));
OAI21X1 OAI21X1_1268 ( .A(alu__abc_38674_new_n1460_), .B(alu__abc_38674_new_n1459_), .C(alu__abc_38674_new_n1463_), .Y(alu__abc_38674_new_n1464_));
OAI21X1 OAI21X1_1269 ( .A(alu__abc_38674_new_n408_), .B(alu__abc_38674_new_n710_), .C(alu__abc_38674_new_n1465_), .Y(alu__abc_38674_new_n1466_));
OAI21X1 OAI21X1_127 ( .A(_abc_40298_new_n1245_), .B(_abc_40298_new_n1071_), .C(_abc_40298_new_n1248_), .Y(_abc_40298_new_n1249_));
OAI21X1 OAI21X1_1270 ( .A(alu__abc_38674_new_n382_), .B(alu__abc_38674_new_n1447_), .C(alu__abc_38674_new_n1468_), .Y(alu_p_o_21_));
OAI21X1 OAI21X1_1271 ( .A(alu_a_i_22_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n676_), .Y(alu__abc_38674_new_n1475_));
OAI21X1 OAI21X1_1272 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n1426_), .C(alu__abc_38674_new_n1476_), .Y(alu__abc_38674_new_n1477_));
OAI21X1 OAI21X1_1273 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n1372_), .C(alu__abc_38674_new_n1478_), .Y(alu__abc_38674_new_n1479_));
OAI21X1 OAI21X1_1274 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n1474_), .C(alu__abc_38674_new_n1480_), .Y(alu__abc_38674_new_n1481_));
OAI21X1 OAI21X1_1275 ( .A(alu_b_i_4_), .B(alu__abc_38674_new_n1481_), .C(alu__abc_38674_new_n1482_), .Y(alu__abc_38674_new_n1483_));
OAI21X1 OAI21X1_1276 ( .A(alu__abc_38674_new_n1473_), .B(alu__abc_38674_new_n1470_), .C(alu__abc_38674_new_n1485_), .Y(alu__abc_38674_new_n1486_));
OAI21X1 OAI21X1_1277 ( .A(alu__abc_38674_new_n131_), .B(alu__abc_38674_new_n1422_), .C(alu__abc_38674_new_n320_), .Y(alu__abc_38674_new_n1487_));
OAI21X1 OAI21X1_1278 ( .A(alu__abc_38674_new_n115_), .B(alu__abc_38674_new_n1487_), .C(alu__abc_38674_new_n1489_), .Y(alu__abc_38674_new_n1490_));
OAI21X1 OAI21X1_1279 ( .A(alu__abc_38674_new_n111_), .B(alu__abc_38674_new_n713_), .C(alu__abc_38674_new_n1495_), .Y(alu_p_o_22_));
OAI21X1 OAI21X1_128 ( .A(epc_q_3_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n1250_));
OAI21X1 OAI21X1_1280 ( .A(alu__abc_38674_new_n1498_), .B(alu__abc_38674_new_n1445_), .C(alu__abc_38674_new_n624_), .Y(alu__abc_38674_new_n1499_));
OAI21X1 OAI21X1_1281 ( .A(alu__abc_38674_new_n382_), .B(alu__abc_38674_new_n1501_), .C(alu__abc_38674_new_n1497_), .Y(alu__abc_38674_new_n1502_));
OAI21X1 OAI21X1_1282 ( .A(alu__abc_38674_new_n321_), .B(alu__abc_38674_new_n1503_), .C(alu__abc_38674_new_n706_), .Y(alu__abc_38674_new_n1505_));
OAI21X1 OAI21X1_1283 ( .A(alu_a_i_23_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n745_), .Y(alu__abc_38674_new_n1507_));
OAI21X1 OAI21X1_1284 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n1454_), .C(alu__abc_38674_new_n1508_), .Y(alu__abc_38674_new_n1509_));
OAI21X1 OAI21X1_1285 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n1506_), .C(alu__abc_38674_new_n1510_), .Y(alu__abc_38674_new_n1511_));
OAI21X1 OAI21X1_1286 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n1511_), .C(alu__abc_38674_new_n1513_), .Y(alu__abc_38674_new_n1514_));
OAI21X1 OAI21X1_1287 ( .A(alu__abc_38674_new_n117_), .B(alu__abc_38674_new_n713_), .C(alu__abc_38674_new_n1518_), .Y(alu__abc_38674_new_n1519_));
OAI21X1 OAI21X1_1288 ( .A(alu__abc_38674_new_n1504_), .B(alu__abc_38674_new_n1505_), .C(alu__abc_38674_new_n1521_), .Y(alu__abc_38674_new_n1522_));
OAI21X1 OAI21X1_1289 ( .A(alu__abc_38674_new_n508_), .B(alu__abc_38674_new_n1524_), .C(alu__abc_38674_new_n1526_), .Y(alu__abc_38674_new_n1527_));
OAI21X1 OAI21X1_129 ( .A(_abc_40298_new_n992_), .B(_abc_40298_new_n1185_), .C(_abc_40298_new_n1252_), .Y(_abc_40298_new_n1253_));
OAI21X1 OAI21X1_1290 ( .A(alu__abc_38674_new_n471_), .B(alu__abc_38674_new_n1529_), .C(alu__abc_38674_new_n1530_), .Y(alu__abc_38674_new_n1531_));
OAI21X1 OAI21X1_1291 ( .A(alu_a_i_24_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n1533_), .Y(alu__abc_38674_new_n1534_));
OAI21X1 OAI21X1_1292 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n1535_), .C(alu__abc_38674_new_n1536_), .Y(alu__abc_38674_new_n1537_));
OAI21X1 OAI21X1_1293 ( .A(alu_b_i_3_), .B(alu__abc_38674_new_n1537_), .C(alu__abc_38674_new_n1538_), .Y(alu__abc_38674_new_n1539_));
OAI21X1 OAI21X1_1294 ( .A(alu__abc_38674_new_n178_), .B(alu__abc_38674_new_n713_), .C(alu__abc_38674_new_n1541_), .Y(alu__abc_38674_new_n1542_));
OAI21X1 OAI21X1_1295 ( .A(alu__abc_38674_new_n1067_), .B(alu__abc_38674_new_n1318_), .C(alu__abc_38674_new_n1543_), .Y(alu__abc_38674_new_n1544_));
OAI21X1 OAI21X1_1296 ( .A(alu__abc_38674_new_n503_), .B(alu__abc_38674_new_n1525_), .C(alu__abc_38674_new_n1548_), .Y(alu__abc_38674_new_n1549_));
OAI21X1 OAI21X1_1297 ( .A(alu_a_i_25_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n742_), .Y(alu__abc_38674_new_n1552_));
OAI21X1 OAI21X1_1298 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n1551_), .C(alu__abc_38674_new_n1553_), .Y(alu__abc_38674_new_n1554_));
OAI21X1 OAI21X1_1299 ( .A(alu__abc_38674_new_n471_), .B(alu__abc_38674_new_n1529_), .C(alu__abc_38674_new_n1560_), .Y(alu__abc_38674_new_n1561_));
OAI21X1 OAI21X1_13 ( .A(_abc_40298_new_n694_), .B(_abc_40298_new_n699_), .C(_abc_40298_new_n700_), .Y(_abc_40298_new_n701_));
OAI21X1 OAI21X1_130 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_4_), .B(_abc_40298_new_n1187_), .C(_abc_40298_new_n1253_), .Y(_abc_40298_new_n1254_));
OAI21X1 OAI21X1_1300 ( .A(alu__abc_38674_new_n182_), .B(alu__abc_38674_new_n787_), .C(alu__abc_38674_new_n1564_), .Y(alu__abc_38674_new_n1565_));
OAI21X1 OAI21X1_1301 ( .A(alu__abc_38674_new_n1318_), .B(alu__abc_38674_new_n1093_), .C(alu__abc_38674_new_n1566_), .Y(alu__abc_38674_new_n1567_));
OAI21X1 OAI21X1_1302 ( .A(alu__abc_38674_new_n1559_), .B(alu__abc_38674_new_n1562_), .C(alu__abc_38674_new_n1568_), .Y(alu__abc_38674_new_n1569_));
OAI21X1 OAI21X1_1303 ( .A(alu__abc_38674_new_n185_), .B(alu__abc_38674_new_n1529_), .C(alu__abc_38674_new_n299_), .Y(alu__abc_38674_new_n1579_));
OAI21X1 OAI21X1_1304 ( .A(alu__abc_38674_new_n191_), .B(alu__abc_38674_new_n1579_), .C(alu__abc_38674_new_n1581_), .Y(alu__abc_38674_new_n1582_));
OAI21X1 OAI21X1_1305 ( .A(alu_a_i_26_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n668_), .Y(alu__abc_38674_new_n1585_));
OAI21X1 OAI21X1_1306 ( .A(alu_b_i_1_), .B(alu__abc_38674_new_n1586_), .C(alu__abc_38674_new_n1587_), .Y(alu__abc_38674_new_n1588_));
OAI21X1 OAI21X1_1307 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n1584_), .C(alu__abc_38674_new_n1589_), .Y(alu__abc_38674_new_n1590_));
OAI21X1 OAI21X1_1308 ( .A(alu__abc_38674_new_n1591_), .B(alu__abc_38674_new_n1592_), .C(alu__abc_38674_new_n701_), .Y(alu__abc_38674_new_n1593_));
OAI21X1 OAI21X1_1309 ( .A(alu__abc_38674_new_n189_), .B(alu__abc_38674_new_n787_), .C(alu__abc_38674_new_n1595_), .Y(alu__abc_38674_new_n1596_));
OAI21X1 OAI21X1_131 ( .A(_abc_40298_new_n1215_), .B(_abc_40298_new_n1255_), .C(_abc_40298_new_n1256_), .Y(_abc_40298_new_n1257_));
OAI21X1 OAI21X1_1310 ( .A(alu__abc_38674_new_n620_), .B(alu__abc_38674_new_n1602_), .C(alu__abc_38674_new_n381_), .Y(alu__abc_38674_new_n1603_));
OAI21X1 OAI21X1_1311 ( .A(alu__abc_38674_new_n395_), .B(alu__abc_38674_new_n1604_), .C(alu__abc_38674_new_n706_), .Y(alu__abc_38674_new_n1606_));
OAI21X1 OAI21X1_1312 ( .A(alu_a_i_27_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n760_), .Y(alu__abc_38674_new_n1607_));
OAI21X1 OAI21X1_1313 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n1552_), .C(alu__abc_38674_new_n1609_), .Y(alu__abc_38674_new_n1610_));
OAI21X1 OAI21X1_1314 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n1610_), .C(alu__abc_38674_new_n1611_), .Y(alu__abc_38674_new_n1612_));
OAI21X1 OAI21X1_1315 ( .A(alu_b_i_4_), .B(alu__abc_38674_new_n1148_), .C(alu__abc_38674_new_n1306_), .Y(alu__abc_38674_new_n1614_));
OAI21X1 OAI21X1_1316 ( .A(alu__abc_38674_new_n195_), .B(alu__abc_38674_new_n787_), .C(alu__abc_38674_new_n1616_), .Y(alu__abc_38674_new_n1617_));
OAI21X1 OAI21X1_1317 ( .A(alu__abc_38674_new_n1605_), .B(alu__abc_38674_new_n1606_), .C(alu__abc_38674_new_n1620_), .Y(alu__abc_38674_new_n1621_));
OAI21X1 OAI21X1_1318 ( .A(alu__abc_38674_new_n1601_), .B(alu__abc_38674_new_n1603_), .C(alu__abc_38674_new_n1622_), .Y(alu_p_o_27_));
OAI21X1 OAI21X1_1319 ( .A(alu__abc_38674_new_n620_), .B(alu__abc_38674_new_n1602_), .C(alu__abc_38674_new_n1624_), .Y(alu__abc_38674_new_n1626_));
OAI21X1 OAI21X1_132 ( .A(_abc_40298_new_n909_), .B(_abc_40298_new_n1255_), .C(_abc_40298_new_n1236_), .Y(_abc_40298_new_n1261_));
OAI21X1 OAI21X1_1320 ( .A(alu__abc_38674_new_n305_), .B(alu__abc_38674_new_n371_), .C(alu__abc_38674_new_n390_), .Y(alu__abc_38674_new_n1629_));
OAI21X1 OAI21X1_1321 ( .A(alu_b_i_4_), .B(alu__abc_38674_new_n1192_), .C(alu__abc_38674_new_n1306_), .Y(alu__abc_38674_new_n1632_));
OAI21X1 OAI21X1_1322 ( .A(alu_a_i_28_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n665_), .Y(alu__abc_38674_new_n1634_));
OAI21X1 OAI21X1_1323 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n1585_), .C(alu__abc_38674_new_n338_), .Y(alu__abc_38674_new_n1636_));
OAI21X1 OAI21X1_1324 ( .A(alu__abc_38674_new_n390_), .B(alu__abc_38674_new_n788_), .C(alu__abc_38674_new_n1640_), .Y(alu__abc_38674_new_n1641_));
OAI21X1 OAI21X1_1325 ( .A(alu__abc_38674_new_n1318_), .B(alu__abc_38674_new_n1187_), .C(alu__abc_38674_new_n1642_), .Y(alu__abc_38674_new_n1643_));
OAI21X1 OAI21X1_1326 ( .A(alu__abc_38674_new_n1625_), .B(alu__abc_38674_new_n1627_), .C(alu__abc_38674_new_n1647_), .Y(alu_p_o_28_));
OAI21X1 OAI21X1_1327 ( .A(alu_b_i_28_), .B(alu__abc_38674_new_n171_), .C(alu__abc_38674_new_n1629_), .Y(alu__abc_38674_new_n1652_));
OAI21X1 OAI21X1_1328 ( .A(alu__abc_38674_new_n169_), .B(alu__abc_38674_new_n1652_), .C(alu__abc_38674_new_n1653_), .Y(alu__abc_38674_new_n1654_));
OAI21X1 OAI21X1_1329 ( .A(alu_a_i_29_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n757_), .Y(alu__abc_38674_new_n1656_));
OAI21X1 OAI21X1_133 ( .A(_abc_40298_new_n1261_), .B(_abc_40298_new_n1264_), .C(_abc_40298_new_n1266_), .Y(_abc_40298_new_n1267_));
OAI21X1 OAI21X1_1330 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n1608_), .C(alu__abc_38674_new_n1657_), .Y(alu__abc_38674_new_n1658_));
OAI21X1 OAI21X1_1331 ( .A(alu__abc_38674_new_n519_), .B(alu__abc_38674_new_n1655_), .C(alu__abc_38674_new_n1661_), .Y(alu__abc_38674_new_n1662_));
OAI21X1 OAI21X1_1332 ( .A(alu__abc_38674_new_n165_), .B(alu__abc_38674_new_n713_), .C(alu__abc_38674_new_n1665_), .Y(alu__abc_38674_new_n1666_));
OAI21X1 OAI21X1_1333 ( .A(alu__abc_38674_new_n382_), .B(alu__abc_38674_new_n1651_), .C(alu__abc_38674_new_n1669_), .Y(alu_p_o_29_));
OAI21X1 OAI21X1_1334 ( .A(alu__abc_38674_new_n1649_), .B(alu__abc_38674_new_n1650_), .C(alu__abc_38674_new_n1671_), .Y(alu__abc_38674_new_n1672_));
OAI21X1 OAI21X1_1335 ( .A(alu__abc_38674_new_n383_), .B(alu__abc_38674_new_n376_), .C(alu__abc_38674_new_n1676_), .Y(alu__abc_38674_new_n1677_));
OAI21X1 OAI21X1_1336 ( .A(alu_b_i_4_), .B(alu__abc_38674_new_n1241_), .C(alu__abc_38674_new_n1306_), .Y(alu__abc_38674_new_n1679_));
OAI21X1 OAI21X1_1337 ( .A(alu_b_i_1_), .B(alu__abc_38674_new_n1680_), .C(alu__abc_38674_new_n1681_), .Y(alu__abc_38674_new_n1682_));
OAI21X1 OAI21X1_1338 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n1479_), .C(alu__abc_38674_new_n519_), .Y(alu__abc_38674_new_n1684_));
OAI21X1 OAI21X1_1339 ( .A(alu__abc_38674_new_n158_), .B(alu__abc_38674_new_n787_), .C(alu__abc_38674_new_n1688_), .Y(alu__abc_38674_new_n1689_));
OAI21X1 OAI21X1_134 ( .A(_abc_40298_new_n1213_), .B(_abc_40298_new_n1259_), .C(_abc_40298_new_n1270_), .Y(_abc_40298_new_n1271_));
OAI21X1 OAI21X1_1340 ( .A(alu__abc_38674_new_n626_), .B(alu__abc_38674_new_n609_), .C(alu__abc_38674_new_n381_), .Y(alu__abc_38674_new_n1698_));
OAI21X1 OAI21X1_1341 ( .A(alu__abc_38674_new_n1699_), .B(alu__abc_38674_new_n1675_), .C(alu__abc_38674_new_n384_), .Y(alu__abc_38674_new_n1702_));
OAI21X1 OAI21X1_1342 ( .A(alu_a_i_31_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n768_), .Y(alu__abc_38674_new_n1706_));
OAI21X1 OAI21X1_1343 ( .A(alu__abc_38674_new_n1708_), .B(alu__abc_38674_new_n1709_), .C(alu__abc_38674_new_n340_), .Y(alu__abc_38674_new_n1710_));
OAI21X1 OAI21X1_1344 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n1705_), .C(alu__abc_38674_new_n1710_), .Y(alu__abc_38674_new_n1711_));
OAI21X1 OAI21X1_1345 ( .A(alu__abc_38674_new_n161_), .B(alu__abc_38674_new_n787_), .C(alu__abc_38674_new_n1712_), .Y(alu__abc_38674_new_n1713_));
OAI21X1 OAI21X1_1346 ( .A(alu__abc_38674_new_n294_), .B(alu__abc_38674_new_n713_), .C(alu__abc_38674_new_n1714_), .Y(alu__abc_38674_new_n1715_));
OAI21X1 OAI21X1_1347 ( .A(alu__abc_38674_new_n702_), .B(alu__abc_38674_new_n1711_), .C(alu__abc_38674_new_n1716_), .Y(alu__abc_38674_new_n1717_));
OAI21X1 OAI21X1_1348 ( .A(alu__abc_38674_new_n782_), .B(alu__abc_38674_new_n1703_), .C(alu__abc_38674_new_n1718_), .Y(alu__abc_38674_new_n1719_));
OAI21X1 OAI21X1_1349 ( .A(alu__abc_38674_new_n1698_), .B(alu__abc_38674_new_n1697_), .C(alu__abc_38674_new_n1720_), .Y(alu_p_o_31_));
OAI21X1 OAI21X1_135 ( .A(_abc_40298_new_n1070_), .B(_abc_40298_new_n1173_), .C(_abc_40298_new_n1271_), .Y(_abc_40298_new_n1272_));
OAI21X1 OAI21X1_1350 ( .A(alu__abc_38674_new_n326_), .B(alu__abc_38674_new_n316_), .C(alu__abc_38674_new_n199_), .Y(alu__abc_38674_new_n1724_));
OAI21X1 OAI21X1_1351 ( .A(alu__abc_38674_new_n161_), .B(alu__abc_38674_new_n160_), .C(alu__abc_38674_new_n1699_), .Y(alu__abc_38674_new_n1727_));
OAI21X1 OAI21X1_1352 ( .A(alu_b_i_31_), .B(alu__abc_38674_new_n294_), .C(alu__abc_38674_new_n1727_), .Y(alu__abc_38674_new_n1728_));
OAI21X1 OAI21X1_136 ( .A(_abc_40298_new_n1134_), .B(_abc_40298_new_n1254_), .C(_abc_40298_new_n1272_), .Y(_abc_40298_new_n1273_));
OAI21X1 OAI21X1_137 ( .A(_abc_40298_new_n888_), .B(_abc_40298_new_n1027_), .C(_abc_40298_new_n1259_), .Y(_abc_40298_new_n1274_));
OAI21X1 OAI21X1_138 ( .A(_abc_40298_new_n1273_), .B(_abc_40298_new_n1071_), .C(_abc_40298_new_n1274_), .Y(_abc_40298_new_n1275_));
OAI21X1 OAI21X1_139 ( .A(epc_q_4_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n1276_));
OAI21X1 OAI21X1_14 ( .A(_abc_40298_new_n631_), .B(_abc_40298_new_n704_), .C(_abc_40298_new_n693_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_1_));
OAI21X1 OAI21X1_140 ( .A(_abc_40298_new_n1000_), .B(_abc_40298_new_n1177_), .C(REGFILE_SIM_reg_bank_reg_rb_o_5_), .Y(_abc_40298_new_n1285_));
OAI21X1 OAI21X1_141 ( .A(_abc_40298_new_n1176_), .B(_abc_40298_new_n1284_), .C(_abc_40298_new_n1285_), .Y(_abc_40298_new_n1286_));
OAI21X1 OAI21X1_142 ( .A(_abc_40298_new_n1232_), .B(_abc_40298_new_n1286_), .C(_abc_40298_new_n1291_), .Y(_abc_40298_new_n1292_));
OAI21X1 OAI21X1_143 ( .A(_abc_40298_new_n992_), .B(_abc_40298_new_n1185_), .C(epc_q_5_), .Y(_abc_40298_new_n1294_));
OAI21X1 OAI21X1_144 ( .A(_abc_40298_new_n1293_), .B(_abc_40298_new_n1187_), .C(_abc_40298_new_n1294_), .Y(_abc_40298_new_n1295_));
OAI21X1 OAI21X1_145 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1292_), .C(_abc_40298_new_n1296_), .Y(_abc_40298_new_n1297_));
OAI21X1 OAI21X1_146 ( .A(_abc_40298_new_n888_), .B(_abc_40298_new_n1027_), .C(_abc_40298_new_n1290_), .Y(_abc_40298_new_n1298_));
OAI21X1 OAI21X1_147 ( .A(_abc_40298_new_n1297_), .B(_abc_40298_new_n1071_), .C(_abc_40298_new_n1298_), .Y(_abc_40298_new_n1299_));
OAI21X1 OAI21X1_148 ( .A(epc_q_5_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n1300_));
OAI21X1 OAI21X1_149 ( .A(_abc_40298_new_n1287_), .B(_abc_40298_new_n1258_), .C(_abc_40298_new_n1302_), .Y(_abc_40298_new_n1303_));
OAI21X1 OAI21X1_15 ( .A(_abc_40298_new_n707_), .B(_abc_40298_new_n695_), .C(_abc_40298_new_n708_), .Y(_abc_40298_new_n709_));
OAI21X1 OAI21X1_150 ( .A(_abc_40298_new_n1138_), .B(_abc_40298_new_n1306_), .C(_abc_40298_new_n1169_), .Y(_abc_40298_new_n1307_));
OAI21X1 OAI21X1_151 ( .A(_abc_40298_new_n1313_), .B(_abc_40298_new_n1318_), .C(_abc_40298_new_n1319_), .Y(_abc_40298_new_n1320_));
OAI21X1 OAI21X1_152 ( .A(_abc_40298_new_n1309_), .B(_abc_40298_new_n1066_), .C(_abc_40298_new_n1320_), .Y(_abc_40298_new_n1321_));
OAI21X1 OAI21X1_153 ( .A(_abc_40298_new_n1322_), .B(_abc_40298_new_n1175_), .C(_abc_40298_new_n1213_), .Y(_abc_40298_new_n1323_));
OAI21X1 OAI21X1_154 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1325_), .C(_abc_40298_new_n1327_), .Y(_abc_40298_new_n1328_));
OAI21X1 OAI21X1_155 ( .A(epc_q_6_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n1329_));
OAI21X1 OAI21X1_156 ( .A(_abc_40298_new_n1138_), .B(_abc_40298_new_n1334_), .C(_abc_40298_new_n1169_), .Y(_abc_40298_new_n1335_));
OAI21X1 OAI21X1_157 ( .A(_abc_40298_new_n1314_), .B(_abc_40298_new_n1344_), .C(_abc_40298_new_n1345_), .Y(_abc_40298_new_n1346_));
OAI21X1 OAI21X1_158 ( .A(_abc_40298_new_n1350_), .B(_abc_40298_new_n1344_), .C(_abc_40298_new_n1351_), .Y(_abc_40298_new_n1352_));
OAI21X1 OAI21X1_159 ( .A(_abc_40298_new_n1338_), .B(_abc_40298_new_n1175_), .C(_abc_40298_new_n1354_), .Y(_abc_40298_new_n1355_));
OAI21X1 OAI21X1_16 ( .A(_abc_40298_new_n707_), .B(_abc_40298_new_n699_), .C(_abc_40298_new_n711_), .Y(_abc_40298_new_n712_));
OAI21X1 OAI21X1_160 ( .A(_abc_40298_new_n1331_), .B(_abc_40298_new_n1333_), .C(_abc_40298_new_n1232_), .Y(_abc_40298_new_n1356_));
OAI21X1 OAI21X1_161 ( .A(_abc_40298_new_n1232_), .B(_abc_40298_new_n1355_), .C(_abc_40298_new_n1356_), .Y(_abc_40298_new_n1357_));
OAI21X1 OAI21X1_162 ( .A(_abc_40298_new_n1337_), .B(_abc_40298_new_n1358_), .C(_abc_40298_new_n1028_), .Y(_abc_40298_new_n1359_));
OAI21X1 OAI21X1_163 ( .A(epc_q_7_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n1360_));
OAI21X1 OAI21X1_164 ( .A(_abc_40298_new_n1332_), .B(_abc_40298_new_n1305_), .C(_abc_40298_new_n1362_), .Y(_abc_40298_new_n1363_));
OAI21X1 OAI21X1_165 ( .A(_abc_40298_new_n1365_), .B(_abc_40298_new_n1028_), .C(REGFILE_SIM_reg_bank_wr_i), .Y(_abc_40298_new_n1366_));
OAI21X1 OAI21X1_166 ( .A(_abc_40298_new_n1340_), .B(_abc_40298_new_n1345_), .C(_abc_40298_new_n1370_), .Y(_abc_40298_new_n1371_));
OAI21X1 OAI21X1_167 ( .A(_abc_40298_new_n1373_), .B(_abc_40298_new_n1376_), .C(_abc_40298_new_n1378_), .Y(_abc_40298_new_n1379_));
OAI21X1 OAI21X1_168 ( .A(_abc_40298_new_n1369_), .B(_abc_40298_new_n1066_), .C(_abc_40298_new_n1379_), .Y(_abc_40298_new_n1380_));
OAI21X1 OAI21X1_169 ( .A(_abc_40298_new_n1368_), .B(_abc_40298_new_n1175_), .C(_abc_40298_new_n1381_), .Y(_abc_40298_new_n1382_));
OAI21X1 OAI21X1_17 ( .A(_abc_40298_new_n631_), .B(_abc_40298_new_n715_), .C(_abc_40298_new_n706_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_2_));
OAI21X1 OAI21X1_170 ( .A(_abc_40298_new_n1232_), .B(_abc_40298_new_n1382_), .C(_abc_40298_new_n1383_), .Y(_abc_40298_new_n1384_));
OAI21X1 OAI21X1_171 ( .A(_abc_40298_new_n1070_), .B(_abc_40298_new_n1173_), .C(_abc_40298_new_n1385_), .Y(_abc_40298_new_n1386_));
OAI21X1 OAI21X1_172 ( .A(_abc_40298_new_n1134_), .B(_abc_40298_new_n1367_), .C(_abc_40298_new_n1386_), .Y(_abc_40298_new_n1387_));
OAI21X1 OAI21X1_173 ( .A(epc_q_8_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n1389_));
OAI21X1 OAI21X1_174 ( .A(_abc_40298_new_n1138_), .B(_abc_40298_new_n1391_), .C(_abc_40298_new_n1169_), .Y(_abc_40298_new_n1392_));
OAI21X1 OAI21X1_175 ( .A(_abc_40298_new_n983_), .B(_abc_40298_new_n1396_), .C(_abc_40298_new_n1066_), .Y(_abc_40298_new_n1397_));
OAI21X1 OAI21X1_176 ( .A(_abc_40298_new_n1398_), .B(_abc_40298_new_n1400_), .C(_abc_40298_new_n1401_), .Y(_abc_40298_new_n1402_));
OAI21X1 OAI21X1_177 ( .A(_abc_40298_new_n1375_), .B(_abc_40298_new_n1377_), .C(_abc_40298_new_n1403_), .Y(_abc_40298_new_n1404_));
OAI21X1 OAI21X1_178 ( .A(_abc_40298_new_n1140_), .B(_abc_40298_new_n1175_), .C(_abc_40298_new_n1213_), .Y(_abc_40298_new_n1408_));
OAI21X1 OAI21X1_179 ( .A(_abc_40298_new_n1394_), .B(_abc_40298_new_n1410_), .C(_abc_40298_new_n1028_), .Y(_abc_40298_new_n1411_));
OAI21X1 OAI21X1_18 ( .A(_abc_40298_new_n718_), .B(_abc_40298_new_n695_), .C(_abc_40298_new_n719_), .Y(_abc_40298_new_n720_));
OAI21X1 OAI21X1_180 ( .A(epc_q_9_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n1412_));
OAI21X1 OAI21X1_181 ( .A(_abc_40298_new_n1399_), .B(_abc_40298_new_n1364_), .C(_abc_40298_new_n1414_), .Y(_abc_40298_new_n1415_));
OAI21X1 OAI21X1_182 ( .A(_abc_40298_new_n1138_), .B(_abc_40298_new_n1419_), .C(_abc_40298_new_n1169_), .Y(_abc_40298_new_n1420_));
OAI21X1 OAI21X1_183 ( .A(_abc_40298_new_n973_), .B(_abc_40298_new_n1399_), .C(_abc_40298_new_n1425_), .Y(_abc_40298_new_n1426_));
OAI21X1 OAI21X1_184 ( .A(_abc_40298_new_n1426_), .B(_abc_40298_new_n1424_), .C(_abc_40298_new_n1430_), .Y(_abc_40298_new_n1431_));
OAI21X1 OAI21X1_185 ( .A(_abc_40298_new_n1432_), .B(_abc_40298_new_n1435_), .C(_abc_40298_new_n985_), .Y(_abc_40298_new_n1436_));
OAI21X1 OAI21X1_186 ( .A(_abc_40298_new_n1213_), .B(_abc_40298_new_n1419_), .C(_abc_40298_new_n1440_), .Y(_abc_40298_new_n1441_));
OAI21X1 OAI21X1_187 ( .A(_abc_40298_new_n1422_), .B(_abc_40298_new_n1442_), .C(_abc_40298_new_n1028_), .Y(_abc_40298_new_n1443_));
OAI21X1 OAI21X1_188 ( .A(epc_q_10_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n1444_));
OAI21X1 OAI21X1_189 ( .A(_abc_40298_new_n1138_), .B(_abc_40298_new_n1450_), .C(_abc_40298_new_n1169_), .Y(_abc_40298_new_n1451_));
OAI21X1 OAI21X1_19 ( .A(_abc_40298_new_n718_), .B(_abc_40298_new_n699_), .C(_abc_40298_new_n722_), .Y(_abc_40298_new_n723_));
OAI21X1 OAI21X1_190 ( .A(_abc_40298_new_n1455_), .B(_abc_40298_new_n1414_), .C(_abc_40298_new_n1431_), .Y(_abc_40298_new_n1456_));
OAI21X1 OAI21X1_191 ( .A(_abc_40298_new_n1456_), .B(_abc_40298_new_n1461_), .C(_abc_40298_new_n1462_), .Y(_abc_40298_new_n1463_));
OAI21X1 OAI21X1_192 ( .A(_abc_40298_new_n1454_), .B(_abc_40298_new_n1066_), .C(_abc_40298_new_n1463_), .Y(_abc_40298_new_n1464_));
OAI21X1 OAI21X1_193 ( .A(_abc_40298_new_n1466_), .B(_abc_40298_new_n1175_), .C(_abc_40298_new_n1213_), .Y(_abc_40298_new_n1467_));
OAI21X1 OAI21X1_194 ( .A(_abc_40298_new_n1453_), .B(_abc_40298_new_n1469_), .C(_abc_40298_new_n1028_), .Y(_abc_40298_new_n1470_));
OAI21X1 OAI21X1_195 ( .A(epc_q_11_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n1471_));
OAI21X1 OAI21X1_196 ( .A(_abc_40298_new_n1447_), .B(_abc_40298_new_n1417_), .C(_abc_40298_new_n1473_), .Y(_abc_40298_new_n1474_));
OAI21X1 OAI21X1_197 ( .A(_abc_40298_new_n1138_), .B(_abc_40298_new_n1476_), .C(_abc_40298_new_n1169_), .Y(_abc_40298_new_n1477_));
OAI21X1 OAI21X1_198 ( .A(_abc_40298_new_n1484_), .B(_abc_40298_new_n1488_), .C(_abc_40298_new_n1493_), .Y(_abc_40298_new_n1494_));
OAI21X1 OAI21X1_199 ( .A(_abc_40298_new_n1489_), .B(_abc_40298_new_n1493_), .C(_abc_40298_new_n1496_), .Y(_abc_40298_new_n1497_));
OAI21X1 OAI21X1_2 ( .A(_abc_40298_new_n630_), .B(_abc_40298_new_n631_), .C(_abc_40298_new_n632_), .Y(_abc_27663_auto_fsm_map_cc_170_map_fsm_2376_3_));
OAI21X1 OAI21X1_20 ( .A(_abc_40298_new_n631_), .B(_abc_40298_new_n726_), .C(_abc_40298_new_n717_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_3_));
OAI21X1 OAI21X1_200 ( .A(_abc_40298_new_n1479_), .B(_abc_40298_new_n1066_), .C(_abc_40298_new_n1497_), .Y(_abc_40298_new_n1498_));
OAI21X1 OAI21X1_201 ( .A(_abc_40298_new_n1478_), .B(_abc_40298_new_n1175_), .C(_abc_40298_new_n1499_), .Y(_abc_40298_new_n1500_));
OAI21X1 OAI21X1_202 ( .A(_abc_40298_new_n1232_), .B(_abc_40298_new_n1500_), .C(_abc_40298_new_n1501_), .Y(_abc_40298_new_n1502_));
OAI21X1 OAI21X1_203 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1503_), .C(_abc_40298_new_n1505_), .Y(_abc_40298_new_n1506_));
OAI21X1 OAI21X1_204 ( .A(epc_q_12_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n1507_));
OAI21X1 OAI21X1_205 ( .A(_abc_40298_new_n1138_), .B(_abc_40298_new_n1509_), .C(_abc_40298_new_n1169_), .Y(_abc_40298_new_n1510_));
OAI21X1 OAI21X1_206 ( .A(_abc_40298_new_n1484_), .B(_abc_40298_new_n1488_), .C(_abc_40298_new_n1516_), .Y(_abc_40298_new_n1517_));
OAI21X1 OAI21X1_207 ( .A(_abc_40298_new_n1491_), .B(_abc_40298_new_n1519_), .C(_abc_40298_new_n985_), .Y(_abc_40298_new_n1520_));
OAI21X1 OAI21X1_208 ( .A(_abc_40298_new_n1232_), .B(_abc_40298_new_n1524_), .C(_abc_40298_new_n1525_), .Y(_abc_40298_new_n1526_));
OAI21X1 OAI21X1_209 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1526_), .C(_abc_40298_new_n1528_), .Y(_abc_40298_new_n1529_));
OAI21X1 OAI21X1_21 ( .A(_abc_40298_new_n655_), .B(_abc_40298_new_n732_), .C(_abc_40298_new_n734_), .Y(_abc_40298_new_n735_));
OAI21X1 OAI21X1_210 ( .A(epc_q_13_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n1530_));
OAI21X1 OAI21X1_211 ( .A(_abc_40298_new_n1512_), .B(_abc_40298_new_n1475_), .C(_abc_40298_new_n1532_), .Y(_abc_40298_new_n1533_));
OAI21X1 OAI21X1_212 ( .A(_abc_40298_new_n1138_), .B(_abc_40298_new_n1537_), .C(_abc_40298_new_n1169_), .Y(_abc_40298_new_n1538_));
OAI21X1 OAI21X1_213 ( .A(_abc_40298_new_n1491_), .B(_abc_40298_new_n1511_), .C(_abc_40298_new_n1541_), .Y(_abc_40298_new_n1542_));
OAI21X1 OAI21X1_214 ( .A(_abc_40298_new_n1542_), .B(_abc_40298_new_n1540_), .C(_abc_40298_new_n1546_), .Y(_abc_40298_new_n1547_));
OAI21X1 OAI21X1_215 ( .A(_abc_40298_new_n1519_), .B(_abc_40298_new_n1494_), .C(_abc_40298_new_n1549_), .Y(_abc_40298_new_n1550_));
OAI21X1 OAI21X1_216 ( .A(_abc_40298_new_n1546_), .B(_abc_40298_new_n1550_), .C(_abc_40298_new_n985_), .Y(_abc_40298_new_n1551_));
OAI21X1 OAI21X1_217 ( .A(_abc_40298_new_n1551_), .B(_abc_40298_new_n1548_), .C(_abc_40298_new_n1539_), .Y(_abc_40298_new_n1552_));
OAI21X1 OAI21X1_218 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1555_), .C(_abc_40298_new_n1557_), .Y(_abc_40298_new_n1558_));
OAI21X1 OAI21X1_219 ( .A(epc_q_14_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n1559_));
OAI21X1 OAI21X1_22 ( .A(state_q_1_), .B(_abc_40298_new_n728_), .C(_abc_40298_new_n735_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_4_));
OAI21X1 OAI21X1_220 ( .A(_abc_40298_new_n1532_), .B(_abc_40298_new_n1562_), .C(_abc_40298_new_n1561_), .Y(_abc_40298_new_n1563_));
OAI21X1 OAI21X1_221 ( .A(_abc_40298_new_n1138_), .B(_abc_40298_new_n1566_), .C(_abc_40298_new_n1169_), .Y(_abc_40298_new_n1567_));
OAI21X1 OAI21X1_222 ( .A(_abc_40298_new_n1545_), .B(_abc_40298_new_n1548_), .C(_abc_40298_new_n1573_), .Y(_abc_40298_new_n1576_));
OAI21X1 OAI21X1_223 ( .A(_abc_40298_new_n1569_), .B(_abc_40298_new_n1066_), .C(_abc_40298_new_n1577_), .Y(_abc_40298_new_n1578_));
OAI21X1 OAI21X1_224 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1581_), .C(_abc_40298_new_n1583_), .Y(_abc_40298_new_n1584_));
OAI21X1 OAI21X1_225 ( .A(epc_q_15_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n1585_));
OAI21X1 OAI21X1_226 ( .A(_abc_40298_new_n1561_), .B(_abc_40298_new_n1535_), .C(_abc_40298_new_n1587_), .Y(_abc_40298_new_n1588_));
OAI21X1 OAI21X1_227 ( .A(_abc_40298_new_n1138_), .B(_abc_40298_new_n1590_), .C(_abc_40298_new_n1169_), .Y(_abc_40298_new_n1591_));
OAI21X1 OAI21X1_228 ( .A(_abc_40298_new_n1000_), .B(_abc_40298_new_n1177_), .C(REGFILE_SIM_reg_bank_reg_rb_o_16_), .Y(_abc_40298_new_n1592_));
OAI21X1 OAI21X1_229 ( .A(_abc_40298_new_n1596_), .B(_abc_40298_new_n1549_), .C(_abc_40298_new_n1597_), .Y(_abc_40298_new_n1598_));
OAI21X1 OAI21X1_23 ( .A(_abc_40298_new_n655_), .B(_abc_40298_new_n741_), .C(_abc_40298_new_n743_), .Y(_abc_40298_new_n744_));
OAI21X1 OAI21X1_230 ( .A(_abc_40298_new_n1607_), .B(_abc_40298_new_n1602_), .C(_abc_40298_new_n985_), .Y(_abc_40298_new_n1608_));
OAI21X1 OAI21X1_231 ( .A(_abc_40298_new_n1176_), .B(_abc_40298_new_n1610_), .C(_abc_40298_new_n1592_), .Y(_abc_40298_new_n1611_));
OAI21X1 OAI21X1_232 ( .A(_abc_40298_new_n1232_), .B(_abc_40298_new_n1611_), .C(_abc_40298_new_n1612_), .Y(_abc_40298_new_n1613_));
OAI21X1 OAI21X1_233 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1614_), .C(_abc_40298_new_n1616_), .Y(_abc_40298_new_n1617_));
OAI21X1 OAI21X1_234 ( .A(epc_q_16_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n1618_));
OAI21X1 OAI21X1_235 ( .A(_abc_40298_new_n1587_), .B(_abc_40298_new_n1565_), .C(_abc_40298_new_n1620_), .Y(_abc_40298_new_n1621_));
OAI21X1 OAI21X1_236 ( .A(_abc_40298_new_n1138_), .B(_abc_40298_new_n1623_), .C(_abc_40298_new_n1169_), .Y(_abc_40298_new_n1624_));
OAI21X1 OAI21X1_237 ( .A(_abc_40298_new_n984_), .B(_abc_40298_new_n1634_), .C(_abc_40298_new_n1626_), .Y(_abc_40298_new_n1635_));
OAI21X1 OAI21X1_238 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1638_), .C(_abc_40298_new_n1640_), .Y(_abc_40298_new_n1641_));
OAI21X1 OAI21X1_239 ( .A(epc_q_17_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n1642_));
OAI21X1 OAI21X1_24 ( .A(state_q_1_), .B(_abc_40298_new_n737_), .C(_abc_40298_new_n744_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_5_));
OAI21X1 OAI21X1_240 ( .A(_abc_40298_new_n1620_), .B(_abc_40298_new_n1589_), .C(_abc_40298_new_n1644_), .Y(_abc_40298_new_n1645_));
OAI21X1 OAI21X1_241 ( .A(_abc_40298_new_n1138_), .B(_abc_40298_new_n1649_), .C(_abc_40298_new_n1169_), .Y(_abc_40298_new_n1650_));
OAI21X1 OAI21X1_242 ( .A(_abc_40298_new_n1660_), .B(_abc_40298_new_n1663_), .C(_abc_40298_new_n985_), .Y(_abc_40298_new_n1664_));
OAI21X1 OAI21X1_243 ( .A(_abc_40298_new_n1662_), .B(_abc_40298_new_n1664_), .C(_abc_40298_new_n1651_), .Y(_abc_40298_new_n1665_));
OAI21X1 OAI21X1_244 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1668_), .C(_abc_40298_new_n1670_), .Y(_abc_40298_new_n1671_));
OAI21X1 OAI21X1_245 ( .A(epc_q_18_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n1672_));
OAI21X1 OAI21X1_246 ( .A(_abc_40298_new_n1138_), .B(_abc_40298_new_n1677_), .C(_abc_40298_new_n1169_), .Y(_abc_40298_new_n1678_));
OAI21X1 OAI21X1_247 ( .A(_abc_40298_new_n1685_), .B(_abc_40298_new_n1681_), .C(_abc_40298_new_n985_), .Y(_abc_40298_new_n1687_));
OAI21X1 OAI21X1_248 ( .A(_abc_40298_new_n1686_), .B(_abc_40298_new_n1687_), .C(_abc_40298_new_n1680_), .Y(_abc_40298_new_n1688_));
OAI21X1 OAI21X1_249 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1691_), .C(_abc_40298_new_n1693_), .Y(_abc_40298_new_n1694_));
OAI21X1 OAI21X1_25 ( .A(_abc_40298_new_n747_), .B(_abc_40298_new_n695_), .C(_abc_40298_new_n748_), .Y(_abc_40298_new_n749_));
OAI21X1 OAI21X1_250 ( .A(epc_q_19_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n1695_));
OAI21X1 OAI21X1_251 ( .A(_abc_40298_new_n1675_), .B(_abc_40298_new_n1647_), .C(_abc_40298_new_n1697_), .Y(_abc_40298_new_n1698_));
OAI21X1 OAI21X1_252 ( .A(_abc_40298_new_n1138_), .B(_abc_40298_new_n1701_), .C(_abc_40298_new_n1169_), .Y(_abc_40298_new_n1702_));
OAI21X1 OAI21X1_253 ( .A(_abc_40298_new_n1704_), .B(_abc_40298_new_n1654_), .C(_abc_40298_new_n1705_), .Y(_abc_40298_new_n1706_));
OAI21X1 OAI21X1_254 ( .A(_abc_40298_new_n1709_), .B(_abc_40298_new_n1602_), .C(_abc_40298_new_n1707_), .Y(_abc_40298_new_n1710_));
OAI21X1 OAI21X1_255 ( .A(_abc_40298_new_n1714_), .B(_abc_40298_new_n1710_), .C(_abc_40298_new_n985_), .Y(_abc_40298_new_n1716_));
OAI21X1 OAI21X1_256 ( .A(_abc_40298_new_n1715_), .B(_abc_40298_new_n1716_), .C(_abc_40298_new_n1703_), .Y(_abc_40298_new_n1717_));
OAI21X1 OAI21X1_257 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1720_), .C(_abc_40298_new_n1722_), .Y(_abc_40298_new_n1723_));
OAI21X1 OAI21X1_258 ( .A(epc_q_20_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n1724_));
OAI21X1 OAI21X1_259 ( .A(_abc_40298_new_n1138_), .B(_abc_40298_new_n1729_), .C(_abc_40298_new_n1169_), .Y(_abc_40298_new_n1730_));
OAI21X1 OAI21X1_26 ( .A(_abc_40298_new_n631_), .B(_abc_40298_new_n753_), .C(_abc_40298_new_n746_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_6_));
OAI21X1 OAI21X1_260 ( .A(_abc_40298_new_n1734_), .B(_abc_40298_new_n1736_), .C(_abc_40298_new_n1733_), .Y(_abc_40298_new_n1737_));
OAI21X1 OAI21X1_261 ( .A(_abc_40298_new_n1741_), .B(_abc_40298_new_n1739_), .C(_abc_40298_new_n1742_), .Y(_abc_40298_new_n1743_));
OAI21X1 OAI21X1_262 ( .A(_abc_40298_new_n1743_), .B(_abc_40298_new_n1738_), .C(_abc_40298_new_n1732_), .Y(_abc_40298_new_n1744_));
OAI21X1 OAI21X1_263 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1747_), .C(_abc_40298_new_n1749_), .Y(_abc_40298_new_n1750_));
OAI21X1 OAI21X1_264 ( .A(epc_q_21_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n1751_));
OAI21X1 OAI21X1_265 ( .A(_abc_40298_new_n1726_), .B(_abc_40298_new_n1699_), .C(_abc_40298_new_n1753_), .Y(_abc_40298_new_n1754_));
OAI21X1 OAI21X1_266 ( .A(_abc_40298_new_n1138_), .B(_abc_40298_new_n1758_), .C(_abc_40298_new_n1169_), .Y(_abc_40298_new_n1759_));
OAI21X1 OAI21X1_267 ( .A(_abc_40298_new_n1726_), .B(_abc_40298_new_n1735_), .C(_abc_40298_new_n1762_), .Y(_abc_40298_new_n1763_));
OAI21X1 OAI21X1_268 ( .A(_abc_40298_new_n1768_), .B(_abc_40298_new_n1771_), .C(_abc_40298_new_n985_), .Y(_abc_40298_new_n1772_));
OAI21X1 OAI21X1_269 ( .A(_abc_40298_new_n1770_), .B(_abc_40298_new_n1772_), .C(_abc_40298_new_n1760_), .Y(_abc_40298_new_n1773_));
OAI21X1 OAI21X1_27 ( .A(_abc_40298_new_n655_), .B(_abc_40298_new_n757_), .C(_abc_40298_new_n759_), .Y(_abc_40298_new_n760_));
OAI21X1 OAI21X1_270 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1776_), .C(_abc_40298_new_n1778_), .Y(_abc_40298_new_n1779_));
OAI21X1 OAI21X1_271 ( .A(epc_q_22_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n1780_));
OAI21X1 OAI21X1_272 ( .A(_abc_40298_new_n1138_), .B(_abc_40298_new_n1785_), .C(_abc_40298_new_n1169_), .Y(_abc_40298_new_n1786_));
OAI21X1 OAI21X1_273 ( .A(_abc_40298_new_n1793_), .B(_abc_40298_new_n1789_), .C(_abc_40298_new_n985_), .Y(_abc_40298_new_n1795_));
OAI21X1 OAI21X1_274 ( .A(_abc_40298_new_n1794_), .B(_abc_40298_new_n1795_), .C(_abc_40298_new_n1788_), .Y(_abc_40298_new_n1796_));
OAI21X1 OAI21X1_275 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1799_), .C(_abc_40298_new_n1801_), .Y(_abc_40298_new_n1802_));
OAI21X1 OAI21X1_276 ( .A(epc_q_23_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n1803_));
OAI21X1 OAI21X1_277 ( .A(_abc_40298_new_n1783_), .B(_abc_40298_new_n1756_), .C(_abc_40298_new_n1805_), .Y(_abc_40298_new_n1806_));
OAI21X1 OAI21X1_278 ( .A(_abc_40298_new_n1138_), .B(_abc_40298_new_n1809_), .C(_abc_40298_new_n1169_), .Y(_abc_40298_new_n1810_));
OAI21X1 OAI21X1_279 ( .A(_abc_40298_new_n1812_), .B(_abc_40298_new_n1814_), .C(_abc_40298_new_n1815_), .Y(_abc_40298_new_n1816_));
OAI21X1 OAI21X1_28 ( .A(_abc_40298_new_n631_), .B(_abc_40298_new_n760_), .C(_abc_40298_new_n761_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_7_));
OAI21X1 OAI21X1_280 ( .A(_abc_40298_new_n1601_), .B(_abc_40298_new_n1599_), .C(_abc_40298_new_n1819_), .Y(_abc_40298_new_n1820_));
OAI21X1 OAI21X1_281 ( .A(_abc_40298_new_n1827_), .B(_abc_40298_new_n1826_), .C(_abc_40298_new_n985_), .Y(_abc_40298_new_n1828_));
OAI21X1 OAI21X1_282 ( .A(_abc_40298_new_n1825_), .B(_abc_40298_new_n1828_), .C(_abc_40298_new_n1829_), .Y(_abc_40298_new_n1830_));
OAI21X1 OAI21X1_283 ( .A(_abc_40298_new_n1811_), .B(_abc_40298_new_n1175_), .C(_abc_40298_new_n1831_), .Y(_abc_40298_new_n1832_));
OAI21X1 OAI21X1_284 ( .A(_abc_40298_new_n1232_), .B(_abc_40298_new_n1832_), .C(_abc_40298_new_n1833_), .Y(_abc_40298_new_n1834_));
OAI21X1 OAI21X1_285 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1835_), .C(_abc_40298_new_n1837_), .Y(_abc_40298_new_n1838_));
OAI21X1 OAI21X1_286 ( .A(epc_q_24_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n1839_));
OAI21X1 OAI21X1_287 ( .A(_abc_40298_new_n1138_), .B(_abc_40298_new_n1841_), .C(_abc_40298_new_n1169_), .Y(_abc_40298_new_n1842_));
OAI21X1 OAI21X1_288 ( .A(_abc_40298_new_n1822_), .B(_abc_40298_new_n1826_), .C(_abc_40298_new_n1847_), .Y(_abc_40298_new_n1848_));
OAI21X1 OAI21X1_289 ( .A(_abc_40298_new_n984_), .B(_abc_40298_new_n1849_), .C(_abc_40298_new_n1851_), .Y(_abc_40298_new_n1852_));
OAI21X1 OAI21X1_29 ( .A(\mem_dat_i[8] ), .B(_abc_40298_new_n686_), .C(_abc_40298_new_n764_), .Y(_abc_40298_new_n765_));
OAI21X1 OAI21X1_290 ( .A(_abc_40298_new_n1070_), .B(_abc_40298_new_n1173_), .C(_abc_40298_new_n1855_), .Y(_abc_40298_new_n1856_));
OAI21X1 OAI21X1_291 ( .A(epc_q_25_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n1860_));
OAI21X1 OAI21X1_292 ( .A(_abc_40298_new_n1844_), .B(_abc_40298_new_n1807_), .C(_abc_40298_new_n1862_), .Y(_abc_40298_new_n1863_));
OAI21X1 OAI21X1_293 ( .A(_abc_40298_new_n1138_), .B(_abc_40298_new_n1866_), .C(_abc_40298_new_n1169_), .Y(_abc_40298_new_n1867_));
OAI21X1 OAI21X1_294 ( .A(_abc_40298_new_n1878_), .B(_abc_40298_new_n1874_), .C(_abc_40298_new_n985_), .Y(_abc_40298_new_n1879_));
OAI21X1 OAI21X1_295 ( .A(_abc_40298_new_n1881_), .B(_abc_40298_new_n1880_), .C(_abc_40298_new_n1175_), .Y(_abc_40298_new_n1882_));
OAI21X1 OAI21X1_296 ( .A(_abc_40298_new_n1868_), .B(_abc_40298_new_n1175_), .C(_abc_40298_new_n1882_), .Y(_abc_40298_new_n1883_));
OAI21X1 OAI21X1_297 ( .A(_abc_40298_new_n1070_), .B(_abc_40298_new_n1173_), .C(_abc_40298_new_n1884_), .Y(_abc_40298_new_n1885_));
OAI21X1 OAI21X1_298 ( .A(epc_q_26_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n1889_));
OAI21X1 OAI21X1_299 ( .A(_abc_40298_new_n1138_), .B(_abc_40298_new_n1892_), .C(_abc_40298_new_n1169_), .Y(_abc_40298_new_n1893_));
OAI21X1 OAI21X1_3 ( .A(inst_r_1_), .B(inst_r_0_), .C(_abc_40298_new_n641_), .Y(_abc_40298_new_n642_));
OAI21X1 OAI21X1_30 ( .A(\mem_dat_i[12] ), .B(_abc_40298_new_n686_), .C(_abc_40298_new_n786_), .Y(_abc_40298_new_n787_));
OAI21X1 OAI21X1_300 ( .A(_abc_40298_new_n1875_), .B(_abc_40298_new_n1874_), .C(_abc_40298_new_n1898_), .Y(_abc_40298_new_n1899_));
OAI21X1 OAI21X1_301 ( .A(_abc_40298_new_n984_), .B(_abc_40298_new_n1900_), .C(_abc_40298_new_n1901_), .Y(_abc_40298_new_n1902_));
OAI21X1 OAI21X1_302 ( .A(_abc_40298_new_n1232_), .B(_abc_40298_new_n1903_), .C(_abc_40298_new_n1904_), .Y(_abc_40298_new_n1905_));
OAI21X1 OAI21X1_303 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1905_), .C(_abc_40298_new_n1907_), .Y(_abc_40298_new_n1908_));
OAI21X1 OAI21X1_304 ( .A(epc_q_27_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n1909_));
OAI21X1 OAI21X1_305 ( .A(_abc_40298_new_n1895_), .B(_abc_40298_new_n1865_), .C(_abc_40298_new_n1911_), .Y(_abc_40298_new_n1912_));
OAI21X1 OAI21X1_306 ( .A(_abc_40298_new_n1138_), .B(_abc_40298_new_n1914_), .C(_abc_40298_new_n1169_), .Y(_abc_40298_new_n1915_));
OAI21X1 OAI21X1_307 ( .A(_abc_40298_new_n1922_), .B(_abc_40298_new_n1872_), .C(_abc_40298_new_n1923_), .Y(_abc_40298_new_n1924_));
OAI21X1 OAI21X1_308 ( .A(_abc_40298_new_n1232_), .B(_abc_40298_new_n1933_), .C(_abc_40298_new_n1934_), .Y(_abc_40298_new_n1935_));
OAI21X1 OAI21X1_309 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1935_), .C(_abc_40298_new_n1937_), .Y(_abc_40298_new_n1938_));
OAI21X1 OAI21X1_31 ( .A(\mem_dat_i[13] ), .B(_abc_40298_new_n686_), .C(_abc_40298_new_n790_), .Y(_abc_40298_new_n791_));
OAI21X1 OAI21X1_310 ( .A(epc_q_28_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n1939_));
OAI21X1 OAI21X1_311 ( .A(_abc_40298_new_n1138_), .B(_abc_40298_new_n1941_), .C(_abc_40298_new_n1169_), .Y(_abc_40298_new_n1942_));
OAI21X1 OAI21X1_312 ( .A(_abc_40298_new_n1945_), .B(_abc_40298_new_n1943_), .C(_abc_40298_new_n985_), .Y(_abc_40298_new_n1947_));
OAI21X1 OAI21X1_313 ( .A(_abc_40298_new_n1946_), .B(_abc_40298_new_n1947_), .C(_abc_40298_new_n1948_), .Y(_abc_40298_new_n1949_));
OAI21X1 OAI21X1_314 ( .A(_abc_40298_new_n1000_), .B(_abc_40298_new_n1177_), .C(_abc_40298_new_n1950_), .Y(_abc_40298_new_n1951_));
OAI21X1 OAI21X1_315 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1954_), .C(_abc_40298_new_n1956_), .Y(_abc_40298_new_n1957_));
OAI21X1 OAI21X1_316 ( .A(epc_q_29_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n1958_));
OAI21X1 OAI21X1_317 ( .A(_abc_40298_new_n1960_), .B(_abc_40298_new_n1913_), .C(_abc_40298_new_n1961_), .Y(_abc_40298_new_n1962_));
OAI21X1 OAI21X1_318 ( .A(_abc_40298_new_n1138_), .B(_abc_40298_new_n1965_), .C(_abc_40298_new_n1169_), .Y(_abc_40298_new_n1966_));
OAI21X1 OAI21X1_319 ( .A(_abc_40298_new_n1924_), .B(_abc_40298_new_n1921_), .C(_abc_40298_new_n1968_), .Y(_abc_40298_new_n1969_));
OAI21X1 OAI21X1_32 ( .A(\mem_dat_i[15] ), .B(_abc_40298_new_n686_), .C(_abc_40298_new_n800_), .Y(_abc_40298_new_n801_));
OAI21X1 OAI21X1_320 ( .A(pc_q_28_), .B(pc_q_29_), .C(opcode_q_25_), .Y(_abc_40298_new_n1970_));
OAI21X1 OAI21X1_321 ( .A(_abc_40298_new_n1975_), .B(_abc_40298_new_n1971_), .C(_abc_40298_new_n985_), .Y(_abc_40298_new_n1976_));
OAI21X1 OAI21X1_322 ( .A(_abc_40298_new_n1978_), .B(_abc_40298_new_n1977_), .C(_abc_40298_new_n1175_), .Y(_abc_40298_new_n1979_));
OAI21X1 OAI21X1_323 ( .A(_abc_40298_new_n1967_), .B(_abc_40298_new_n1175_), .C(_abc_40298_new_n1979_), .Y(_abc_40298_new_n1980_));
OAI21X1 OAI21X1_324 ( .A(_abc_40298_new_n1168_), .B(_abc_40298_new_n1983_), .C(_abc_40298_new_n1985_), .Y(_abc_40298_new_n1986_));
OAI21X1 OAI21X1_325 ( .A(epc_q_30_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n1987_));
OAI21X1 OAI21X1_326 ( .A(pc_q_31_), .B(_abc_40298_new_n1991_), .C(_abc_40298_new_n985_), .Y(_abc_40298_new_n1993_));
OAI21X1 OAI21X1_327 ( .A(_abc_40298_new_n1992_), .B(_abc_40298_new_n1993_), .C(_abc_40298_new_n1994_), .Y(_abc_40298_new_n1995_));
OAI21X1 OAI21X1_328 ( .A(_abc_40298_new_n1000_), .B(_abc_40298_new_n1177_), .C(_abc_40298_new_n1996_), .Y(_abc_40298_new_n1997_));
OAI21X1 OAI21X1_329 ( .A(_abc_40298_new_n1961_), .B(_abc_40298_new_n2002_), .C(_abc_40298_new_n1999_), .Y(_abc_40298_new_n2003_));
OAI21X1 OAI21X1_33 ( .A(_abc_40298_new_n804_), .B(_abc_40298_new_n806_), .C(_abc_40298_new_n655_), .Y(_abc_40298_new_n807_));
OAI21X1 OAI21X1_330 ( .A(epc_q_31_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n2012_));
OAI21X1 OAI21X1_331 ( .A(next_pc_r_0_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n2016_));
OAI21X1 OAI21X1_332 ( .A(next_pc_r_1_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n2019_));
OAI21X1 OAI21X1_333 ( .A(pc_q_2_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n2022_));
OAI21X1 OAI21X1_334 ( .A(_abc_40298_new_n1244_), .B(_abc_40298_new_n2024_), .C(REGFILE_SIM_reg_bank_wr_i), .Y(_abc_40298_new_n2025_));
OAI21X1 OAI21X1_335 ( .A(pc_q_3_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n2025_), .Y(_abc_40298_new_n2026_));
OAI21X1 OAI21X1_336 ( .A(pc_q_4_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n2029_));
OAI21X1 OAI21X1_337 ( .A(_abc_40298_new_n1292_), .B(_abc_40298_new_n2024_), .C(REGFILE_SIM_reg_bank_wr_i), .Y(_abc_40298_new_n2031_));
OAI21X1 OAI21X1_338 ( .A(pc_q_5_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n2031_), .Y(_abc_40298_new_n2032_));
OAI21X1 OAI21X1_339 ( .A(pc_q_6_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n2035_));
OAI21X1 OAI21X1_34 ( .A(_abc_40298_new_n804_), .B(_abc_40298_new_n811_), .C(_abc_40298_new_n655_), .Y(_abc_40298_new_n812_));
OAI21X1 OAI21X1_340 ( .A(_abc_40298_new_n1357_), .B(_abc_40298_new_n2024_), .C(REGFILE_SIM_reg_bank_wr_i), .Y(_abc_40298_new_n2037_));
OAI21X1 OAI21X1_341 ( .A(pc_q_7_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n2037_), .Y(_abc_40298_new_n2038_));
OAI21X1 OAI21X1_342 ( .A(_abc_40298_new_n1134_), .B(_abc_40298_new_n1385_), .C(_abc_40298_new_n1170_), .Y(_abc_40298_new_n2040_));
OAI21X1 OAI21X1_343 ( .A(_abc_40298_new_n1362_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n2041_), .Y(_0pc_q_31_0__8_));
OAI21X1 OAI21X1_344 ( .A(inst_trap_w), .B(_abc_40298_new_n2044_), .C(_abc_40298_new_n2043_), .Y(_abc_40298_new_n2045_));
OAI21X1 OAI21X1_345 ( .A(pc_q_9_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n2047_));
OAI21X1 OAI21X1_346 ( .A(_abc_40298_new_n1173_), .B(_abc_40298_new_n1441_), .C(_abc_40298_new_n885_), .Y(_abc_40298_new_n2049_));
OAI21X1 OAI21X1_347 ( .A(_abc_40298_new_n888_), .B(_abc_40298_new_n2049_), .C(_abc_40298_new_n2043_), .Y(_abc_40298_new_n2050_));
OAI21X1 OAI21X1_348 ( .A(pc_q_10_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n2051_), .Y(_abc_40298_new_n2052_));
OAI21X1 OAI21X1_349 ( .A(_abc_40298_new_n1134_), .B(_abc_40298_new_n1468_), .C(_abc_40298_new_n2043_), .Y(_abc_40298_new_n2054_));
OAI21X1 OAI21X1_35 ( .A(_abc_40298_new_n804_), .B(_abc_40298_new_n816_), .C(_abc_40298_new_n655_), .Y(_abc_40298_new_n817_));
OAI21X1 OAI21X1_350 ( .A(pc_q_11_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n2056_));
OAI21X1 OAI21X1_351 ( .A(_abc_40298_new_n2024_), .B(_abc_40298_new_n1502_), .C(REGFILE_SIM_reg_bank_wr_i), .Y(_abc_40298_new_n2058_));
OAI21X1 OAI21X1_352 ( .A(pc_q_12_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n2058_), .Y(_abc_40298_new_n2059_));
OAI21X1 OAI21X1_353 ( .A(pc_q_13_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n2062_));
OAI21X1 OAI21X1_354 ( .A(pc_q_14_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n2065_));
OAI21X1 OAI21X1_355 ( .A(pc_q_15_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n2068_));
OAI21X1 OAI21X1_356 ( .A(_abc_40298_new_n2024_), .B(_abc_40298_new_n1613_), .C(REGFILE_SIM_reg_bank_wr_i), .Y(_abc_40298_new_n2070_));
OAI21X1 OAI21X1_357 ( .A(pc_q_16_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n2070_), .Y(_abc_40298_new_n2071_));
OAI21X1 OAI21X1_358 ( .A(pc_q_17_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n2074_));
OAI21X1 OAI21X1_359 ( .A(pc_q_18_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n2077_));
OAI21X1 OAI21X1_36 ( .A(_abc_40298_new_n804_), .B(_abc_40298_new_n821_), .C(_abc_40298_new_n655_), .Y(_abc_40298_new_n822_));
OAI21X1 OAI21X1_360 ( .A(pc_q_19_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n2080_));
OAI21X1 OAI21X1_361 ( .A(pc_q_20_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n2083_));
OAI21X1 OAI21X1_362 ( .A(pc_q_21_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n2086_));
OAI21X1 OAI21X1_363 ( .A(pc_q_22_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n2089_));
OAI21X1 OAI21X1_364 ( .A(pc_q_23_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n2092_));
OAI21X1 OAI21X1_365 ( .A(_abc_40298_new_n2024_), .B(_abc_40298_new_n1834_), .C(REGFILE_SIM_reg_bank_wr_i), .Y(_abc_40298_new_n2094_));
OAI21X1 OAI21X1_366 ( .A(pc_q_24_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n2094_), .Y(_abc_40298_new_n2095_));
OAI21X1 OAI21X1_367 ( .A(_abc_40298_new_n2024_), .B(_abc_40298_new_n1855_), .C(REGFILE_SIM_reg_bank_wr_i), .Y(_abc_40298_new_n2097_));
OAI21X1 OAI21X1_368 ( .A(pc_q_25_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n2097_), .Y(_abc_40298_new_n2098_));
OAI21X1 OAI21X1_369 ( .A(_abc_40298_new_n2024_), .B(_abc_40298_new_n1884_), .C(REGFILE_SIM_reg_bank_wr_i), .Y(_abc_40298_new_n2100_));
OAI21X1 OAI21X1_37 ( .A(_abc_40298_new_n804_), .B(_abc_40298_new_n826_), .C(_abc_40298_new_n655_), .Y(_abc_40298_new_n827_));
OAI21X1 OAI21X1_370 ( .A(pc_q_26_), .B(REGFILE_SIM_reg_bank_wr_i), .C(_abc_40298_new_n2100_), .Y(_abc_40298_new_n2101_));
OAI21X1 OAI21X1_371 ( .A(pc_q_27_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n2104_));
OAI21X1 OAI21X1_372 ( .A(pc_q_28_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n2107_));
OAI21X1 OAI21X1_373 ( .A(pc_q_29_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n2110_));
OAI21X1 OAI21X1_374 ( .A(pc_q_30_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n2113_));
OAI21X1 OAI21X1_375 ( .A(pc_q_31_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n2117_));
OAI21X1 OAI21X1_376 ( .A(_abc_40298_new_n923_), .B(_abc_40298_new_n925_), .C(_abc_40298_new_n2122_), .Y(_abc_40298_new_n2123_));
OAI21X1 OAI21X1_377 ( .A(_abc_40298_new_n949_), .B(_abc_40298_new_n2130_), .C(_abc_40298_new_n1013_), .Y(_0ex_rd_q_4_0__0_));
OAI21X1 OAI21X1_378 ( .A(_abc_40298_new_n623_), .B(_abc_40298_new_n2130_), .C(_abc_40298_new_n1013_), .Y(_0ex_rd_q_4_0__3_));
OAI21X1 OAI21X1_379 ( .A(_abc_40298_new_n646_), .B(_abc_40298_new_n929_), .C(_abc_40298_new_n982_), .Y(_abc_40298_new_n2140_));
OAI21X1 OAI21X1_38 ( .A(_abc_40298_new_n804_), .B(_abc_40298_new_n831_), .C(_abc_40298_new_n655_), .Y(_abc_40298_new_n832_));
OAI21X1 OAI21X1_380 ( .A(_abc_40298_new_n918_), .B(_abc_40298_new_n974_), .C(_abc_40298_new_n955_), .Y(_abc_40298_new_n2144_));
OAI21X1 OAI21X1_381 ( .A(_abc_40298_new_n921_), .B(_abc_40298_new_n976_), .C(_abc_40298_new_n897_), .Y(_abc_40298_new_n2148_));
OAI21X1 OAI21X1_382 ( .A(_abc_40298_new_n659_), .B(_abc_40298_new_n958_), .C(_abc_40298_new_n2141_), .Y(_abc_40298_new_n2159_));
OAI21X1 OAI21X1_383 ( .A(_abc_40298_new_n2165_), .B(_abc_40298_new_n2167_), .C(_abc_40298_new_n897_), .Y(_abc_40298_new_n2168_));
OAI21X1 OAI21X1_384 ( .A(_abc_40298_new_n906_), .B(_abc_40298_new_n2163_), .C(_abc_40298_new_n2171_), .Y(_abc_40298_new_n2172_));
OAI21X1 OAI21X1_385 ( .A(_abc_40298_new_n2174_), .B(_abc_40298_new_n906_), .C(_abc_40298_new_n2173_), .Y(_abc_40298_new_n2175_));
OAI21X1 OAI21X1_386 ( .A(_abc_40298_new_n1322_), .B(_abc_40298_new_n2176_), .C(_abc_40298_new_n2161_), .Y(alu_input_b_r_6_));
OAI21X1 OAI21X1_387 ( .A(_abc_40298_new_n1338_), .B(_abc_40298_new_n2176_), .C(_abc_40298_new_n2178_), .Y(alu_input_b_r_7_));
OAI21X1 OAI21X1_388 ( .A(_abc_40298_new_n1368_), .B(_abc_40298_new_n2176_), .C(_abc_40298_new_n2180_), .Y(alu_input_b_r_8_));
OAI21X1 OAI21X1_389 ( .A(_abc_40298_new_n1140_), .B(_abc_40298_new_n2176_), .C(_abc_40298_new_n2182_), .Y(alu_input_b_r_9_));
OAI21X1 OAI21X1_39 ( .A(_abc_40298_new_n804_), .B(_abc_40298_new_n836_), .C(_abc_40298_new_n655_), .Y(_abc_40298_new_n837_));
OAI21X1 OAI21X1_390 ( .A(_abc_40298_new_n1154_), .B(_abc_40298_new_n2176_), .C(_abc_40298_new_n2184_), .Y(alu_input_b_r_10_));
OAI21X1 OAI21X1_391 ( .A(_abc_40298_new_n1466_), .B(_abc_40298_new_n2176_), .C(_abc_40298_new_n2186_), .Y(alu_input_b_r_11_));
OAI21X1 OAI21X1_392 ( .A(_abc_40298_new_n1478_), .B(_abc_40298_new_n2176_), .C(_abc_40298_new_n2188_), .Y(alu_input_b_r_12_));
OAI21X1 OAI21X1_393 ( .A(_abc_40298_new_n2190_), .B(_abc_40298_new_n2176_), .C(_abc_40298_new_n2191_), .Y(alu_input_b_r_13_));
OAI21X1 OAI21X1_394 ( .A(_abc_40298_new_n2193_), .B(_abc_40298_new_n2176_), .C(_abc_40298_new_n2194_), .Y(alu_input_b_r_14_));
OAI21X1 OAI21X1_395 ( .A(_abc_40298_new_n2159_), .B(_abc_40298_new_n2198_), .C(_abc_40298_new_n2199_), .Y(_abc_40298_new_n2200_));
OAI21X1 OAI21X1_396 ( .A(_abc_40298_new_n2196_), .B(_abc_40298_new_n2176_), .C(_abc_40298_new_n2200_), .Y(alu_input_b_r_15_));
OAI21X1 OAI21X1_397 ( .A(_abc_40298_new_n2206_), .B(_abc_40298_new_n2197_), .C(_abc_40298_new_n2205_), .Y(_abc_40298_new_n2207_));
OAI21X1 OAI21X1_398 ( .A(_abc_40298_new_n2175_), .B(_abc_40298_new_n2172_), .C(REGFILE_SIM_reg_bank_reg_rb_o_16_), .Y(_abc_40298_new_n2209_));
OAI21X1 OAI21X1_399 ( .A(_abc_40298_new_n2202_), .B(_abc_40298_new_n2208_), .C(_abc_40298_new_n2209_), .Y(alu_input_b_r_16_));
OAI21X1 OAI21X1_4 ( .A(_abc_40298_new_n645_), .B(_abc_40298_new_n650_), .C(_abc_40298_new_n653_), .Y(_abc_40298_new_n654_));
OAI21X1 OAI21X1_40 ( .A(_abc_40298_new_n804_), .B(_abc_40298_new_n841_), .C(_abc_40298_new_n655_), .Y(_abc_40298_new_n842_));
OAI21X1 OAI21X1_400 ( .A(_abc_40298_new_n2211_), .B(_abc_40298_new_n2197_), .C(_abc_40298_new_n2205_), .Y(_abc_40298_new_n2212_));
OAI21X1 OAI21X1_401 ( .A(_abc_40298_new_n2175_), .B(_abc_40298_new_n2172_), .C(REGFILE_SIM_reg_bank_reg_rb_o_17_), .Y(_abc_40298_new_n2214_));
OAI21X1 OAI21X1_402 ( .A(_abc_40298_new_n2202_), .B(_abc_40298_new_n2213_), .C(_abc_40298_new_n2214_), .Y(alu_input_b_r_17_));
OAI21X1 OAI21X1_403 ( .A(_abc_40298_new_n2216_), .B(_abc_40298_new_n2197_), .C(_abc_40298_new_n2205_), .Y(_abc_40298_new_n2217_));
OAI21X1 OAI21X1_404 ( .A(_abc_40298_new_n2175_), .B(_abc_40298_new_n2172_), .C(REGFILE_SIM_reg_bank_reg_rb_o_18_), .Y(_abc_40298_new_n2219_));
OAI21X1 OAI21X1_405 ( .A(_abc_40298_new_n2202_), .B(_abc_40298_new_n2218_), .C(_abc_40298_new_n2219_), .Y(alu_input_b_r_18_));
OAI21X1 OAI21X1_406 ( .A(_abc_40298_new_n2221_), .B(_abc_40298_new_n2197_), .C(_abc_40298_new_n2205_), .Y(_abc_40298_new_n2222_));
OAI21X1 OAI21X1_407 ( .A(_abc_40298_new_n2175_), .B(_abc_40298_new_n2172_), .C(REGFILE_SIM_reg_bank_reg_rb_o_19_), .Y(_abc_40298_new_n2224_));
OAI21X1 OAI21X1_408 ( .A(_abc_40298_new_n2202_), .B(_abc_40298_new_n2223_), .C(_abc_40298_new_n2224_), .Y(alu_input_b_r_19_));
OAI21X1 OAI21X1_409 ( .A(_abc_40298_new_n2226_), .B(_abc_40298_new_n2197_), .C(_abc_40298_new_n2205_), .Y(_abc_40298_new_n2227_));
OAI21X1 OAI21X1_41 ( .A(_abc_40298_new_n804_), .B(_abc_40298_new_n846_), .C(_abc_40298_new_n655_), .Y(_abc_40298_new_n847_));
OAI21X1 OAI21X1_410 ( .A(_abc_40298_new_n2175_), .B(_abc_40298_new_n2172_), .C(REGFILE_SIM_reg_bank_reg_rb_o_20_), .Y(_abc_40298_new_n2229_));
OAI21X1 OAI21X1_411 ( .A(_abc_40298_new_n2202_), .B(_abc_40298_new_n2228_), .C(_abc_40298_new_n2229_), .Y(alu_input_b_r_20_));
OAI21X1 OAI21X1_412 ( .A(_abc_40298_new_n2231_), .B(_abc_40298_new_n2197_), .C(_abc_40298_new_n2205_), .Y(_abc_40298_new_n2232_));
OAI21X1 OAI21X1_413 ( .A(_abc_40298_new_n2175_), .B(_abc_40298_new_n2172_), .C(REGFILE_SIM_reg_bank_reg_rb_o_21_), .Y(_abc_40298_new_n2234_));
OAI21X1 OAI21X1_414 ( .A(_abc_40298_new_n2202_), .B(_abc_40298_new_n2233_), .C(_abc_40298_new_n2234_), .Y(alu_input_b_r_21_));
OAI21X1 OAI21X1_415 ( .A(_abc_40298_new_n2236_), .B(_abc_40298_new_n2197_), .C(_abc_40298_new_n2205_), .Y(_abc_40298_new_n2237_));
OAI21X1 OAI21X1_416 ( .A(_abc_40298_new_n2175_), .B(_abc_40298_new_n2172_), .C(REGFILE_SIM_reg_bank_reg_rb_o_22_), .Y(_abc_40298_new_n2239_));
OAI21X1 OAI21X1_417 ( .A(_abc_40298_new_n2202_), .B(_abc_40298_new_n2238_), .C(_abc_40298_new_n2239_), .Y(alu_input_b_r_22_));
OAI21X1 OAI21X1_418 ( .A(_abc_40298_new_n2241_), .B(_abc_40298_new_n2197_), .C(_abc_40298_new_n2205_), .Y(_abc_40298_new_n2242_));
OAI21X1 OAI21X1_419 ( .A(_abc_40298_new_n2175_), .B(_abc_40298_new_n2172_), .C(REGFILE_SIM_reg_bank_reg_rb_o_23_), .Y(_abc_40298_new_n2244_));
OAI21X1 OAI21X1_42 ( .A(_abc_40298_new_n804_), .B(_abc_40298_new_n851_), .C(_abc_40298_new_n655_), .Y(_abc_40298_new_n852_));
OAI21X1 OAI21X1_420 ( .A(_abc_40298_new_n2202_), .B(_abc_40298_new_n2243_), .C(_abc_40298_new_n2244_), .Y(alu_input_b_r_23_));
OAI21X1 OAI21X1_421 ( .A(_abc_40298_new_n2246_), .B(_abc_40298_new_n2197_), .C(_abc_40298_new_n2205_), .Y(_abc_40298_new_n2247_));
OAI21X1 OAI21X1_422 ( .A(_abc_40298_new_n2250_), .B(_abc_40298_new_n2197_), .C(_abc_40298_new_n2205_), .Y(_abc_40298_new_n2251_));
OAI21X1 OAI21X1_423 ( .A(_abc_40298_new_n2254_), .B(_abc_40298_new_n2197_), .C(_abc_40298_new_n2205_), .Y(_abc_40298_new_n2255_));
OAI21X1 OAI21X1_424 ( .A(_abc_40298_new_n2258_), .B(_abc_40298_new_n2197_), .C(_abc_40298_new_n2205_), .Y(_abc_40298_new_n2259_));
OAI21X1 OAI21X1_425 ( .A(_abc_40298_new_n2175_), .B(_abc_40298_new_n2172_), .C(REGFILE_SIM_reg_bank_reg_rb_o_27_), .Y(_abc_40298_new_n2261_));
OAI21X1 OAI21X1_426 ( .A(_abc_40298_new_n2202_), .B(_abc_40298_new_n2260_), .C(_abc_40298_new_n2261_), .Y(alu_input_b_r_27_));
OAI21X1 OAI21X1_427 ( .A(_abc_40298_new_n2263_), .B(_abc_40298_new_n2197_), .C(_abc_40298_new_n2205_), .Y(_abc_40298_new_n2264_));
OAI21X1 OAI21X1_428 ( .A(_abc_40298_new_n2175_), .B(_abc_40298_new_n2172_), .C(REGFILE_SIM_reg_bank_reg_rb_o_28_), .Y(_abc_40298_new_n2266_));
OAI21X1 OAI21X1_429 ( .A(_abc_40298_new_n2202_), .B(_abc_40298_new_n2265_), .C(_abc_40298_new_n2266_), .Y(alu_input_b_r_28_));
OAI21X1 OAI21X1_43 ( .A(_abc_40298_new_n804_), .B(_abc_40298_new_n856_), .C(_abc_40298_new_n655_), .Y(_abc_40298_new_n857_));
OAI21X1 OAI21X1_430 ( .A(_abc_40298_new_n2268_), .B(_abc_40298_new_n2197_), .C(_abc_40298_new_n2205_), .Y(_abc_40298_new_n2269_));
OAI21X1 OAI21X1_431 ( .A(_abc_40298_new_n2272_), .B(_abc_40298_new_n2197_), .C(_abc_40298_new_n2205_), .Y(_abc_40298_new_n2273_));
OAI21X1 OAI21X1_432 ( .A(_abc_40298_new_n2276_), .B(_abc_40298_new_n2197_), .C(_abc_40298_new_n2205_), .Y(_abc_40298_new_n2277_));
OAI21X1 OAI21X1_433 ( .A(_abc_40298_new_n918_), .B(_abc_40298_new_n974_), .C(_abc_40298_new_n955_), .Y(_abc_40298_new_n2282_));
OAI21X1 OAI21X1_434 ( .A(_abc_40298_new_n646_), .B(_abc_40298_new_n958_), .C(_abc_40298_new_n932_), .Y(_abc_40298_new_n2284_));
OAI21X1 OAI21X1_435 ( .A(_abc_40298_new_n2281_), .B(_abc_40298_new_n1013_), .C(_abc_40298_new_n2288_), .Y(_abc_40298_new_n2289_));
OAI21X1 OAI21X1_436 ( .A(_abc_40298_new_n2280_), .B(_abc_40298_new_n2120_), .C(_abc_40298_new_n2290_), .Y(alu_input_a_r_0_));
OAI21X1 OAI21X1_437 ( .A(_abc_40298_new_n2293_), .B(_abc_40298_new_n1013_), .C(_abc_40298_new_n2295_), .Y(_abc_40298_new_n2296_));
OAI21X1 OAI21X1_438 ( .A(_abc_40298_new_n2292_), .B(_abc_40298_new_n2120_), .C(_abc_40298_new_n2297_), .Y(alu_input_a_r_1_));
OAI21X1 OAI21X1_439 ( .A(_abc_40298_new_n1061_), .B(_abc_40298_new_n1069_), .C(_abc_40298_new_n2300_), .Y(_abc_40298_new_n2301_));
OAI21X1 OAI21X1_44 ( .A(_abc_40298_new_n804_), .B(_abc_40298_new_n861_), .C(_abc_40298_new_n655_), .Y(_abc_40298_new_n862_));
OAI21X1 OAI21X1_440 ( .A(_abc_40298_new_n2299_), .B(_abc_40298_new_n2302_), .C(_abc_40298_new_n1013_), .Y(_abc_40298_new_n2303_));
OAI21X1 OAI21X1_441 ( .A(_abc_40298_new_n1215_), .B(_abc_40298_new_n1013_), .C(_abc_40298_new_n982_), .Y(_abc_40298_new_n2305_));
OAI21X1 OAI21X1_442 ( .A(_abc_40298_new_n2307_), .B(_abc_40298_new_n2302_), .C(_abc_40298_new_n1002_), .Y(_abc_40298_new_n2308_));
OAI21X1 OAI21X1_443 ( .A(_abc_40298_new_n1229_), .B(_abc_40298_new_n1185_), .C(_abc_40298_new_n1001_), .Y(_abc_40298_new_n2309_));
OAI21X1 OAI21X1_444 ( .A(_abc_40298_new_n1013_), .B(_abc_40298_new_n1247_), .C(_abc_40298_new_n2310_), .Y(_abc_40298_new_n2311_));
OAI21X1 OAI21X1_445 ( .A(_abc_40298_new_n2307_), .B(_abc_40298_new_n2120_), .C(_abc_40298_new_n2312_), .Y(alu_input_a_r_3_));
OAI21X1 OAI21X1_446 ( .A(_abc_40298_new_n2314_), .B(_abc_40298_new_n2302_), .C(_abc_40298_new_n1002_), .Y(_abc_40298_new_n2315_));
OAI21X1 OAI21X1_447 ( .A(_abc_40298_new_n1252_), .B(_abc_40298_new_n1185_), .C(_abc_40298_new_n1001_), .Y(_abc_40298_new_n2316_));
OAI21X1 OAI21X1_448 ( .A(_abc_40298_new_n1013_), .B(_abc_40298_new_n1259_), .C(_abc_40298_new_n2317_), .Y(_abc_40298_new_n2318_));
OAI21X1 OAI21X1_449 ( .A(_abc_40298_new_n2314_), .B(_abc_40298_new_n2120_), .C(_abc_40298_new_n2319_), .Y(alu_input_a_r_4_));
OAI21X1 OAI21X1_45 ( .A(_abc_40298_new_n804_), .B(_abc_40298_new_n866_), .C(_abc_40298_new_n655_), .Y(_abc_40298_new_n867_));
OAI21X1 OAI21X1_450 ( .A(_abc_40298_new_n2321_), .B(_abc_40298_new_n2120_), .C(_abc_40298_new_n2325_), .Y(alu_input_a_r_5_));
OAI21X1 OAI21X1_451 ( .A(_abc_40298_new_n2327_), .B(_abc_40298_new_n2302_), .C(_abc_40298_new_n1002_), .Y(_abc_40298_new_n2328_));
OAI21X1 OAI21X1_452 ( .A(_abc_40298_new_n1309_), .B(_abc_40298_new_n1185_), .C(_abc_40298_new_n1001_), .Y(_abc_40298_new_n2329_));
OAI21X1 OAI21X1_453 ( .A(_abc_40298_new_n1013_), .B(_abc_40298_new_n1308_), .C(_abc_40298_new_n2330_), .Y(_abc_40298_new_n2331_));
OAI21X1 OAI21X1_454 ( .A(_abc_40298_new_n2327_), .B(_abc_40298_new_n2120_), .C(_abc_40298_new_n2332_), .Y(alu_input_a_r_6_));
OAI21X1 OAI21X1_455 ( .A(_abc_40298_new_n2334_), .B(_abc_40298_new_n2302_), .C(_abc_40298_new_n1002_), .Y(_abc_40298_new_n2336_));
OAI21X1 OAI21X1_456 ( .A(_abc_40298_new_n1339_), .B(_abc_40298_new_n1185_), .C(_abc_40298_new_n1001_), .Y(_abc_40298_new_n2337_));
OAI21X1 OAI21X1_457 ( .A(_abc_40298_new_n1013_), .B(_abc_40298_new_n2335_), .C(_abc_40298_new_n2338_), .Y(_abc_40298_new_n2339_));
OAI21X1 OAI21X1_458 ( .A(_abc_40298_new_n2334_), .B(_abc_40298_new_n2120_), .C(_abc_40298_new_n2340_), .Y(alu_input_a_r_7_));
OAI21X1 OAI21X1_459 ( .A(_abc_40298_new_n2342_), .B(_abc_40298_new_n2302_), .C(_abc_40298_new_n1002_), .Y(_abc_40298_new_n2343_));
OAI21X1 OAI21X1_46 ( .A(_abc_40298_new_n804_), .B(_abc_40298_new_n871_), .C(_abc_40298_new_n655_), .Y(_abc_40298_new_n872_));
OAI21X1 OAI21X1_460 ( .A(_abc_40298_new_n1369_), .B(_abc_40298_new_n1185_), .C(_abc_40298_new_n1001_), .Y(_abc_40298_new_n2344_));
OAI21X1 OAI21X1_461 ( .A(_abc_40298_new_n1013_), .B(_abc_40298_new_n1365_), .C(_abc_40298_new_n2345_), .Y(_abc_40298_new_n2346_));
OAI21X1 OAI21X1_462 ( .A(_abc_40298_new_n2342_), .B(_abc_40298_new_n2120_), .C(_abc_40298_new_n2347_), .Y(alu_input_a_r_8_));
OAI21X1 OAI21X1_463 ( .A(_abc_40298_new_n1395_), .B(_abc_40298_new_n1185_), .C(_abc_40298_new_n2349_), .Y(_abc_40298_new_n2350_));
OAI21X1 OAI21X1_464 ( .A(_abc_40298_new_n2352_), .B(_abc_40298_new_n2302_), .C(_abc_40298_new_n1002_), .Y(_abc_40298_new_n2353_));
OAI21X1 OAI21X1_465 ( .A(_abc_40298_new_n2350_), .B(_abc_40298_new_n2351_), .C(_abc_40298_new_n2353_), .Y(_abc_40298_new_n2354_));
OAI21X1 OAI21X1_466 ( .A(_abc_40298_new_n916_), .B(_abc_40298_new_n2119_), .C(REGFILE_SIM_reg_bank_reg_ra_o_9_), .Y(_abc_40298_new_n2356_));
OAI21X1 OAI21X1_467 ( .A(_abc_40298_new_n2358_), .B(_abc_40298_new_n2120_), .C(_abc_40298_new_n2362_), .Y(alu_input_a_r_10_));
OAI21X1 OAI21X1_468 ( .A(_abc_40298_new_n2364_), .B(_abc_40298_new_n2365_), .C(_abc_40298_new_n1013_), .Y(_abc_40298_new_n2366_));
OAI21X1 OAI21X1_469 ( .A(_abc_40298_new_n1013_), .B(_abc_40298_new_n1450_), .C(_abc_40298_new_n2366_), .Y(_abc_40298_new_n2367_));
OAI21X1 OAI21X1_47 ( .A(_abc_40298_new_n804_), .B(_abc_40298_new_n876_), .C(_abc_40298_new_n655_), .Y(_abc_40298_new_n877_));
OAI21X1 OAI21X1_470 ( .A(_abc_40298_new_n1038_), .B(_abc_40298_new_n2120_), .C(_abc_40298_new_n2367_), .Y(alu_input_a_r_11_));
OAI21X1 OAI21X1_471 ( .A(_abc_40298_new_n1034_), .B(_abc_40298_new_n2302_), .C(_abc_40298_new_n1002_), .Y(_abc_40298_new_n2369_));
OAI21X1 OAI21X1_472 ( .A(_abc_40298_new_n1479_), .B(_abc_40298_new_n1185_), .C(_abc_40298_new_n1001_), .Y(_abc_40298_new_n2370_));
OAI21X1 OAI21X1_473 ( .A(_abc_40298_new_n1034_), .B(_abc_40298_new_n2120_), .C(_abc_40298_new_n2371_), .Y(alu_input_a_r_12_));
OAI21X1 OAI21X1_474 ( .A(_abc_40298_new_n1039_), .B(_abc_40298_new_n2302_), .C(_abc_40298_new_n2373_), .Y(_abc_40298_new_n2374_));
OAI21X1 OAI21X1_475 ( .A(_abc_40298_new_n1039_), .B(_abc_40298_new_n2120_), .C(_abc_40298_new_n2375_), .Y(alu_input_a_r_13_));
OAI21X1 OAI21X1_476 ( .A(_abc_40298_new_n1036_), .B(_abc_40298_new_n2302_), .C(_abc_40298_new_n2377_), .Y(_abc_40298_new_n2378_));
OAI21X1 OAI21X1_477 ( .A(_abc_40298_new_n1036_), .B(_abc_40298_new_n2120_), .C(_abc_40298_new_n2379_), .Y(alu_input_a_r_14_));
OAI21X1 OAI21X1_478 ( .A(_abc_40298_new_n1035_), .B(_abc_40298_new_n2302_), .C(_abc_40298_new_n1002_), .Y(_abc_40298_new_n2381_));
OAI21X1 OAI21X1_479 ( .A(_abc_40298_new_n1569_), .B(_abc_40298_new_n1185_), .C(_abc_40298_new_n1001_), .Y(_abc_40298_new_n2382_));
OAI21X1 OAI21X1_48 ( .A(_abc_40298_new_n804_), .B(_abc_40298_new_n881_), .C(_abc_40298_new_n655_), .Y(_abc_40298_new_n882_));
OAI21X1 OAI21X1_480 ( .A(_abc_40298_new_n1035_), .B(_abc_40298_new_n2120_), .C(_abc_40298_new_n2383_), .Y(alu_input_a_r_15_));
OAI21X1 OAI21X1_481 ( .A(_abc_40298_new_n911_), .B(_abc_40298_new_n1014_), .C(_abc_40298_new_n2386_), .Y(_abc_40298_new_n2387_));
OAI21X1 OAI21X1_482 ( .A(_abc_40298_new_n2388_), .B(_abc_40298_new_n1185_), .C(_abc_40298_new_n1013_), .Y(_abc_40298_new_n2389_));
OAI21X1 OAI21X1_483 ( .A(_abc_40298_new_n2385_), .B(_abc_40298_new_n2120_), .C(_abc_40298_new_n2390_), .Y(alu_input_a_r_16_));
OAI21X1 OAI21X1_484 ( .A(_abc_40298_new_n909_), .B(_abc_40298_new_n1014_), .C(_abc_40298_new_n2393_), .Y(_abc_40298_new_n2394_));
OAI21X1 OAI21X1_485 ( .A(_abc_40298_new_n2395_), .B(_abc_40298_new_n1185_), .C(_abc_40298_new_n1013_), .Y(_abc_40298_new_n2396_));
OAI21X1 OAI21X1_486 ( .A(_abc_40298_new_n2392_), .B(_abc_40298_new_n2120_), .C(_abc_40298_new_n2397_), .Y(alu_input_a_r_17_));
OAI21X1 OAI21X1_487 ( .A(_abc_40298_new_n898_), .B(_abc_40298_new_n1014_), .C(_abc_40298_new_n2400_), .Y(_abc_40298_new_n2401_));
OAI21X1 OAI21X1_488 ( .A(_abc_40298_new_n2402_), .B(_abc_40298_new_n1185_), .C(_abc_40298_new_n1013_), .Y(_abc_40298_new_n2403_));
OAI21X1 OAI21X1_489 ( .A(_abc_40298_new_n2399_), .B(_abc_40298_new_n2120_), .C(_abc_40298_new_n2404_), .Y(alu_input_a_r_18_));
OAI21X1 OAI21X1_49 ( .A(_abc_40298_new_n630_), .B(_abc_40298_new_n631_), .C(_abc_40298_new_n634_), .Y(REGFILE_SIM_reg_bank_wr_i));
OAI21X1 OAI21X1_490 ( .A(_abc_40298_new_n903_), .B(_abc_40298_new_n1014_), .C(_abc_40298_new_n2407_), .Y(_abc_40298_new_n2408_));
OAI21X1 OAI21X1_491 ( .A(_abc_40298_new_n2409_), .B(_abc_40298_new_n1185_), .C(_abc_40298_new_n1013_), .Y(_abc_40298_new_n2410_));
OAI21X1 OAI21X1_492 ( .A(_abc_40298_new_n2406_), .B(_abc_40298_new_n2120_), .C(_abc_40298_new_n2411_), .Y(alu_input_a_r_19_));
OAI21X1 OAI21X1_493 ( .A(_abc_40298_new_n1315_), .B(_abc_40298_new_n1014_), .C(_abc_40298_new_n2414_), .Y(_abc_40298_new_n2415_));
OAI21X1 OAI21X1_494 ( .A(_abc_40298_new_n2416_), .B(_abc_40298_new_n1185_), .C(_abc_40298_new_n1013_), .Y(_abc_40298_new_n2417_));
OAI21X1 OAI21X1_495 ( .A(_abc_40298_new_n2413_), .B(_abc_40298_new_n2120_), .C(_abc_40298_new_n2418_), .Y(alu_input_a_r_20_));
OAI21X1 OAI21X1_496 ( .A(_abc_40298_new_n1341_), .B(_abc_40298_new_n1014_), .C(_abc_40298_new_n2421_), .Y(_abc_40298_new_n2422_));
OAI21X1 OAI21X1_497 ( .A(_abc_40298_new_n2423_), .B(_abc_40298_new_n1185_), .C(_abc_40298_new_n1013_), .Y(_abc_40298_new_n2424_));
OAI21X1 OAI21X1_498 ( .A(_abc_40298_new_n2420_), .B(_abc_40298_new_n2120_), .C(_abc_40298_new_n2425_), .Y(alu_input_a_r_21_));
OAI21X1 OAI21X1_499 ( .A(_abc_40298_new_n917_), .B(_abc_40298_new_n1014_), .C(_abc_40298_new_n2428_), .Y(_abc_40298_new_n2429_));
OAI21X1 OAI21X1_5 ( .A(mem_ack_i), .B(_abc_40298_new_n666_), .C(_abc_40298_new_n667_), .Y(_abc_27663_auto_fsm_map_cc_170_map_fsm_2376_2_));
OAI21X1 OAI21X1_50 ( .A(_abc_40298_new_n627_), .B(_abc_40298_new_n886_), .C(_abc_40298_new_n622_), .Y(_abc_40298_new_n887_));
OAI21X1 OAI21X1_500 ( .A(_abc_40298_new_n2430_), .B(_abc_40298_new_n1185_), .C(_abc_40298_new_n1013_), .Y(_abc_40298_new_n2431_));
OAI21X1 OAI21X1_501 ( .A(_abc_40298_new_n2427_), .B(_abc_40298_new_n2120_), .C(_abc_40298_new_n2432_), .Y(alu_input_a_r_22_));
OAI21X1 OAI21X1_502 ( .A(_abc_40298_new_n973_), .B(_abc_40298_new_n1014_), .C(_abc_40298_new_n2435_), .Y(_abc_40298_new_n2436_));
OAI21X1 OAI21X1_503 ( .A(_abc_40298_new_n2437_), .B(_abc_40298_new_n1185_), .C(_abc_40298_new_n1013_), .Y(_abc_40298_new_n2438_));
OAI21X1 OAI21X1_504 ( .A(_abc_40298_new_n2434_), .B(_abc_40298_new_n2120_), .C(_abc_40298_new_n2439_), .Y(alu_input_a_r_23_));
OAI21X1 OAI21X1_505 ( .A(_abc_40298_new_n1455_), .B(_abc_40298_new_n1014_), .C(_abc_40298_new_n2442_), .Y(_abc_40298_new_n2443_));
OAI21X1 OAI21X1_506 ( .A(_abc_40298_new_n2444_), .B(_abc_40298_new_n1185_), .C(_abc_40298_new_n1013_), .Y(_abc_40298_new_n2445_));
OAI21X1 OAI21X1_507 ( .A(_abc_40298_new_n2441_), .B(_abc_40298_new_n2120_), .C(_abc_40298_new_n2446_), .Y(alu_input_a_r_24_));
OAI21X1 OAI21X1_508 ( .A(_abc_40298_new_n1457_), .B(_abc_40298_new_n1014_), .C(_abc_40298_new_n2449_), .Y(_abc_40298_new_n2450_));
OAI21X1 OAI21X1_509 ( .A(_abc_40298_new_n2451_), .B(_abc_40298_new_n1185_), .C(_abc_40298_new_n1013_), .Y(_abc_40298_new_n2452_));
OAI21X1 OAI21X1_51 ( .A(_abc_40298_new_n908_), .B(_abc_40298_new_n910_), .C(_abc_40298_new_n913_), .Y(_abc_40298_new_n914_));
OAI21X1 OAI21X1_510 ( .A(_abc_40298_new_n2448_), .B(_abc_40298_new_n2120_), .C(_abc_40298_new_n2453_), .Y(alu_input_a_r_25_));
OAI21X1 OAI21X1_511 ( .A(_abc_40298_new_n2456_), .B(_abc_40298_new_n1014_), .C(_abc_40298_new_n2457_), .Y(_abc_40298_new_n2458_));
OAI21X1 OAI21X1_512 ( .A(_abc_40298_new_n2459_), .B(_abc_40298_new_n1185_), .C(_abc_40298_new_n1013_), .Y(_abc_40298_new_n2460_));
OAI21X1 OAI21X1_513 ( .A(_abc_40298_new_n2455_), .B(_abc_40298_new_n2120_), .C(_abc_40298_new_n2461_), .Y(alu_input_a_r_26_));
OAI21X1 OAI21X1_514 ( .A(_abc_40298_new_n1513_), .B(_abc_40298_new_n1014_), .C(_abc_40298_new_n2464_), .Y(_abc_40298_new_n2465_));
OAI21X1 OAI21X1_515 ( .A(_abc_40298_new_n2466_), .B(_abc_40298_new_n1185_), .C(_abc_40298_new_n1013_), .Y(_abc_40298_new_n2467_));
OAI21X1 OAI21X1_516 ( .A(_abc_40298_new_n2463_), .B(_abc_40298_new_n2120_), .C(_abc_40298_new_n2468_), .Y(alu_input_a_r_27_));
OAI21X1 OAI21X1_517 ( .A(_abc_40298_new_n2471_), .B(_abc_40298_new_n1014_), .C(_abc_40298_new_n2472_), .Y(_abc_40298_new_n2473_));
OAI21X1 OAI21X1_518 ( .A(_abc_40298_new_n2474_), .B(_abc_40298_new_n1185_), .C(_abc_40298_new_n1013_), .Y(_abc_40298_new_n2475_));
OAI21X1 OAI21X1_519 ( .A(_abc_40298_new_n2470_), .B(_abc_40298_new_n2120_), .C(_abc_40298_new_n2476_), .Y(alu_input_a_r_28_));
OAI21X1 OAI21X1_52 ( .A(_abc_40298_new_n905_), .B(_abc_40298_new_n914_), .C(_abc_40298_new_n907_), .Y(_abc_40298_new_n915_));
OAI21X1 OAI21X1_520 ( .A(_abc_40298_new_n2479_), .B(_abc_40298_new_n1014_), .C(_abc_40298_new_n2480_), .Y(_abc_40298_new_n2481_));
OAI21X1 OAI21X1_521 ( .A(_abc_40298_new_n2482_), .B(_abc_40298_new_n1185_), .C(_abc_40298_new_n1013_), .Y(_abc_40298_new_n2483_));
OAI21X1 OAI21X1_522 ( .A(_abc_40298_new_n2478_), .B(_abc_40298_new_n2120_), .C(_abc_40298_new_n2484_), .Y(alu_input_a_r_29_));
OAI21X1 OAI21X1_523 ( .A(_abc_40298_new_n1604_), .B(_abc_40298_new_n1014_), .C(_abc_40298_new_n2487_), .Y(_abc_40298_new_n2488_));
OAI21X1 OAI21X1_524 ( .A(_abc_40298_new_n2489_), .B(_abc_40298_new_n1185_), .C(_abc_40298_new_n1013_), .Y(_abc_40298_new_n2490_));
OAI21X1 OAI21X1_525 ( .A(_abc_40298_new_n2486_), .B(_abc_40298_new_n2120_), .C(_abc_40298_new_n2491_), .Y(alu_input_a_r_30_));
OAI21X1 OAI21X1_526 ( .A(_abc_40298_new_n1628_), .B(_abc_40298_new_n1014_), .C(_abc_40298_new_n2494_), .Y(_abc_40298_new_n2495_));
OAI21X1 OAI21X1_527 ( .A(_abc_40298_new_n2496_), .B(_abc_40298_new_n1185_), .C(_abc_40298_new_n1013_), .Y(_abc_40298_new_n2497_));
OAI21X1 OAI21X1_528 ( .A(_abc_40298_new_n2493_), .B(_abc_40298_new_n2120_), .C(_abc_40298_new_n2498_), .Y(alu_input_a_r_31_));
OAI21X1 OAI21X1_529 ( .A(_abc_40298_new_n914_), .B(_abc_40298_new_n926_), .C(_abc_40298_new_n907_), .Y(_abc_40298_new_n2502_));
OAI21X1 OAI21X1_53 ( .A(_abc_40298_new_n924_), .B(_abc_40298_new_n926_), .C(_abc_40298_new_n907_), .Y(_abc_40298_new_n927_));
OAI21X1 OAI21X1_530 ( .A(_abc_40298_new_n2515_), .B(_abc_40298_new_n2522_), .C(_abc_40298_new_n2571_), .Y(_abc_40298_new_n2572_));
OAI21X1 OAI21X1_531 ( .A(\mem_sel_o[0] ), .B(_abc_40298_new_n2570_), .C(_abc_40298_new_n2572_), .Y(_abc_40298_new_n2573_));
OAI21X1 OAI21X1_532 ( .A(_abc_40298_new_n2567_), .B(_abc_40298_new_n2516_), .C(_abc_40298_new_n2573_), .Y(_abc_40298_new_n2574_));
OAI21X1 OAI21X1_533 ( .A(_abc_40298_new_n2568_), .B(_abc_40298_new_n659_), .C(_abc_40298_new_n2574_), .Y(_abc_40298_new_n2575_));
OAI21X1 OAI21X1_534 ( .A(_abc_40298_new_n1046_), .B(_abc_40298_new_n2514_), .C(_abc_40298_new_n2521_), .Y(_abc_40298_new_n2585_));
OAI21X1 OAI21X1_535 ( .A(_abc_40298_new_n642_), .B(_abc_40298_new_n2587_), .C(_abc_40298_new_n2584_), .Y(_abc_40298_new_n2588_));
OAI21X1 OAI21X1_536 ( .A(_abc_40298_new_n2586_), .B(_abc_40298_new_n2589_), .C(_abc_40298_new_n2588_), .Y(_abc_40298_new_n2590_));
OAI21X1 OAI21X1_537 ( .A(_abc_40298_new_n2515_), .B(_abc_40298_new_n2521_), .C(_abc_40298_new_n2571_), .Y(_abc_40298_new_n2593_));
OAI21X1 OAI21X1_538 ( .A(\mem_sel_o[2] ), .B(_abc_40298_new_n2570_), .C(_abc_40298_new_n2593_), .Y(_abc_40298_new_n2594_));
OAI21X1 OAI21X1_539 ( .A(_abc_40298_new_n2592_), .B(_abc_40298_new_n2516_), .C(_abc_40298_new_n2594_), .Y(_abc_40298_new_n2595_));
OAI21X1 OAI21X1_54 ( .A(_abc_40298_new_n948_), .B(_abc_40298_new_n951_), .C(_abc_40298_new_n933_), .Y(_abc_40298_new_n952_));
OAI21X1 OAI21X1_540 ( .A(_abc_40298_new_n2568_), .B(_abc_40298_new_n659_), .C(_abc_40298_new_n2595_), .Y(_abc_40298_new_n2596_));
OAI21X1 OAI21X1_541 ( .A(_abc_40298_new_n1046_), .B(_abc_40298_new_n2514_), .C(_abc_40298_new_n2522_), .Y(_abc_40298_new_n2601_));
OAI21X1 OAI21X1_542 ( .A(_abc_40298_new_n642_), .B(_abc_40298_new_n2603_), .C(_abc_40298_new_n2600_), .Y(_abc_40298_new_n2604_));
OAI21X1 OAI21X1_543 ( .A(_abc_40298_new_n2589_), .B(_abc_40298_new_n2602_), .C(_abc_40298_new_n2604_), .Y(_abc_40298_new_n2605_));
OAI21X1 OAI21X1_544 ( .A(_abc_40298_new_n2139_), .B(_abc_40298_new_n2585_), .C(_abc_40298_new_n2609_), .Y(_abc_40298_new_n2610_));
OAI21X1 OAI21X1_545 ( .A(_abc_40298_new_n640_), .B(_abc_40298_new_n683_), .C(_abc_40298_new_n2607_), .Y(_abc_40298_new_n2613_));
OAI21X1 OAI21X1_546 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_0_), .B(_abc_40298_new_n2612_), .C(_abc_40298_new_n2613_), .Y(_abc_40298_new_n2614_));
OAI21X1 OAI21X1_547 ( .A(_abc_40298_new_n2153_), .B(_abc_40298_new_n2585_), .C(_abc_40298_new_n2619_), .Y(_abc_40298_new_n2620_));
OAI21X1 OAI21X1_548 ( .A(_abc_40298_new_n640_), .B(_abc_40298_new_n683_), .C(_abc_40298_new_n2618_), .Y(_abc_40298_new_n2621_));
OAI21X1 OAI21X1_549 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_1_), .B(_abc_40298_new_n2612_), .C(_abc_40298_new_n2621_), .Y(_abc_40298_new_n2622_));
OAI21X1 OAI21X1_55 ( .A(alu_op_r_4_), .B(_abc_40298_new_n956_), .C(_abc_40298_new_n960_), .Y(_abc_40298_new_n961_));
OAI21X1 OAI21X1_550 ( .A(_abc_40298_new_n1030_), .B(_abc_40298_new_n2585_), .C(_abc_40298_new_n2627_), .Y(_abc_40298_new_n2628_));
OAI21X1 OAI21X1_551 ( .A(_abc_40298_new_n640_), .B(_abc_40298_new_n683_), .C(_abc_40298_new_n2626_), .Y(_abc_40298_new_n2629_));
OAI21X1 OAI21X1_552 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_2_), .B(_abc_40298_new_n2612_), .C(_abc_40298_new_n2629_), .Y(_abc_40298_new_n2630_));
OAI21X1 OAI21X1_553 ( .A(_abc_40298_new_n1233_), .B(_abc_40298_new_n2585_), .C(_abc_40298_new_n2635_), .Y(_abc_40298_new_n2636_));
OAI21X1 OAI21X1_554 ( .A(_abc_40298_new_n640_), .B(_abc_40298_new_n683_), .C(_abc_40298_new_n2634_), .Y(_abc_40298_new_n2637_));
OAI21X1 OAI21X1_555 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_3_), .B(_abc_40298_new_n2612_), .C(_abc_40298_new_n2637_), .Y(_abc_40298_new_n2638_));
OAI21X1 OAI21X1_556 ( .A(_abc_40298_new_n1260_), .B(_abc_40298_new_n2585_), .C(_abc_40298_new_n2643_), .Y(_abc_40298_new_n2644_));
OAI21X1 OAI21X1_557 ( .A(_abc_40298_new_n640_), .B(_abc_40298_new_n683_), .C(_abc_40298_new_n2642_), .Y(_abc_40298_new_n2645_));
OAI21X1 OAI21X1_558 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_4_), .B(_abc_40298_new_n2612_), .C(_abc_40298_new_n2645_), .Y(_abc_40298_new_n2646_));
OAI21X1 OAI21X1_559 ( .A(_abc_40298_new_n1293_), .B(_abc_40298_new_n2585_), .C(_abc_40298_new_n2651_), .Y(_abc_40298_new_n2652_));
OAI21X1 OAI21X1_56 ( .A(_abc_40298_new_n931_), .B(_abc_40298_new_n930_), .C(_abc_40298_new_n968_), .Y(_abc_40298_new_n969_));
OAI21X1 OAI21X1_560 ( .A(_abc_40298_new_n640_), .B(_abc_40298_new_n683_), .C(_abc_40298_new_n2650_), .Y(_abc_40298_new_n2653_));
OAI21X1 OAI21X1_561 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_5_), .B(_abc_40298_new_n2612_), .C(_abc_40298_new_n2653_), .Y(_abc_40298_new_n2654_));
OAI21X1 OAI21X1_562 ( .A(_abc_40298_new_n1322_), .B(_abc_40298_new_n2585_), .C(_abc_40298_new_n2659_), .Y(_abc_40298_new_n2660_));
OAI21X1 OAI21X1_563 ( .A(_abc_40298_new_n640_), .B(_abc_40298_new_n683_), .C(_abc_40298_new_n2658_), .Y(_abc_40298_new_n2661_));
OAI21X1 OAI21X1_564 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_6_), .B(_abc_40298_new_n2612_), .C(_abc_40298_new_n2661_), .Y(_abc_40298_new_n2662_));
OAI21X1 OAI21X1_565 ( .A(_abc_40298_new_n1338_), .B(_abc_40298_new_n2585_), .C(_abc_40298_new_n2667_), .Y(_abc_40298_new_n2668_));
OAI21X1 OAI21X1_566 ( .A(_abc_40298_new_n640_), .B(_abc_40298_new_n683_), .C(_abc_40298_new_n2666_), .Y(_abc_40298_new_n2669_));
OAI21X1 OAI21X1_567 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_7_), .B(_abc_40298_new_n2612_), .C(_abc_40298_new_n2669_), .Y(_abc_40298_new_n2670_));
OAI21X1 OAI21X1_568 ( .A(inst_r_1_), .B(REGFILE_SIM_reg_bank_reg_rb_o_8_), .C(_abc_40298_new_n2570_), .Y(_abc_40298_new_n2675_));
OAI21X1 OAI21X1_569 ( .A(_abc_40298_new_n2674_), .B(_abc_40298_new_n2611_), .C(_abc_40298_new_n2675_), .Y(_abc_40298_new_n2676_));
OAI21X1 OAI21X1_57 ( .A(_abc_40298_new_n657_), .B(_abc_40298_new_n958_), .C(_abc_40298_new_n980_), .Y(_abc_40298_new_n981_));
OAI21X1 OAI21X1_570 ( .A(_abc_40298_new_n1368_), .B(_abc_40298_new_n2585_), .C(_abc_40298_new_n2677_), .Y(_abc_40298_new_n2678_));
OAI21X1 OAI21X1_571 ( .A(_abc_40298_new_n2139_), .B(_abc_40298_new_n2585_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2680_));
OAI21X1 OAI21X1_572 ( .A(inst_r_1_), .B(REGFILE_SIM_reg_bank_reg_rb_o_9_), .C(_abc_40298_new_n2570_), .Y(_abc_40298_new_n2684_));
OAI21X1 OAI21X1_573 ( .A(_abc_40298_new_n2683_), .B(_abc_40298_new_n2611_), .C(_abc_40298_new_n2684_), .Y(_abc_40298_new_n2685_));
OAI21X1 OAI21X1_574 ( .A(_abc_40298_new_n1140_), .B(_abc_40298_new_n2585_), .C(_abc_40298_new_n2686_), .Y(_abc_40298_new_n2687_));
OAI21X1 OAI21X1_575 ( .A(_abc_40298_new_n2153_), .B(_abc_40298_new_n2585_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2689_));
OAI21X1 OAI21X1_576 ( .A(inst_r_1_), .B(REGFILE_SIM_reg_bank_reg_rb_o_10_), .C(_abc_40298_new_n2570_), .Y(_abc_40298_new_n2693_));
OAI21X1 OAI21X1_577 ( .A(_abc_40298_new_n2692_), .B(_abc_40298_new_n2611_), .C(_abc_40298_new_n2693_), .Y(_abc_40298_new_n2694_));
OAI21X1 OAI21X1_578 ( .A(_abc_40298_new_n1154_), .B(_abc_40298_new_n2585_), .C(_abc_40298_new_n2695_), .Y(_abc_40298_new_n2696_));
OAI21X1 OAI21X1_579 ( .A(_abc_40298_new_n1030_), .B(_abc_40298_new_n2585_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2698_));
OAI21X1 OAI21X1_58 ( .A(_abc_40298_new_n657_), .B(_abc_40298_new_n983_), .C(_abc_40298_new_n887_), .Y(_abc_40298_new_n984_));
OAI21X1 OAI21X1_580 ( .A(inst_r_1_), .B(REGFILE_SIM_reg_bank_reg_rb_o_11_), .C(_abc_40298_new_n2570_), .Y(_abc_40298_new_n2702_));
OAI21X1 OAI21X1_581 ( .A(_abc_40298_new_n2701_), .B(_abc_40298_new_n2611_), .C(_abc_40298_new_n2702_), .Y(_abc_40298_new_n2703_));
OAI21X1 OAI21X1_582 ( .A(_abc_40298_new_n1466_), .B(_abc_40298_new_n2585_), .C(_abc_40298_new_n2704_), .Y(_abc_40298_new_n2705_));
OAI21X1 OAI21X1_583 ( .A(_abc_40298_new_n1233_), .B(_abc_40298_new_n2585_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2707_));
OAI21X1 OAI21X1_584 ( .A(inst_r_1_), .B(REGFILE_SIM_reg_bank_reg_rb_o_12_), .C(_abc_40298_new_n2570_), .Y(_abc_40298_new_n2711_));
OAI21X1 OAI21X1_585 ( .A(_abc_40298_new_n2710_), .B(_abc_40298_new_n2611_), .C(_abc_40298_new_n2711_), .Y(_abc_40298_new_n2712_));
OAI21X1 OAI21X1_586 ( .A(_abc_40298_new_n1478_), .B(_abc_40298_new_n2585_), .C(_abc_40298_new_n2713_), .Y(_abc_40298_new_n2714_));
OAI21X1 OAI21X1_587 ( .A(_abc_40298_new_n1260_), .B(_abc_40298_new_n2585_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2716_));
OAI21X1 OAI21X1_588 ( .A(inst_r_1_), .B(REGFILE_SIM_reg_bank_reg_rb_o_13_), .C(_abc_40298_new_n2570_), .Y(_abc_40298_new_n2720_));
OAI21X1 OAI21X1_589 ( .A(_abc_40298_new_n2719_), .B(_abc_40298_new_n2611_), .C(_abc_40298_new_n2720_), .Y(_abc_40298_new_n2721_));
OAI21X1 OAI21X1_59 ( .A(_abc_40298_new_n987_), .B(_abc_40298_new_n969_), .C(_abc_40298_new_n988_), .Y(_abc_40298_new_n989_));
OAI21X1 OAI21X1_590 ( .A(_abc_40298_new_n2190_), .B(_abc_40298_new_n2585_), .C(_abc_40298_new_n2722_), .Y(_abc_40298_new_n2723_));
OAI21X1 OAI21X1_591 ( .A(_abc_40298_new_n1293_), .B(_abc_40298_new_n2585_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2725_));
OAI21X1 OAI21X1_592 ( .A(inst_r_1_), .B(REGFILE_SIM_reg_bank_reg_rb_o_14_), .C(_abc_40298_new_n2570_), .Y(_abc_40298_new_n2729_));
OAI21X1 OAI21X1_593 ( .A(_abc_40298_new_n2728_), .B(_abc_40298_new_n2611_), .C(_abc_40298_new_n2729_), .Y(_abc_40298_new_n2730_));
OAI21X1 OAI21X1_594 ( .A(_abc_40298_new_n2193_), .B(_abc_40298_new_n2585_), .C(_abc_40298_new_n2731_), .Y(_abc_40298_new_n2732_));
OAI21X1 OAI21X1_595 ( .A(_abc_40298_new_n1322_), .B(_abc_40298_new_n2585_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2734_));
OAI21X1 OAI21X1_596 ( .A(inst_r_1_), .B(REGFILE_SIM_reg_bank_reg_rb_o_15_), .C(_abc_40298_new_n2570_), .Y(_abc_40298_new_n2738_));
OAI21X1 OAI21X1_597 ( .A(_abc_40298_new_n2737_), .B(_abc_40298_new_n2611_), .C(_abc_40298_new_n2738_), .Y(_abc_40298_new_n2739_));
OAI21X1 OAI21X1_598 ( .A(_abc_40298_new_n2196_), .B(_abc_40298_new_n2585_), .C(_abc_40298_new_n2740_), .Y(_abc_40298_new_n2741_));
OAI21X1 OAI21X1_599 ( .A(_abc_40298_new_n1338_), .B(_abc_40298_new_n2585_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2743_));
OAI21X1 OAI21X1_6 ( .A(_abc_40298_new_n643_), .B(_abc_40298_new_n662_), .C(state_q_5_), .Y(_abc_40298_new_n669_));
OAI21X1 OAI21X1_60 ( .A(inst_r_1_), .B(_abc_40298_new_n1003_), .C(_abc_40298_new_n1002_), .Y(_abc_40298_new_n1004_));
OAI21X1 OAI21X1_600 ( .A(_abc_40298_new_n2139_), .B(_abc_40298_new_n2601_), .C(_abc_40298_new_n2747_), .Y(_abc_40298_new_n2748_));
OAI21X1 OAI21X1_601 ( .A(_abc_40298_new_n640_), .B(_abc_40298_new_n683_), .C(_abc_40298_new_n2746_), .Y(_abc_40298_new_n2749_));
OAI21X1 OAI21X1_602 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_16_), .B(_abc_40298_new_n2612_), .C(_abc_40298_new_n2749_), .Y(_abc_40298_new_n2750_));
OAI21X1 OAI21X1_603 ( .A(_abc_40298_new_n2153_), .B(_abc_40298_new_n2601_), .C(_abc_40298_new_n2755_), .Y(_abc_40298_new_n2756_));
OAI21X1 OAI21X1_604 ( .A(_abc_40298_new_n640_), .B(_abc_40298_new_n683_), .C(_abc_40298_new_n2754_), .Y(_abc_40298_new_n2757_));
OAI21X1 OAI21X1_605 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_17_), .B(_abc_40298_new_n2612_), .C(_abc_40298_new_n2757_), .Y(_abc_40298_new_n2758_));
OAI21X1 OAI21X1_606 ( .A(_abc_40298_new_n1030_), .B(_abc_40298_new_n2601_), .C(_abc_40298_new_n2763_), .Y(_abc_40298_new_n2764_));
OAI21X1 OAI21X1_607 ( .A(_abc_40298_new_n640_), .B(_abc_40298_new_n683_), .C(_abc_40298_new_n2762_), .Y(_abc_40298_new_n2765_));
OAI21X1 OAI21X1_608 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_18_), .B(_abc_40298_new_n2612_), .C(_abc_40298_new_n2765_), .Y(_abc_40298_new_n2766_));
OAI21X1 OAI21X1_609 ( .A(_abc_40298_new_n1233_), .B(_abc_40298_new_n2601_), .C(_abc_40298_new_n2771_), .Y(_abc_40298_new_n2772_));
OAI21X1 OAI21X1_61 ( .A(_abc_40298_new_n618_), .B(_abc_40298_new_n1009_), .C(_abc_40298_new_n1011_), .Y(_abc_40298_new_n1012_));
OAI21X1 OAI21X1_610 ( .A(_abc_40298_new_n640_), .B(_abc_40298_new_n683_), .C(_abc_40298_new_n2770_), .Y(_abc_40298_new_n2773_));
OAI21X1 OAI21X1_611 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_19_), .B(_abc_40298_new_n2612_), .C(_abc_40298_new_n2773_), .Y(_abc_40298_new_n2774_));
OAI21X1 OAI21X1_612 ( .A(_abc_40298_new_n1260_), .B(_abc_40298_new_n2601_), .C(_abc_40298_new_n2779_), .Y(_abc_40298_new_n2780_));
OAI21X1 OAI21X1_613 ( .A(_abc_40298_new_n640_), .B(_abc_40298_new_n683_), .C(_abc_40298_new_n2778_), .Y(_abc_40298_new_n2781_));
OAI21X1 OAI21X1_614 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_20_), .B(_abc_40298_new_n2612_), .C(_abc_40298_new_n2781_), .Y(_abc_40298_new_n2782_));
OAI21X1 OAI21X1_615 ( .A(_abc_40298_new_n1293_), .B(_abc_40298_new_n2601_), .C(_abc_40298_new_n2787_), .Y(_abc_40298_new_n2788_));
OAI21X1 OAI21X1_616 ( .A(_abc_40298_new_n640_), .B(_abc_40298_new_n683_), .C(_abc_40298_new_n2786_), .Y(_abc_40298_new_n2789_));
OAI21X1 OAI21X1_617 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_21_), .B(_abc_40298_new_n2612_), .C(_abc_40298_new_n2789_), .Y(_abc_40298_new_n2790_));
OAI21X1 OAI21X1_618 ( .A(_abc_40298_new_n1322_), .B(_abc_40298_new_n2601_), .C(_abc_40298_new_n2795_), .Y(_abc_40298_new_n2796_));
OAI21X1 OAI21X1_619 ( .A(_abc_40298_new_n640_), .B(_abc_40298_new_n683_), .C(_abc_40298_new_n2794_), .Y(_abc_40298_new_n2797_));
OAI21X1 OAI21X1_62 ( .A(_abc_40298_new_n1043_), .B(_abc_40298_new_n1059_), .C(sr_q_2_), .Y(_abc_40298_new_n1062_));
OAI21X1 OAI21X1_620 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_22_), .B(_abc_40298_new_n2612_), .C(_abc_40298_new_n2797_), .Y(_abc_40298_new_n2798_));
OAI21X1 OAI21X1_621 ( .A(_abc_40298_new_n1338_), .B(_abc_40298_new_n2601_), .C(_abc_40298_new_n2803_), .Y(_abc_40298_new_n2804_));
OAI21X1 OAI21X1_622 ( .A(_abc_40298_new_n640_), .B(_abc_40298_new_n683_), .C(_abc_40298_new_n2802_), .Y(_abc_40298_new_n2805_));
OAI21X1 OAI21X1_623 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_23_), .B(_abc_40298_new_n2612_), .C(_abc_40298_new_n2805_), .Y(_abc_40298_new_n2806_));
OAI21X1 OAI21X1_624 ( .A(inst_r_1_), .B(REGFILE_SIM_reg_bank_reg_rb_o_24_), .C(_abc_40298_new_n2570_), .Y(_abc_40298_new_n2811_));
OAI21X1 OAI21X1_625 ( .A(_abc_40298_new_n2810_), .B(_abc_40298_new_n2611_), .C(_abc_40298_new_n2811_), .Y(_abc_40298_new_n2812_));
OAI21X1 OAI21X1_626 ( .A(_abc_40298_new_n1368_), .B(_abc_40298_new_n2601_), .C(_abc_40298_new_n2813_), .Y(_abc_40298_new_n2814_));
OAI21X1 OAI21X1_627 ( .A(_abc_40298_new_n2139_), .B(_abc_40298_new_n2601_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2816_));
OAI21X1 OAI21X1_628 ( .A(inst_r_1_), .B(REGFILE_SIM_reg_bank_reg_rb_o_25_), .C(_abc_40298_new_n2570_), .Y(_abc_40298_new_n2820_));
OAI21X1 OAI21X1_629 ( .A(_abc_40298_new_n2819_), .B(_abc_40298_new_n2611_), .C(_abc_40298_new_n2820_), .Y(_abc_40298_new_n2821_));
OAI21X1 OAI21X1_63 ( .A(_abc_40298_new_n1030_), .B(_abc_40298_new_n1061_), .C(_abc_40298_new_n1062_), .Y(_abc_40298_new_n1063_));
OAI21X1 OAI21X1_630 ( .A(_abc_40298_new_n1140_), .B(_abc_40298_new_n2601_), .C(_abc_40298_new_n2822_), .Y(_abc_40298_new_n2823_));
OAI21X1 OAI21X1_631 ( .A(_abc_40298_new_n2153_), .B(_abc_40298_new_n2601_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2825_));
OAI21X1 OAI21X1_632 ( .A(inst_r_1_), .B(REGFILE_SIM_reg_bank_reg_rb_o_26_), .C(_abc_40298_new_n2570_), .Y(_abc_40298_new_n2829_));
OAI21X1 OAI21X1_633 ( .A(_abc_40298_new_n2828_), .B(_abc_40298_new_n2611_), .C(_abc_40298_new_n2829_), .Y(_abc_40298_new_n2830_));
OAI21X1 OAI21X1_634 ( .A(_abc_40298_new_n1154_), .B(_abc_40298_new_n2601_), .C(_abc_40298_new_n2831_), .Y(_abc_40298_new_n2832_));
OAI21X1 OAI21X1_635 ( .A(_abc_40298_new_n1030_), .B(_abc_40298_new_n2601_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2834_));
OAI21X1 OAI21X1_636 ( .A(inst_r_1_), .B(REGFILE_SIM_reg_bank_reg_rb_o_27_), .C(_abc_40298_new_n2570_), .Y(_abc_40298_new_n2838_));
OAI21X1 OAI21X1_637 ( .A(_abc_40298_new_n2837_), .B(_abc_40298_new_n2611_), .C(_abc_40298_new_n2838_), .Y(_abc_40298_new_n2839_));
OAI21X1 OAI21X1_638 ( .A(_abc_40298_new_n1466_), .B(_abc_40298_new_n2601_), .C(_abc_40298_new_n2840_), .Y(_abc_40298_new_n2841_));
OAI21X1 OAI21X1_639 ( .A(_abc_40298_new_n1233_), .B(_abc_40298_new_n2601_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2843_));
OAI21X1 OAI21X1_64 ( .A(_abc_40298_new_n1064_), .B(_abc_40298_new_n1066_), .C(_abc_40298_new_n1067_), .Y(_abc_40298_new_n1068_));
OAI21X1 OAI21X1_640 ( .A(inst_r_1_), .B(REGFILE_SIM_reg_bank_reg_rb_o_28_), .C(_abc_40298_new_n2570_), .Y(_abc_40298_new_n2847_));
OAI21X1 OAI21X1_641 ( .A(_abc_40298_new_n2846_), .B(_abc_40298_new_n2611_), .C(_abc_40298_new_n2847_), .Y(_abc_40298_new_n2848_));
OAI21X1 OAI21X1_642 ( .A(_abc_40298_new_n1478_), .B(_abc_40298_new_n2601_), .C(_abc_40298_new_n2849_), .Y(_abc_40298_new_n2850_));
OAI21X1 OAI21X1_643 ( .A(_abc_40298_new_n1260_), .B(_abc_40298_new_n2601_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2852_));
OAI21X1 OAI21X1_644 ( .A(inst_r_1_), .B(REGFILE_SIM_reg_bank_reg_rb_o_29_), .C(_abc_40298_new_n2570_), .Y(_abc_40298_new_n2856_));
OAI21X1 OAI21X1_645 ( .A(_abc_40298_new_n2855_), .B(_abc_40298_new_n2611_), .C(_abc_40298_new_n2856_), .Y(_abc_40298_new_n2857_));
OAI21X1 OAI21X1_646 ( .A(_abc_40298_new_n2190_), .B(_abc_40298_new_n2601_), .C(_abc_40298_new_n2858_), .Y(_abc_40298_new_n2859_));
OAI21X1 OAI21X1_647 ( .A(_abc_40298_new_n1293_), .B(_abc_40298_new_n2601_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2861_));
OAI21X1 OAI21X1_648 ( .A(inst_r_1_), .B(REGFILE_SIM_reg_bank_reg_rb_o_30_), .C(_abc_40298_new_n2570_), .Y(_abc_40298_new_n2865_));
OAI21X1 OAI21X1_649 ( .A(_abc_40298_new_n2864_), .B(_abc_40298_new_n2611_), .C(_abc_40298_new_n2865_), .Y(_abc_40298_new_n2866_));
OAI21X1 OAI21X1_65 ( .A(_abc_40298_new_n992_), .B(_abc_40298_new_n1063_), .C(_abc_40298_new_n1068_), .Y(_abc_40298_new_n1069_));
OAI21X1 OAI21X1_650 ( .A(_abc_40298_new_n2193_), .B(_abc_40298_new_n2601_), .C(_abc_40298_new_n2867_), .Y(_abc_40298_new_n2868_));
OAI21X1 OAI21X1_651 ( .A(_abc_40298_new_n1322_), .B(_abc_40298_new_n2601_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2870_));
OAI21X1 OAI21X1_652 ( .A(inst_r_1_), .B(REGFILE_SIM_reg_bank_reg_rb_o_31_), .C(_abc_40298_new_n2570_), .Y(_abc_40298_new_n2874_));
OAI21X1 OAI21X1_653 ( .A(_abc_40298_new_n2873_), .B(_abc_40298_new_n2611_), .C(_abc_40298_new_n2874_), .Y(_abc_40298_new_n2875_));
OAI21X1 OAI21X1_654 ( .A(_abc_40298_new_n2196_), .B(_abc_40298_new_n2601_), .C(_abc_40298_new_n2876_), .Y(_abc_40298_new_n2877_));
OAI21X1 OAI21X1_655 ( .A(_abc_40298_new_n1338_), .B(_abc_40298_new_n2601_), .C(_abc_40298_new_n2578_), .Y(_abc_40298_new_n2879_));
OAI21X1 OAI21X1_656 ( .A(_abc_40298_new_n2568_), .B(_abc_40298_new_n657_), .C(_abc_40298_new_n2589_), .Y(_abc_40298_new_n2885_));
OAI21X1 OAI21X1_657 ( .A(mem_we_o), .B(_abc_40298_new_n2885_), .C(_abc_40298_new_n2576_), .Y(_abc_40298_new_n2886_));
OAI21X1 OAI21X1_658 ( .A(_abc_40298_new_n2882_), .B(_abc_40298_new_n2884_), .C(_abc_40298_new_n2886_), .Y(_0mem_we_o_0_0_));
OAI21X1 OAI21X1_659 ( .A(_abc_40298_new_n662_), .B(_abc_40298_new_n2885_), .C(state_q_5_), .Y(_abc_40298_new_n2888_));
OAI21X1 OAI21X1_66 ( .A(_abc_40298_new_n1070_), .B(_abc_40298_new_n1071_), .C(_abc_40298_new_n1069_), .Y(_abc_40298_new_n1072_));
OAI21X1 OAI21X1_660 ( .A(state_q_1_), .B(state_q_2_), .C(_abc_40298_new_n2891_), .Y(_abc_40298_new_n2892_));
OAI21X1 OAI21X1_661 ( .A(_abc_40298_new_n635_), .B(_abc_40298_new_n664_), .C(_abc_40298_new_n2884_), .Y(_abc_40298_new_n2895_));
OAI21X1 OAI21X1_662 ( .A(_abc_40298_new_n667_), .B(_abc_40298_new_n2281_), .C(_abc_40298_new_n2896_), .Y(_0mem_addr_o_31_0__0_));
OAI21X1 OAI21X1_663 ( .A(_abc_40298_new_n667_), .B(_abc_40298_new_n2293_), .C(_abc_40298_new_n2898_), .Y(_0mem_addr_o_31_0__1_));
OAI21X1 OAI21X1_664 ( .A(_abc_40298_new_n2513_), .B(_abc_40298_new_n1050_), .C(_abc_40298_new_n2518_), .Y(_abc_40298_new_n2903_));
OAI21X1 OAI21X1_665 ( .A(_abc_40298_new_n1055_), .B(_abc_40298_new_n2912_), .C(_abc_40298_new_n2911_), .Y(_abc_40298_new_n2913_));
OAI21X1 OAI21X1_666 ( .A(_abc_40298_new_n2904_), .B(_abc_40298_new_n2907_), .C(_abc_40298_new_n2914_), .Y(_abc_40298_new_n2915_));
OAI21X1 OAI21X1_667 ( .A(\mem_addr_o[3] ), .B(_abc_40298_new_n664_), .C(state_q_5_), .Y(_abc_40298_new_n2917_));
OAI21X1 OAI21X1_668 ( .A(_abc_40298_new_n2916_), .B(_abc_40298_new_n2917_), .C(_abc_40298_new_n2918_), .Y(_0mem_addr_o_31_0__3_));
OAI21X1 OAI21X1_669 ( .A(_abc_40298_new_n1055_), .B(_abc_40298_new_n2911_), .C(_abc_40298_new_n2922_), .Y(_abc_40298_new_n2923_));
OAI21X1 OAI21X1_67 ( .A(_abc_40298_new_n992_), .B(_abc_40298_new_n1080_), .C(_abc_40298_new_n1064_), .Y(_abc_40298_new_n1083_));
OAI21X1 OAI21X1_670 ( .A(_abc_40298_new_n669_), .B(_abc_40298_new_n2924_), .C(_abc_40298_new_n2925_), .Y(_0mem_addr_o_31_0__4_));
OAI21X1 OAI21X1_671 ( .A(_abc_40298_new_n2314_), .B(_abc_40298_new_n1315_), .C(_abc_40298_new_n2927_), .Y(_abc_40298_new_n2928_));
OAI21X1 OAI21X1_672 ( .A(\mem_addr_o[5] ), .B(_abc_40298_new_n664_), .C(state_q_5_), .Y(_abc_40298_new_n2937_));
OAI21X1 OAI21X1_673 ( .A(_abc_40298_new_n2937_), .B(_abc_40298_new_n2936_), .C(_abc_40298_new_n2938_), .Y(_0mem_addr_o_31_0__5_));
OAI21X1 OAI21X1_674 ( .A(_abc_40298_new_n1053_), .B(_abc_40298_new_n2941_), .C(_abc_40298_new_n2940_), .Y(_abc_40298_new_n2942_));
OAI21X1 OAI21X1_675 ( .A(_abc_40298_new_n2929_), .B(_abc_40298_new_n2934_), .C(_abc_40298_new_n2943_), .Y(_abc_40298_new_n2944_));
OAI21X1 OAI21X1_676 ( .A(_abc_40298_new_n669_), .B(_abc_40298_new_n2945_), .C(_abc_40298_new_n2946_), .Y(_0mem_addr_o_31_0__6_));
OAI21X1 OAI21X1_677 ( .A(_abc_40298_new_n2327_), .B(_abc_40298_new_n917_), .C(_abc_40298_new_n2944_), .Y(_abc_40298_new_n2950_));
OAI21X1 OAI21X1_678 ( .A(_abc_40298_new_n2941_), .B(_abc_40298_new_n2951_), .C(_abc_40298_new_n2949_), .Y(_abc_40298_new_n2952_));
OAI21X1 OAI21X1_679 ( .A(_abc_40298_new_n2949_), .B(_abc_40298_new_n2950_), .C(_abc_40298_new_n2953_), .Y(_abc_40298_new_n2954_));
OAI21X1 OAI21X1_68 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_2_), .B(_abc_40298_new_n1082_), .C(_abc_40298_new_n1083_), .Y(_abc_40298_new_n1084_));
OAI21X1 OAI21X1_680 ( .A(_abc_40298_new_n2958_), .B(_abc_40298_new_n2940_), .C(_abc_40298_new_n2959_), .Y(_abc_40298_new_n2960_));
OAI21X1 OAI21X1_681 ( .A(_abc_40298_new_n2963_), .B(_abc_40298_new_n2965_), .C(_abc_40298_new_n2966_), .Y(_0mem_addr_o_31_0__8_));
OAI21X1 OAI21X1_682 ( .A(_abc_40298_new_n2342_), .B(_abc_40298_new_n1455_), .C(_abc_40298_new_n2964_), .Y(_abc_40298_new_n2968_));
OAI21X1 OAI21X1_683 ( .A(\mem_addr_o[9] ), .B(_abc_40298_new_n664_), .C(state_q_5_), .Y(_abc_40298_new_n2973_));
OAI21X1 OAI21X1_684 ( .A(_abc_40298_new_n2973_), .B(_abc_40298_new_n2972_), .C(_abc_40298_new_n2974_), .Y(_0mem_addr_o_31_0__9_));
OAI21X1 OAI21X1_685 ( .A(\mem_addr_o[10] ), .B(_abc_40298_new_n664_), .C(state_q_5_), .Y(_abc_40298_new_n2983_));
OAI21X1 OAI21X1_686 ( .A(_abc_40298_new_n2983_), .B(_abc_40298_new_n2982_), .C(_abc_40298_new_n2984_), .Y(_0mem_addr_o_31_0__10_));
OAI21X1 OAI21X1_687 ( .A(_abc_40298_new_n2358_), .B(_abc_40298_new_n2456_), .C(_abc_40298_new_n2980_), .Y(_abc_40298_new_n2986_));
OAI21X1 OAI21X1_688 ( .A(_abc_40298_new_n625_), .B(_abc_40298_new_n2568_), .C(_abc_40298_new_n1513_), .Y(_abc_40298_new_n2987_));
OAI21X1 OAI21X1_689 ( .A(opcode_q_21_), .B(_abc_40298_new_n642_), .C(_abc_40298_new_n2987_), .Y(_abc_40298_new_n2988_));
OAI21X1 OAI21X1_69 ( .A(_abc_40298_new_n1073_), .B(_abc_40298_new_n1069_), .C(_abc_40298_new_n1084_), .Y(_abc_40298_new_n1085_));
OAI21X1 OAI21X1_690 ( .A(_abc_40298_new_n2989_), .B(_abc_40298_new_n2986_), .C(_abc_40298_new_n2902_), .Y(_abc_40298_new_n2991_));
OAI21X1 OAI21X1_691 ( .A(_abc_40298_new_n2990_), .B(_abc_40298_new_n2991_), .C(_abc_40298_new_n2992_), .Y(_0mem_addr_o_31_0__11_));
OAI21X1 OAI21X1_692 ( .A(_abc_40298_new_n2997_), .B(_abc_40298_new_n2995_), .C(_abc_40298_new_n2999_), .Y(_abc_40298_new_n3000_));
OAI21X1 OAI21X1_693 ( .A(_abc_40298_new_n625_), .B(_abc_40298_new_n2568_), .C(REGFILE_SIM_reg_bank_rb_i_1_), .Y(_abc_40298_new_n3002_));
OAI21X1 OAI21X1_694 ( .A(_abc_40298_new_n944_), .B(_abc_40298_new_n642_), .C(_abc_40298_new_n3002_), .Y(_abc_40298_new_n3003_));
OAI21X1 OAI21X1_695 ( .A(_abc_40298_new_n669_), .B(_abc_40298_new_n3007_), .C(_abc_40298_new_n3008_), .Y(_0mem_addr_o_31_0__12_));
OAI21X1 OAI21X1_696 ( .A(_abc_40298_new_n625_), .B(_abc_40298_new_n2568_), .C(_abc_40298_new_n2479_), .Y(_abc_40298_new_n3011_));
OAI21X1 OAI21X1_697 ( .A(opcode_q_23_), .B(_abc_40298_new_n642_), .C(_abc_40298_new_n3011_), .Y(_abc_40298_new_n3012_));
OAI21X1 OAI21X1_698 ( .A(_abc_40298_new_n3004_), .B(_abc_40298_new_n3001_), .C(_abc_40298_new_n3010_), .Y(_abc_40298_new_n3017_));
OAI21X1 OAI21X1_699 ( .A(_abc_40298_new_n1039_), .B(_abc_40298_new_n3012_), .C(_abc_40298_new_n3018_), .Y(_abc_40298_new_n3023_));
OAI21X1 OAI21X1_7 ( .A(mem_ack_i), .B(_abc_40298_new_n631_), .C(_abc_40298_new_n669_), .Y(_abc_27663_auto_fsm_map_cc_170_map_fsm_2376_1_));
OAI21X1 OAI21X1_70 ( .A(_abc_40298_new_n1085_), .B(_abc_40298_new_n1029_), .C(_abc_40298_new_n1072_), .Y(_abc_40298_new_n1086_));
OAI21X1 OAI21X1_700 ( .A(_abc_40298_new_n625_), .B(_abc_40298_new_n2568_), .C(REGFILE_SIM_reg_bank_rb_i_3_), .Y(_abc_40298_new_n3024_));
OAI21X1 OAI21X1_701 ( .A(_abc_40298_new_n623_), .B(_abc_40298_new_n642_), .C(_abc_40298_new_n3024_), .Y(_abc_40298_new_n3025_));
OAI21X1 OAI21X1_702 ( .A(\mem_addr_o[14] ), .B(_abc_40298_new_n664_), .C(state_q_5_), .Y(_abc_40298_new_n3029_));
OAI21X1 OAI21X1_703 ( .A(_abc_40298_new_n3029_), .B(_abc_40298_new_n3028_), .C(_abc_40298_new_n3030_), .Y(_0mem_addr_o_31_0__14_));
OAI21X1 OAI21X1_704 ( .A(_abc_40298_new_n3026_), .B(_abc_40298_new_n3032_), .C(_abc_40298_new_n3033_), .Y(_abc_40298_new_n3034_));
OAI21X1 OAI21X1_705 ( .A(_abc_40298_new_n625_), .B(_abc_40298_new_n2568_), .C(REGFILE_SIM_reg_bank_rb_i_4_), .Y(_abc_40298_new_n3035_));
OAI21X1 OAI21X1_706 ( .A(_abc_40298_new_n624_), .B(_abc_40298_new_n642_), .C(_abc_40298_new_n3035_), .Y(_abc_40298_new_n3036_));
OAI21X1 OAI21X1_707 ( .A(_abc_40298_new_n625_), .B(_abc_40298_new_n2568_), .C(_abc_40298_new_n1628_), .Y(_abc_40298_new_n3038_));
OAI21X1 OAI21X1_708 ( .A(opcode_q_25_), .B(_abc_40298_new_n642_), .C(_abc_40298_new_n3038_), .Y(_abc_40298_new_n3039_));
OAI21X1 OAI21X1_709 ( .A(_abc_40298_new_n669_), .B(_abc_40298_new_n3042_), .C(_abc_40298_new_n3043_), .Y(_0mem_addr_o_31_0__15_));
OAI21X1 OAI21X1_71 ( .A(esr_q_2_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n1087_));
OAI21X1 OAI21X1_710 ( .A(_abc_40298_new_n3010_), .B(_abc_40298_new_n3015_), .C(_abc_40298_new_n3013_), .Y(_abc_40298_new_n3045_));
OAI21X1 OAI21X1_711 ( .A(_abc_40298_new_n3033_), .B(_abc_40298_new_n3041_), .C(_abc_40298_new_n3037_), .Y(_abc_40298_new_n3047_));
OAI21X1 OAI21X1_712 ( .A(_abc_40298_new_n3050_), .B(_abc_40298_new_n3001_), .C(_abc_40298_new_n3048_), .Y(_abc_40298_new_n3051_));
OAI21X1 OAI21X1_713 ( .A(_abc_40298_new_n3054_), .B(_abc_40298_new_n3057_), .C(_abc_40298_new_n2902_), .Y(_abc_40298_new_n3058_));
OAI21X1 OAI21X1_714 ( .A(_abc_40298_new_n3056_), .B(_abc_40298_new_n3058_), .C(_abc_40298_new_n3059_), .Y(_0mem_addr_o_31_0__16_));
OAI21X1 OAI21X1_715 ( .A(_abc_40298_new_n3054_), .B(_abc_40298_new_n3057_), .C(_abc_40298_new_n3052_), .Y(_abc_40298_new_n3061_));
OAI21X1 OAI21X1_716 ( .A(_abc_40298_new_n669_), .B(_abc_40298_new_n3063_), .C(_abc_40298_new_n3064_), .Y(_0mem_addr_o_31_0__17_));
OAI21X1 OAI21X1_717 ( .A(_abc_40298_new_n2392_), .B(_abc_40298_new_n3039_), .C(_abc_40298_new_n3052_), .Y(_abc_40298_new_n3067_));
OAI21X1 OAI21X1_718 ( .A(_abc_40298_new_n669_), .B(_abc_40298_new_n3072_), .C(_abc_40298_new_n3073_), .Y(_0mem_addr_o_31_0__18_));
OAI21X1 OAI21X1_719 ( .A(_abc_40298_new_n2399_), .B(_abc_40298_new_n3039_), .C(_abc_40298_new_n3071_), .Y(_abc_40298_new_n3075_));
OAI21X1 OAI21X1_72 ( .A(_abc_40298_new_n931_), .B(_abc_40298_new_n930_), .C(_abc_40298_new_n950_), .Y(_abc_40298_new_n1090_));
OAI21X1 OAI21X1_720 ( .A(_abc_40298_new_n3076_), .B(_abc_40298_new_n3075_), .C(_abc_40298_new_n664_), .Y(_abc_40298_new_n3077_));
OAI21X1 OAI21X1_721 ( .A(\mem_addr_o[19] ), .B(_abc_40298_new_n664_), .C(state_q_5_), .Y(_abc_40298_new_n3079_));
OAI21X1 OAI21X1_722 ( .A(_abc_40298_new_n3079_), .B(_abc_40298_new_n3078_), .C(_abc_40298_new_n3080_), .Y(_0mem_addr_o_31_0__19_));
OAI21X1 OAI21X1_723 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_18_), .B(REGFILE_SIM_reg_bank_reg_ra_o_19_), .C(_abc_40298_new_n3036_), .Y(_abc_40298_new_n3086_));
OAI21X1 OAI21X1_724 ( .A(_abc_40298_new_n3092_), .B(_abc_40298_new_n3089_), .C(_abc_40298_new_n2902_), .Y(_abc_40298_new_n3094_));
OAI21X1 OAI21X1_725 ( .A(_abc_40298_new_n3093_), .B(_abc_40298_new_n3094_), .C(_abc_40298_new_n3095_), .Y(_0mem_addr_o_31_0__20_));
OAI21X1 OAI21X1_726 ( .A(_abc_40298_new_n3092_), .B(_abc_40298_new_n3089_), .C(_abc_40298_new_n3090_), .Y(_abc_40298_new_n3097_));
OAI21X1 OAI21X1_727 ( .A(_abc_40298_new_n3098_), .B(_abc_40298_new_n3097_), .C(_abc_40298_new_n664_), .Y(_abc_40298_new_n3099_));
OAI21X1 OAI21X1_728 ( .A(\mem_addr_o[21] ), .B(_abc_40298_new_n664_), .C(state_q_5_), .Y(_abc_40298_new_n3101_));
OAI21X1 OAI21X1_729 ( .A(_abc_40298_new_n3101_), .B(_abc_40298_new_n3100_), .C(_abc_40298_new_n3102_), .Y(_0mem_addr_o_31_0__21_));
OAI21X1 OAI21X1_73 ( .A(_abc_40298_new_n987_), .B(_abc_40298_new_n969_), .C(_abc_40298_new_n1093_), .Y(_abc_40298_new_n1094_));
OAI21X1 OAI21X1_730 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_20_), .B(REGFILE_SIM_reg_bank_reg_ra_o_21_), .C(_abc_40298_new_n3036_), .Y(_abc_40298_new_n3105_));
OAI21X1 OAI21X1_731 ( .A(_abc_40298_new_n3107_), .B(_abc_40298_new_n3089_), .C(_abc_40298_new_n3105_), .Y(_abc_40298_new_n3108_));
OAI21X1 OAI21X1_732 ( .A(_abc_40298_new_n3109_), .B(_abc_40298_new_n3111_), .C(_abc_40298_new_n3112_), .Y(_0mem_addr_o_31_0__22_));
OAI21X1 OAI21X1_733 ( .A(_abc_40298_new_n2427_), .B(_abc_40298_new_n3039_), .C(_abc_40298_new_n3110_), .Y(_abc_40298_new_n3118_));
OAI21X1 OAI21X1_734 ( .A(_abc_40298_new_n3115_), .B(_abc_40298_new_n3118_), .C(_abc_40298_new_n2902_), .Y(_abc_40298_new_n3119_));
OAI21X1 OAI21X1_735 ( .A(_abc_40298_new_n3117_), .B(_abc_40298_new_n3119_), .C(_abc_40298_new_n3120_), .Y(_0mem_addr_o_31_0__23_));
OAI21X1 OAI21X1_736 ( .A(_abc_40298_new_n3105_), .B(_abc_40298_new_n3122_), .C(_abc_40298_new_n3114_), .Y(_abc_40298_new_n3123_));
OAI21X1 OAI21X1_737 ( .A(_abc_40298_new_n3125_), .B(_abc_40298_new_n3087_), .C(_abc_40298_new_n3124_), .Y(_abc_40298_new_n3126_));
OAI21X1 OAI21X1_738 ( .A(_abc_40298_new_n3130_), .B(_abc_40298_new_n3128_), .C(_abc_40298_new_n2902_), .Y(_abc_40298_new_n3132_));
OAI21X1 OAI21X1_739 ( .A(_abc_40298_new_n3131_), .B(_abc_40298_new_n3132_), .C(_abc_40298_new_n3133_), .Y(_0mem_addr_o_31_0__24_));
OAI21X1 OAI21X1_74 ( .A(_abc_40298_new_n1098_), .B(_abc_40298_new_n942_), .C(_abc_40298_new_n971_), .Y(_abc_40298_new_n1099_));
OAI21X1 OAI21X1_740 ( .A(_abc_40298_new_n3130_), .B(_abc_40298_new_n3128_), .C(_abc_40298_new_n3135_), .Y(_abc_40298_new_n3136_));
OAI21X1 OAI21X1_741 ( .A(_abc_40298_new_n3138_), .B(_abc_40298_new_n3136_), .C(_abc_40298_new_n664_), .Y(_abc_40298_new_n3140_));
OAI21X1 OAI21X1_742 ( .A(\mem_addr_o[25] ), .B(_abc_40298_new_n664_), .C(state_q_5_), .Y(_abc_40298_new_n3142_));
OAI21X1 OAI21X1_743 ( .A(_abc_40298_new_n3142_), .B(_abc_40298_new_n3141_), .C(_abc_40298_new_n3143_), .Y(_0mem_addr_o_31_0__25_));
OAI21X1 OAI21X1_744 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_24_), .B(REGFILE_SIM_reg_bank_reg_ra_o_25_), .C(_abc_40298_new_n3036_), .Y(_abc_40298_new_n3147_));
OAI21X1 OAI21X1_745 ( .A(_abc_40298_new_n3146_), .B(_abc_40298_new_n3128_), .C(_abc_40298_new_n3147_), .Y(_abc_40298_new_n3148_));
OAI21X1 OAI21X1_746 ( .A(_abc_40298_new_n3148_), .B(_abc_40298_new_n3149_), .C(_abc_40298_new_n3150_), .Y(_abc_40298_new_n3151_));
OAI21X1 OAI21X1_747 ( .A(_abc_40298_new_n2455_), .B(_abc_40298_new_n3039_), .C(_abc_40298_new_n3155_), .Y(_abc_40298_new_n3156_));
OAI21X1 OAI21X1_748 ( .A(_abc_40298_new_n669_), .B(_abc_40298_new_n3158_), .C(_abc_40298_new_n3159_), .Y(_0mem_addr_o_31_0__27_));
OAI21X1 OAI21X1_749 ( .A(_abc_40298_new_n3162_), .B(_abc_40298_new_n3128_), .C(_abc_40298_new_n3164_), .Y(_abc_40298_new_n3165_));
OAI21X1 OAI21X1_75 ( .A(alu_equal_o), .B(alu_less_than_signed_o), .C(_abc_40298_new_n1091_), .Y(_abc_40298_new_n1104_));
OAI21X1 OAI21X1_750 ( .A(_abc_40298_new_n3167_), .B(_abc_40298_new_n3169_), .C(_abc_40298_new_n3170_), .Y(_0mem_addr_o_31_0__28_));
OAI21X1 OAI21X1_751 ( .A(_abc_40298_new_n2470_), .B(_abc_40298_new_n3039_), .C(_abc_40298_new_n3168_), .Y(_abc_40298_new_n3172_));
OAI21X1 OAI21X1_752 ( .A(_abc_40298_new_n669_), .B(_abc_40298_new_n3174_), .C(_abc_40298_new_n3175_), .Y(_0mem_addr_o_31_0__29_));
OAI21X1 OAI21X1_753 ( .A(\mem_addr_o[30] ), .B(_abc_40298_new_n664_), .C(state_q_5_), .Y(_abc_40298_new_n3187_));
OAI21X1 OAI21X1_754 ( .A(_abc_40298_new_n3187_), .B(_abc_40298_new_n3186_), .C(_abc_40298_new_n3188_), .Y(_0mem_addr_o_31_0__30_));
OAI21X1 OAI21X1_755 ( .A(_abc_40298_new_n3179_), .B(_abc_40298_new_n3183_), .C(_abc_40298_new_n3177_), .Y(_abc_40298_new_n3190_));
OAI21X1 OAI21X1_756 ( .A(_abc_40298_new_n3191_), .B(_abc_40298_new_n3190_), .C(_abc_40298_new_n664_), .Y(_abc_40298_new_n3192_));
OAI21X1 OAI21X1_757 ( .A(\mem_addr_o[31] ), .B(_abc_40298_new_n664_), .C(state_q_5_), .Y(_abc_40298_new_n3194_));
OAI21X1 OAI21X1_758 ( .A(_abc_40298_new_n3194_), .B(_abc_40298_new_n3193_), .C(_abc_40298_new_n3195_), .Y(_0mem_addr_o_31_0__31_));
OAI21X1 OAI21X1_759 ( .A(nmi_q), .B(nmi_i), .C(enable_i), .Y(_abc_40298_new_n3198_));
OAI21X1 OAI21X1_76 ( .A(_abc_40298_new_n930_), .B(_abc_40298_new_n931_), .C(_abc_40298_new_n948_), .Y(_abc_40298_new_n1106_));
OAI21X1 OAI21X1_760 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2269_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4180_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4185_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4186_));
OAI21X1 OAI21X1_761 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3264_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4211_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4210_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4212_));
OAI21X1 OAI21X1_762 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2274_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4180_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4256_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4257_));
OAI21X1 OAI21X1_763 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3267_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4211_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4265_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4266_));
OAI21X1 OAI21X1_764 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2276_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4180_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4288_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4289_));
OAI21X1 OAI21X1_765 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3269_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4211_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4297_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4298_));
OAI21X1 OAI21X1_766 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2278_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4180_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4320_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4321_));
OAI21X1 OAI21X1_767 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3271_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4211_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4329_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4330_));
OAI21X1 OAI21X1_768 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2280_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4180_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4352_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4353_));
OAI21X1 OAI21X1_769 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3273_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4211_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4361_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4362_));
OAI21X1 OAI21X1_77 ( .A(_abc_40298_new_n1105_), .B(_abc_40298_new_n1103_), .C(_abc_40298_new_n1109_), .Y(_abc_40298_new_n1110_));
OAI21X1 OAI21X1_770 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2282_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4180_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4384_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4385_));
OAI21X1 OAI21X1_771 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3275_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4211_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4393_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4394_));
OAI21X1 OAI21X1_772 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2284_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4180_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4416_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4417_));
OAI21X1 OAI21X1_773 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3277_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4211_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4425_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4426_));
OAI21X1 OAI21X1_774 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2286_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4180_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4448_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4449_));
OAI21X1 OAI21X1_775 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3279_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4211_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4457_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4458_));
OAI21X1 OAI21X1_776 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2288_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4180_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4480_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4481_));
OAI21X1 OAI21X1_777 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3281_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4211_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4489_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4490_));
OAI21X1 OAI21X1_778 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2290_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4180_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4512_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4513_));
OAI21X1 OAI21X1_779 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3283_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4211_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4521_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4522_));
OAI21X1 OAI21X1_78 ( .A(_abc_40298_new_n930_), .B(_abc_40298_new_n931_), .C(_abc_40298_new_n1008_), .Y(_abc_40298_new_n1112_));
OAI21X1 OAI21X1_780 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2292_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4180_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4544_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4545_));
OAI21X1 OAI21X1_781 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3285_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4211_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4553_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4554_));
OAI21X1 OAI21X1_782 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2294_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4180_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4576_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4577_));
OAI21X1 OAI21X1_783 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3287_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4211_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4585_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4586_));
OAI21X1 OAI21X1_784 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2296_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4180_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4608_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4609_));
OAI21X1 OAI21X1_785 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3289_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4211_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4617_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4618_));
OAI21X1 OAI21X1_786 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2298_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4180_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4640_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4641_));
OAI21X1 OAI21X1_787 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3291_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4211_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4649_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4650_));
OAI21X1 OAI21X1_788 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2300_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4180_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4672_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4673_));
OAI21X1 OAI21X1_789 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3293_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4211_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4681_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4682_));
OAI21X1 OAI21X1_79 ( .A(_abc_40298_new_n1115_), .B(_abc_40298_new_n1113_), .C(_abc_40298_new_n1112_), .Y(_abc_40298_new_n1116_));
OAI21X1 OAI21X1_790 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2302_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4180_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4704_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4705_));
OAI21X1 OAI21X1_791 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3295_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4211_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4713_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4714_));
OAI21X1 OAI21X1_792 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2304_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4180_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4736_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4737_));
OAI21X1 OAI21X1_793 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3297_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4211_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4745_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4746_));
OAI21X1 OAI21X1_794 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2306_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4180_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4768_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4769_));
OAI21X1 OAI21X1_795 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3299_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4211_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4777_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4778_));
OAI21X1 OAI21X1_796 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2308_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4180_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4800_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4801_));
OAI21X1 OAI21X1_797 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3301_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4211_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4809_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4810_));
OAI21X1 OAI21X1_798 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2310_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4180_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4832_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4833_));
OAI21X1 OAI21X1_799 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3303_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4211_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4841_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4842_));
OAI21X1 OAI21X1_8 ( .A(_abc_40298_new_n683_), .B(_abc_40298_new_n645_), .C(_abc_40298_new_n685_), .Y(_abc_40298_new_n686_));
OAI21X1 OAI21X1_80 ( .A(_abc_40298_new_n1119_), .B(_abc_40298_new_n1117_), .C(alu_flag_update_o), .Y(_abc_40298_new_n1120_));
OAI21X1 OAI21X1_800 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2312_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4180_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4864_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4865_));
OAI21X1 OAI21X1_801 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3305_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4211_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4873_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4874_));
OAI21X1 OAI21X1_802 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2314_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4180_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4896_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4897_));
OAI21X1 OAI21X1_803 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3307_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4211_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4905_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4906_));
OAI21X1 OAI21X1_804 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2316_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4180_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4928_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4929_));
OAI21X1 OAI21X1_805 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3309_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4211_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4937_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4938_));
OAI21X1 OAI21X1_806 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2318_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4180_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4960_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4961_));
OAI21X1 OAI21X1_807 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3311_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4211_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4969_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4970_));
OAI21X1 OAI21X1_808 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2320_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4180_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4992_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4993_));
OAI21X1 OAI21X1_809 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3313_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4211_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5001_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5002_));
OAI21X1 OAI21X1_81 ( .A(_abc_40298_new_n1089_), .B(alu_flag_update_o), .C(_abc_40298_new_n1120_), .Y(_abc_40298_new_n1121_));
OAI21X1 OAI21X1_810 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2322_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4180_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5024_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5025_));
OAI21X1 OAI21X1_811 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3315_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4211_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5033_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5034_));
OAI21X1 OAI21X1_812 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2324_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4180_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5056_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5057_));
OAI21X1 OAI21X1_813 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3317_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4211_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5065_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5066_));
OAI21X1 OAI21X1_814 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2326_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4180_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5088_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5089_));
OAI21X1 OAI21X1_815 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3319_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4211_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5097_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5098_));
OAI21X1 OAI21X1_816 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2328_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4180_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5120_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5121_));
OAI21X1 OAI21X1_817 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3321_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4211_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5129_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5130_));
OAI21X1 OAI21X1_818 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2330_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4180_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5152_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5153_));
OAI21X1 OAI21X1_819 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3323_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4211_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5161_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5162_));
OAI21X1 OAI21X1_82 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_9_), .B(_abc_40298_new_n1061_), .C(_abc_40298_new_n993_), .Y(_abc_40298_new_n1122_));
OAI21X1 OAI21X1_820 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2332_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4180_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5184_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5185_));
OAI21X1 OAI21X1_821 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3325_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4211_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5193_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5194_));
OAI21X1 OAI21X1_822 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2334_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4180_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5216_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5217_));
OAI21X1 OAI21X1_823 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3327_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4211_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5225_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5226_));
OAI21X1 OAI21X1_824 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2269_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5252_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5257_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5258_));
OAI21X1 OAI21X1_825 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3264_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5283_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5282_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5284_));
OAI21X1 OAI21X1_826 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2274_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5252_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5328_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5329_));
OAI21X1 OAI21X1_827 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3267_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5283_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5337_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5338_));
OAI21X1 OAI21X1_828 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2276_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5252_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5360_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5361_));
OAI21X1 OAI21X1_829 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3269_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5283_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5369_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5370_));
OAI21X1 OAI21X1_83 ( .A(_abc_40298_new_n1060_), .B(_abc_40298_new_n1121_), .C(_abc_40298_new_n1123_), .Y(_abc_40298_new_n1124_));
OAI21X1 OAI21X1_830 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2278_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5252_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5392_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5393_));
OAI21X1 OAI21X1_831 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3271_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5283_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5401_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5402_));
OAI21X1 OAI21X1_832 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2280_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5252_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5424_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5425_));
OAI21X1 OAI21X1_833 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3273_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5283_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5433_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5434_));
OAI21X1 OAI21X1_834 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2282_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5252_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5456_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5457_));
OAI21X1 OAI21X1_835 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3275_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5283_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5465_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5466_));
OAI21X1 OAI21X1_836 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2284_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5252_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5488_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5489_));
OAI21X1 OAI21X1_837 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3277_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5283_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5497_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5498_));
OAI21X1 OAI21X1_838 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2286_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5252_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5520_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5521_));
OAI21X1 OAI21X1_839 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3279_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5283_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5529_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5530_));
OAI21X1 OAI21X1_84 ( .A(_abc_40298_new_n1119_), .B(_abc_40298_new_n1117_), .C(_abc_40298_new_n933_), .Y(_abc_40298_new_n1128_));
OAI21X1 OAI21X1_840 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2288_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5252_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5552_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5553_));
OAI21X1 OAI21X1_841 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3281_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5283_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5561_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5562_));
OAI21X1 OAI21X1_842 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2290_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5252_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5584_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5585_));
OAI21X1 OAI21X1_843 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3283_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5283_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5593_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5594_));
OAI21X1 OAI21X1_844 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2292_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5252_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5616_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5617_));
OAI21X1 OAI21X1_845 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3285_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5283_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5625_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5626_));
OAI21X1 OAI21X1_846 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2294_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5252_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5648_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5649_));
OAI21X1 OAI21X1_847 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3287_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5283_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5657_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5658_));
OAI21X1 OAI21X1_848 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2296_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5252_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5680_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5681_));
OAI21X1 OAI21X1_849 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3289_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5283_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5689_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5690_));
OAI21X1 OAI21X1_85 ( .A(_abc_40298_new_n983_), .B(_abc_40298_new_n657_), .C(_abc_40298_new_n1128_), .Y(_abc_40298_new_n1129_));
OAI21X1 OAI21X1_850 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2298_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5252_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5712_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5713_));
OAI21X1 OAI21X1_851 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3291_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5283_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5721_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5722_));
OAI21X1 OAI21X1_852 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2300_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5252_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5744_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5745_));
OAI21X1 OAI21X1_853 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3293_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5283_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5753_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5754_));
OAI21X1 OAI21X1_854 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2302_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5252_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5776_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5777_));
OAI21X1 OAI21X1_855 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3295_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5283_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5785_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5786_));
OAI21X1 OAI21X1_856 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2304_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5252_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5808_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5809_));
OAI21X1 OAI21X1_857 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3297_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5283_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5817_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5818_));
OAI21X1 OAI21X1_858 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2306_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5252_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5840_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5841_));
OAI21X1 OAI21X1_859 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3299_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5283_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5849_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5850_));
OAI21X1 OAI21X1_86 ( .A(esr_q_9_), .B(_abc_40298_new_n1066_), .C(_abc_40298_new_n992_), .Y(_abc_40298_new_n1130_));
OAI21X1 OAI21X1_860 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2308_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5252_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5872_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5873_));
OAI21X1 OAI21X1_861 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3301_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5283_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5881_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5882_));
OAI21X1 OAI21X1_862 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2310_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5252_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5904_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5905_));
OAI21X1 OAI21X1_863 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3303_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5283_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5913_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5914_));
OAI21X1 OAI21X1_864 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2312_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5252_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5936_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5937_));
OAI21X1 OAI21X1_865 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3305_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5283_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5945_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5946_));
OAI21X1 OAI21X1_866 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2314_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5252_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5968_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5969_));
OAI21X1 OAI21X1_867 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3307_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5283_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n5977_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5978_));
OAI21X1 OAI21X1_868 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2316_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5252_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n6000_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6001_));
OAI21X1 OAI21X1_869 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3309_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5283_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n6009_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6010_));
OAI21X1 OAI21X1_87 ( .A(_abc_40298_new_n1129_), .B(_abc_40298_new_n1127_), .C(_abc_40298_new_n1131_), .Y(_abc_40298_new_n1132_));
OAI21X1 OAI21X1_870 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2318_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5252_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n6032_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6033_));
OAI21X1 OAI21X1_871 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3311_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5283_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n6041_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6042_));
OAI21X1 OAI21X1_872 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2320_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5252_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n6064_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6065_));
OAI21X1 OAI21X1_873 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3313_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5283_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n6073_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6074_));
OAI21X1 OAI21X1_874 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2322_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5252_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n6096_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6097_));
OAI21X1 OAI21X1_875 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3315_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5283_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n6105_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6106_));
OAI21X1 OAI21X1_876 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2324_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5252_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n6128_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6129_));
OAI21X1 OAI21X1_877 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3317_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5283_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n6137_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6138_));
OAI21X1 OAI21X1_878 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2326_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5252_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n6160_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6161_));
OAI21X1 OAI21X1_879 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3319_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5283_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n6169_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6170_));
OAI21X1 OAI21X1_88 ( .A(_abc_40298_new_n1073_), .B(_abc_40298_new_n1069_), .C(_abc_40298_new_n885_), .Y(_abc_40298_new_n1134_));
OAI21X1 OAI21X1_880 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2328_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5252_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n6192_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6193_));
OAI21X1 OAI21X1_881 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3321_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5283_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n6201_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6202_));
OAI21X1 OAI21X1_882 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2330_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5252_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n6224_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6225_));
OAI21X1 OAI21X1_883 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3323_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5283_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n6233_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6234_));
OAI21X1 OAI21X1_884 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2332_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5252_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n6256_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6257_));
OAI21X1 OAI21X1_885 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3325_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5283_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n6265_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6266_));
OAI21X1 OAI21X1_886 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2334_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5252_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n6288_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6289_));
OAI21X1 OAI21X1_887 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3327_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5283_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n6297_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6298_));
OAI21X1 OAI21X1_888 ( .A(alu__abc_38674_new_n118_), .B(alu__abc_38674_new_n119_), .C(alu__abc_38674_new_n115_), .Y(alu__abc_38674_new_n120_));
OAI21X1 OAI21X1_889 ( .A(alu__abc_38674_new_n129_), .B(alu__abc_38674_new_n130_), .C(alu__abc_38674_new_n126_), .Y(alu__abc_38674_new_n131_));
OAI21X1 OAI21X1_89 ( .A(_abc_40298_new_n1125_), .B(_abc_40298_new_n1133_), .C(_abc_40298_new_n1136_), .Y(_abc_40298_new_n1137_));
OAI21X1 OAI21X1_890 ( .A(alu__abc_38674_new_n136_), .B(alu__abc_38674_new_n137_), .C(alu__abc_38674_new_n141_), .Y(alu__abc_38674_new_n142_));
OAI21X1 OAI21X1_891 ( .A(alu__abc_38674_new_n145_), .B(alu__abc_38674_new_n146_), .C(alu__abc_38674_new_n150_), .Y(alu__abc_38674_new_n151_));
OAI21X1 OAI21X1_892 ( .A(alu__abc_38674_new_n172_), .B(alu__abc_38674_new_n173_), .C(alu__abc_38674_new_n169_), .Y(alu__abc_38674_new_n174_));
OAI21X1 OAI21X1_893 ( .A(alu__abc_38674_new_n179_), .B(alu__abc_38674_new_n180_), .C(alu__abc_38674_new_n184_), .Y(alu__abc_38674_new_n185_));
OAI21X1 OAI21X1_894 ( .A(alu__abc_38674_new_n194_), .B(alu__abc_38674_new_n195_), .C(alu__abc_38674_new_n191_), .Y(alu__abc_38674_new_n196_));
OAI21X1 OAI21X1_895 ( .A(alu__abc_38674_new_n203_), .B(alu__abc_38674_new_n204_), .C(alu__abc_38674_new_n208_), .Y(alu__abc_38674_new_n209_));
OAI21X1 OAI21X1_896 ( .A(alu__abc_38674_new_n218_), .B(alu__abc_38674_new_n219_), .C(alu__abc_38674_new_n215_), .Y(alu__abc_38674_new_n220_));
OAI21X1 OAI21X1_897 ( .A(alu__abc_38674_new_n248_), .B(alu__abc_38674_new_n249_), .C(alu__abc_38674_new_n247_), .Y(alu__abc_38674_new_n250_));
OAI21X1 OAI21X1_898 ( .A(alu__abc_38674_new_n254_), .B(alu__abc_38674_new_n255_), .C(alu__abc_38674_new_n253_), .Y(alu__abc_38674_new_n256_));
OAI21X1 OAI21X1_899 ( .A(alu__abc_38674_new_n262_), .B(alu__abc_38674_new_n261_), .C(alu__abc_38674_new_n263_), .Y(alu__abc_38674_new_n264_));
OAI21X1 OAI21X1_9 ( .A(_abc_40298_new_n672_), .B(mem_offset_q_0_), .C(_abc_40298_new_n686_), .Y(_abc_40298_new_n687_));
OAI21X1 OAI21X1_90 ( .A(esr_q_9_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n1143_));
OAI21X1 OAI21X1_900 ( .A(alu__abc_38674_new_n279_), .B(alu__abc_38674_new_n286_), .C(alu__abc_38674_new_n283_), .Y(alu_c_update_o));
OAI21X1 OAI21X1_901 ( .A(alu__abc_38674_new_n182_), .B(alu__abc_38674_new_n181_), .C(alu__abc_38674_new_n296_), .Y(alu__abc_38674_new_n297_));
OAI21X1 OAI21X1_902 ( .A(alu_b_i_25_), .B(alu__abc_38674_new_n295_), .C(alu__abc_38674_new_n297_), .Y(alu__abc_38674_new_n298_));
OAI21X1 OAI21X1_903 ( .A(alu__abc_38674_new_n195_), .B(alu__abc_38674_new_n194_), .C(alu__abc_38674_new_n301_), .Y(alu__abc_38674_new_n302_));
OAI21X1 OAI21X1_904 ( .A(alu_b_i_27_), .B(alu__abc_38674_new_n193_), .C(alu__abc_38674_new_n302_), .Y(alu__abc_38674_new_n303_));
OAI21X1 OAI21X1_905 ( .A(alu_b_i_17_), .B(alu__abc_38674_new_n308_), .C(alu__abc_38674_new_n309_), .Y(alu__abc_38674_new_n310_));
OAI21X1 OAI21X1_906 ( .A(alu__abc_38674_new_n130_), .B(alu__abc_38674_new_n129_), .C(alu__abc_38674_new_n317_), .Y(alu__abc_38674_new_n318_));
OAI21X1 OAI21X1_907 ( .A(alu_b_i_21_), .B(alu__abc_38674_new_n128_), .C(alu__abc_38674_new_n318_), .Y(alu__abc_38674_new_n319_));
OAI21X1 OAI21X1_908 ( .A(alu__abc_38674_new_n120_), .B(alu__abc_38674_new_n320_), .C(alu__abc_38674_new_n325_), .Y(alu__abc_38674_new_n326_));
OAI21X1 OAI21X1_909 ( .A(alu__abc_38674_new_n248_), .B(alu__abc_38674_new_n249_), .C(alu__abc_38674_new_n331_), .Y(alu__abc_38674_new_n332_));
OAI21X1 OAI21X1_91 ( .A(_abc_40298_new_n657_), .B(_abc_40298_new_n983_), .C(_abc_40298_new_n1145_), .Y(_abc_40298_new_n1146_));
OAI21X1 OAI21X1_910 ( .A(alu_b_i_7_), .B(alu__abc_38674_new_n329_), .C(alu__abc_38674_new_n332_), .Y(alu__abc_38674_new_n333_));
OAI21X1 OAI21X1_911 ( .A(alu__abc_38674_new_n336_), .B(alu_b_i_1_), .C(alu__abc_38674_new_n264_), .Y(alu__abc_38674_new_n337_));
OAI21X1 OAI21X1_912 ( .A(alu__abc_38674_new_n339_), .B(alu__abc_38674_new_n271_), .C(alu__abc_38674_new_n341_), .Y(alu__abc_38674_new_n342_));
OAI21X1 OAI21X1_913 ( .A(alu__abc_38674_new_n346_), .B(alu__abc_38674_new_n344_), .C(alu__abc_38674_new_n253_), .Y(alu__abc_38674_new_n347_));
OAI21X1 OAI21X1_914 ( .A(alu_b_i_5_), .B(alu__abc_38674_new_n334_), .C(alu__abc_38674_new_n347_), .Y(alu__abc_38674_new_n348_));
OAI21X1 OAI21X1_915 ( .A(alu_b_i_9_), .B(alu__abc_38674_new_n228_), .C(alu__abc_38674_new_n353_), .Y(alu__abc_38674_new_n354_));
OAI21X1 OAI21X1_916 ( .A(alu_b_i_11_), .B(alu__abc_38674_new_n356_), .C(alu__abc_38674_new_n357_), .Y(alu__abc_38674_new_n358_));
OAI21X1 OAI21X1_917 ( .A(alu__abc_38674_new_n219_), .B(alu__abc_38674_new_n218_), .C(alu__abc_38674_new_n361_), .Y(alu__abc_38674_new_n362_));
OAI21X1 OAI21X1_918 ( .A(alu_b_i_13_), .B(alu__abc_38674_new_n217_), .C(alu__abc_38674_new_n362_), .Y(alu__abc_38674_new_n363_));
OAI21X1 OAI21X1_919 ( .A(alu__abc_38674_new_n366_), .B(alu__abc_38674_new_n207_), .C(alu__abc_38674_new_n365_), .Y(alu__abc_38674_new_n367_));
OAI21X1 OAI21X1_92 ( .A(esr_q_10_), .B(_abc_40298_new_n1066_), .C(_abc_40298_new_n1146_), .Y(_abc_40298_new_n1147_));
OAI21X1 OAI21X1_920 ( .A(alu__abc_38674_new_n222_), .B(alu__abc_38674_new_n359_), .C(alu__abc_38674_new_n368_), .Y(alu__abc_38674_new_n369_));
OAI21X1 OAI21X1_921 ( .A(alu__abc_38674_new_n369_), .B(alu__abc_38674_new_n350_), .C(alu__abc_38674_new_n154_), .Y(alu__abc_38674_new_n370_));
OAI21X1 OAI21X1_922 ( .A(alu__abc_38674_new_n174_), .B(alu__abc_38674_new_n372_), .C(alu__abc_38674_new_n375_), .Y(alu__abc_38674_new_n376_));
OAI21X1 OAI21X1_923 ( .A(alu__abc_38674_new_n157_), .B(alu__abc_38674_new_n158_), .C(alu__abc_38674_new_n376_), .Y(alu__abc_38674_new_n377_));
OAI21X1 OAI21X1_924 ( .A(alu_b_i_30_), .B(alu__abc_38674_new_n156_), .C(alu__abc_38674_new_n377_), .Y(alu__abc_38674_new_n378_));
OAI21X1 OAI21X1_925 ( .A(alu_b_i_31_), .B(alu__abc_38674_new_n294_), .C(alu__abc_38674_new_n379_), .Y(alu_less_than_signed_o));
OAI21X1 OAI21X1_926 ( .A(alu__abc_38674_new_n167_), .B(alu__abc_38674_new_n387_), .C(alu__abc_38674_new_n386_), .Y(alu__abc_38674_new_n388_));
OAI21X1 OAI21X1_927 ( .A(alu__abc_38674_new_n393_), .B(alu__abc_38674_new_n396_), .C(alu__abc_38674_new_n394_), .Y(alu__abc_38674_new_n397_));
OAI21X1 OAI21X1_928 ( .A(alu__abc_38674_new_n392_), .B(alu__abc_38674_new_n401_), .C(alu__abc_38674_new_n402_), .Y(alu__abc_38674_new_n403_));
OAI21X1 OAI21X1_929 ( .A(alu__abc_38674_new_n130_), .B(alu__abc_38674_new_n407_), .C(alu__abc_38674_new_n408_), .Y(alu__abc_38674_new_n409_));
OAI21X1 OAI21X1_93 ( .A(_abc_40298_new_n1150_), .B(_abc_40298_new_n1149_), .C(_abc_40298_new_n993_), .Y(_abc_40298_new_n1151_));
OAI21X1 OAI21X1_930 ( .A(alu__abc_38674_new_n414_), .B(alu__abc_38674_new_n413_), .C(alu__abc_38674_new_n416_), .Y(alu__abc_38674_new_n417_));
OAI21X1 OAI21X1_931 ( .A(alu__abc_38674_new_n420_), .B(alu__abc_38674_new_n262_), .C(alu__abc_38674_new_n260_), .Y(alu__abc_38674_new_n421_));
OAI21X1 OAI21X1_932 ( .A(alu__abc_38674_new_n436_), .B(alu__abc_38674_new_n432_), .C(alu__abc_38674_new_n251_), .Y(alu__abc_38674_new_n437_));
OAI21X1 OAI21X1_933 ( .A(alu__abc_38674_new_n438_), .B(alu__abc_38674_new_n430_), .C(alu__abc_38674_new_n440_), .Y(alu__abc_38674_new_n441_));
OAI21X1 OAI21X1_934 ( .A(alu__abc_38674_new_n227_), .B(alu__abc_38674_new_n228_), .C(alu__abc_38674_new_n223_), .Y(alu__abc_38674_new_n444_));
OAI21X1 OAI21X1_935 ( .A(alu_b_i_9_), .B(alu_a_i_9_), .C(alu__abc_38674_new_n444_), .Y(alu__abc_38674_new_n445_));
OAI21X1 OAI21X1_936 ( .A(alu_b_i_11_), .B(alu_a_i_11_), .C(alu__abc_38674_new_n446_), .Y(alu__abc_38674_new_n447_));
OAI21X1 OAI21X1_937 ( .A(alu__abc_38674_new_n445_), .B(alu__abc_38674_new_n443_), .C(alu__abc_38674_new_n448_), .Y(alu__abc_38674_new_n449_));
OAI21X1 OAI21X1_938 ( .A(alu__abc_38674_new_n454_), .B(alu__abc_38674_new_n452_), .C(alu__abc_38674_new_n450_), .Y(alu__abc_38674_new_n455_));
OAI21X1 OAI21X1_939 ( .A(alu__abc_38674_new_n442_), .B(alu__abc_38674_new_n463_), .C(alu__abc_38674_new_n458_), .Y(alu__abc_38674_new_n464_));
OAI21X1 OAI21X1_94 ( .A(esr_q_10_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n1157_));
OAI21X1 OAI21X1_940 ( .A(alu__abc_38674_new_n476_), .B(alu__abc_38674_new_n475_), .C(alu__abc_38674_new_n404_), .Y(alu__abc_38674_new_n477_));
OAI21X1 OAI21X1_941 ( .A(alu__abc_38674_new_n282_), .B(alu__abc_38674_new_n381_), .C(alu__abc_38674_new_n477_), .Y(alu__abc_38674_new_n478_));
OAI21X1 OAI21X1_942 ( .A(alu__abc_38674_new_n479_), .B(alu__abc_38674_new_n470_), .C(alu__abc_38674_new_n401_), .Y(alu__abc_38674_new_n480_));
OAI21X1 OAI21X1_943 ( .A(alu__abc_38674_new_n170_), .B(alu__abc_38674_new_n171_), .C(alu__abc_38674_new_n481_), .Y(alu__abc_38674_new_n482_));
OAI21X1 OAI21X1_944 ( .A(alu__abc_38674_new_n146_), .B(alu__abc_38674_new_n488_), .C(alu__abc_38674_new_n485_), .Y(alu__abc_38674_new_n489_));
OAI21X1 OAI21X1_945 ( .A(alu__abc_38674_new_n126_), .B(alu__abc_38674_new_n491_), .C(alu__abc_38674_new_n407_), .Y(alu__abc_38674_new_n492_));
OAI21X1 OAI21X1_946 ( .A(alu__abc_38674_new_n411_), .B(alu__abc_38674_new_n491_), .C(alu__abc_38674_new_n494_), .Y(alu__abc_38674_new_n495_));
OAI21X1 OAI21X1_947 ( .A(alu__abc_38674_new_n474_), .B(alu__abc_38674_new_n470_), .C(alu__abc_38674_new_n399_), .Y(alu__abc_38674_new_n498_));
OAI21X1 OAI21X1_948 ( .A(alu__abc_38674_new_n180_), .B(alu__abc_38674_new_n470_), .C(alu__abc_38674_new_n501_), .Y(alu__abc_38674_new_n502_));
OAI21X1 OAI21X1_949 ( .A(alu__abc_38674_new_n179_), .B(alu__abc_38674_new_n180_), .C(alu__abc_38674_new_n470_), .Y(alu__abc_38674_new_n506_));
OAI21X1 OAI21X1_95 ( .A(sr_q_2_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n1161_));
OAI21X1 OAI21X1_950 ( .A(alu__abc_38674_new_n441_), .B(alu__abc_38674_new_n524_), .C(alu__abc_38674_new_n462_), .Y(alu__abc_38674_new_n525_));
OAI21X1 OAI21X1_951 ( .A(alu__abc_38674_new_n513_), .B(alu__abc_38674_new_n526_), .C(alu__abc_38674_new_n453_), .Y(alu__abc_38674_new_n527_));
OAI21X1 OAI21X1_952 ( .A(alu__abc_38674_new_n461_), .B(alu__abc_38674_new_n442_), .C(alu__abc_38674_new_n515_), .Y(alu__abc_38674_new_n531_));
OAI21X1 OAI21X1_953 ( .A(alu__abc_38674_new_n529_), .B(alu__abc_38674_new_n532_), .C(alu__abc_38674_new_n512_), .Y(alu__abc_38674_new_n533_));
OAI21X1 OAI21X1_954 ( .A(alu__abc_38674_new_n225_), .B(alu__abc_38674_new_n442_), .C(alu__abc_38674_new_n223_), .Y(alu__abc_38674_new_n536_));
OAI21X1 OAI21X1_955 ( .A(alu__abc_38674_new_n437_), .B(alu__abc_38674_new_n541_), .C(alu__abc_38674_new_n428_), .Y(alu__abc_38674_new_n542_));
OAI21X1 OAI21X1_956 ( .A(alu__abc_38674_new_n254_), .B(alu__abc_38674_new_n550_), .C(alu__abc_38674_new_n433_), .Y(alu__abc_38674_new_n551_));
OAI21X1 OAI21X1_957 ( .A(alu__abc_38674_new_n266_), .B(alu__abc_38674_new_n556_), .C(alu__abc_38674_new_n555_), .Y(alu__abc_38674_new_n557_));
OAI21X1 OAI21X1_958 ( .A(alu__abc_38674_new_n203_), .B(alu__abc_38674_new_n204_), .C(alu__abc_38674_new_n532_), .Y(alu__abc_38674_new_n575_));
OAI21X1 OAI21X1_959 ( .A(alu__abc_38674_new_n212_), .B(alu__abc_38674_new_n582_), .C(alu__abc_38674_new_n451_), .Y(alu__abc_38674_new_n583_));
OAI21X1 OAI21X1_96 ( .A(_abc_40298_new_n1125_), .B(_abc_40298_new_n1133_), .C(_abc_40298_new_n1135_), .Y(_abc_40298_new_n1163_));
OAI21X1 OAI21X1_960 ( .A(alu__abc_38674_new_n585_), .B(alu__abc_38674_new_n442_), .C(alu__abc_38674_new_n445_), .Y(alu__abc_38674_new_n586_));
OAI21X1 OAI21X1_961 ( .A(alu__abc_38674_new_n441_), .B(alu__abc_38674_new_n524_), .C(alu__abc_38674_new_n460_), .Y(alu__abc_38674_new_n589_));
OAI21X1 OAI21X1_962 ( .A(alu__abc_38674_new_n446_), .B(alu__abc_38674_new_n590_), .C(alu__abc_38674_new_n240_), .Y(alu__abc_38674_new_n591_));
OAI21X1 OAI21X1_963 ( .A(alu__abc_38674_new_n134_), .B(alu__abc_38674_new_n135_), .C(alu__abc_38674_new_n601_), .Y(alu__abc_38674_new_n602_));
OAI21X1 OAI21X1_964 ( .A(alu__abc_38674_new_n383_), .B(alu__abc_38674_new_n611_), .C(alu__abc_38674_new_n610_), .Y(alu__abc_38674_new_n612_));
OAI21X1 OAI21X1_965 ( .A(alu__abc_38674_new_n186_), .B(alu__abc_38674_new_n187_), .C(alu__abc_38674_new_n617_), .Y(alu__abc_38674_new_n618_));
OAI21X1 OAI21X1_966 ( .A(alu__abc_38674_new_n110_), .B(alu__abc_38674_new_n111_), .C(alu__abc_38674_new_n621_), .Y(alu__abc_38674_new_n622_));
OAI21X1 OAI21X1_967 ( .A(alu__abc_38674_new_n382_), .B(alu__abc_38674_new_n627_), .C(alu__abc_38674_new_n478_), .Y(alu_c_o));
OAI21X1 OAI21X1_968 ( .A(alu_a_i_10_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n629_), .Y(alu__abc_38674_new_n630_));
OAI21X1 OAI21X1_969 ( .A(alu_a_i_8_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n631_), .Y(alu__abc_38674_new_n632_));
OAI21X1 OAI21X1_97 ( .A(sr_q_9_), .B(REGFILE_SIM_reg_bank_wr_i), .C(enable_i), .Y(_abc_40298_new_n1164_));
OAI21X1 OAI21X1_970 ( .A(alu_a_i_12_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n635_), .Y(alu__abc_38674_new_n636_));
OAI21X1 OAI21X1_971 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n634_), .C(alu__abc_38674_new_n637_), .Y(alu__abc_38674_new_n638_));
OAI21X1 OAI21X1_972 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n633_), .C(alu__abc_38674_new_n639_), .Y(alu__abc_38674_new_n640_));
OAI21X1 OAI21X1_973 ( .A(alu_a_i_2_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n642_), .Y(alu__abc_38674_new_n643_));
OAI21X1 OAI21X1_974 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n643_), .C(alu__abc_38674_new_n646_), .Y(alu__abc_38674_new_n647_));
OAI21X1 OAI21X1_975 ( .A(alu_a_i_4_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n649_), .Y(alu__abc_38674_new_n650_));
OAI21X1 OAI21X1_976 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n648_), .C(alu__abc_38674_new_n651_), .Y(alu__abc_38674_new_n652_));
OAI21X1 OAI21X1_977 ( .A(alu_b_i_2_), .B(alu__abc_38674_new_n647_), .C(alu__abc_38674_new_n653_), .Y(alu__abc_38674_new_n654_));
OAI21X1 OAI21X1_978 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n640_), .C(alu__abc_38674_new_n654_), .Y(alu__abc_38674_new_n655_));
OAI21X1 OAI21X1_979 ( .A(alu__abc_38674_new_n289_), .B(alu__abc_38674_new_n657_), .C(alu__abc_38674_new_n656_), .Y(alu__abc_38674_new_n658_));
OAI21X1 OAI21X1_98 ( .A(_abc_40298_new_n998_), .B(_abc_40298_new_n1010_), .C(_abc_40298_new_n999_), .Y(_abc_40298_new_n1175_));
OAI21X1 OAI21X1_980 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n661_), .C(alu__abc_38674_new_n663_), .Y(alu__abc_38674_new_n664_));
OAI21X1 OAI21X1_981 ( .A(alu_a_i_26_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n665_), .Y(alu__abc_38674_new_n666_));
OAI21X1 OAI21X1_982 ( .A(alu_a_i_24_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n668_), .Y(alu__abc_38674_new_n669_));
OAI21X1 OAI21X1_983 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n667_), .C(alu__abc_38674_new_n670_), .Y(alu__abc_38674_new_n671_));
OAI21X1 OAI21X1_984 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n664_), .C(alu__abc_38674_new_n672_), .Y(alu__abc_38674_new_n673_));
OAI21X1 OAI21X1_985 ( .A(alu_a_i_20_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n676_), .Y(alu__abc_38674_new_n677_));
OAI21X1 OAI21X1_986 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n675_), .C(alu__abc_38674_new_n678_), .Y(alu__abc_38674_new_n679_));
OAI21X1 OAI21X1_987 ( .A(alu_a_i_18_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n682_), .Y(alu__abc_38674_new_n683_));
OAI21X1 OAI21X1_988 ( .A(alu_b_i_1_), .B(alu__abc_38674_new_n681_), .C(alu__abc_38674_new_n684_), .Y(alu__abc_38674_new_n685_));
OAI21X1 OAI21X1_989 ( .A(alu__abc_38674_new_n338_), .B(alu__abc_38674_new_n680_), .C(alu__abc_38674_new_n686_), .Y(alu__abc_38674_new_n687_));
OAI21X1 OAI21X1_99 ( .A(_abc_40298_new_n1000_), .B(_abc_40298_new_n1177_), .C(REGFILE_SIM_reg_bank_reg_rb_o_0_), .Y(_abc_40298_new_n1178_));
OAI21X1 OAI21X1_990 ( .A(alu__abc_38674_new_n340_), .B(alu__abc_38674_new_n674_), .C(alu__abc_38674_new_n688_), .Y(alu__abc_38674_new_n689_));
OAI21X1 OAI21X1_991 ( .A(alu_b_i_4_), .B(alu__abc_38674_new_n655_), .C(alu__abc_38674_new_n690_), .Y(alu__abc_38674_new_n691_));
OAI21X1 OAI21X1_992 ( .A(alu_c_i), .B(alu__abc_38674_new_n692_), .C(alu__abc_38674_new_n693_), .Y(alu__abc_38674_new_n694_));
OAI21X1 OAI21X1_993 ( .A(alu__abc_38674_new_n706_), .B(alu__abc_38674_new_n705_), .C(alu__abc_38674_new_n692_), .Y(alu__abc_38674_new_n707_));
OAI21X1 OAI21X1_994 ( .A(alu__abc_38674_new_n697_), .B(alu__abc_38674_new_n702_), .C(alu__abc_38674_new_n708_), .Y(alu__abc_38674_new_n709_));
OAI21X1 OAI21X1_995 ( .A(alu_op_i_1_), .B(alu_op_i_2_), .C(alu_op_i_3_), .Y(alu__abc_38674_new_n711_));
OAI21X1 OAI21X1_996 ( .A(alu__abc_38674_new_n281_), .B(alu__abc_38674_new_n698_), .C(alu__abc_38674_new_n711_), .Y(alu__abc_38674_new_n712_));
OAI21X1 OAI21X1_997 ( .A(alu__abc_38674_new_n719_), .B(alu__abc_38674_new_n718_), .C(alu__abc_38674_new_n559_), .Y(alu__abc_38674_new_n720_));
OAI21X1 OAI21X1_998 ( .A(alu__abc_38674_new_n559_), .B(alu__abc_38674_new_n717_), .C(alu__abc_38674_new_n720_), .Y(alu__abc_38674_new_n721_));
OAI21X1 OAI21X1_999 ( .A(alu_a_i_15_), .B(alu_b_i_0_), .C(alu__abc_38674_new_n727_), .Y(alu__abc_38674_new_n728_));
OAI22X1 OAI22X1_1 ( .A(_abc_40298_new_n634_), .B(enable_i), .C(_abc_40298_new_n635_), .D(_abc_40298_new_n664_), .Y(_abc_27663_auto_fsm_map_cc_170_map_fsm_2376_4_));
OAI22X1 OAI22X1_10 ( .A(_abc_40298_new_n1213_), .B(_abc_40298_new_n1450_), .C(_abc_40298_new_n1467_), .D(_abc_40298_new_n1465_), .Y(_abc_40298_new_n1468_));
OAI22X1 OAI22X1_100 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3724_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4243_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3659_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4242_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4280_));
OAI22X1 OAI22X1_101 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4049_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4247_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4114_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4246_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4282_));
OAI22X1 OAI22X1_102 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2207_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4250_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3789_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4249_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4283_));
OAI22X1 OAI22X1_103 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2477_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4190_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2543_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4187_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4290_));
OAI22X1 OAI22X1_104 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2675_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4198_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2807_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4195_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4292_));
OAI22X1 OAI22X1_105 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3006_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4202_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3072_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4201_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4293_));
OAI22X1 OAI22X1_106 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3465_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4207_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3530_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4206_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4296_));
OAI22X1 OAI22X1_107 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3986_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4216_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3596_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4214_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4300_));
OAI22X1 OAI22X1_108 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3856_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4218_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3921_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4219_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4301_));
OAI22X1 OAI22X1_109 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3137_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4226_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2411_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4224_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4305_));
OAI22X1 OAI22X1_11 ( .A(_abc_40298_new_n1916_), .B(_abc_40298_new_n1066_), .C(_abc_40298_new_n1929_), .D(_abc_40298_new_n1931_), .Y(_abc_40298_new_n1932_));
OAI22X1 OAI22X1_110 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2343_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4229_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2111_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4228_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4306_));
OAI22X1 OAI22X1_111 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2940_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4235_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2872_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4234_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4308_));
OAI22X1 OAI22X1_112 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3400_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4239_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3334_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4240_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4311_));
OAI22X1 OAI22X1_113 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3726_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4243_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3661_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4242_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4312_));
OAI22X1 OAI22X1_114 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4051_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4247_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4116_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4246_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4314_));
OAI22X1 OAI22X1_115 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2209_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4250_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3791_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4249_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4315_));
OAI22X1 OAI22X1_116 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2479_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4190_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2545_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4187_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4322_));
OAI22X1 OAI22X1_117 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2677_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4198_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2809_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4195_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4324_));
OAI22X1 OAI22X1_118 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3008_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4202_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3074_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4201_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4325_));
OAI22X1 OAI22X1_119 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3467_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4207_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3532_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4206_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4328_));
OAI22X1 OAI22X1_12 ( .A(_abc_40298_new_n2139_), .B(_abc_40298_new_n2151_), .C(_abc_40298_new_n911_), .D(_abc_40298_new_n2146_), .Y(alu_input_b_r_0_));
OAI22X1 OAI22X1_120 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3988_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4216_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3598_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4214_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4332_));
OAI22X1 OAI22X1_121 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3858_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4218_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3923_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4219_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4333_));
OAI22X1 OAI22X1_122 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3139_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4226_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2413_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4224_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4337_));
OAI22X1 OAI22X1_123 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2345_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4229_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2114_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4228_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4338_));
OAI22X1 OAI22X1_124 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2942_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4235_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2874_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4234_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4340_));
OAI22X1 OAI22X1_125 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3402_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4239_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3336_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4240_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4343_));
OAI22X1 OAI22X1_126 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3728_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4243_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3663_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4242_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4344_));
OAI22X1 OAI22X1_127 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4053_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4247_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4118_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4246_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4346_));
OAI22X1 OAI22X1_128 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2211_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4250_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3793_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4249_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4347_));
OAI22X1 OAI22X1_129 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2481_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4190_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2547_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4187_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4354_));
OAI22X1 OAI22X1_13 ( .A(_abc_40298_new_n2153_), .B(_abc_40298_new_n2151_), .C(_abc_40298_new_n909_), .D(_abc_40298_new_n2146_), .Y(alu_input_b_r_1_));
OAI22X1 OAI22X1_130 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2679_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4198_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2811_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4195_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4356_));
OAI22X1 OAI22X1_131 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3010_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4202_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3076_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4201_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4357_));
OAI22X1 OAI22X1_132 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3469_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4207_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3534_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4206_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4360_));
OAI22X1 OAI22X1_133 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3990_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4216_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3600_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4214_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4364_));
OAI22X1 OAI22X1_134 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3860_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4218_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3925_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4219_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4365_));
OAI22X1 OAI22X1_135 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3141_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4226_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2415_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4224_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4369_));
OAI22X1 OAI22X1_136 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2347_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4229_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2117_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4228_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4370_));
OAI22X1 OAI22X1_137 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2944_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4235_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2876_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4234_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4372_));
OAI22X1 OAI22X1_138 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3404_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4239_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3338_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4240_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4375_));
OAI22X1 OAI22X1_139 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3730_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4243_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3665_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4242_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4376_));
OAI22X1 OAI22X1_14 ( .A(_abc_40298_new_n1030_), .B(_abc_40298_new_n2151_), .C(_abc_40298_new_n898_), .D(_abc_40298_new_n2146_), .Y(alu_input_b_r_2_));
OAI22X1 OAI22X1_140 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4055_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4247_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4120_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4246_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4378_));
OAI22X1 OAI22X1_141 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2213_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4250_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3795_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4249_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4379_));
OAI22X1 OAI22X1_142 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2483_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4190_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2549_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4187_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4386_));
OAI22X1 OAI22X1_143 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2681_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4198_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2813_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4195_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4388_));
OAI22X1 OAI22X1_144 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3012_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4202_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3078_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4201_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4389_));
OAI22X1 OAI22X1_145 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3471_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4207_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3536_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4206_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4392_));
OAI22X1 OAI22X1_146 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3992_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4216_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3602_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4214_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4396_));
OAI22X1 OAI22X1_147 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3862_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4218_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3927_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4219_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4397_));
OAI22X1 OAI22X1_148 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3143_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4226_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2417_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4224_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4401_));
OAI22X1 OAI22X1_149 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2349_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4229_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2120_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4228_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4402_));
OAI22X1 OAI22X1_15 ( .A(_abc_40298_new_n1233_), .B(_abc_40298_new_n2151_), .C(_abc_40298_new_n903_), .D(_abc_40298_new_n2146_), .Y(alu_input_b_r_3_));
OAI22X1 OAI22X1_150 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2946_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4235_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2878_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4234_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4404_));
OAI22X1 OAI22X1_151 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3406_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4239_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3340_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4240_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4407_));
OAI22X1 OAI22X1_152 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3732_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4243_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3667_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4242_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4408_));
OAI22X1 OAI22X1_153 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4057_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4247_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4122_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4246_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4410_));
OAI22X1 OAI22X1_154 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2215_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4250_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3797_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4249_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4411_));
OAI22X1 OAI22X1_155 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2485_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4190_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2551_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4187_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4418_));
OAI22X1 OAI22X1_156 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2683_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4198_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2815_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4195_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4420_));
OAI22X1 OAI22X1_157 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3014_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4202_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3080_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4201_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4421_));
OAI22X1 OAI22X1_158 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3473_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4207_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3538_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4206_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4424_));
OAI22X1 OAI22X1_159 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3994_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4216_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3604_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4214_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4428_));
OAI22X1 OAI22X1_16 ( .A(_abc_40298_new_n1260_), .B(_abc_40298_new_n2151_), .C(_abc_40298_new_n1315_), .D(_abc_40298_new_n2146_), .Y(alu_input_b_r_4_));
OAI22X1 OAI22X1_160 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3864_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4218_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3929_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4219_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4429_));
OAI22X1 OAI22X1_161 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3145_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4226_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2419_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4224_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4433_));
OAI22X1 OAI22X1_162 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2351_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4229_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2123_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4228_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4434_));
OAI22X1 OAI22X1_163 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2948_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4235_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2880_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4234_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4436_));
OAI22X1 OAI22X1_164 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3408_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4239_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3342_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4240_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4439_));
OAI22X1 OAI22X1_165 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3734_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4243_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3669_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4242_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4440_));
OAI22X1 OAI22X1_166 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4059_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4247_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4124_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4246_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4442_));
OAI22X1 OAI22X1_167 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2217_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4250_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3799_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4249_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4443_));
OAI22X1 OAI22X1_168 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2487_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4190_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2553_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4187_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4450_));
OAI22X1 OAI22X1_169 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2685_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4198_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2817_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4195_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4452_));
OAI22X1 OAI22X1_17 ( .A(_abc_40298_new_n1293_), .B(_abc_40298_new_n2151_), .C(_abc_40298_new_n1341_), .D(_abc_40298_new_n2146_), .Y(alu_input_b_r_5_));
OAI22X1 OAI22X1_170 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3016_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4202_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3082_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4201_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4453_));
OAI22X1 OAI22X1_171 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3475_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4207_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3540_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4206_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4456_));
OAI22X1 OAI22X1_172 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3996_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4216_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3606_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4214_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4460_));
OAI22X1 OAI22X1_173 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3866_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4218_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3931_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4219_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4461_));
OAI22X1 OAI22X1_174 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3147_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4226_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2421_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4224_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4465_));
OAI22X1 OAI22X1_175 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2353_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4229_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2126_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4228_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4466_));
OAI22X1 OAI22X1_176 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2950_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4235_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2882_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4234_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4468_));
OAI22X1 OAI22X1_177 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3410_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4239_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3344_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4240_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4471_));
OAI22X1 OAI22X1_178 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3736_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4243_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3671_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4242_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4472_));
OAI22X1 OAI22X1_179 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4061_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4247_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4126_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4246_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4474_));
OAI22X1 OAI22X1_18 ( .A(_abc_40298_new_n1811_), .B(_abc_40298_new_n2176_), .C(_abc_40298_new_n2202_), .D(_abc_40298_new_n2248_), .Y(alu_input_b_r_24_));
OAI22X1 OAI22X1_180 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2219_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4250_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3801_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4249_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4475_));
OAI22X1 OAI22X1_181 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2489_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4190_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2555_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4187_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4482_));
OAI22X1 OAI22X1_182 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2687_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4198_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2819_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4195_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4484_));
OAI22X1 OAI22X1_183 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3018_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4202_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3084_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4201_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4485_));
OAI22X1 OAI22X1_184 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3477_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4207_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3542_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4206_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4488_));
OAI22X1 OAI22X1_185 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3998_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4216_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3608_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4214_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4492_));
OAI22X1 OAI22X1_186 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3868_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4218_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3933_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4219_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4493_));
OAI22X1 OAI22X1_187 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3149_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4226_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2423_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4224_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4497_));
OAI22X1 OAI22X1_188 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2355_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4229_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2129_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4228_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4498_));
OAI22X1 OAI22X1_189 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2952_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4235_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2884_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4234_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4500_));
OAI22X1 OAI22X1_19 ( .A(_abc_40298_new_n1853_), .B(_abc_40298_new_n2176_), .C(_abc_40298_new_n2202_), .D(_abc_40298_new_n2252_), .Y(alu_input_b_r_25_));
OAI22X1 OAI22X1_190 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3412_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4239_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3346_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4240_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4503_));
OAI22X1 OAI22X1_191 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3738_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4243_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3673_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4242_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4504_));
OAI22X1 OAI22X1_192 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4063_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4247_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4128_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4246_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4506_));
OAI22X1 OAI22X1_193 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2221_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4250_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3803_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4249_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4507_));
OAI22X1 OAI22X1_194 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2491_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4190_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2557_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4187_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4514_));
OAI22X1 OAI22X1_195 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2689_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4198_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2821_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4195_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4516_));
OAI22X1 OAI22X1_196 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3020_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4202_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3086_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4201_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4517_));
OAI22X1 OAI22X1_197 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3479_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4207_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3544_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4206_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4520_));
OAI22X1 OAI22X1_198 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4000_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4216_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3610_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4214_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4524_));
OAI22X1 OAI22X1_199 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3870_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4218_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3935_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4219_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4525_));
OAI22X1 OAI22X1_2 ( .A(_abc_40298_new_n771_), .B(_abc_40298_new_n698_), .C(_abc_40298_new_n770_), .D(_abc_40298_new_n695_), .Y(_abc_40298_new_n772_));
OAI22X1 OAI22X1_20 ( .A(_abc_40298_new_n1868_), .B(_abc_40298_new_n2176_), .C(_abc_40298_new_n2202_), .D(_abc_40298_new_n2256_), .Y(alu_input_b_r_26_));
OAI22X1 OAI22X1_200 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3151_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4226_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2425_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4224_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4529_));
OAI22X1 OAI22X1_201 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2357_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4229_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2132_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4228_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4530_));
OAI22X1 OAI22X1_202 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2954_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4235_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2886_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4234_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4532_));
OAI22X1 OAI22X1_203 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3414_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4239_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3348_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4240_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4535_));
OAI22X1 OAI22X1_204 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3740_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4243_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3675_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4242_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4536_));
OAI22X1 OAI22X1_205 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4065_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4247_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4130_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4246_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4538_));
OAI22X1 OAI22X1_206 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2223_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4250_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3805_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4249_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4539_));
OAI22X1 OAI22X1_207 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2493_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4190_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2559_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4187_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4546_));
OAI22X1 OAI22X1_208 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2691_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4198_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2823_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4195_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4548_));
OAI22X1 OAI22X1_209 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3022_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4202_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3088_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4201_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4549_));
OAI22X1 OAI22X1_21 ( .A(_abc_40298_new_n1950_), .B(_abc_40298_new_n2176_), .C(_abc_40298_new_n2202_), .D(_abc_40298_new_n2270_), .Y(alu_input_b_r_29_));
OAI22X1 OAI22X1_210 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3481_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4207_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3546_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4206_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4552_));
OAI22X1 OAI22X1_211 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4002_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4216_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3612_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4214_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4556_));
OAI22X1 OAI22X1_212 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3872_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4218_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3937_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4219_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4557_));
OAI22X1 OAI22X1_213 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3153_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4226_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2427_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4224_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4561_));
OAI22X1 OAI22X1_214 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2359_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4229_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2135_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4228_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4562_));
OAI22X1 OAI22X1_215 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2956_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4235_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2888_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4234_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4564_));
OAI22X1 OAI22X1_216 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3416_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4239_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3350_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4240_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4567_));
OAI22X1 OAI22X1_217 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3742_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4243_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3677_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4242_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4568_));
OAI22X1 OAI22X1_218 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4067_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4247_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4132_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4246_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4570_));
OAI22X1 OAI22X1_219 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2225_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4250_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3807_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4249_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4571_));
OAI22X1 OAI22X1_22 ( .A(_abc_40298_new_n1967_), .B(_abc_40298_new_n2176_), .C(_abc_40298_new_n2202_), .D(_abc_40298_new_n2274_), .Y(alu_input_b_r_30_));
OAI22X1 OAI22X1_220 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2495_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4190_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2561_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4187_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4578_));
OAI22X1 OAI22X1_221 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2693_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4198_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2825_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4195_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4580_));
OAI22X1 OAI22X1_222 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3024_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4202_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3090_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4201_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4581_));
OAI22X1 OAI22X1_223 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3483_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4207_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3548_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4206_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4584_));
OAI22X1 OAI22X1_224 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4004_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4216_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3614_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4214_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4588_));
OAI22X1 OAI22X1_225 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3874_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4218_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3939_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4219_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4589_));
OAI22X1 OAI22X1_226 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3155_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4226_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2429_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4224_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4593_));
OAI22X1 OAI22X1_227 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2361_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4229_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2138_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4228_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4594_));
OAI22X1 OAI22X1_228 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2958_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4235_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2890_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4234_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4596_));
OAI22X1 OAI22X1_229 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3418_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4239_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3352_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4240_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4599_));
OAI22X1 OAI22X1_23 ( .A(_abc_40298_new_n1996_), .B(_abc_40298_new_n2176_), .C(_abc_40298_new_n2202_), .D(_abc_40298_new_n2278_), .Y(alu_input_b_r_31_));
OAI22X1 OAI22X1_230 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3744_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4243_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3679_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4242_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4600_));
OAI22X1 OAI22X1_231 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4069_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4247_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4134_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4246_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4602_));
OAI22X1 OAI22X1_232 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2227_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4250_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3809_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4249_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4603_));
OAI22X1 OAI22X1_233 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2497_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4190_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2563_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4187_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4610_));
OAI22X1 OAI22X1_234 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2695_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4198_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2827_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4195_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4612_));
OAI22X1 OAI22X1_235 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3026_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4202_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3092_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4201_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4613_));
OAI22X1 OAI22X1_236 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3485_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4207_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3550_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4206_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4616_));
OAI22X1 OAI22X1_237 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4006_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4216_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3616_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4214_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4620_));
OAI22X1 OAI22X1_238 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3876_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4218_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3941_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4219_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4621_));
OAI22X1 OAI22X1_239 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3157_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4226_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2431_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4224_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4625_));
OAI22X1 OAI22X1_24 ( .A(_abc_40298_new_n2299_), .B(_abc_40298_new_n2120_), .C(_abc_40298_new_n2305_), .D(_abc_40298_new_n2304_), .Y(alu_input_a_r_2_));
OAI22X1 OAI22X1_240 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2363_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4229_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2141_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4228_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4626_));
OAI22X1 OAI22X1_241 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2960_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4235_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2892_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4234_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4628_));
OAI22X1 OAI22X1_242 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3420_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4239_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3354_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4240_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4631_));
OAI22X1 OAI22X1_243 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3746_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4243_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3681_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4242_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4632_));
OAI22X1 OAI22X1_244 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4071_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4247_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4136_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4246_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4634_));
OAI22X1 OAI22X1_245 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2229_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4250_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3811_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4249_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4635_));
OAI22X1 OAI22X1_246 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2499_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4190_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2565_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4187_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4642_));
OAI22X1 OAI22X1_247 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2697_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4198_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2829_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4195_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4644_));
OAI22X1 OAI22X1_248 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3028_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4202_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3094_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4201_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4645_));
OAI22X1 OAI22X1_249 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3487_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4207_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3552_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4206_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4648_));
OAI22X1 OAI22X1_25 ( .A(_abc_40298_new_n1013_), .B(_abc_40298_new_n1290_), .C(_abc_40298_new_n2323_), .D(_abc_40298_new_n2322_), .Y(_abc_40298_new_n2324_));
OAI22X1 OAI22X1_250 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4008_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4216_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3618_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4214_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4652_));
OAI22X1 OAI22X1_251 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3878_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4218_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3943_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4219_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4653_));
OAI22X1 OAI22X1_252 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3159_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4226_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2433_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4224_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4657_));
OAI22X1 OAI22X1_253 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2365_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4229_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2144_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4228_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4658_));
OAI22X1 OAI22X1_254 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2962_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4235_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2894_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4234_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4660_));
OAI22X1 OAI22X1_255 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3422_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4239_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3356_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4240_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4663_));
OAI22X1 OAI22X1_256 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3748_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4243_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3683_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4242_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4664_));
OAI22X1 OAI22X1_257 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4073_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4247_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4138_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4246_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4666_));
OAI22X1 OAI22X1_258 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2231_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4250_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3813_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4249_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4667_));
OAI22X1 OAI22X1_259 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2501_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4190_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2567_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4187_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4674_));
OAI22X1 OAI22X1_26 ( .A(_abc_40298_new_n1153_), .B(_abc_40298_new_n1080_), .C(_abc_40298_new_n1437_), .D(_abc_40298_new_n1185_), .Y(_abc_40298_new_n2359_));
OAI22X1 OAI22X1_260 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2699_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4198_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2831_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4195_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4676_));
OAI22X1 OAI22X1_261 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3030_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4202_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3096_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4201_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4677_));
OAI22X1 OAI22X1_262 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3489_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4207_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3554_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4206_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4680_));
OAI22X1 OAI22X1_263 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4010_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4216_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3620_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4214_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4684_));
OAI22X1 OAI22X1_264 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3880_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4218_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3945_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4219_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4685_));
OAI22X1 OAI22X1_265 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3161_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4226_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2435_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4224_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4689_));
OAI22X1 OAI22X1_266 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2367_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4229_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2147_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4228_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4690_));
OAI22X1 OAI22X1_267 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2964_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4235_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2896_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4234_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4692_));
OAI22X1 OAI22X1_268 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3424_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4239_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3358_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4240_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4695_));
OAI22X1 OAI22X1_269 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3750_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4243_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3685_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4242_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4696_));
OAI22X1 OAI22X1_27 ( .A(_abc_40298_new_n2358_), .B(_abc_40298_new_n2302_), .C(_abc_40298_new_n1002_), .D(_abc_40298_new_n2360_), .Y(_abc_40298_new_n2361_));
OAI22X1 OAI22X1_270 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4075_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4247_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4140_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4246_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4698_));
OAI22X1 OAI22X1_271 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2233_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4250_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3815_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4249_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4699_));
OAI22X1 OAI22X1_272 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2503_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4190_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2569_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4187_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4706_));
OAI22X1 OAI22X1_273 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2701_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4198_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2833_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4195_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4708_));
OAI22X1 OAI22X1_274 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3032_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4202_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3098_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4201_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4709_));
OAI22X1 OAI22X1_275 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3491_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4207_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3556_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4206_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4712_));
OAI22X1 OAI22X1_276 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4012_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4216_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3622_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4214_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4716_));
OAI22X1 OAI22X1_277 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3882_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4218_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3947_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4219_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4717_));
OAI22X1 OAI22X1_278 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3163_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4226_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2437_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4224_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4721_));
OAI22X1 OAI22X1_279 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2369_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4229_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2150_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4228_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4722_));
OAI22X1 OAI22X1_28 ( .A(_abc_40298_new_n2387_), .B(_abc_40298_new_n2389_), .C(_abc_40298_new_n1013_), .D(_abc_40298_new_n1590_), .Y(_abc_40298_new_n2390_));
OAI22X1 OAI22X1_280 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2966_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4235_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2898_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4234_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4724_));
OAI22X1 OAI22X1_281 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3426_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4239_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3360_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4240_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4727_));
OAI22X1 OAI22X1_282 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3752_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4243_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3687_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4242_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4728_));
OAI22X1 OAI22X1_283 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4077_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4247_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4142_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4246_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4730_));
OAI22X1 OAI22X1_284 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2235_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4250_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3817_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4249_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4731_));
OAI22X1 OAI22X1_285 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2505_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4190_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2571_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4187_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4738_));
OAI22X1 OAI22X1_286 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2703_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4198_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2835_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4195_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4740_));
OAI22X1 OAI22X1_287 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3034_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4202_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3100_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4201_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4741_));
OAI22X1 OAI22X1_288 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3493_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4207_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3558_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4206_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4744_));
OAI22X1 OAI22X1_289 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4014_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4216_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3624_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4214_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4748_));
OAI22X1 OAI22X1_29 ( .A(_abc_40298_new_n2394_), .B(_abc_40298_new_n2396_), .C(_abc_40298_new_n1013_), .D(_abc_40298_new_n1623_), .Y(_abc_40298_new_n2397_));
OAI22X1 OAI22X1_290 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3884_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4218_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3949_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4219_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4749_));
OAI22X1 OAI22X1_291 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3165_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4226_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2439_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4224_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4753_));
OAI22X1 OAI22X1_292 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2371_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4229_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2153_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4228_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4754_));
OAI22X1 OAI22X1_293 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2968_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4235_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2900_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4234_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4756_));
OAI22X1 OAI22X1_294 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3428_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4239_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3362_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4240_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4759_));
OAI22X1 OAI22X1_295 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3754_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4243_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3689_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4242_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4760_));
OAI22X1 OAI22X1_296 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4079_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4247_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4144_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4246_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4762_));
OAI22X1 OAI22X1_297 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2237_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4250_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3819_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4249_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4763_));
OAI22X1 OAI22X1_298 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2507_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4190_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2573_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4187_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4770_));
OAI22X1 OAI22X1_299 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2705_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4198_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2837_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4195_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4772_));
OAI22X1 OAI22X1_3 ( .A(_abc_40298_new_n771_), .B(_abc_40298_new_n710_), .C(_abc_40298_new_n776_), .D(_abc_40298_new_n695_), .Y(_abc_40298_new_n777_));
OAI22X1 OAI22X1_30 ( .A(_abc_40298_new_n2401_), .B(_abc_40298_new_n2403_), .C(_abc_40298_new_n1013_), .D(_abc_40298_new_n1649_), .Y(_abc_40298_new_n2404_));
OAI22X1 OAI22X1_300 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3036_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4202_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3102_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4201_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4773_));
OAI22X1 OAI22X1_301 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3495_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4207_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3560_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4206_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4776_));
OAI22X1 OAI22X1_302 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4016_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4216_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3626_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4214_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4780_));
OAI22X1 OAI22X1_303 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3886_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4218_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3951_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4219_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4781_));
OAI22X1 OAI22X1_304 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3167_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4226_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2441_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4224_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4785_));
OAI22X1 OAI22X1_305 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2373_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4229_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2156_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4228_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4786_));
OAI22X1 OAI22X1_306 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2970_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4235_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2902_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4234_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4788_));
OAI22X1 OAI22X1_307 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3430_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4239_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3364_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4240_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4791_));
OAI22X1 OAI22X1_308 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3756_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4243_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3691_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4242_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4792_));
OAI22X1 OAI22X1_309 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4081_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4247_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4146_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4246_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4794_));
OAI22X1 OAI22X1_31 ( .A(_abc_40298_new_n2408_), .B(_abc_40298_new_n2410_), .C(_abc_40298_new_n1013_), .D(_abc_40298_new_n1677_), .Y(_abc_40298_new_n2411_));
OAI22X1 OAI22X1_310 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2239_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4250_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3821_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4249_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4795_));
OAI22X1 OAI22X1_311 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2509_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4190_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2575_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4187_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4802_));
OAI22X1 OAI22X1_312 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2707_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4198_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2839_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4195_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4804_));
OAI22X1 OAI22X1_313 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3038_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4202_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3104_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4201_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4805_));
OAI22X1 OAI22X1_314 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3497_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4207_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3562_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4206_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4808_));
OAI22X1 OAI22X1_315 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4018_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4216_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3628_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4214_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4812_));
OAI22X1 OAI22X1_316 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3888_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4218_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3953_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4219_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4813_));
OAI22X1 OAI22X1_317 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3169_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4226_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2443_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4224_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4817_));
OAI22X1 OAI22X1_318 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2375_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4229_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2159_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4228_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4818_));
OAI22X1 OAI22X1_319 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2972_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4235_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2904_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4234_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4820_));
OAI22X1 OAI22X1_32 ( .A(_abc_40298_new_n2415_), .B(_abc_40298_new_n2417_), .C(_abc_40298_new_n1013_), .D(_abc_40298_new_n1701_), .Y(_abc_40298_new_n2418_));
OAI22X1 OAI22X1_320 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3432_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4239_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3366_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4240_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4823_));
OAI22X1 OAI22X1_321 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3758_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4243_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3693_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4242_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4824_));
OAI22X1 OAI22X1_322 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4083_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4247_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4148_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4246_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4826_));
OAI22X1 OAI22X1_323 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2241_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4250_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3823_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4249_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4827_));
OAI22X1 OAI22X1_324 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2511_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4190_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2577_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4187_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4834_));
OAI22X1 OAI22X1_325 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2709_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4198_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2841_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4195_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4836_));
OAI22X1 OAI22X1_326 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3040_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4202_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3106_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4201_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4837_));
OAI22X1 OAI22X1_327 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3499_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4207_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3564_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4206_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4840_));
OAI22X1 OAI22X1_328 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4020_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4216_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3630_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4214_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4844_));
OAI22X1 OAI22X1_329 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3890_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4218_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3955_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4219_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4845_));
OAI22X1 OAI22X1_33 ( .A(_abc_40298_new_n2422_), .B(_abc_40298_new_n2424_), .C(_abc_40298_new_n1013_), .D(_abc_40298_new_n1729_), .Y(_abc_40298_new_n2425_));
OAI22X1 OAI22X1_330 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3171_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4226_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2445_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4224_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4849_));
OAI22X1 OAI22X1_331 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2377_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4229_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2162_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4228_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4850_));
OAI22X1 OAI22X1_332 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2974_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4235_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2906_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4234_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4852_));
OAI22X1 OAI22X1_333 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3434_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4239_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3368_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4240_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4855_));
OAI22X1 OAI22X1_334 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3760_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4243_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3695_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4242_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4856_));
OAI22X1 OAI22X1_335 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4085_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4247_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4150_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4246_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4858_));
OAI22X1 OAI22X1_336 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2243_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4250_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3825_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4249_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4859_));
OAI22X1 OAI22X1_337 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2513_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4190_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2579_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4187_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4866_));
OAI22X1 OAI22X1_338 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2711_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4198_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2843_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4195_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4868_));
OAI22X1 OAI22X1_339 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3042_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4202_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3108_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4201_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4869_));
OAI22X1 OAI22X1_34 ( .A(_abc_40298_new_n2429_), .B(_abc_40298_new_n2431_), .C(_abc_40298_new_n1013_), .D(_abc_40298_new_n1758_), .Y(_abc_40298_new_n2432_));
OAI22X1 OAI22X1_340 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3501_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4207_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3566_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4206_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4872_));
OAI22X1 OAI22X1_341 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4022_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4216_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3632_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4214_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4876_));
OAI22X1 OAI22X1_342 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3892_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4218_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3957_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4219_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4877_));
OAI22X1 OAI22X1_343 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3173_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4226_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2447_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4224_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4881_));
OAI22X1 OAI22X1_344 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2379_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4229_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2165_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4228_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4882_));
OAI22X1 OAI22X1_345 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2976_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4235_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2908_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4234_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4884_));
OAI22X1 OAI22X1_346 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3436_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4239_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3370_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4240_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4887_));
OAI22X1 OAI22X1_347 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3762_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4243_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3697_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4242_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4888_));
OAI22X1 OAI22X1_348 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4087_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4247_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4152_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4246_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4890_));
OAI22X1 OAI22X1_349 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2245_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4250_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3827_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4249_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4891_));
OAI22X1 OAI22X1_35 ( .A(_abc_40298_new_n2436_), .B(_abc_40298_new_n2438_), .C(_abc_40298_new_n1013_), .D(_abc_40298_new_n1785_), .Y(_abc_40298_new_n2439_));
OAI22X1 OAI22X1_350 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2515_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4190_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2581_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4187_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4898_));
OAI22X1 OAI22X1_351 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2713_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4198_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2845_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4195_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4900_));
OAI22X1 OAI22X1_352 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3044_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4202_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3110_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4201_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4901_));
OAI22X1 OAI22X1_353 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3503_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4207_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3568_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4206_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4904_));
OAI22X1 OAI22X1_354 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4024_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4216_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3634_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4214_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4908_));
OAI22X1 OAI22X1_355 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3894_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4218_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3959_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4219_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4909_));
OAI22X1 OAI22X1_356 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3175_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4226_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2449_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4224_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4913_));
OAI22X1 OAI22X1_357 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2381_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4229_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2168_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4228_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4914_));
OAI22X1 OAI22X1_358 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2978_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4235_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2910_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4234_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4916_));
OAI22X1 OAI22X1_359 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3438_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4239_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3372_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4240_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4919_));
OAI22X1 OAI22X1_36 ( .A(_abc_40298_new_n2443_), .B(_abc_40298_new_n2445_), .C(_abc_40298_new_n1013_), .D(_abc_40298_new_n1809_), .Y(_abc_40298_new_n2446_));
OAI22X1 OAI22X1_360 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3764_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4243_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3699_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4242_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4920_));
OAI22X1 OAI22X1_361 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4089_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4247_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4154_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4246_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4922_));
OAI22X1 OAI22X1_362 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2247_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4250_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3829_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4249_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4923_));
OAI22X1 OAI22X1_363 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2517_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4190_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2583_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4187_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4930_));
OAI22X1 OAI22X1_364 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2715_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4198_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2847_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4195_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4932_));
OAI22X1 OAI22X1_365 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3046_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4202_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3112_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4201_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4933_));
OAI22X1 OAI22X1_366 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3505_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4207_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3570_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4206_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4936_));
OAI22X1 OAI22X1_367 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4026_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4216_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3636_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4214_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4940_));
OAI22X1 OAI22X1_368 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3896_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4218_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3961_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4219_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4941_));
OAI22X1 OAI22X1_369 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3177_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4226_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2451_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4224_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4945_));
OAI22X1 OAI22X1_37 ( .A(_abc_40298_new_n2450_), .B(_abc_40298_new_n2452_), .C(_abc_40298_new_n1013_), .D(_abc_40298_new_n1841_), .Y(_abc_40298_new_n2453_));
OAI22X1 OAI22X1_370 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2383_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4229_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2171_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4228_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4946_));
OAI22X1 OAI22X1_371 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2980_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4235_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2912_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4234_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4948_));
OAI22X1 OAI22X1_372 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3440_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4239_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3374_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4240_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4951_));
OAI22X1 OAI22X1_373 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3766_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4243_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3701_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4242_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4952_));
OAI22X1 OAI22X1_374 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4091_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4247_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4156_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4246_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4954_));
OAI22X1 OAI22X1_375 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2249_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4250_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3831_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4249_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4955_));
OAI22X1 OAI22X1_376 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2519_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4190_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2585_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4187_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4962_));
OAI22X1 OAI22X1_377 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2717_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4198_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2849_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4195_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4964_));
OAI22X1 OAI22X1_378 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3048_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4202_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3114_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4201_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4965_));
OAI22X1 OAI22X1_379 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3507_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4207_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3572_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4206_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4968_));
OAI22X1 OAI22X1_38 ( .A(_abc_40298_new_n2458_), .B(_abc_40298_new_n2460_), .C(_abc_40298_new_n1013_), .D(_abc_40298_new_n1866_), .Y(_abc_40298_new_n2461_));
OAI22X1 OAI22X1_380 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4028_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4216_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3638_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4214_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4972_));
OAI22X1 OAI22X1_381 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3898_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4218_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3963_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4219_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4973_));
OAI22X1 OAI22X1_382 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3179_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4226_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2453_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4224_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4977_));
OAI22X1 OAI22X1_383 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2385_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4229_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2174_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4228_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4978_));
OAI22X1 OAI22X1_384 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2982_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4235_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2914_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4234_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4980_));
OAI22X1 OAI22X1_385 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3442_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4239_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3376_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4240_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4983_));
OAI22X1 OAI22X1_386 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3768_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4243_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3703_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4242_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4984_));
OAI22X1 OAI22X1_387 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4093_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4247_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4158_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4246_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4986_));
OAI22X1 OAI22X1_388 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2251_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4250_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3833_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4249_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4987_));
OAI22X1 OAI22X1_389 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2521_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4190_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2587_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4187_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4994_));
OAI22X1 OAI22X1_39 ( .A(_abc_40298_new_n2465_), .B(_abc_40298_new_n2467_), .C(_abc_40298_new_n1013_), .D(_abc_40298_new_n1892_), .Y(_abc_40298_new_n2468_));
OAI22X1 OAI22X1_390 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2719_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4198_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2851_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4195_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4996_));
OAI22X1 OAI22X1_391 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3050_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4202_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3116_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4201_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4997_));
OAI22X1 OAI22X1_392 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3509_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4207_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3574_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4206_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5000_));
OAI22X1 OAI22X1_393 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4030_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4216_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3640_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4214_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5004_));
OAI22X1 OAI22X1_394 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3900_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4218_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3965_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4219_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5005_));
OAI22X1 OAI22X1_395 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3181_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4226_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2455_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4224_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5009_));
OAI22X1 OAI22X1_396 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2387_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4229_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2177_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4228_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5010_));
OAI22X1 OAI22X1_397 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2984_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4235_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2916_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4234_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5012_));
OAI22X1 OAI22X1_398 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3444_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4239_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3378_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4240_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5015_));
OAI22X1 OAI22X1_399 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3770_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4243_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3705_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4242_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5016_));
OAI22X1 OAI22X1_4 ( .A(_abc_40298_new_n771_), .B(_abc_40298_new_n721_), .C(_abc_40298_new_n781_), .D(_abc_40298_new_n695_), .Y(_abc_40298_new_n782_));
OAI22X1 OAI22X1_40 ( .A(_abc_40298_new_n2473_), .B(_abc_40298_new_n2475_), .C(_abc_40298_new_n1013_), .D(_abc_40298_new_n1914_), .Y(_abc_40298_new_n2476_));
OAI22X1 OAI22X1_400 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4095_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4247_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4160_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4246_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5018_));
OAI22X1 OAI22X1_401 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2253_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4250_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3835_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4249_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5019_));
OAI22X1 OAI22X1_402 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2523_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4190_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2589_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4187_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5026_));
OAI22X1 OAI22X1_403 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2721_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4198_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2853_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4195_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5028_));
OAI22X1 OAI22X1_404 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3052_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4202_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3118_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4201_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5029_));
OAI22X1 OAI22X1_405 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3511_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4207_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3576_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4206_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5032_));
OAI22X1 OAI22X1_406 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4032_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4216_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3642_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4214_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5036_));
OAI22X1 OAI22X1_407 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3902_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4218_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3967_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4219_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5037_));
OAI22X1 OAI22X1_408 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3183_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4226_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2457_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4224_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5041_));
OAI22X1 OAI22X1_409 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2389_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4229_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2180_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4228_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5042_));
OAI22X1 OAI22X1_41 ( .A(_abc_40298_new_n2481_), .B(_abc_40298_new_n2483_), .C(_abc_40298_new_n1013_), .D(_abc_40298_new_n1941_), .Y(_abc_40298_new_n2484_));
OAI22X1 OAI22X1_410 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2986_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4235_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2918_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4234_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5044_));
OAI22X1 OAI22X1_411 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3446_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4239_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3380_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4240_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5047_));
OAI22X1 OAI22X1_412 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3772_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4243_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3707_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4242_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5048_));
OAI22X1 OAI22X1_413 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4097_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4247_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4162_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4246_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5050_));
OAI22X1 OAI22X1_414 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2255_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4250_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3837_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4249_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5051_));
OAI22X1 OAI22X1_415 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2525_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4190_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2591_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4187_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5058_));
OAI22X1 OAI22X1_416 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2723_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4198_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2855_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4195_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5060_));
OAI22X1 OAI22X1_417 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3054_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4202_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3120_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4201_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5061_));
OAI22X1 OAI22X1_418 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3513_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4207_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3578_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4206_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5064_));
OAI22X1 OAI22X1_419 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4034_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4216_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3644_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4214_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5068_));
OAI22X1 OAI22X1_42 ( .A(_abc_40298_new_n2488_), .B(_abc_40298_new_n2490_), .C(_abc_40298_new_n1013_), .D(_abc_40298_new_n1965_), .Y(_abc_40298_new_n2491_));
OAI22X1 OAI22X1_420 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3904_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4218_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3969_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4219_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5069_));
OAI22X1 OAI22X1_421 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3185_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4226_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2459_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4224_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5073_));
OAI22X1 OAI22X1_422 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2391_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4229_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2183_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4228_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5074_));
OAI22X1 OAI22X1_423 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2988_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4235_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2920_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4234_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5076_));
OAI22X1 OAI22X1_424 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3448_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4239_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3382_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4240_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5079_));
OAI22X1 OAI22X1_425 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3774_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4243_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3709_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4242_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5080_));
OAI22X1 OAI22X1_426 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4099_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4247_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4164_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4246_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5082_));
OAI22X1 OAI22X1_427 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2257_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4250_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3839_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4249_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5083_));
OAI22X1 OAI22X1_428 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2527_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4190_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2593_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4187_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5090_));
OAI22X1 OAI22X1_429 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2725_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4198_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2857_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4195_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5092_));
OAI22X1 OAI22X1_43 ( .A(_abc_40298_new_n2495_), .B(_abc_40298_new_n2497_), .C(_abc_40298_new_n1013_), .D(_abc_40298_new_n2010_), .Y(_abc_40298_new_n2498_));
OAI22X1 OAI22X1_430 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3056_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4202_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3122_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4201_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5093_));
OAI22X1 OAI22X1_431 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3515_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4207_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3580_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4206_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5096_));
OAI22X1 OAI22X1_432 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4036_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4216_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3646_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4214_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5100_));
OAI22X1 OAI22X1_433 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3906_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4218_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3971_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4219_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5101_));
OAI22X1 OAI22X1_434 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3187_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4226_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2461_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4224_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5105_));
OAI22X1 OAI22X1_435 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2393_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4229_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2186_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4228_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5106_));
OAI22X1 OAI22X1_436 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2990_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4235_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2922_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4234_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5108_));
OAI22X1 OAI22X1_437 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3450_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4239_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3384_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4240_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5111_));
OAI22X1 OAI22X1_438 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3776_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4243_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3711_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4242_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5112_));
OAI22X1 OAI22X1_439 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4101_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4247_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4166_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4246_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5114_));
OAI22X1 OAI22X1_44 ( .A(state_q_5_), .B(_abc_40298_new_n2607_), .C(_abc_40298_new_n2577_), .D(_abc_40298_new_n2616_), .Y(_0mem_dat_o_31_0__0_));
OAI22X1 OAI22X1_440 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2259_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4250_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3841_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4249_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5115_));
OAI22X1 OAI22X1_441 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2529_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4190_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2595_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4187_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5122_));
OAI22X1 OAI22X1_442 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2727_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4198_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2859_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4195_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5124_));
OAI22X1 OAI22X1_443 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3058_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4202_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3124_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4201_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5125_));
OAI22X1 OAI22X1_444 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3517_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4207_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3582_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4206_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5128_));
OAI22X1 OAI22X1_445 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4038_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4216_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3648_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4214_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5132_));
OAI22X1 OAI22X1_446 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3908_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4218_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3973_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4219_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5133_));
OAI22X1 OAI22X1_447 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3189_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4226_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2463_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4224_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5137_));
OAI22X1 OAI22X1_448 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2395_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4229_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2189_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4228_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5138_));
OAI22X1 OAI22X1_449 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2992_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4235_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2924_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4234_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5140_));
OAI22X1 OAI22X1_45 ( .A(state_q_5_), .B(_abc_40298_new_n2618_), .C(_abc_40298_new_n2577_), .D(_abc_40298_new_n2624_), .Y(_0mem_dat_o_31_0__1_));
OAI22X1 OAI22X1_450 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3452_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4239_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3386_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4240_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5143_));
OAI22X1 OAI22X1_451 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3778_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4243_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3713_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4242_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5144_));
OAI22X1 OAI22X1_452 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4103_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4247_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4168_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4246_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5146_));
OAI22X1 OAI22X1_453 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2261_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4250_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3843_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4249_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5147_));
OAI22X1 OAI22X1_454 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2531_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4190_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2597_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4187_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5154_));
OAI22X1 OAI22X1_455 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2729_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4198_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2861_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4195_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5156_));
OAI22X1 OAI22X1_456 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3060_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4202_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3126_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4201_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5157_));
OAI22X1 OAI22X1_457 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3519_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4207_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3584_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4206_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5160_));
OAI22X1 OAI22X1_458 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4040_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4216_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3650_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4214_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5164_));
OAI22X1 OAI22X1_459 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3910_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4218_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3975_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4219_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5165_));
OAI22X1 OAI22X1_46 ( .A(state_q_5_), .B(_abc_40298_new_n2626_), .C(_abc_40298_new_n2577_), .D(_abc_40298_new_n2632_), .Y(_0mem_dat_o_31_0__2_));
OAI22X1 OAI22X1_460 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3191_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4226_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2465_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4224_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5169_));
OAI22X1 OAI22X1_461 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2397_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4229_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2192_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4228_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5170_));
OAI22X1 OAI22X1_462 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2994_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4235_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2926_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4234_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5172_));
OAI22X1 OAI22X1_463 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3454_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4239_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3388_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4240_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5175_));
OAI22X1 OAI22X1_464 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3780_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4243_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3715_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4242_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5176_));
OAI22X1 OAI22X1_465 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4105_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4247_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4170_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4246_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5178_));
OAI22X1 OAI22X1_466 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2263_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4250_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3845_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4249_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5179_));
OAI22X1 OAI22X1_467 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2533_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4190_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2599_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4187_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5186_));
OAI22X1 OAI22X1_468 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2731_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4198_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2863_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4195_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5188_));
OAI22X1 OAI22X1_469 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3062_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4202_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3128_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4201_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5189_));
OAI22X1 OAI22X1_47 ( .A(state_q_5_), .B(_abc_40298_new_n2634_), .C(_abc_40298_new_n2577_), .D(_abc_40298_new_n2640_), .Y(_0mem_dat_o_31_0__3_));
OAI22X1 OAI22X1_470 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3521_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4207_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3586_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4206_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5192_));
OAI22X1 OAI22X1_471 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4042_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4216_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3652_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4214_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5196_));
OAI22X1 OAI22X1_472 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3912_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4218_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3977_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4219_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5197_));
OAI22X1 OAI22X1_473 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3193_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4226_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2467_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4224_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5201_));
OAI22X1 OAI22X1_474 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2399_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4229_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2195_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4228_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5202_));
OAI22X1 OAI22X1_475 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2996_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4235_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2928_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4234_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5204_));
OAI22X1 OAI22X1_476 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3456_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4239_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3390_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4240_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5207_));
OAI22X1 OAI22X1_477 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3782_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4243_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3717_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4242_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5208_));
OAI22X1 OAI22X1_478 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4107_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4247_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4172_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4246_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5210_));
OAI22X1 OAI22X1_479 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2265_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4250_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3847_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4249_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5211_));
OAI22X1 OAI22X1_48 ( .A(state_q_5_), .B(_abc_40298_new_n2642_), .C(_abc_40298_new_n2577_), .D(_abc_40298_new_n2648_), .Y(_0mem_dat_o_31_0__4_));
OAI22X1 OAI22X1_480 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2535_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4190_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2601_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4187_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5218_));
OAI22X1 OAI22X1_481 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2733_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4198_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2865_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4195_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5220_));
OAI22X1 OAI22X1_482 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3064_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4202_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3130_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4201_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5221_));
OAI22X1 OAI22X1_483 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3523_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4207_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3588_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4206_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5224_));
OAI22X1 OAI22X1_484 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4044_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4216_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3654_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4214_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5228_));
OAI22X1 OAI22X1_485 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3914_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4218_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3979_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4219_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5229_));
OAI22X1 OAI22X1_486 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3195_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4226_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2469_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4224_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5233_));
OAI22X1 OAI22X1_487 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2401_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4229_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2198_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4228_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5234_));
OAI22X1 OAI22X1_488 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2998_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4235_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2930_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4234_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5236_));
OAI22X1 OAI22X1_489 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3458_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4239_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3392_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4240_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5239_));
OAI22X1 OAI22X1_49 ( .A(state_q_5_), .B(_abc_40298_new_n2650_), .C(_abc_40298_new_n2577_), .D(_abc_40298_new_n2656_), .Y(_0mem_dat_o_31_0__5_));
OAI22X1 OAI22X1_490 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3784_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4243_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3719_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4242_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5240_));
OAI22X1 OAI22X1_491 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4109_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4247_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4174_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4246_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5242_));
OAI22X1 OAI22X1_492 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2267_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4250_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3849_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4249_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5243_));
OAI22X1 OAI22X1_493 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2471_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5262_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2537_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5259_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5263_));
OAI22X1 OAI22X1_494 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2668_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5270_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2801_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5267_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5271_));
OAI22X1 OAI22X1_495 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3000_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5274_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3066_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5273_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5275_));
OAI22X1 OAI22X1_496 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3460_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5279_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3525_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5278_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5280_));
OAI22X1 OAI22X1_497 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3981_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5288_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3590_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5286_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5289_));
OAI22X1 OAI22X1_498 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3851_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5290_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3916_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5291_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5292_));
OAI22X1 OAI22X1_499 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3132_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5298_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2403_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5296_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5299_));
OAI22X1 OAI22X1_5 ( .A(_abc_40298_new_n771_), .B(_abc_40298_new_n795_), .C(_abc_40298_new_n794_), .D(_abc_40298_new_n695_), .Y(_abc_40298_new_n796_));
OAI22X1 OAI22X1_50 ( .A(state_q_5_), .B(_abc_40298_new_n2658_), .C(_abc_40298_new_n2577_), .D(_abc_40298_new_n2664_), .Y(_0mem_dat_o_31_0__6_));
OAI22X1 OAI22X1_500 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2336_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5301_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2099_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5300_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5302_));
OAI22X1 OAI22X1_501 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2932_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5307_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2867_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5306_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5308_));
OAI22X1 OAI22X1_502 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3394_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5311_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3329_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5312_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5313_));
OAI22X1 OAI22X1_503 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3721_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5315_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3656_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5314_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5316_));
OAI22X1 OAI22X1_504 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4046_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5319_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4111_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5318_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5320_));
OAI22X1 OAI22X1_505 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2201_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5322_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3786_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5321_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5323_));
OAI22X1 OAI22X1_506 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2475_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5262_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2541_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5259_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5330_));
OAI22X1 OAI22X1_507 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2673_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5270_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2805_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5267_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5332_));
OAI22X1 OAI22X1_508 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3004_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5274_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3070_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5273_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5333_));
OAI22X1 OAI22X1_509 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3463_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5279_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3528_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5278_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5336_));
OAI22X1 OAI22X1_51 ( .A(state_q_5_), .B(_abc_40298_new_n2666_), .C(_abc_40298_new_n2577_), .D(_abc_40298_new_n2672_), .Y(_0mem_dat_o_31_0__7_));
OAI22X1 OAI22X1_510 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3984_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5288_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3594_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5286_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5340_));
OAI22X1 OAI22X1_511 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3854_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5290_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3919_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5291_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5341_));
OAI22X1 OAI22X1_512 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3135_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5298_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2409_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5296_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5345_));
OAI22X1 OAI22X1_513 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2341_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5301_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2108_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5300_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5346_));
OAI22X1 OAI22X1_514 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2938_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5307_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2870_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5306_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5348_));
OAI22X1 OAI22X1_515 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3398_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5311_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3332_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5312_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5351_));
OAI22X1 OAI22X1_516 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3724_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5315_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3659_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5314_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5352_));
OAI22X1 OAI22X1_517 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4049_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5319_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4114_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5318_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5354_));
OAI22X1 OAI22X1_518 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2207_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5322_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3789_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5321_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5355_));
OAI22X1 OAI22X1_519 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2477_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5262_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2543_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5259_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5362_));
OAI22X1 OAI22X1_52 ( .A(state_q_5_), .B(_abc_40298_new_n2674_), .C(_abc_40298_new_n2681_), .D(_abc_40298_new_n2679_), .Y(_0mem_dat_o_31_0__8_));
OAI22X1 OAI22X1_520 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2675_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5270_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2807_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5267_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5364_));
OAI22X1 OAI22X1_521 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3006_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5274_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3072_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5273_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5365_));
OAI22X1 OAI22X1_522 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3465_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5279_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3530_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5278_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5368_));
OAI22X1 OAI22X1_523 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3986_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5288_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3596_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5286_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5372_));
OAI22X1 OAI22X1_524 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3856_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5290_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3921_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5291_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5373_));
OAI22X1 OAI22X1_525 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3137_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5298_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2411_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5296_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5377_));
OAI22X1 OAI22X1_526 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2343_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5301_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2111_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5300_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5378_));
OAI22X1 OAI22X1_527 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2940_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5307_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2872_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5306_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5380_));
OAI22X1 OAI22X1_528 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3400_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5311_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3334_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5312_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5383_));
OAI22X1 OAI22X1_529 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3726_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5315_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3661_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5314_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5384_));
OAI22X1 OAI22X1_53 ( .A(state_q_5_), .B(_abc_40298_new_n2683_), .C(_abc_40298_new_n2690_), .D(_abc_40298_new_n2688_), .Y(_0mem_dat_o_31_0__9_));
OAI22X1 OAI22X1_530 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4051_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5319_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4116_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5318_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5386_));
OAI22X1 OAI22X1_531 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2209_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5322_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3791_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5321_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5387_));
OAI22X1 OAI22X1_532 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2479_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5262_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2545_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5259_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5394_));
OAI22X1 OAI22X1_533 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2677_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5270_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2809_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5267_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5396_));
OAI22X1 OAI22X1_534 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3008_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5274_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3074_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5273_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5397_));
OAI22X1 OAI22X1_535 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3467_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5279_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3532_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5278_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5400_));
OAI22X1 OAI22X1_536 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3988_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5288_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3598_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5286_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5404_));
OAI22X1 OAI22X1_537 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3858_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5290_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3923_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5291_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5405_));
OAI22X1 OAI22X1_538 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3139_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5298_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2413_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5296_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5409_));
OAI22X1 OAI22X1_539 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2345_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5301_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2114_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5300_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5410_));
OAI22X1 OAI22X1_54 ( .A(state_q_5_), .B(_abc_40298_new_n2692_), .C(_abc_40298_new_n2699_), .D(_abc_40298_new_n2697_), .Y(_0mem_dat_o_31_0__10_));
OAI22X1 OAI22X1_540 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2942_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5307_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2874_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5306_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5412_));
OAI22X1 OAI22X1_541 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3402_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5311_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3336_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5312_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5415_));
OAI22X1 OAI22X1_542 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3728_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5315_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3663_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5314_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5416_));
OAI22X1 OAI22X1_543 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4053_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5319_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4118_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5318_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5418_));
OAI22X1 OAI22X1_544 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2211_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5322_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3793_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5321_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5419_));
OAI22X1 OAI22X1_545 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2481_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5262_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2547_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5259_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5426_));
OAI22X1 OAI22X1_546 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2679_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5270_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2811_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5267_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5428_));
OAI22X1 OAI22X1_547 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3010_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5274_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3076_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5273_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5429_));
OAI22X1 OAI22X1_548 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3469_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5279_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3534_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5278_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5432_));
OAI22X1 OAI22X1_549 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3990_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5288_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3600_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5286_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5436_));
OAI22X1 OAI22X1_55 ( .A(state_q_5_), .B(_abc_40298_new_n2701_), .C(_abc_40298_new_n2708_), .D(_abc_40298_new_n2706_), .Y(_0mem_dat_o_31_0__11_));
OAI22X1 OAI22X1_550 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3860_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5290_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3925_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5291_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5437_));
OAI22X1 OAI22X1_551 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3141_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5298_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2415_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5296_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5441_));
OAI22X1 OAI22X1_552 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2347_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5301_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2117_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5300_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5442_));
OAI22X1 OAI22X1_553 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2944_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5307_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2876_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5306_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5444_));
OAI22X1 OAI22X1_554 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3404_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5311_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3338_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5312_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5447_));
OAI22X1 OAI22X1_555 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3730_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5315_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3665_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5314_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5448_));
OAI22X1 OAI22X1_556 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4055_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5319_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4120_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5318_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5450_));
OAI22X1 OAI22X1_557 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2213_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5322_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3795_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5321_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5451_));
OAI22X1 OAI22X1_558 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2483_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5262_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2549_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5259_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5458_));
OAI22X1 OAI22X1_559 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2681_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5270_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2813_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5267_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5460_));
OAI22X1 OAI22X1_56 ( .A(state_q_5_), .B(_abc_40298_new_n2710_), .C(_abc_40298_new_n2717_), .D(_abc_40298_new_n2715_), .Y(_0mem_dat_o_31_0__12_));
OAI22X1 OAI22X1_560 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3012_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5274_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3078_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5273_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5461_));
OAI22X1 OAI22X1_561 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3471_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5279_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3536_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5278_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5464_));
OAI22X1 OAI22X1_562 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3992_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5288_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3602_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5286_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5468_));
OAI22X1 OAI22X1_563 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3862_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5290_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3927_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5291_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5469_));
OAI22X1 OAI22X1_564 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3143_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5298_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2417_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5296_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5473_));
OAI22X1 OAI22X1_565 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2349_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5301_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2120_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5300_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5474_));
OAI22X1 OAI22X1_566 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2946_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5307_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2878_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5306_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5476_));
OAI22X1 OAI22X1_567 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3406_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5311_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3340_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5312_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5479_));
OAI22X1 OAI22X1_568 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3732_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5315_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3667_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5314_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5480_));
OAI22X1 OAI22X1_569 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4057_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5319_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4122_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5318_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5482_));
OAI22X1 OAI22X1_57 ( .A(state_q_5_), .B(_abc_40298_new_n2719_), .C(_abc_40298_new_n2726_), .D(_abc_40298_new_n2724_), .Y(_0mem_dat_o_31_0__13_));
OAI22X1 OAI22X1_570 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2215_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5322_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3797_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5321_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5483_));
OAI22X1 OAI22X1_571 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2485_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5262_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2551_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5259_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5490_));
OAI22X1 OAI22X1_572 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2683_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5270_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2815_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5267_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5492_));
OAI22X1 OAI22X1_573 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3014_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5274_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3080_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5273_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5493_));
OAI22X1 OAI22X1_574 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3473_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5279_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3538_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5278_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5496_));
OAI22X1 OAI22X1_575 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3994_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5288_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3604_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5286_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5500_));
OAI22X1 OAI22X1_576 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3864_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5290_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3929_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5291_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5501_));
OAI22X1 OAI22X1_577 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3145_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5298_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2419_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5296_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5505_));
OAI22X1 OAI22X1_578 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2351_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5301_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2123_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5300_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5506_));
OAI22X1 OAI22X1_579 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2948_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5307_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2880_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5306_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5508_));
OAI22X1 OAI22X1_58 ( .A(state_q_5_), .B(_abc_40298_new_n2728_), .C(_abc_40298_new_n2735_), .D(_abc_40298_new_n2733_), .Y(_0mem_dat_o_31_0__14_));
OAI22X1 OAI22X1_580 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3408_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5311_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3342_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5312_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5511_));
OAI22X1 OAI22X1_581 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3734_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5315_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3669_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5314_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5512_));
OAI22X1 OAI22X1_582 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4059_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5319_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4124_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5318_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5514_));
OAI22X1 OAI22X1_583 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2217_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5322_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3799_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5321_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5515_));
OAI22X1 OAI22X1_584 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2487_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5262_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2553_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5259_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5522_));
OAI22X1 OAI22X1_585 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2685_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5270_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2817_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5267_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5524_));
OAI22X1 OAI22X1_586 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3016_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5274_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3082_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5273_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5525_));
OAI22X1 OAI22X1_587 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3475_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5279_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3540_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5278_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5528_));
OAI22X1 OAI22X1_588 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3996_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5288_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3606_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5286_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5532_));
OAI22X1 OAI22X1_589 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3866_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5290_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3931_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5291_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5533_));
OAI22X1 OAI22X1_59 ( .A(state_q_5_), .B(_abc_40298_new_n2737_), .C(_abc_40298_new_n2744_), .D(_abc_40298_new_n2742_), .Y(_0mem_dat_o_31_0__15_));
OAI22X1 OAI22X1_590 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3147_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5298_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2421_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5296_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5537_));
OAI22X1 OAI22X1_591 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2353_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5301_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2126_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5300_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5538_));
OAI22X1 OAI22X1_592 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2950_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5307_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2882_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5306_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5540_));
OAI22X1 OAI22X1_593 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3410_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5311_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3344_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5312_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5543_));
OAI22X1 OAI22X1_594 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3736_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5315_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3671_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5314_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5544_));
OAI22X1 OAI22X1_595 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4061_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5319_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4126_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5318_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5546_));
OAI22X1 OAI22X1_596 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2219_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5322_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3801_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5321_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5547_));
OAI22X1 OAI22X1_597 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2489_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5262_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2555_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5259_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5554_));
OAI22X1 OAI22X1_598 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2687_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5270_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2819_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5267_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5556_));
OAI22X1 OAI22X1_599 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3018_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5274_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3084_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5273_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5557_));
OAI22X1 OAI22X1_6 ( .A(_abc_40298_new_n1089_), .B(_abc_40298_new_n1209_), .C(_abc_40298_new_n984_), .D(_abc_40298_new_n1210_), .Y(_abc_40298_new_n1211_));
OAI22X1 OAI22X1_60 ( .A(state_q_5_), .B(_abc_40298_new_n2746_), .C(_abc_40298_new_n2577_), .D(_abc_40298_new_n2752_), .Y(_0mem_dat_o_31_0__16_));
OAI22X1 OAI22X1_600 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3477_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5279_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3542_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5278_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5560_));
OAI22X1 OAI22X1_601 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3998_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5288_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3608_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5286_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5564_));
OAI22X1 OAI22X1_602 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3868_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5290_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3933_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5291_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5565_));
OAI22X1 OAI22X1_603 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3149_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5298_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2423_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5296_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5569_));
OAI22X1 OAI22X1_604 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2355_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5301_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2129_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5300_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5570_));
OAI22X1 OAI22X1_605 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2952_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5307_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2884_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5306_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5572_));
OAI22X1 OAI22X1_606 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3412_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5311_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3346_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5312_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5575_));
OAI22X1 OAI22X1_607 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3738_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5315_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3673_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5314_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5576_));
OAI22X1 OAI22X1_608 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4063_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5319_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4128_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5318_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5578_));
OAI22X1 OAI22X1_609 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2221_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5322_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3803_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5321_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5579_));
OAI22X1 OAI22X1_61 ( .A(state_q_5_), .B(_abc_40298_new_n2754_), .C(_abc_40298_new_n2577_), .D(_abc_40298_new_n2760_), .Y(_0mem_dat_o_31_0__17_));
OAI22X1 OAI22X1_610 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2491_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5262_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2557_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5259_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5586_));
OAI22X1 OAI22X1_611 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2689_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5270_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2821_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5267_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5588_));
OAI22X1 OAI22X1_612 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3020_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5274_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3086_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5273_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5589_));
OAI22X1 OAI22X1_613 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3479_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5279_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3544_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5278_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5592_));
OAI22X1 OAI22X1_614 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4000_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5288_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3610_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5286_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5596_));
OAI22X1 OAI22X1_615 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3870_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5290_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3935_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5291_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5597_));
OAI22X1 OAI22X1_616 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3151_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5298_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2425_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5296_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5601_));
OAI22X1 OAI22X1_617 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2357_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5301_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2132_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5300_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5602_));
OAI22X1 OAI22X1_618 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2954_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5307_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2886_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5306_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5604_));
OAI22X1 OAI22X1_619 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3414_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5311_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3348_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5312_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5607_));
OAI22X1 OAI22X1_62 ( .A(state_q_5_), .B(_abc_40298_new_n2762_), .C(_abc_40298_new_n2577_), .D(_abc_40298_new_n2768_), .Y(_0mem_dat_o_31_0__18_));
OAI22X1 OAI22X1_620 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3740_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5315_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3675_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5314_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5608_));
OAI22X1 OAI22X1_621 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4065_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5319_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4130_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5318_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5610_));
OAI22X1 OAI22X1_622 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2223_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5322_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3805_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5321_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5611_));
OAI22X1 OAI22X1_623 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2493_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5262_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2559_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5259_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5618_));
OAI22X1 OAI22X1_624 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2691_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5270_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2823_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5267_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5620_));
OAI22X1 OAI22X1_625 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3022_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5274_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3088_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5273_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5621_));
OAI22X1 OAI22X1_626 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3481_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5279_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3546_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5278_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5624_));
OAI22X1 OAI22X1_627 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4002_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5288_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3612_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5286_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5628_));
OAI22X1 OAI22X1_628 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3872_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5290_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3937_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5291_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5629_));
OAI22X1 OAI22X1_629 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3153_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5298_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2427_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5296_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5633_));
OAI22X1 OAI22X1_63 ( .A(state_q_5_), .B(_abc_40298_new_n2770_), .C(_abc_40298_new_n2577_), .D(_abc_40298_new_n2776_), .Y(_0mem_dat_o_31_0__19_));
OAI22X1 OAI22X1_630 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2359_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5301_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2135_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5300_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5634_));
OAI22X1 OAI22X1_631 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2956_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5307_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2888_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5306_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5636_));
OAI22X1 OAI22X1_632 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3416_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5311_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3350_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5312_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5639_));
OAI22X1 OAI22X1_633 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3742_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5315_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3677_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5314_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5640_));
OAI22X1 OAI22X1_634 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4067_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5319_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4132_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5318_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5642_));
OAI22X1 OAI22X1_635 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2225_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5322_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3807_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5321_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5643_));
OAI22X1 OAI22X1_636 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2495_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5262_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2561_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5259_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5650_));
OAI22X1 OAI22X1_637 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2693_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5270_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2825_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5267_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5652_));
OAI22X1 OAI22X1_638 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3024_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5274_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3090_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5273_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5653_));
OAI22X1 OAI22X1_639 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3483_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5279_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3548_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5278_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5656_));
OAI22X1 OAI22X1_64 ( .A(state_q_5_), .B(_abc_40298_new_n2778_), .C(_abc_40298_new_n2577_), .D(_abc_40298_new_n2784_), .Y(_0mem_dat_o_31_0__20_));
OAI22X1 OAI22X1_640 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4004_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5288_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3614_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5286_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5660_));
OAI22X1 OAI22X1_641 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3874_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5290_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3939_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5291_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5661_));
OAI22X1 OAI22X1_642 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3155_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5298_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2429_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5296_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5665_));
OAI22X1 OAI22X1_643 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2361_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5301_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2138_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5300_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5666_));
OAI22X1 OAI22X1_644 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2958_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5307_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2890_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5306_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5668_));
OAI22X1 OAI22X1_645 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3418_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5311_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3352_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5312_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5671_));
OAI22X1 OAI22X1_646 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3744_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5315_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3679_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5314_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5672_));
OAI22X1 OAI22X1_647 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4069_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5319_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4134_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5318_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5674_));
OAI22X1 OAI22X1_648 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2227_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5322_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3809_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5321_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5675_));
OAI22X1 OAI22X1_649 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2497_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5262_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2563_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5259_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5682_));
OAI22X1 OAI22X1_65 ( .A(state_q_5_), .B(_abc_40298_new_n2786_), .C(_abc_40298_new_n2577_), .D(_abc_40298_new_n2792_), .Y(_0mem_dat_o_31_0__21_));
OAI22X1 OAI22X1_650 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2695_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5270_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2827_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5267_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5684_));
OAI22X1 OAI22X1_651 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3026_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5274_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3092_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5273_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5685_));
OAI22X1 OAI22X1_652 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3485_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5279_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3550_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5278_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5688_));
OAI22X1 OAI22X1_653 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4006_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5288_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3616_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5286_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5692_));
OAI22X1 OAI22X1_654 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3876_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5290_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3941_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5291_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5693_));
OAI22X1 OAI22X1_655 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3157_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5298_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2431_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5296_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5697_));
OAI22X1 OAI22X1_656 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2363_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5301_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2141_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5300_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5698_));
OAI22X1 OAI22X1_657 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2960_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5307_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2892_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5306_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5700_));
OAI22X1 OAI22X1_658 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3420_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5311_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3354_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5312_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5703_));
OAI22X1 OAI22X1_659 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3746_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5315_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3681_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5314_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5704_));
OAI22X1 OAI22X1_66 ( .A(state_q_5_), .B(_abc_40298_new_n2794_), .C(_abc_40298_new_n2577_), .D(_abc_40298_new_n2800_), .Y(_0mem_dat_o_31_0__22_));
OAI22X1 OAI22X1_660 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4071_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5319_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4136_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5318_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5706_));
OAI22X1 OAI22X1_661 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2229_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5322_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3811_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5321_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5707_));
OAI22X1 OAI22X1_662 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2499_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5262_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2565_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5259_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5714_));
OAI22X1 OAI22X1_663 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2697_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5270_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2829_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5267_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5716_));
OAI22X1 OAI22X1_664 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3028_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5274_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3094_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5273_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5717_));
OAI22X1 OAI22X1_665 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3487_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5279_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3552_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5278_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5720_));
OAI22X1 OAI22X1_666 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4008_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5288_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3618_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5286_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5724_));
OAI22X1 OAI22X1_667 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3878_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5290_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3943_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5291_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5725_));
OAI22X1 OAI22X1_668 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3159_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5298_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2433_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5296_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5729_));
OAI22X1 OAI22X1_669 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2365_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5301_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2144_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5300_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5730_));
OAI22X1 OAI22X1_67 ( .A(state_q_5_), .B(_abc_40298_new_n2802_), .C(_abc_40298_new_n2577_), .D(_abc_40298_new_n2808_), .Y(_0mem_dat_o_31_0__23_));
OAI22X1 OAI22X1_670 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2962_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5307_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2894_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5306_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5732_));
OAI22X1 OAI22X1_671 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3422_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5311_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3356_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5312_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5735_));
OAI22X1 OAI22X1_672 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3748_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5315_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3683_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5314_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5736_));
OAI22X1 OAI22X1_673 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4073_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5319_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4138_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5318_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5738_));
OAI22X1 OAI22X1_674 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2231_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5322_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3813_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5321_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5739_));
OAI22X1 OAI22X1_675 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2501_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5262_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2567_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5259_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5746_));
OAI22X1 OAI22X1_676 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2699_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5270_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2831_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5267_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5748_));
OAI22X1 OAI22X1_677 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3030_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5274_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3096_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5273_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5749_));
OAI22X1 OAI22X1_678 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3489_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5279_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3554_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5278_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5752_));
OAI22X1 OAI22X1_679 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4010_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5288_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3620_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5286_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5756_));
OAI22X1 OAI22X1_68 ( .A(state_q_5_), .B(_abc_40298_new_n2810_), .C(_abc_40298_new_n2817_), .D(_abc_40298_new_n2815_), .Y(_0mem_dat_o_31_0__24_));
OAI22X1 OAI22X1_680 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3880_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5290_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3945_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5291_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5757_));
OAI22X1 OAI22X1_681 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3161_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5298_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2435_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5296_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5761_));
OAI22X1 OAI22X1_682 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2367_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5301_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2147_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5300_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5762_));
OAI22X1 OAI22X1_683 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2964_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5307_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2896_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5306_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5764_));
OAI22X1 OAI22X1_684 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3424_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5311_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3358_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5312_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5767_));
OAI22X1 OAI22X1_685 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3750_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5315_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3685_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5314_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5768_));
OAI22X1 OAI22X1_686 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4075_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5319_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4140_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5318_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5770_));
OAI22X1 OAI22X1_687 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2233_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5322_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3815_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5321_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5771_));
OAI22X1 OAI22X1_688 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2503_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5262_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2569_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5259_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5778_));
OAI22X1 OAI22X1_689 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2701_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5270_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2833_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5267_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5780_));
OAI22X1 OAI22X1_69 ( .A(state_q_5_), .B(_abc_40298_new_n2819_), .C(_abc_40298_new_n2826_), .D(_abc_40298_new_n2824_), .Y(_0mem_dat_o_31_0__25_));
OAI22X1 OAI22X1_690 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3032_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5274_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3098_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5273_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5781_));
OAI22X1 OAI22X1_691 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3491_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5279_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3556_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5278_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5784_));
OAI22X1 OAI22X1_692 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4012_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5288_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3622_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5286_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5788_));
OAI22X1 OAI22X1_693 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3882_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5290_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3947_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5291_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5789_));
OAI22X1 OAI22X1_694 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3163_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5298_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2437_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5296_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5793_));
OAI22X1 OAI22X1_695 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2369_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5301_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2150_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5300_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5794_));
OAI22X1 OAI22X1_696 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2966_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5307_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2898_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5306_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5796_));
OAI22X1 OAI22X1_697 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3426_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5311_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3360_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5312_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5799_));
OAI22X1 OAI22X1_698 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3752_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5315_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3687_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5314_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5800_));
OAI22X1 OAI22X1_699 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4077_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5319_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4142_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5318_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5802_));
OAI22X1 OAI22X1_7 ( .A(_abc_40298_new_n1339_), .B(_abc_40298_new_n1066_), .C(_abc_40298_new_n1352_), .D(_abc_40298_new_n1347_), .Y(_abc_40298_new_n1353_));
OAI22X1 OAI22X1_70 ( .A(state_q_5_), .B(_abc_40298_new_n2828_), .C(_abc_40298_new_n2835_), .D(_abc_40298_new_n2833_), .Y(_0mem_dat_o_31_0__26_));
OAI22X1 OAI22X1_700 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2235_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5322_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3817_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5321_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5803_));
OAI22X1 OAI22X1_701 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2505_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5262_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2571_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5259_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5810_));
OAI22X1 OAI22X1_702 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2703_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5270_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2835_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5267_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5812_));
OAI22X1 OAI22X1_703 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3034_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5274_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3100_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5273_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5813_));
OAI22X1 OAI22X1_704 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3493_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5279_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3558_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5278_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5816_));
OAI22X1 OAI22X1_705 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4014_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5288_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3624_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5286_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5820_));
OAI22X1 OAI22X1_706 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3884_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5290_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3949_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5291_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5821_));
OAI22X1 OAI22X1_707 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3165_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5298_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2439_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5296_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5825_));
OAI22X1 OAI22X1_708 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2371_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5301_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2153_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5300_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5826_));
OAI22X1 OAI22X1_709 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2968_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5307_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2900_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5306_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5828_));
OAI22X1 OAI22X1_71 ( .A(state_q_5_), .B(_abc_40298_new_n2837_), .C(_abc_40298_new_n2844_), .D(_abc_40298_new_n2842_), .Y(_0mem_dat_o_31_0__27_));
OAI22X1 OAI22X1_710 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3428_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5311_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3362_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5312_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5831_));
OAI22X1 OAI22X1_711 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3754_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5315_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3689_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5314_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5832_));
OAI22X1 OAI22X1_712 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4079_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5319_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4144_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5318_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5834_));
OAI22X1 OAI22X1_713 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2237_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5322_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3819_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5321_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5835_));
OAI22X1 OAI22X1_714 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2507_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5262_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2573_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5259_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5842_));
OAI22X1 OAI22X1_715 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2705_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5270_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2837_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5267_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5844_));
OAI22X1 OAI22X1_716 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3036_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5274_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3102_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5273_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5845_));
OAI22X1 OAI22X1_717 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3495_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5279_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3560_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5278_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5848_));
OAI22X1 OAI22X1_718 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4016_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5288_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3626_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5286_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5852_));
OAI22X1 OAI22X1_719 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3886_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5290_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3951_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5291_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5853_));
OAI22X1 OAI22X1_72 ( .A(state_q_5_), .B(_abc_40298_new_n2846_), .C(_abc_40298_new_n2853_), .D(_abc_40298_new_n2851_), .Y(_0mem_dat_o_31_0__28_));
OAI22X1 OAI22X1_720 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3167_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5298_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2441_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5296_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5857_));
OAI22X1 OAI22X1_721 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2373_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5301_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2156_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5300_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5858_));
OAI22X1 OAI22X1_722 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2970_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5307_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2902_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5306_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5860_));
OAI22X1 OAI22X1_723 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3430_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5311_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3364_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5312_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5863_));
OAI22X1 OAI22X1_724 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3756_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5315_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3691_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5314_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5864_));
OAI22X1 OAI22X1_725 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4081_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5319_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4146_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5318_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5866_));
OAI22X1 OAI22X1_726 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2239_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5322_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3821_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5321_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5867_));
OAI22X1 OAI22X1_727 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2509_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5262_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2575_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5259_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5874_));
OAI22X1 OAI22X1_728 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2707_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5270_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2839_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5267_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5876_));
OAI22X1 OAI22X1_729 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3038_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5274_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3104_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5273_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5877_));
OAI22X1 OAI22X1_73 ( .A(state_q_5_), .B(_abc_40298_new_n2855_), .C(_abc_40298_new_n2862_), .D(_abc_40298_new_n2860_), .Y(_0mem_dat_o_31_0__29_));
OAI22X1 OAI22X1_730 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3497_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5279_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3562_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5278_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5880_));
OAI22X1 OAI22X1_731 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4018_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5288_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3628_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5286_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5884_));
OAI22X1 OAI22X1_732 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3888_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5290_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3953_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5291_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5885_));
OAI22X1 OAI22X1_733 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3169_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5298_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2443_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5296_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5889_));
OAI22X1 OAI22X1_734 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2375_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5301_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2159_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5300_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5890_));
OAI22X1 OAI22X1_735 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2972_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5307_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2904_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5306_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5892_));
OAI22X1 OAI22X1_736 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3432_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5311_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3366_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5312_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5895_));
OAI22X1 OAI22X1_737 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3758_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5315_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3693_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5314_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5896_));
OAI22X1 OAI22X1_738 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4083_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5319_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4148_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5318_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5898_));
OAI22X1 OAI22X1_739 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2241_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5322_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3823_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5321_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5899_));
OAI22X1 OAI22X1_74 ( .A(state_q_5_), .B(_abc_40298_new_n2864_), .C(_abc_40298_new_n2871_), .D(_abc_40298_new_n2869_), .Y(_0mem_dat_o_31_0__30_));
OAI22X1 OAI22X1_740 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2511_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5262_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2577_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5259_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5906_));
OAI22X1 OAI22X1_741 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2709_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5270_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2841_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5267_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5908_));
OAI22X1 OAI22X1_742 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3040_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5274_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3106_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5273_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5909_));
OAI22X1 OAI22X1_743 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3499_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5279_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3564_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5278_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5912_));
OAI22X1 OAI22X1_744 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4020_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5288_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3630_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5286_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5916_));
OAI22X1 OAI22X1_745 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3890_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5290_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3955_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5291_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5917_));
OAI22X1 OAI22X1_746 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3171_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5298_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2445_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5296_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5921_));
OAI22X1 OAI22X1_747 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2377_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5301_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2162_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5300_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5922_));
OAI22X1 OAI22X1_748 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2974_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5307_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2906_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5306_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5924_));
OAI22X1 OAI22X1_749 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3434_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5311_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3368_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5312_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5927_));
OAI22X1 OAI22X1_75 ( .A(state_q_5_), .B(_abc_40298_new_n2873_), .C(_abc_40298_new_n2880_), .D(_abc_40298_new_n2878_), .Y(_0mem_dat_o_31_0__31_));
OAI22X1 OAI22X1_750 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3760_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5315_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3695_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5314_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5928_));
OAI22X1 OAI22X1_751 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4085_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5319_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4150_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5318_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5930_));
OAI22X1 OAI22X1_752 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2243_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5322_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3825_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5321_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5931_));
OAI22X1 OAI22X1_753 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2513_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5262_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2579_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5259_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5938_));
OAI22X1 OAI22X1_754 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2711_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5270_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2843_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5267_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5940_));
OAI22X1 OAI22X1_755 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3042_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5274_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3108_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5273_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5941_));
OAI22X1 OAI22X1_756 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3501_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5279_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3566_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5278_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5944_));
OAI22X1 OAI22X1_757 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4022_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5288_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3632_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5286_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5948_));
OAI22X1 OAI22X1_758 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3892_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5290_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3957_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5291_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5949_));
OAI22X1 OAI22X1_759 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3173_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5298_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2447_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5296_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5953_));
OAI22X1 OAI22X1_76 ( .A(_abc_40298_new_n2455_), .B(_abc_40298_new_n3039_), .C(_abc_40298_new_n3147_), .D(_abc_40298_new_n3161_), .Y(_abc_40298_new_n3163_));
OAI22X1 OAI22X1_760 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2379_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5301_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2165_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5300_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5954_));
OAI22X1 OAI22X1_761 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2976_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5307_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2908_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5306_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5956_));
OAI22X1 OAI22X1_762 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3436_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5311_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3370_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5312_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5959_));
OAI22X1 OAI22X1_763 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3762_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5315_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3697_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5314_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5960_));
OAI22X1 OAI22X1_764 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4087_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5319_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4152_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5318_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5962_));
OAI22X1 OAI22X1_765 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2245_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5322_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3827_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5321_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5963_));
OAI22X1 OAI22X1_766 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2515_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5262_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2581_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5259_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5970_));
OAI22X1 OAI22X1_767 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2713_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5270_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2845_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5267_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5972_));
OAI22X1 OAI22X1_768 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3044_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5274_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3110_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5273_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5973_));
OAI22X1 OAI22X1_769 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3503_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5279_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3568_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5278_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5976_));
OAI22X1 OAI22X1_77 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2471_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4190_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2537_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4187_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4191_));
OAI22X1 OAI22X1_770 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4024_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5288_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3634_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5286_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5980_));
OAI22X1 OAI22X1_771 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3894_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5290_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3959_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5291_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5981_));
OAI22X1 OAI22X1_772 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3175_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5298_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2449_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5296_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5985_));
OAI22X1 OAI22X1_773 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2381_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5301_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2168_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5300_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5986_));
OAI22X1 OAI22X1_774 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2978_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5307_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2910_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5306_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5988_));
OAI22X1 OAI22X1_775 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3438_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5311_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3372_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5312_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5991_));
OAI22X1 OAI22X1_776 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3764_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5315_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3699_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5314_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5992_));
OAI22X1 OAI22X1_777 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4089_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5319_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4154_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5318_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5994_));
OAI22X1 OAI22X1_778 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2247_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5322_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3829_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5321_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n5995_));
OAI22X1 OAI22X1_779 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2517_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5262_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2583_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5259_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6002_));
OAI22X1 OAI22X1_78 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2668_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4198_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2801_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4195_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4199_));
OAI22X1 OAI22X1_780 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2715_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5270_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2847_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5267_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6004_));
OAI22X1 OAI22X1_781 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3046_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5274_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3112_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5273_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6005_));
OAI22X1 OAI22X1_782 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3505_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5279_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3570_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5278_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6008_));
OAI22X1 OAI22X1_783 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4026_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5288_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3636_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5286_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6012_));
OAI22X1 OAI22X1_784 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3896_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5290_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3961_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5291_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6013_));
OAI22X1 OAI22X1_785 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3177_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5298_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2451_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5296_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6017_));
OAI22X1 OAI22X1_786 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2383_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5301_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2171_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5300_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6018_));
OAI22X1 OAI22X1_787 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2980_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5307_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2912_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5306_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6020_));
OAI22X1 OAI22X1_788 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3440_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5311_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3374_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5312_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6023_));
OAI22X1 OAI22X1_789 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3766_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5315_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3701_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5314_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6024_));
OAI22X1 OAI22X1_79 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3000_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4202_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3066_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4201_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4203_));
OAI22X1 OAI22X1_790 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4091_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5319_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4156_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5318_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6026_));
OAI22X1 OAI22X1_791 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2249_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5322_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3831_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5321_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6027_));
OAI22X1 OAI22X1_792 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2519_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5262_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2585_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5259_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6034_));
OAI22X1 OAI22X1_793 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2717_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5270_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2849_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5267_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6036_));
OAI22X1 OAI22X1_794 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3048_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5274_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3114_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5273_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6037_));
OAI22X1 OAI22X1_795 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3507_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5279_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3572_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5278_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6040_));
OAI22X1 OAI22X1_796 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4028_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5288_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3638_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5286_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6044_));
OAI22X1 OAI22X1_797 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3898_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5290_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3963_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5291_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6045_));
OAI22X1 OAI22X1_798 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3179_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5298_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2453_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5296_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6049_));
OAI22X1 OAI22X1_799 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2385_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5301_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2174_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5300_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6050_));
OAI22X1 OAI22X1_8 ( .A(_abc_40298_new_n1395_), .B(_abc_40298_new_n1066_), .C(_abc_40298_new_n1397_), .D(_abc_40298_new_n1405_), .Y(_abc_40298_new_n1406_));
OAI22X1 OAI22X1_80 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3460_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4207_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3525_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4206_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4208_));
OAI22X1 OAI22X1_800 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2982_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5307_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2914_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5306_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6052_));
OAI22X1 OAI22X1_801 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3442_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5311_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3376_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5312_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6055_));
OAI22X1 OAI22X1_802 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3768_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5315_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3703_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5314_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6056_));
OAI22X1 OAI22X1_803 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4093_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5319_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4158_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5318_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6058_));
OAI22X1 OAI22X1_804 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2251_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5322_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3833_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5321_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6059_));
OAI22X1 OAI22X1_805 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2521_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5262_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2587_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5259_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6066_));
OAI22X1 OAI22X1_806 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2719_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5270_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2851_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5267_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6068_));
OAI22X1 OAI22X1_807 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3050_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5274_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3116_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5273_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6069_));
OAI22X1 OAI22X1_808 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3509_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5279_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3574_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5278_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6072_));
OAI22X1 OAI22X1_809 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4030_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5288_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3640_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5286_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6076_));
OAI22X1 OAI22X1_81 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3981_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4216_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3590_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4214_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4217_));
OAI22X1 OAI22X1_810 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3900_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5290_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3965_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5291_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6077_));
OAI22X1 OAI22X1_811 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3181_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5298_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2455_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5296_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6081_));
OAI22X1 OAI22X1_812 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2387_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5301_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2177_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5300_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6082_));
OAI22X1 OAI22X1_813 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2984_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5307_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2916_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5306_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6084_));
OAI22X1 OAI22X1_814 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3444_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5311_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3378_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5312_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6087_));
OAI22X1 OAI22X1_815 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3770_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5315_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3705_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5314_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6088_));
OAI22X1 OAI22X1_816 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4095_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5319_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4160_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5318_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6090_));
OAI22X1 OAI22X1_817 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2253_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5322_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3835_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5321_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6091_));
OAI22X1 OAI22X1_818 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2523_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5262_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2589_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5259_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6098_));
OAI22X1 OAI22X1_819 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2721_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5270_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2853_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5267_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6100_));
OAI22X1 OAI22X1_82 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3851_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4218_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3916_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4219_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4220_));
OAI22X1 OAI22X1_820 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3052_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5274_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3118_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5273_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6101_));
OAI22X1 OAI22X1_821 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3511_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5279_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3576_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5278_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6104_));
OAI22X1 OAI22X1_822 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4032_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5288_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3642_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5286_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6108_));
OAI22X1 OAI22X1_823 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3902_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5290_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3967_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5291_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6109_));
OAI22X1 OAI22X1_824 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3183_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5298_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2457_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5296_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6113_));
OAI22X1 OAI22X1_825 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2389_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5301_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2180_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5300_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6114_));
OAI22X1 OAI22X1_826 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2986_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5307_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2918_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5306_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6116_));
OAI22X1 OAI22X1_827 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3446_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5311_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3380_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5312_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6119_));
OAI22X1 OAI22X1_828 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3772_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5315_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3707_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5314_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6120_));
OAI22X1 OAI22X1_829 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4097_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5319_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4162_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5318_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6122_));
OAI22X1 OAI22X1_83 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3132_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4226_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2403_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4224_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4227_));
OAI22X1 OAI22X1_830 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2255_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5322_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3837_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5321_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6123_));
OAI22X1 OAI22X1_831 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2525_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5262_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2591_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5259_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6130_));
OAI22X1 OAI22X1_832 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2723_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5270_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2855_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5267_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6132_));
OAI22X1 OAI22X1_833 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3054_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5274_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3120_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5273_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6133_));
OAI22X1 OAI22X1_834 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3513_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5279_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3578_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5278_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6136_));
OAI22X1 OAI22X1_835 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4034_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5288_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3644_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5286_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6140_));
OAI22X1 OAI22X1_836 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3904_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5290_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3969_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5291_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6141_));
OAI22X1 OAI22X1_837 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3185_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5298_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2459_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5296_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6145_));
OAI22X1 OAI22X1_838 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2391_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5301_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2183_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5300_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6146_));
OAI22X1 OAI22X1_839 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2988_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5307_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2920_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5306_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6148_));
OAI22X1 OAI22X1_84 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2336_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4229_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2099_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4228_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4230_));
OAI22X1 OAI22X1_840 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3448_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5311_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3382_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5312_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6151_));
OAI22X1 OAI22X1_841 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3774_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5315_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3709_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5314_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6152_));
OAI22X1 OAI22X1_842 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4099_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5319_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4164_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5318_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6154_));
OAI22X1 OAI22X1_843 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2257_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5322_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3839_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5321_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6155_));
OAI22X1 OAI22X1_844 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2527_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5262_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2593_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5259_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6162_));
OAI22X1 OAI22X1_845 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2725_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5270_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2857_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5267_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6164_));
OAI22X1 OAI22X1_846 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3056_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5274_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3122_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5273_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6165_));
OAI22X1 OAI22X1_847 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3515_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5279_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3580_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5278_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6168_));
OAI22X1 OAI22X1_848 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4036_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5288_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3646_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5286_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6172_));
OAI22X1 OAI22X1_849 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3906_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5290_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3971_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5291_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6173_));
OAI22X1 OAI22X1_85 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2932_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4235_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2867_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4234_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4236_));
OAI22X1 OAI22X1_850 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3187_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5298_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2461_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5296_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6177_));
OAI22X1 OAI22X1_851 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2393_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5301_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2186_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5300_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6178_));
OAI22X1 OAI22X1_852 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2990_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5307_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2922_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5306_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6180_));
OAI22X1 OAI22X1_853 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3450_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5311_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3384_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5312_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6183_));
OAI22X1 OAI22X1_854 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3776_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5315_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3711_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5314_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6184_));
OAI22X1 OAI22X1_855 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4101_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5319_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4166_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5318_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6186_));
OAI22X1 OAI22X1_856 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2259_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5322_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3841_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5321_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6187_));
OAI22X1 OAI22X1_857 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2529_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5262_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2595_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5259_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6194_));
OAI22X1 OAI22X1_858 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2727_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5270_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2859_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5267_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6196_));
OAI22X1 OAI22X1_859 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3058_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5274_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3124_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5273_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6197_));
OAI22X1 OAI22X1_86 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3394_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4239_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3329_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4240_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4241_));
OAI22X1 OAI22X1_860 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3517_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5279_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3582_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5278_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6200_));
OAI22X1 OAI22X1_861 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4038_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5288_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3648_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5286_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6204_));
OAI22X1 OAI22X1_862 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3908_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5290_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3973_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5291_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6205_));
OAI22X1 OAI22X1_863 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3189_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5298_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2463_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5296_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6209_));
OAI22X1 OAI22X1_864 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2395_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5301_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2189_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5300_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6210_));
OAI22X1 OAI22X1_865 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2992_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5307_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2924_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5306_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6212_));
OAI22X1 OAI22X1_866 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3452_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5311_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3386_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5312_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6215_));
OAI22X1 OAI22X1_867 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3778_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5315_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3713_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5314_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6216_));
OAI22X1 OAI22X1_868 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4103_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5319_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4168_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5318_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6218_));
OAI22X1 OAI22X1_869 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2261_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5322_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3843_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5321_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6219_));
OAI22X1 OAI22X1_87 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3721_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4243_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3656_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4242_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4244_));
OAI22X1 OAI22X1_870 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2531_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5262_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2597_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5259_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6226_));
OAI22X1 OAI22X1_871 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2729_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5270_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2861_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5267_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6228_));
OAI22X1 OAI22X1_872 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3060_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5274_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3126_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5273_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6229_));
OAI22X1 OAI22X1_873 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3519_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5279_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3584_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5278_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6232_));
OAI22X1 OAI22X1_874 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4040_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5288_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3650_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5286_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6236_));
OAI22X1 OAI22X1_875 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3910_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5290_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3975_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5291_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6237_));
OAI22X1 OAI22X1_876 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3191_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5298_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2465_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5296_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6241_));
OAI22X1 OAI22X1_877 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2397_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5301_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2192_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5300_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6242_));
OAI22X1 OAI22X1_878 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2994_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5307_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2926_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5306_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6244_));
OAI22X1 OAI22X1_879 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3454_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5311_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3388_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5312_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6247_));
OAI22X1 OAI22X1_88 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4046_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4247_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4111_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4246_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4248_));
OAI22X1 OAI22X1_880 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3780_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5315_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3715_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5314_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6248_));
OAI22X1 OAI22X1_881 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4105_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5319_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4170_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5318_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6250_));
OAI22X1 OAI22X1_882 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2263_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5322_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3845_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5321_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6251_));
OAI22X1 OAI22X1_883 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2533_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5262_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2599_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5259_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6258_));
OAI22X1 OAI22X1_884 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2731_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5270_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2863_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5267_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6260_));
OAI22X1 OAI22X1_885 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3062_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5274_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3128_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5273_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6261_));
OAI22X1 OAI22X1_886 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3521_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5279_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3586_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5278_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6264_));
OAI22X1 OAI22X1_887 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4042_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5288_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3652_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5286_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6268_));
OAI22X1 OAI22X1_888 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3912_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5290_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3977_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5291_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6269_));
OAI22X1 OAI22X1_889 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3193_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5298_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2467_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5296_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6273_));
OAI22X1 OAI22X1_89 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2201_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4250_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3786_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4249_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4251_));
OAI22X1 OAI22X1_890 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2399_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5301_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2195_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5300_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6274_));
OAI22X1 OAI22X1_891 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2996_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5307_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2928_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5306_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6276_));
OAI22X1 OAI22X1_892 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3456_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5311_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3390_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5312_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6279_));
OAI22X1 OAI22X1_893 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3782_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5315_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3717_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5314_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6280_));
OAI22X1 OAI22X1_894 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4107_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5319_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4172_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5318_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6282_));
OAI22X1 OAI22X1_895 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2265_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5322_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3847_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5321_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6283_));
OAI22X1 OAI22X1_896 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2535_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5262_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2601_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5259_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6290_));
OAI22X1 OAI22X1_897 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2733_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5270_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2865_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5267_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6292_));
OAI22X1 OAI22X1_898 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3064_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5274_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3130_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5273_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6293_));
OAI22X1 OAI22X1_899 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3523_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5279_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3588_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5278_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6296_));
OAI22X1 OAI22X1_9 ( .A(_abc_40298_new_n1213_), .B(_abc_40298_new_n1391_), .C(_abc_40298_new_n1408_), .D(_abc_40298_new_n1407_), .Y(_abc_40298_new_n1409_));
OAI22X1 OAI22X1_90 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2475_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4190_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2541_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4187_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4258_));
OAI22X1 OAI22X1_900 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4044_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5288_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3654_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5286_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6300_));
OAI22X1 OAI22X1_901 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3914_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5290_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3979_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5291_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6301_));
OAI22X1 OAI22X1_902 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3195_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5298_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2469_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5296_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6305_));
OAI22X1 OAI22X1_903 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2401_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5301_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2198_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5300_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6306_));
OAI22X1 OAI22X1_904 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2998_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5307_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2930_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5306_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6308_));
OAI22X1 OAI22X1_905 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3458_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5311_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3392_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5312_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6311_));
OAI22X1 OAI22X1_906 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3784_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5315_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3719_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5314_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6312_));
OAI22X1 OAI22X1_907 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n4109_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5319_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n4174_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5318_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6314_));
OAI22X1 OAI22X1_908 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2267_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n5322_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3849_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n5321_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n6315_));
OAI22X1 OAI22X1_909 ( .A(alu__abc_38674_new_n420_), .B(alu__abc_38674_new_n710_), .C(alu__abc_38674_new_n258_), .D(alu__abc_38674_new_n713_), .Y(alu__abc_38674_new_n714_));
OAI22X1 OAI22X1_91 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2673_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4198_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2805_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4195_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4260_));
OAI22X1 OAI22X1_910 ( .A(alu__abc_38674_new_n267_), .B(alu__abc_38674_new_n787_), .C(alu__abc_38674_new_n834_), .D(alu__abc_38674_new_n788_), .Y(alu__abc_38674_new_n845_));
OAI22X1 OAI22X1_911 ( .A(alu__abc_38674_new_n245_), .B(alu__abc_38674_new_n710_), .C(alu__abc_38674_new_n247_), .D(alu__abc_38674_new_n788_), .Y(alu__abc_38674_new_n1000_));
OAI22X1 OAI22X1_912 ( .A(alu__abc_38674_new_n249_), .B(alu__abc_38674_new_n787_), .C(alu__abc_38674_new_n517_), .D(alu__abc_38674_new_n788_), .Y(alu__abc_38674_new_n1034_));
OAI22X1 OAI22X1_913 ( .A(alu__abc_38674_new_n283_), .B(alu__abc_38674_new_n538_), .C(alu__abc_38674_new_n1075_), .D(alu__abc_38674_new_n1077_), .Y(alu__abc_38674_new_n1078_));
OAI22X1 OAI22X1_914 ( .A(alu__abc_38674_new_n702_), .B(alu__abc_38674_new_n1093_), .C(alu__abc_38674_new_n658_), .D(alu__abc_38674_new_n1084_), .Y(alu__abc_38674_new_n1094_));
OAI22X1 OAI22X1_915 ( .A(alu__abc_38674_new_n1146_), .B(alu__abc_38674_new_n1149_), .C(alu__abc_38674_new_n519_), .D(alu__abc_38674_new_n1148_), .Y(alu__abc_38674_new_n1150_));
OAI22X1 OAI22X1_916 ( .A(alu__abc_38674_new_n213_), .B(alu__abc_38674_new_n787_), .C(alu__abc_38674_new_n215_), .D(alu__abc_38674_new_n788_), .Y(alu__abc_38674_new_n1188_));
OAI22X1 OAI22X1_917 ( .A(alu__abc_38674_new_n1193_), .B(alu__abc_38674_new_n1194_), .C(alu__abc_38674_new_n519_), .D(alu__abc_38674_new_n1192_), .Y(alu__abc_38674_new_n1195_));
OAI22X1 OAI22X1_918 ( .A(alu__abc_38674_new_n578_), .B(alu__abc_38674_new_n710_), .C(alu__abc_38674_new_n658_), .D(alu__abc_38674_new_n1195_), .Y(alu__abc_38674_new_n1196_));
OAI22X1 OAI22X1_919 ( .A(alu__abc_38674_new_n283_), .B(alu__abc_38674_new_n584_), .C(alu__abc_38674_new_n382_), .D(alu__abc_38674_new_n1205_), .Y(alu__abc_38674_new_n1206_));
OAI22X1 OAI22X1_92 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3004_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4202_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3070_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4201_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4261_));
OAI22X1 OAI22X1_920 ( .A(alu__abc_38674_new_n512_), .B(alu__abc_38674_new_n710_), .C(alu__abc_38674_new_n204_), .D(alu__abc_38674_new_n787_), .Y(alu__abc_38674_new_n1256_));
OAI22X1 OAI22X1_921 ( .A(alu__abc_38674_new_n283_), .B(alu__abc_38674_new_n1266_), .C(alu__abc_38674_new_n382_), .D(alu__abc_38674_new_n1270_), .Y(alu__abc_38674_new_n1271_));
OAI22X1 OAI22X1_922 ( .A(alu__abc_38674_new_n206_), .B(alu__abc_38674_new_n787_), .C(alu__abc_38674_new_n208_), .D(alu__abc_38674_new_n788_), .Y(alu__abc_38674_new_n1289_));
OAI22X1 OAI22X1_923 ( .A(alu__abc_38674_new_n485_), .B(alu__abc_38674_new_n710_), .C(alu__abc_38674_new_n307_), .D(alu__abc_38674_new_n788_), .Y(alu__abc_38674_new_n1379_));
OAI22X1 OAI22X1_924 ( .A(alu__abc_38674_new_n283_), .B(alu__abc_38674_new_n1412_), .C(alu__abc_38674_new_n382_), .D(alu__abc_38674_new_n1417_), .Y(alu__abc_38674_new_n1418_));
OAI22X1 OAI22X1_925 ( .A(alu__abc_38674_new_n124_), .B(alu__abc_38674_new_n787_), .C(alu__abc_38674_new_n126_), .D(alu__abc_38674_new_n788_), .Y(alu__abc_38674_new_n1434_));
OAI22X1 OAI22X1_926 ( .A(alu__abc_38674_new_n130_), .B(alu__abc_38674_new_n787_), .C(alu__abc_38674_new_n1461_), .D(alu__abc_38674_new_n788_), .Y(alu__abc_38674_new_n1462_));
OAI22X1 OAI22X1_927 ( .A(alu__abc_38674_new_n119_), .B(alu__abc_38674_new_n787_), .C(alu__abc_38674_new_n322_), .D(alu__abc_38674_new_n788_), .Y(alu__abc_38674_new_n1517_));
OAI22X1 OAI22X1_928 ( .A(alu__abc_38674_new_n283_), .B(alu__abc_38674_new_n507_), .C(alu__abc_38674_new_n382_), .D(alu__abc_38674_new_n1525_), .Y(alu__abc_38674_new_n1526_));
OAI22X1 OAI22X1_929 ( .A(alu__abc_38674_new_n501_), .B(alu__abc_38674_new_n710_), .C(alu__abc_38674_new_n180_), .D(alu__abc_38674_new_n787_), .Y(alu__abc_38674_new_n1540_));
OAI22X1 OAI22X1_93 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3463_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4207_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3528_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4206_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4264_));
OAI22X1 OAI22X1_930 ( .A(alu__abc_38674_new_n394_), .B(alu__abc_38674_new_n710_), .C(alu__abc_38674_new_n396_), .D(alu__abc_38674_new_n788_), .Y(alu__abc_38674_new_n1615_));
OAI22X1 OAI22X1_931 ( .A(alu__abc_38674_new_n1635_), .B(alu__abc_38674_new_n1636_), .C(alu__abc_38674_new_n338_), .D(alu__abc_38674_new_n1535_), .Y(alu__abc_38674_new_n1637_));
OAI22X1 OAI22X1_932 ( .A(alu__abc_38674_new_n386_), .B(alu__abc_38674_new_n710_), .C(alu__abc_38674_new_n167_), .D(alu__abc_38674_new_n787_), .Y(alu__abc_38674_new_n1664_));
OAI22X1 OAI22X1_933 ( .A(alu__abc_38674_new_n610_), .B(alu__abc_38674_new_n710_), .C(alu__abc_38674_new_n383_), .D(alu__abc_38674_new_n788_), .Y(alu__abc_38674_new_n1687_));
OAI22X1 OAI22X1_94 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3984_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4216_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3594_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4214_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4268_));
OAI22X1 OAI22X1_95 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3854_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4218_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3919_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4219_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4269_));
OAI22X1 OAI22X1_96 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3135_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4226_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2409_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4224_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4273_));
OAI22X1 OAI22X1_97 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2341_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4229_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2108_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4228_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4274_));
OAI22X1 OAI22X1_98 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2938_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4235_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n2870_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4234_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4276_));
OAI22X1 OAI22X1_99 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n3398_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n4239_), .C(REGFILE_SIM_reg_bank__abc_34451_new_n3332_), .D(REGFILE_SIM_reg_bank__abc_34451_new_n4240_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n4279_));
OR2X2 OR2X2_1 ( .A(_abc_40298_new_n618_), .B(_abc_40298_new_n636_), .Y(_abc_40298_new_n1003_));
OR2X2 OR2X2_10 ( .A(_abc_40298_new_n1708_), .B(_abc_40298_new_n1704_), .Y(_abc_40298_new_n1709_));
OR2X2 OR2X2_11 ( .A(_abc_40298_new_n1921_), .B(_abc_40298_new_n1924_), .Y(_abc_40298_new_n1925_));
OR2X2 OR2X2_12 ( .A(_abc_40298_new_n1930_), .B(_abc_40298_new_n984_), .Y(_abc_40298_new_n1931_));
OR2X2 OR2X2_13 ( .A(_abc_40298_new_n2159_), .B(_abc_40298_new_n959_), .Y(_abc_40298_new_n2160_));
OR2X2 OR2X2_14 ( .A(_abc_40298_new_n2162_), .B(_abc_40298_new_n891_), .Y(_abc_40298_new_n2163_));
OR2X2 OR2X2_15 ( .A(_abc_40298_new_n2905_), .B(_abc_40298_new_n2903_), .Y(_abc_40298_new_n2906_));
OR2X2 OR2X2_16 ( .A(_abc_40298_new_n2979_), .B(_abc_40298_new_n2977_), .Y(_abc_40298_new_n2981_));
OR2X2 OR2X2_17 ( .A(_abc_40298_new_n3001_), .B(_abc_40298_new_n3004_), .Y(_abc_40298_new_n3006_));
OR2X2 OR2X2_18 ( .A(_abc_40298_new_n3012_), .B(_abc_40298_new_n1039_), .Y(_abc_40298_new_n3013_));
OR2X2 OR2X2_19 ( .A(_abc_40298_new_n3069_), .B(_abc_40298_new_n3066_), .Y(_abc_40298_new_n3071_));
OR2X2 OR2X2_2 ( .A(_abc_40298_new_n1089_), .B(alu_flag_update_o), .Y(_abc_40298_new_n1126_));
OR2X2 OR2X2_20 ( .A(_abc_40298_new_n3107_), .B(_abc_40298_new_n3122_), .Y(_abc_40298_new_n3125_));
OR2X2 OR2X2_21 ( .A(_abc_40298_new_n3146_), .B(_abc_40298_new_n3161_), .Y(_abc_40298_new_n3162_));
OR2X2 OR2X2_22 ( .A(_abc_40298_new_n3183_), .B(_abc_40298_new_n3179_), .Y(_abc_40298_new_n3184_));
OR2X2 OR2X2_23 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2202_), .B(REGFILE_SIM_reg_bank_rd_i_0_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2203_));
OR2X2 OR2X2_24 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2338_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2101_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2339_));
OR2X2 OR2X2_25 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2404_), .B(REGFILE_SIM_reg_bank_rd_i_2_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n2405_));
OR2X2 OR2X2_26 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2203_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2934_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3001_));
OR2X2 OR2X2_27 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2934_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2270_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3067_));
OR2X2 OR2X2_28 ( .A(REGFILE_SIM_reg_bank__abc_34451_new_n2338_), .B(REGFILE_SIM_reg_bank__abc_34451_new_n2934_), .Y(REGFILE_SIM_reg_bank__abc_34451_new_n3133_));
OR2X2 OR2X2_29 ( .A(alu_b_i_8_), .B(alu_a_i_8_), .Y(alu__abc_38674_new_n224_));
OR2X2 OR2X2_3 ( .A(_abc_40298_new_n1234_), .B(_abc_40298_new_n1216_), .Y(_abc_40298_new_n1235_));
OR2X2 OR2X2_30 ( .A(alu_b_i_11_), .B(alu_a_i_11_), .Y(alu__abc_38674_new_n238_));
OR2X2 OR2X2_31 ( .A(alu__abc_38674_new_n222_), .B(alu__abc_38674_new_n242_), .Y(alu__abc_38674_new_n243_));
OR2X2 OR2X2_32 ( .A(alu_b_i_6_), .B(alu_a_i_6_), .Y(alu__abc_38674_new_n246_));
OR2X2 OR2X2_33 ( .A(alu_b_i_5_), .B(alu_a_i_5_), .Y(alu__abc_38674_new_n252_));
OR2X2 OR2X2_34 ( .A(alu__abc_38674_new_n364_), .B(alu_b_i_15_), .Y(alu__abc_38674_new_n365_));
OR2X2 OR2X2_35 ( .A(alu__abc_38674_new_n378_), .B(alu__abc_38674_new_n162_), .Y(alu__abc_38674_new_n379_));
OR2X2 OR2X2_36 ( .A(alu_b_i_7_), .B(alu_a_i_7_), .Y(alu__abc_38674_new_n439_));
OR2X2 OR2X2_37 ( .A(alu__abc_38674_new_n470_), .B(alu__abc_38674_new_n474_), .Y(alu__abc_38674_new_n475_));
OR2X2 OR2X2_38 ( .A(alu__abc_38674_new_n470_), .B(alu__abc_38674_new_n472_), .Y(alu__abc_38674_new_n505_));
OR2X2 OR2X2_39 ( .A(alu__abc_38674_new_n421_), .B(alu__abc_38674_new_n268_), .Y(alu__abc_38674_new_n568_));
OR2X2 OR2X2_4 ( .A(_abc_40298_new_n1316_), .B(_abc_40298_new_n1314_), .Y(_abc_40298_new_n1317_));
OR2X2 OR2X2_40 ( .A(alu__abc_38674_new_n606_), .B(alu__abc_38674_new_n504_), .Y(alu__abc_38674_new_n607_));
OR2X2 OR2X2_41 ( .A(alu__abc_38674_new_n612_), .B(alu__abc_38674_new_n162_), .Y(alu__abc_38674_new_n613_));
OR2X2 OR2X2_42 ( .A(alu__abc_38674_new_n609_), .B(alu__abc_38674_new_n626_), .Y(alu__abc_38674_new_n627_));
OR2X2 OR2X2_43 ( .A(alu__abc_38674_new_n898_), .B(alu__abc_38674_new_n894_), .Y(alu__abc_38674_new_n899_));
OR2X2 OR2X2_44 ( .A(alu__abc_38674_new_n935_), .B(alu__abc_38674_new_n933_), .Y(alu__abc_38674_new_n936_));
OR2X2 OR2X2_45 ( .A(alu__abc_38674_new_n1067_), .B(alu__abc_38674_new_n702_), .Y(alu__abc_38674_new_n1068_));
OR2X2 OR2X2_46 ( .A(alu__abc_38674_new_n1196_), .B(alu__abc_38674_new_n1190_), .Y(alu__abc_38674_new_n1197_));
OR2X2 OR2X2_47 ( .A(alu__abc_38674_new_n1206_), .B(alu__abc_38674_new_n1232_), .Y(alu_p_o_13_));
OR2X2 OR2X2_48 ( .A(alu__abc_38674_new_n1359_), .B(alu__abc_38674_new_n1384_), .Y(alu__abc_38674_new_n1385_));
OR2X2 OR2X2_49 ( .A(alu__abc_38674_new_n865_), .B(alu_b_i_4_), .Y(alu__abc_38674_new_n1399_));
OR2X2 OR2X2_5 ( .A(_abc_40298_new_n1488_), .B(_abc_40298_new_n1484_), .Y(_abc_40298_new_n1489_));
OR2X2 OR2X2_50 ( .A(alu__abc_38674_new_n533_), .B(alu__abc_38674_new_n208_), .Y(alu__abc_38674_new_n1413_));
OR2X2 OR2X2_51 ( .A(alu__abc_38674_new_n1445_), .B(alu__abc_38674_new_n493_), .Y(alu__abc_38674_new_n1446_));
OR2X2 OR2X2_52 ( .A(alu__abc_38674_new_n1451_), .B(alu__abc_38674_new_n1466_), .Y(alu__abc_38674_new_n1467_));
OR2X2 OR2X2_53 ( .A(alu__abc_38674_new_n496_), .B(alu__abc_38674_new_n493_), .Y(alu__abc_38674_new_n1498_));
OR2X2 OR2X2_54 ( .A(alu__abc_38674_new_n1516_), .B(alu__abc_38674_new_n1519_), .Y(alu__abc_38674_new_n1520_));
OR2X2 OR2X2_55 ( .A(alu__abc_38674_new_n1522_), .B(alu__abc_38674_new_n1502_), .Y(alu_p_o_23_));
OR2X2 OR2X2_56 ( .A(alu__abc_38674_new_n1556_), .B(alu__abc_38674_new_n702_), .Y(alu__abc_38674_new_n1557_));
OR2X2 OR2X2_57 ( .A(alu__abc_38674_new_n1529_), .B(alu__abc_38674_new_n185_), .Y(alu__abc_38674_new_n1558_));
OR2X2 OR2X2_58 ( .A(alu__abc_38674_new_n1080_), .B(alu_b_i_4_), .Y(alu__abc_38674_new_n1563_));
OR2X2 OR2X2_59 ( .A(alu__abc_38674_new_n304_), .B(alu__abc_38674_new_n176_), .Y(alu__abc_38674_new_n1725_));
OR2X2 OR2X2_6 ( .A(_abc_40298_new_n1476_), .B(_abc_40298_new_n1213_), .Y(_abc_40298_new_n1501_));
OR2X2 OR2X2_7 ( .A(_abc_40298_new_n1595_), .B(_abc_40298_new_n1598_), .Y(_abc_40298_new_n1599_));
OR2X2 OR2X2_8 ( .A(_abc_40298_new_n1590_), .B(_abc_40298_new_n1213_), .Y(_abc_40298_new_n1612_));
OR2X2 OR2X2_9 ( .A(_abc_40298_new_n1662_), .B(_abc_40298_new_n1659_), .Y(_abc_40298_new_n1681_));
XNOR2X1 XNOR2X1_1 ( .A(_abc_40298_new_n988_), .B(_abc_40298_new_n1092_), .Y(_abc_40298_new_n1093_));
XNOR2X1 XNOR2X1_10 ( .A(_abc_40298_new_n1913_), .B(pc_q_29_), .Y(_abc_40298_new_n1941_));
XNOR2X1 XNOR2X1_11 ( .A(_abc_40298_new_n2520_), .B(_abc_40298_new_n2513_), .Y(_abc_40298_new_n2521_));
XNOR2X1 XNOR2X1_12 ( .A(_abc_40298_new_n2923_), .B(_abc_40298_new_n2921_), .Y(_abc_40298_new_n2924_));
XNOR2X1 XNOR2X1_13 ( .A(_abc_40298_new_n2988_), .B(REGFILE_SIM_reg_bank_reg_ra_o_11_), .Y(_abc_40298_new_n2989_));
XNOR2X1 XNOR2X1_14 ( .A(_abc_40298_new_n3003_), .B(REGFILE_SIM_reg_bank_reg_ra_o_12_), .Y(_abc_40298_new_n3004_));
XNOR2X1 XNOR2X1_15 ( .A(_abc_40298_new_n3025_), .B(REGFILE_SIM_reg_bank_reg_ra_o_14_), .Y(_abc_40298_new_n3026_));
XNOR2X1 XNOR2X1_16 ( .A(_abc_40298_new_n3023_), .B(_abc_40298_new_n3026_), .Y(_abc_40298_new_n3027_));
XNOR2X1 XNOR2X1_17 ( .A(_abc_40298_new_n3039_), .B(_abc_40298_new_n2392_), .Y(_abc_40298_new_n3062_));
XNOR2X1 XNOR2X1_18 ( .A(_abc_40298_new_n3039_), .B(_abc_40298_new_n2399_), .Y(_abc_40298_new_n3066_));
XNOR2X1 XNOR2X1_19 ( .A(_abc_40298_new_n3039_), .B(_abc_40298_new_n2406_), .Y(_abc_40298_new_n3076_));
XNOR2X1 XNOR2X1_2 ( .A(_abc_40298_new_n1282_), .B(_abc_40298_new_n1281_), .Y(_abc_40298_new_n1283_));
XNOR2X1 XNOR2X1_20 ( .A(_abc_40298_new_n3039_), .B(_abc_40298_new_n2420_), .Y(_abc_40298_new_n3098_));
XNOR2X1 XNOR2X1_21 ( .A(_abc_40298_new_n3036_), .B(_abc_40298_new_n2427_), .Y(_abc_40298_new_n3104_));
XNOR2X1 XNOR2X1_22 ( .A(_abc_40298_new_n3036_), .B(_abc_40298_new_n2434_), .Y(_abc_40298_new_n3115_));
XNOR2X1 XNOR2X1_23 ( .A(_abc_40298_new_n3036_), .B(_abc_40298_new_n2441_), .Y(_abc_40298_new_n3129_));
XNOR2X1 XNOR2X1_24 ( .A(_abc_40298_new_n3036_), .B(_abc_40298_new_n2448_), .Y(_abc_40298_new_n3137_));
XNOR2X1 XNOR2X1_25 ( .A(_abc_40298_new_n3036_), .B(_abc_40298_new_n2455_), .Y(_abc_40298_new_n3149_));
XNOR2X1 XNOR2X1_26 ( .A(_abc_40298_new_n3036_), .B(_abc_40298_new_n2463_), .Y(_abc_40298_new_n3157_));
XNOR2X1 XNOR2X1_27 ( .A(_abc_40298_new_n3156_), .B(_abc_40298_new_n3157_), .Y(_abc_40298_new_n3158_));
XNOR2X1 XNOR2X1_28 ( .A(_abc_40298_new_n3036_), .B(_abc_40298_new_n2470_), .Y(_abc_40298_new_n3166_));
XNOR2X1 XNOR2X1_29 ( .A(_abc_40298_new_n3039_), .B(_abc_40298_new_n2478_), .Y(_abc_40298_new_n3173_));
XNOR2X1 XNOR2X1_3 ( .A(_abc_40298_new_n1364_), .B(pc_q_9_), .Y(_abc_40298_new_n1391_));
XNOR2X1 XNOR2X1_30 ( .A(_abc_40298_new_n3036_), .B(REGFILE_SIM_reg_bank_reg_ra_o_31_), .Y(_abc_40298_new_n3191_));
XNOR2X1 XNOR2X1_31 ( .A(alu__abc_38674_new_n482_), .B(alu__abc_38674_new_n169_), .Y(alu__abc_38674_new_n483_));
XNOR2X1 XNOR2X1_32 ( .A(alu__abc_38674_new_n480_), .B(alu__abc_38674_new_n390_), .Y(alu__abc_38674_new_n484_));
XNOR2X1 XNOR2X1_33 ( .A(alu__abc_38674_new_n489_), .B(alu__abc_38674_new_n150_), .Y(alu__abc_38674_new_n490_));
XNOR2X1 XNOR2X1_34 ( .A(alu__abc_38674_new_n492_), .B(alu__abc_38674_new_n410_), .Y(alu__abc_38674_new_n493_));
XNOR2X1 XNOR2X1_35 ( .A(alu__abc_38674_new_n495_), .B(alu__abc_38674_new_n114_), .Y(alu__abc_38674_new_n496_));
XNOR2X1 XNOR2X1_36 ( .A(alu__abc_38674_new_n498_), .B(alu__abc_38674_new_n191_), .Y(alu__abc_38674_new_n499_));
XNOR2X1 XNOR2X1_37 ( .A(alu__abc_38674_new_n502_), .B(alu__abc_38674_new_n184_), .Y(alu__abc_38674_new_n503_));
XNOR2X1 XNOR2X1_38 ( .A(alu__abc_38674_new_n464_), .B(alu__abc_38674_new_n509_), .Y(alu__abc_38674_new_n510_));
XNOR2X1 XNOR2X1_39 ( .A(alu__abc_38674_new_n536_), .B(alu__abc_38674_new_n230_), .Y(alu__abc_38674_new_n537_));
XNOR2X1 XNOR2X1_4 ( .A(_abc_40298_new_n1475_), .B(pc_q_13_), .Y(_abc_40298_new_n1509_));
XNOR2X1 XNOR2X1_40 ( .A(alu__abc_38674_new_n442_), .B(alu__abc_38674_new_n539_), .Y(alu__abc_38674_new_n540_));
XNOR2X1 XNOR2X1_41 ( .A(alu__abc_38674_new_n543_), .B(alu__abc_38674_new_n517_), .Y(alu__abc_38674_new_n544_));
XNOR2X1 XNOR2X1_42 ( .A(alu__abc_38674_new_n425_), .B(alu__abc_38674_new_n521_), .Y(alu__abc_38674_new_n571_));
XNOR2X1 XNOR2X1_43 ( .A(alu__abc_38674_new_n531_), .B(alu__abc_38674_new_n215_), .Y(alu__abc_38674_new_n595_));
XNOR2X1 XNOR2X1_44 ( .A(alu__abc_38674_new_n491_), .B(alu__abc_38674_new_n125_), .Y(alu__abc_38674_new_n599_));
XNOR2X1 XNOR2X1_45 ( .A(alu__abc_38674_new_n488_), .B(alu__abc_38674_new_n306_), .Y(alu__abc_38674_new_n600_));
XNOR2X1 XNOR2X1_46 ( .A(alu__abc_38674_new_n602_), .B(alu__abc_38674_new_n141_), .Y(alu__abc_38674_new_n603_));
XNOR2X1 XNOR2X1_47 ( .A(alu__abc_38674_new_n611_), .B(alu__abc_38674_new_n159_), .Y(alu__abc_38674_new_n616_));
XNOR2X1 XNOR2X1_48 ( .A(alu__abc_38674_new_n618_), .B(alu__abc_38674_new_n396_), .Y(alu__abc_38674_new_n619_));
XNOR2X1 XNOR2X1_49 ( .A(alu__abc_38674_new_n622_), .B(alu__abc_38674_new_n322_), .Y(alu__abc_38674_new_n623_));
XNOR2X1 XNOR2X1_5 ( .A(_abc_40298_new_n1633_), .B(_abc_40298_new_n1631_), .Y(_abc_40298_new_n1634_));
XNOR2X1 XNOR2X1_50 ( .A(alu__abc_38674_new_n561_), .B(alu__abc_38674_new_n420_), .Y(alu__abc_38674_new_n786_));
XNOR2X1 XNOR2X1_51 ( .A(alu__abc_38674_new_n425_), .B(alu__abc_38674_new_n335_), .Y(alu__abc_38674_new_n903_));
XNOR2X1 XNOR2X1_52 ( .A(alu__abc_38674_new_n531_), .B(alu__abc_38674_new_n214_), .Y(alu__abc_38674_new_n1176_));
XNOR2X1 XNOR2X1_53 ( .A(alu__abc_38674_new_n532_), .B(alu__abc_38674_new_n453_), .Y(alu__abc_38674_new_n1240_));
XNOR2X1 XNOR2X1_54 ( .A(alu__abc_38674_new_n602_), .B(alu__abc_38674_new_n140_), .Y(alu__abc_38674_new_n1327_));
XNOR2X1 XNOR2X1_55 ( .A(alu__abc_38674_new_n488_), .B(alu__abc_38674_new_n307_), .Y(alu__abc_38674_new_n1358_));
XNOR2X1 XNOR2X1_56 ( .A(alu__abc_38674_new_n491_), .B(alu__abc_38674_new_n126_), .Y(alu__abc_38674_new_n1412_));
XNOR2X1 XNOR2X1_57 ( .A(alu__abc_38674_new_n1449_), .B(alu__abc_38674_new_n410_), .Y(alu__abc_38674_new_n1450_));
XNOR2X1 XNOR2X1_58 ( .A(alu__abc_38674_new_n1650_), .B(alu__abc_38674_new_n1649_), .Y(alu__abc_38674_new_n1651_));
XNOR2X1 XNOR2X1_6 ( .A(_abc_40298_new_n1807_), .B(pc_q_25_), .Y(_abc_40298_new_n1841_));
XNOR2X1 XNOR2X1_7 ( .A(_abc_40298_new_n1848_), .B(_abc_40298_new_n1846_), .Y(_abc_40298_new_n1849_));
XNOR2X1 XNOR2X1_8 ( .A(_abc_40298_new_n1864_), .B(pc_q_27_), .Y(_abc_40298_new_n1891_));
XNOR2X1 XNOR2X1_9 ( .A(_abc_40298_new_n1899_), .B(_abc_40298_new_n1897_), .Y(_abc_40298_new_n1900_));
XOR2X1 XOR2X1_1 ( .A(alu_op_r_1_), .B(pc_q_3_), .Y(_abc_40298_new_n1234_));
XOR2X1 XOR2X1_2 ( .A(opcode_q_25_), .B(pc_q_29_), .Y(_abc_40298_new_n1944_));
XOR2X1 XOR2X1_3 ( .A(_abc_40298_new_n2968_), .B(_abc_40298_new_n2970_), .Y(_abc_40298_new_n2971_));
XOR2X1 XOR2X1_4 ( .A(_abc_40298_new_n3034_), .B(_abc_40298_new_n3041_), .Y(_abc_40298_new_n3042_));
XOR2X1 XOR2X1_5 ( .A(_abc_40298_new_n3061_), .B(_abc_40298_new_n3062_), .Y(_abc_40298_new_n3063_));
XOR2X1 XOR2X1_6 ( .A(_abc_40298_new_n3172_), .B(_abc_40298_new_n3173_), .Y(_abc_40298_new_n3174_));

assign \mem_cti_o[0]  = 1'h1;
assign \mem_cti_o[1]  = 1'h1;
assign \mem_cti_o[2]  = 1'h1;

endmodule