module b04_reset(clock, RESET_G, nRESET_G, RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_, DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_, DATA_OUT_REG_7_, DATA_OUT_REG_6_, DATA_OUT_REG_5_, DATA_OUT_REG_4_, DATA_OUT_REG_3_, DATA_OUT_REG_2_, DATA_OUT_REG_1_, DATA_OUT_REG_0_);

input AVERAGE;
input DATA_IN_0_;
input DATA_IN_1_;
input DATA_IN_2_;
input DATA_IN_3_;
input DATA_IN_4_;
input DATA_IN_5_;
input DATA_IN_6_;
input DATA_IN_7_;
output DATA_OUT_REG_0_;
output DATA_OUT_REG_1_;
output DATA_OUT_REG_2_;
output DATA_OUT_REG_3_;
output DATA_OUT_REG_4_;
output DATA_OUT_REG_5_;
output DATA_OUT_REG_6_;
output DATA_OUT_REG_7_;
input ENABLE;
wire REG1_REG_0_; 
wire REG1_REG_1_; 
wire REG1_REG_2_; 
wire REG1_REG_3_; 
wire REG1_REG_4_; 
wire REG1_REG_5_; 
wire REG1_REG_6_; 
wire REG1_REG_7_; 
wire REG2_REG_0_; 
wire REG2_REG_1_; 
wire REG2_REG_2_; 
wire REG2_REG_3_; 
wire REG2_REG_4_; 
wire REG2_REG_5_; 
wire REG2_REG_6_; 
wire REG2_REG_7_; 
wire REG3_REG_0_; 
wire REG3_REG_1_; 
wire REG3_REG_2_; 
wire REG3_REG_3_; 
wire REG3_REG_4_; 
wire REG3_REG_5_; 
wire REG3_REG_6_; 
wire REG3_REG_7_; 
wire REG4_REG_0_; 
wire REG4_REG_1_; 
wire REG4_REG_2_; 
wire REG4_REG_3_; 
wire REG4_REG_4_; 
wire REG4_REG_5_; 
wire REG4_REG_6_; 
wire REG4_REG_7_; 
input RESET_G;
input RESTART;
wire RLAST_REG_0_; 
wire RLAST_REG_1_; 
wire RLAST_REG_2_; 
wire RLAST_REG_3_; 
wire RLAST_REG_4_; 
wire RLAST_REG_5_; 
wire RLAST_REG_6_; 
wire RLAST_REG_7_; 
wire RMAX_REG_0_; 
wire RMAX_REG_1_; 
wire RMAX_REG_2_; 
wire RMAX_REG_3_; 
wire RMAX_REG_4_; 
wire RMAX_REG_5_; 
wire RMAX_REG_6_; 
wire RMAX_REG_7_; 
wire RMIN_REG_0_; 
wire RMIN_REG_1_; 
wire RMIN_REG_2_; 
wire RMIN_REG_3_; 
wire RMIN_REG_4_; 
wire RMIN_REG_5_; 
wire RMIN_REG_6_; 
wire RMIN_REG_7_; 
wire STATO_REG_0_; 
wire STATO_REG_1_; 
wire _abc_3576_new_n146_; 
wire _abc_3576_new_n147_; 
wire _abc_3576_new_n148_; 
wire _abc_3576_new_n149_; 
wire _abc_3576_new_n150_; 
wire _abc_3576_new_n151_; 
wire _abc_3576_new_n153_; 
wire _abc_3576_new_n154_; 
wire _abc_3576_new_n155_; 
wire _abc_3576_new_n156_; 
wire _abc_3576_new_n157_; 
wire _abc_3576_new_n158_; 
wire _abc_3576_new_n159_; 
wire _abc_3576_new_n160_; 
wire _abc_3576_new_n161_; 
wire _abc_3576_new_n162_; 
wire _abc_3576_new_n163_; 
wire _abc_3576_new_n164_; 
wire _abc_3576_new_n165_; 
wire _abc_3576_new_n166_; 
wire _abc_3576_new_n167_; 
wire _abc_3576_new_n168_; 
wire _abc_3576_new_n169_; 
wire _abc_3576_new_n170_; 
wire _abc_3576_new_n171_; 
wire _abc_3576_new_n172_; 
wire _abc_3576_new_n173_; 
wire _abc_3576_new_n174_; 
wire _abc_3576_new_n175_; 
wire _abc_3576_new_n176_; 
wire _abc_3576_new_n177_; 
wire _abc_3576_new_n178_; 
wire _abc_3576_new_n179_; 
wire _abc_3576_new_n180_; 
wire _abc_3576_new_n181_; 
wire _abc_3576_new_n182_; 
wire _abc_3576_new_n183_; 
wire _abc_3576_new_n184_; 
wire _abc_3576_new_n185_; 
wire _abc_3576_new_n186_; 
wire _abc_3576_new_n187_; 
wire _abc_3576_new_n188_; 
wire _abc_3576_new_n189_; 
wire _abc_3576_new_n190_; 
wire _abc_3576_new_n191_; 
wire _abc_3576_new_n192_; 
wire _abc_3576_new_n193_; 
wire _abc_3576_new_n194_; 
wire _abc_3576_new_n195_; 
wire _abc_3576_new_n196_; 
wire _abc_3576_new_n197_; 
wire _abc_3576_new_n198_; 
wire _abc_3576_new_n199_; 
wire _abc_3576_new_n200_; 
wire _abc_3576_new_n201_; 
wire _abc_3576_new_n202_; 
wire _abc_3576_new_n203_; 
wire _abc_3576_new_n204_; 
wire _abc_3576_new_n205_; 
wire _abc_3576_new_n206_; 
wire _abc_3576_new_n207_; 
wire _abc_3576_new_n208_; 
wire _abc_3576_new_n209_; 
wire _abc_3576_new_n210_; 
wire _abc_3576_new_n211_; 
wire _abc_3576_new_n212_; 
wire _abc_3576_new_n213_; 
wire _abc_3576_new_n214_; 
wire _abc_3576_new_n215_; 
wire _abc_3576_new_n216_; 
wire _abc_3576_new_n217_; 
wire _abc_3576_new_n218_; 
wire _abc_3576_new_n219_; 
wire _abc_3576_new_n220_; 
wire _abc_3576_new_n221_; 
wire _abc_3576_new_n222_; 
wire _abc_3576_new_n223_; 
wire _abc_3576_new_n224_; 
wire _abc_3576_new_n225_; 
wire _abc_3576_new_n226_; 
wire _abc_3576_new_n227_; 
wire _abc_3576_new_n228_; 
wire _abc_3576_new_n229_; 
wire _abc_3576_new_n230_; 
wire _abc_3576_new_n231_; 
wire _abc_3576_new_n232_; 
wire _abc_3576_new_n233_; 
wire _abc_3576_new_n234_; 
wire _abc_3576_new_n235_; 
wire _abc_3576_new_n236_; 
wire _abc_3576_new_n237_; 
wire _abc_3576_new_n238_; 
wire _abc_3576_new_n239_; 
wire _abc_3576_new_n240_; 
wire _abc_3576_new_n241_; 
wire _abc_3576_new_n242_; 
wire _abc_3576_new_n243_; 
wire _abc_3576_new_n244_; 
wire _abc_3576_new_n245_; 
wire _abc_3576_new_n246_; 
wire _abc_3576_new_n247_; 
wire _abc_3576_new_n248_; 
wire _abc_3576_new_n249_; 
wire _abc_3576_new_n250_; 
wire _abc_3576_new_n251_; 
wire _abc_3576_new_n252_; 
wire _abc_3576_new_n253_; 
wire _abc_3576_new_n254_; 
wire _abc_3576_new_n255_; 
wire _abc_3576_new_n256_; 
wire _abc_3576_new_n257_; 
wire _abc_3576_new_n258_; 
wire _abc_3576_new_n259_; 
wire _abc_3576_new_n260_; 
wire _abc_3576_new_n261_; 
wire _abc_3576_new_n262_; 
wire _abc_3576_new_n263_; 
wire _abc_3576_new_n264_; 
wire _abc_3576_new_n265_; 
wire _abc_3576_new_n266_; 
wire _abc_3576_new_n267_; 
wire _abc_3576_new_n268_; 
wire _abc_3576_new_n269_; 
wire _abc_3576_new_n270_; 
wire _abc_3576_new_n271_; 
wire _abc_3576_new_n272_; 
wire _abc_3576_new_n273_; 
wire _abc_3576_new_n274_; 
wire _abc_3576_new_n275_; 
wire _abc_3576_new_n276_; 
wire _abc_3576_new_n277_; 
wire _abc_3576_new_n278_; 
wire _abc_3576_new_n279_; 
wire _abc_3576_new_n280_; 
wire _abc_3576_new_n281_; 
wire _abc_3576_new_n282_; 
wire _abc_3576_new_n283_; 
wire _abc_3576_new_n284_; 
wire _abc_3576_new_n285_; 
wire _abc_3576_new_n286_; 
wire _abc_3576_new_n287_; 
wire _abc_3576_new_n288_; 
wire _abc_3576_new_n289_; 
wire _abc_3576_new_n290_; 
wire _abc_3576_new_n291_; 
wire _abc_3576_new_n292_; 
wire _abc_3576_new_n293_; 
wire _abc_3576_new_n294_; 
wire _abc_3576_new_n295_; 
wire _abc_3576_new_n297_; 
wire _abc_3576_new_n298_; 
wire _abc_3576_new_n299_; 
wire _abc_3576_new_n300_; 
wire _abc_3576_new_n301_; 
wire _abc_3576_new_n302_; 
wire _abc_3576_new_n303_; 
wire _abc_3576_new_n304_; 
wire _abc_3576_new_n305_; 
wire _abc_3576_new_n306_; 
wire _abc_3576_new_n307_; 
wire _abc_3576_new_n308_; 
wire _abc_3576_new_n309_; 
wire _abc_3576_new_n310_; 
wire _abc_3576_new_n311_; 
wire _abc_3576_new_n312_; 
wire _abc_3576_new_n313_; 
wire _abc_3576_new_n314_; 
wire _abc_3576_new_n315_; 
wire _abc_3576_new_n316_; 
wire _abc_3576_new_n317_; 
wire _abc_3576_new_n318_; 
wire _abc_3576_new_n319_; 
wire _abc_3576_new_n320_; 
wire _abc_3576_new_n321_; 
wire _abc_3576_new_n322_; 
wire _abc_3576_new_n323_; 
wire _abc_3576_new_n324_; 
wire _abc_3576_new_n325_; 
wire _abc_3576_new_n326_; 
wire _abc_3576_new_n327_; 
wire _abc_3576_new_n328_; 
wire _abc_3576_new_n329_; 
wire _abc_3576_new_n330_; 
wire _abc_3576_new_n331_; 
wire _abc_3576_new_n333_; 
wire _abc_3576_new_n334_; 
wire _abc_3576_new_n335_; 
wire _abc_3576_new_n336_; 
wire _abc_3576_new_n337_; 
wire _abc_3576_new_n338_; 
wire _abc_3576_new_n339_; 
wire _abc_3576_new_n340_; 
wire _abc_3576_new_n341_; 
wire _abc_3576_new_n342_; 
wire _abc_3576_new_n343_; 
wire _abc_3576_new_n344_; 
wire _abc_3576_new_n345_; 
wire _abc_3576_new_n346_; 
wire _abc_3576_new_n347_; 
wire _abc_3576_new_n348_; 
wire _abc_3576_new_n349_; 
wire _abc_3576_new_n350_; 
wire _abc_3576_new_n351_; 
wire _abc_3576_new_n352_; 
wire _abc_3576_new_n353_; 
wire _abc_3576_new_n354_; 
wire _abc_3576_new_n355_; 
wire _abc_3576_new_n356_; 
wire _abc_3576_new_n357_; 
wire _abc_3576_new_n358_; 
wire _abc_3576_new_n359_; 
wire _abc_3576_new_n360_; 
wire _abc_3576_new_n361_; 
wire _abc_3576_new_n362_; 
wire _abc_3576_new_n363_; 
wire _abc_3576_new_n364_; 
wire _abc_3576_new_n365_; 
wire _abc_3576_new_n367_; 
wire _abc_3576_new_n368_; 
wire _abc_3576_new_n369_; 
wire _abc_3576_new_n370_; 
wire _abc_3576_new_n371_; 
wire _abc_3576_new_n372_; 
wire _abc_3576_new_n373_; 
wire _abc_3576_new_n374_; 
wire _abc_3576_new_n375_; 
wire _abc_3576_new_n376_; 
wire _abc_3576_new_n377_; 
wire _abc_3576_new_n378_; 
wire _abc_3576_new_n379_; 
wire _abc_3576_new_n380_; 
wire _abc_3576_new_n381_; 
wire _abc_3576_new_n382_; 
wire _abc_3576_new_n383_; 
wire _abc_3576_new_n384_; 
wire _abc_3576_new_n385_; 
wire _abc_3576_new_n386_; 
wire _abc_3576_new_n387_; 
wire _abc_3576_new_n388_; 
wire _abc_3576_new_n389_; 
wire _abc_3576_new_n390_; 
wire _abc_3576_new_n391_; 
wire _abc_3576_new_n392_; 
wire _abc_3576_new_n393_; 
wire _abc_3576_new_n394_; 
wire _abc_3576_new_n395_; 
wire _abc_3576_new_n396_; 
wire _abc_3576_new_n397_; 
wire _abc_3576_new_n398_; 
wire _abc_3576_new_n399_; 
wire _abc_3576_new_n400_; 
wire _abc_3576_new_n401_; 
wire _abc_3576_new_n402_; 
wire _abc_3576_new_n403_; 
wire _abc_3576_new_n404_; 
wire _abc_3576_new_n405_; 
wire _abc_3576_new_n406_; 
wire _abc_3576_new_n407_; 
wire _abc_3576_new_n408_; 
wire _abc_3576_new_n409_; 
wire _abc_3576_new_n410_; 
wire _abc_3576_new_n412_; 
wire _abc_3576_new_n413_; 
wire _abc_3576_new_n414_; 
wire _abc_3576_new_n415_; 
wire _abc_3576_new_n416_; 
wire _abc_3576_new_n417_; 
wire _abc_3576_new_n418_; 
wire _abc_3576_new_n419_; 
wire _abc_3576_new_n420_; 
wire _abc_3576_new_n421_; 
wire _abc_3576_new_n422_; 
wire _abc_3576_new_n423_; 
wire _abc_3576_new_n424_; 
wire _abc_3576_new_n425_; 
wire _abc_3576_new_n426_; 
wire _abc_3576_new_n427_; 
wire _abc_3576_new_n428_; 
wire _abc_3576_new_n429_; 
wire _abc_3576_new_n430_; 
wire _abc_3576_new_n431_; 
wire _abc_3576_new_n432_; 
wire _abc_3576_new_n433_; 
wire _abc_3576_new_n434_; 
wire _abc_3576_new_n435_; 
wire _abc_3576_new_n436_; 
wire _abc_3576_new_n437_; 
wire _abc_3576_new_n438_; 
wire _abc_3576_new_n439_; 
wire _abc_3576_new_n440_; 
wire _abc_3576_new_n441_; 
wire _abc_3576_new_n442_; 
wire _abc_3576_new_n443_; 
wire _abc_3576_new_n444_; 
wire _abc_3576_new_n445_; 
wire _abc_3576_new_n446_; 
wire _abc_3576_new_n447_; 
wire _abc_3576_new_n448_; 
wire _abc_3576_new_n449_; 
wire _abc_3576_new_n451_; 
wire _abc_3576_new_n452_; 
wire _abc_3576_new_n453_; 
wire _abc_3576_new_n454_; 
wire _abc_3576_new_n455_; 
wire _abc_3576_new_n456_; 
wire _abc_3576_new_n457_; 
wire _abc_3576_new_n458_; 
wire _abc_3576_new_n459_; 
wire _abc_3576_new_n460_; 
wire _abc_3576_new_n461_; 
wire _abc_3576_new_n462_; 
wire _abc_3576_new_n463_; 
wire _abc_3576_new_n464_; 
wire _abc_3576_new_n465_; 
wire _abc_3576_new_n466_; 
wire _abc_3576_new_n467_; 
wire _abc_3576_new_n468_; 
wire _abc_3576_new_n469_; 
wire _abc_3576_new_n470_; 
wire _abc_3576_new_n471_; 
wire _abc_3576_new_n472_; 
wire _abc_3576_new_n473_; 
wire _abc_3576_new_n474_; 
wire _abc_3576_new_n475_; 
wire _abc_3576_new_n476_; 
wire _abc_3576_new_n477_; 
wire _abc_3576_new_n478_; 
wire _abc_3576_new_n479_; 
wire _abc_3576_new_n480_; 
wire _abc_3576_new_n481_; 
wire _abc_3576_new_n482_; 
wire _abc_3576_new_n483_; 
wire _abc_3576_new_n484_; 
wire _abc_3576_new_n485_; 
wire _abc_3576_new_n486_; 
wire _abc_3576_new_n487_; 
wire _abc_3576_new_n488_; 
wire _abc_3576_new_n489_; 
wire _abc_3576_new_n491_; 
wire _abc_3576_new_n492_; 
wire _abc_3576_new_n493_; 
wire _abc_3576_new_n494_; 
wire _abc_3576_new_n495_; 
wire _abc_3576_new_n496_; 
wire _abc_3576_new_n497_; 
wire _abc_3576_new_n498_; 
wire _abc_3576_new_n499_; 
wire _abc_3576_new_n501_; 
wire _abc_3576_new_n502_; 
wire _abc_3576_new_n503_; 
wire _abc_3576_new_n504_; 
wire _abc_3576_new_n505_; 
wire _abc_3576_new_n507_; 
wire _abc_3576_new_n508_; 
wire _abc_3576_new_n509_; 
wire _abc_3576_new_n511_; 
wire _abc_3576_new_n512_; 
wire _abc_3576_new_n513_; 
wire _abc_3576_new_n515_; 
wire _abc_3576_new_n516_; 
wire _abc_3576_new_n517_; 
wire _abc_3576_new_n519_; 
wire _abc_3576_new_n520_; 
wire _abc_3576_new_n521_; 
wire _abc_3576_new_n523_; 
wire _abc_3576_new_n524_; 
wire _abc_3576_new_n525_; 
wire _abc_3576_new_n527_; 
wire _abc_3576_new_n528_; 
wire _abc_3576_new_n529_; 
wire _abc_3576_new_n531_; 
wire _abc_3576_new_n532_; 
wire _abc_3576_new_n533_; 
wire _abc_3576_new_n535_; 
wire _abc_3576_new_n536_; 
wire _abc_3576_new_n537_; 
wire _abc_3576_new_n539_; 
wire _abc_3576_new_n540_; 
wire _abc_3576_new_n541_; 
wire _abc_3576_new_n543_; 
wire _abc_3576_new_n544_; 
wire _abc_3576_new_n545_; 
wire _abc_3576_new_n547_; 
wire _abc_3576_new_n548_; 
wire _abc_3576_new_n549_; 
wire _abc_3576_new_n551_; 
wire _abc_3576_new_n552_; 
wire _abc_3576_new_n553_; 
wire _abc_3576_new_n555_; 
wire _abc_3576_new_n556_; 
wire _abc_3576_new_n557_; 
wire _abc_3576_new_n559_; 
wire _abc_3576_new_n560_; 
wire _abc_3576_new_n561_; 
wire _abc_3576_new_n563_; 
wire _abc_3576_new_n564_; 
wire _abc_3576_new_n565_; 
wire _abc_3576_new_n567_; 
wire _abc_3576_new_n568_; 
wire _abc_3576_new_n569_; 
wire _abc_3576_new_n571_; 
wire _abc_3576_new_n572_; 
wire _abc_3576_new_n573_; 
wire _abc_3576_new_n575_; 
wire _abc_3576_new_n576_; 
wire _abc_3576_new_n577_; 
wire _abc_3576_new_n579_; 
wire _abc_3576_new_n580_; 
wire _abc_3576_new_n581_; 
wire _abc_3576_new_n583_; 
wire _abc_3576_new_n584_; 
wire _abc_3576_new_n585_; 
wire _abc_3576_new_n587_; 
wire _abc_3576_new_n588_; 
wire _abc_3576_new_n589_; 
wire _abc_3576_new_n591_; 
wire _abc_3576_new_n592_; 
wire _abc_3576_new_n593_; 
wire _abc_3576_new_n595_; 
wire _abc_3576_new_n596_; 
wire _abc_3576_new_n597_; 
wire _abc_3576_new_n599_; 
wire _abc_3576_new_n600_; 
wire _abc_3576_new_n601_; 
wire _abc_3576_new_n603_; 
wire _abc_3576_new_n604_; 
wire _abc_3576_new_n605_; 
wire _abc_3576_new_n607_; 
wire _abc_3576_new_n608_; 
wire _abc_3576_new_n609_; 
wire _abc_3576_new_n611_; 
wire _abc_3576_new_n612_; 
wire _abc_3576_new_n613_; 
wire _abc_3576_new_n615_; 
wire _abc_3576_new_n616_; 
wire _abc_3576_new_n617_; 
wire _abc_3576_new_n619_; 
wire _abc_3576_new_n620_; 
wire _abc_3576_new_n621_; 
wire _abc_3576_new_n623_; 
wire _abc_3576_new_n624_; 
wire _abc_3576_new_n625_; 
wire _abc_3576_new_n627_; 
wire _abc_3576_new_n628_; 
wire _abc_3576_new_n629_; 
wire _abc_3576_new_n631_; 
wire _abc_3576_new_n632_; 
wire _abc_3576_new_n633_; 
wire _abc_3576_new_n635_; 
wire _abc_3576_new_n636_; 
wire _abc_3576_new_n637_; 
wire _abc_3576_new_n638_; 
wire _abc_3576_new_n639_; 
wire _abc_3576_new_n640_; 
wire _abc_3576_new_n641_; 
wire _abc_3576_new_n642_; 
wire _abc_3576_new_n644_; 
wire _abc_3576_new_n645_; 
wire _abc_3576_new_n646_; 
wire _abc_3576_new_n648_; 
wire _abc_3576_new_n649_; 
wire _abc_3576_new_n650_; 
wire _abc_3576_new_n652_; 
wire _abc_3576_new_n653_; 
wire _abc_3576_new_n654_; 
wire _abc_3576_new_n656_; 
wire _abc_3576_new_n657_; 
wire _abc_3576_new_n658_; 
wire _abc_3576_new_n660_; 
wire _abc_3576_new_n661_; 
wire _abc_3576_new_n662_; 
wire _abc_3576_new_n664_; 
wire _abc_3576_new_n665_; 
wire _abc_3576_new_n666_; 
wire _abc_3576_new_n668_; 
wire _abc_3576_new_n669_; 
wire _abc_3576_new_n670_; 
wire _abc_3576_new_n672_; 
wire _abc_3576_new_n673_; 
wire _abc_3576_new_n674_; 
wire _abc_3576_new_n675_; 
wire _abc_3576_new_n676_; 
wire _abc_3576_new_n677_; 
wire _abc_3576_new_n678_; 
wire _abc_3576_new_n679_; 
wire _abc_3576_new_n680_; 
wire _abc_3576_new_n681_; 
wire _abc_3576_new_n682_; 
wire _abc_3576_new_n683_; 
wire _abc_3576_new_n684_; 
wire _abc_3576_new_n685_; 
wire _abc_3576_new_n686_; 
wire _abc_3576_new_n687_; 
wire _abc_3576_new_n688_; 
wire _abc_3576_new_n689_; 
wire _abc_3576_new_n690_; 
wire _abc_3576_new_n691_; 
wire _abc_3576_new_n692_; 
wire _abc_3576_new_n693_; 
wire _abc_3576_new_n694_; 
wire _abc_3576_new_n695_; 
wire _abc_3576_new_n696_; 
wire _abc_3576_new_n697_; 
wire _abc_3576_new_n698_; 
wire _abc_3576_new_n699_; 
wire _abc_3576_new_n700_; 
wire _abc_3576_new_n701_; 
wire _abc_3576_new_n702_; 
wire _abc_3576_new_n703_; 
wire _abc_3576_new_n704_; 
wire _abc_3576_new_n705_; 
wire _abc_3576_new_n706_; 
wire _abc_3576_new_n707_; 
wire _abc_3576_new_n708_; 
wire _abc_3576_new_n709_; 
wire _abc_3576_new_n710_; 
wire _abc_3576_new_n711_; 
wire _abc_3576_new_n712_; 
wire _abc_3576_new_n713_; 
wire _abc_3576_new_n714_; 
wire _abc_3576_new_n715_; 
wire _abc_3576_new_n716_; 
wire _abc_3576_new_n717_; 
wire _abc_3576_new_n718_; 
wire _abc_3576_new_n719_; 
wire _abc_3576_new_n720_; 
wire _abc_3576_new_n721_; 
wire _abc_3576_new_n722_; 
wire _abc_3576_new_n723_; 
wire _abc_3576_new_n724_; 
wire _abc_3576_new_n725_; 
wire _abc_3576_new_n726_; 
wire _abc_3576_new_n727_; 
wire _abc_3576_new_n728_; 
wire _abc_3576_new_n729_; 
wire _abc_3576_new_n730_; 
wire _abc_3576_new_n731_; 
wire _abc_3576_new_n732_; 
wire _abc_3576_new_n733_; 
wire _abc_3576_new_n734_; 
wire _abc_3576_new_n735_; 
wire _abc_3576_new_n736_; 
wire _abc_3576_new_n737_; 
wire _abc_3576_new_n738_; 
wire _abc_3576_new_n739_; 
wire _abc_3576_new_n740_; 
wire _abc_3576_new_n741_; 
wire _abc_3576_new_n742_; 
wire _abc_3576_new_n743_; 
wire _abc_3576_new_n744_; 
wire _abc_3576_new_n745_; 
wire _abc_3576_new_n746_; 
wire _abc_3576_new_n747_; 
wire _abc_3576_new_n748_; 
wire _abc_3576_new_n749_; 
wire _abc_3576_new_n750_; 
wire _abc_3576_new_n751_; 
wire _abc_3576_new_n752_; 
wire _abc_3576_new_n753_; 
wire _abc_3576_new_n754_; 
wire _abc_3576_new_n756_; 
wire _abc_3576_new_n757_; 
wire _abc_3576_new_n758_; 
wire _abc_3576_new_n760_; 
wire _abc_3576_new_n761_; 
wire _abc_3576_new_n762_; 
wire _abc_3576_new_n764_; 
wire _abc_3576_new_n765_; 
wire _abc_3576_new_n766_; 
wire _abc_3576_new_n768_; 
wire _abc_3576_new_n769_; 
wire _abc_3576_new_n770_; 
wire _abc_3576_new_n772_; 
wire _abc_3576_new_n773_; 
wire _abc_3576_new_n774_; 
wire _abc_3576_new_n776_; 
wire _abc_3576_new_n777_; 
wire _abc_3576_new_n778_; 
wire _abc_3576_new_n780_; 
wire _abc_3576_new_n781_; 
wire _abc_3576_new_n782_; 
wire _abc_3576_new_n784_; 
wire _abc_3576_new_n785_; 
wire _abc_3576_new_n786_; 
wire _abc_3576_new_n787_; 
wire _abc_3576_new_n788_; 
wire _abc_3576_new_n789_; 
wire _abc_3576_new_n791_; 
wire _abc_3576_new_n792_; 
wire _abc_3576_new_n793_; 
wire _abc_3576_new_n795_; 
wire _abc_3576_new_n796_; 
wire _abc_3576_new_n797_; 
wire _abc_3576_new_n799_; 
wire _abc_3576_new_n800_; 
wire _abc_3576_new_n801_; 
wire _abc_3576_new_n803_; 
wire _abc_3576_new_n804_; 
wire _abc_3576_new_n805_; 
wire _abc_3576_new_n807_; 
wire _abc_3576_new_n808_; 
wire _abc_3576_new_n809_; 
wire _abc_3576_new_n811_; 
wire _abc_3576_new_n812_; 
wire _abc_3576_new_n813_; 
wire _abc_3576_new_n815_; 
wire _abc_3576_new_n816_; 
wire _abc_3576_new_n817_; 
wire _abc_3576_new_n819_; 
input clock;
wire n104; 
wire n109; 
wire n114; 
wire n119; 
wire n124; 
wire n129; 
wire n134; 
wire n139; 
wire n144; 
wire n149; 
wire n154; 
wire n159; 
wire n164; 
wire n169; 
wire n174; 
wire n179; 
wire n184; 
wire n189; 
wire n194; 
wire n199; 
wire n204; 
wire n209; 
wire n214; 
wire n219; 
wire n224; 
wire n229; 
wire n234; 
wire n239; 
wire n244; 
wire n249; 
wire n254; 
wire n259; 
wire n264; 
wire n269; 
wire n274; 
wire n279; 
wire n284; 
wire n289; 
wire n294; 
wire n299; 
wire n304; 
wire n309; 
wire n314; 
wire n319; 
wire n324; 
wire n328; 
wire n332; 
wire n336; 
wire n340; 
wire n344; 
wire n348; 
wire n352; 
wire n356; 
wire n361; 
wire n44; 
wire n49; 
wire n54; 
wire n59; 
wire n64; 
wire n69; 
wire n74; 
wire n79; 
wire n84; 
wire n89; 
wire n94; 
wire n99; 
input nRESET_G;
AND2X2 AND2X2_1 ( .A(_abc_3576_new_n146_), .B(STATO_REG_1_), .Y(_abc_3576_new_n147_));
AND2X2 AND2X2_10 ( .A(_abc_3576_new_n166_), .B(_abc_3576_new_n170_), .Y(_abc_3576_new_n171_));
AND2X2 AND2X2_100 ( .A(_abc_3576_new_n290_), .B(DATA_OUT_REG_2_), .Y(_abc_3576_new_n361_));
AND2X2 AND2X2_101 ( .A(_abc_3576_new_n200_), .B(_abc_3576_new_n317_), .Y(_abc_3576_new_n367_));
AND2X2 AND2X2_102 ( .A(_abc_3576_new_n355_), .B(_abc_3576_new_n367_), .Y(_abc_3576_new_n368_));
AND2X2 AND2X2_103 ( .A(_abc_3576_new_n352_), .B(_abc_3576_new_n319_), .Y(_abc_3576_new_n369_));
AND2X2 AND2X2_104 ( .A(_abc_3576_new_n371_), .B(_abc_3576_new_n344_), .Y(_abc_3576_new_n372_));
AND2X2 AND2X2_105 ( .A(_abc_3576_new_n374_), .B(_abc_3576_new_n373_), .Y(_abc_3576_new_n375_));
AND2X2 AND2X2_106 ( .A(_abc_3576_new_n377_), .B(_abc_3576_new_n376_), .Y(_abc_3576_new_n378_));
AND2X2 AND2X2_107 ( .A(_abc_3576_new_n375_), .B(_abc_3576_new_n378_), .Y(_abc_3576_new_n379_));
AND2X2 AND2X2_108 ( .A(_abc_3576_new_n380_), .B(_abc_3576_new_n381_), .Y(_abc_3576_new_n382_));
AND2X2 AND2X2_109 ( .A(_abc_3576_new_n372_), .B(_abc_3576_new_n383_), .Y(_abc_3576_new_n384_));
AND2X2 AND2X2_11 ( .A(_abc_3576_new_n172_), .B(_abc_3576_new_n161_), .Y(_abc_3576_new_n173_));
AND2X2 AND2X2_110 ( .A(_abc_3576_new_n385_), .B(_abc_3576_new_n172_), .Y(_abc_3576_new_n386_));
AND2X2 AND2X2_111 ( .A(_abc_3576_new_n386_), .B(_abc_3576_new_n308_), .Y(_abc_3576_new_n387_));
AND2X2 AND2X2_112 ( .A(_abc_3576_new_n388_), .B(_abc_3576_new_n342_), .Y(_abc_3576_new_n389_));
AND2X2 AND2X2_113 ( .A(_abc_3576_new_n390_), .B(_abc_3576_new_n382_), .Y(_abc_3576_new_n391_));
AND2X2 AND2X2_114 ( .A(_abc_3576_new_n368_), .B(_abc_3576_new_n392_), .Y(_abc_3576_new_n395_));
AND2X2 AND2X2_115 ( .A(_abc_3576_new_n396_), .B(_abc_3576_new_n393_), .Y(_abc_3576_new_n397_));
AND2X2 AND2X2_116 ( .A(_abc_3576_new_n398_), .B(_abc_3576_new_n370_), .Y(_abc_3576_new_n399_));
AND2X2 AND2X2_117 ( .A(_abc_3576_new_n400_), .B(_abc_3576_new_n394_), .Y(_abc_3576_new_n401_));
AND2X2 AND2X2_118 ( .A(_abc_3576_new_n401_), .B(_abc_3576_new_n275_), .Y(_abc_3576_new_n402_));
AND2X2 AND2X2_119 ( .A(_abc_3576_new_n286_), .B(REG4_REG_3_), .Y(_abc_3576_new_n403_));
AND2X2 AND2X2_12 ( .A(_abc_3576_new_n175_), .B(_abc_3576_new_n174_), .Y(_abc_3576_new_n176_));
AND2X2 AND2X2_120 ( .A(_abc_3576_new_n288_), .B(RLAST_REG_3_), .Y(_abc_3576_new_n404_));
AND2X2 AND2X2_121 ( .A(_abc_3576_new_n290_), .B(DATA_OUT_REG_3_), .Y(_abc_3576_new_n405_));
AND2X2 AND2X2_122 ( .A(_abc_3576_new_n393_), .B(_abc_3576_new_n282_), .Y(_abc_3576_new_n409_));
AND2X2 AND2X2_123 ( .A(_abc_3576_new_n413_), .B(_abc_3576_new_n412_), .Y(_abc_3576_new_n414_));
AND2X2 AND2X2_124 ( .A(_abc_3576_new_n416_), .B(_abc_3576_new_n415_), .Y(_abc_3576_new_n417_));
AND2X2 AND2X2_125 ( .A(_abc_3576_new_n414_), .B(_abc_3576_new_n417_), .Y(_abc_3576_new_n418_));
AND2X2 AND2X2_126 ( .A(_abc_3576_new_n419_), .B(_abc_3576_new_n420_), .Y(_abc_3576_new_n421_));
AND2X2 AND2X2_127 ( .A(_abc_3576_new_n424_), .B(_abc_3576_new_n380_), .Y(_abc_3576_new_n425_));
AND2X2 AND2X2_128 ( .A(_abc_3576_new_n425_), .B(_abc_3576_new_n422_), .Y(_abc_3576_new_n426_));
AND2X2 AND2X2_129 ( .A(_abc_3576_new_n390_), .B(_abc_3576_new_n381_), .Y(_abc_3576_new_n427_));
AND2X2 AND2X2_13 ( .A(_abc_3576_new_n154_), .B(REG4_REG_0_), .Y(_abc_3576_new_n177_));
AND2X2 AND2X2_130 ( .A(_abc_3576_new_n428_), .B(_abc_3576_new_n421_), .Y(_abc_3576_new_n429_));
AND2X2 AND2X2_131 ( .A(_abc_3576_new_n430_), .B(_abc_3576_new_n395_), .Y(_abc_3576_new_n431_));
AND2X2 AND2X2_132 ( .A(_abc_3576_new_n432_), .B(_abc_3576_new_n433_), .Y(_abc_3576_new_n434_));
AND2X2 AND2X2_133 ( .A(_abc_3576_new_n435_), .B(_abc_3576_new_n399_), .Y(_abc_3576_new_n437_));
AND2X2 AND2X2_134 ( .A(_abc_3576_new_n438_), .B(_abc_3576_new_n275_), .Y(_abc_3576_new_n439_));
AND2X2 AND2X2_135 ( .A(_abc_3576_new_n439_), .B(_abc_3576_new_n436_), .Y(_abc_3576_new_n440_));
AND2X2 AND2X2_136 ( .A(_abc_3576_new_n441_), .B(_abc_3576_new_n282_), .Y(_abc_3576_new_n442_));
AND2X2 AND2X2_137 ( .A(_abc_3576_new_n288_), .B(RLAST_REG_4_), .Y(_abc_3576_new_n443_));
AND2X2 AND2X2_138 ( .A(_abc_3576_new_n286_), .B(REG4_REG_4_), .Y(_abc_3576_new_n444_));
AND2X2 AND2X2_139 ( .A(_abc_3576_new_n290_), .B(DATA_OUT_REG_4_), .Y(_abc_3576_new_n445_));
AND2X2 AND2X2_14 ( .A(RMIN_REG_0_), .B(RESTART), .Y(_abc_3576_new_n178_));
AND2X2 AND2X2_140 ( .A(_abc_3576_new_n452_), .B(_abc_3576_new_n419_), .Y(_abc_3576_new_n453_));
AND2X2 AND2X2_141 ( .A(_abc_3576_new_n455_), .B(_abc_3576_new_n454_), .Y(_abc_3576_new_n456_));
AND2X2 AND2X2_142 ( .A(_abc_3576_new_n459_), .B(_abc_3576_new_n458_), .Y(_abc_3576_new_n460_));
AND2X2 AND2X2_143 ( .A(_abc_3576_new_n457_), .B(_abc_3576_new_n460_), .Y(_abc_3576_new_n461_));
AND2X2 AND2X2_144 ( .A(_abc_3576_new_n453_), .B(_abc_3576_new_n465_), .Y(_abc_3576_new_n466_));
AND2X2 AND2X2_145 ( .A(_abc_3576_new_n428_), .B(_abc_3576_new_n420_), .Y(_abc_3576_new_n467_));
AND2X2 AND2X2_146 ( .A(_abc_3576_new_n468_), .B(_abc_3576_new_n464_), .Y(_abc_3576_new_n469_));
AND2X2 AND2X2_147 ( .A(_abc_3576_new_n473_), .B(_abc_3576_new_n472_), .Y(_abc_3576_new_n474_));
AND2X2 AND2X2_148 ( .A(_abc_3576_new_n471_), .B(_abc_3576_new_n475_), .Y(_abc_3576_new_n476_));
AND2X2 AND2X2_149 ( .A(_abc_3576_new_n479_), .B(_abc_3576_new_n275_), .Y(_abc_3576_new_n480_));
AND2X2 AND2X2_15 ( .A(_abc_3576_new_n176_), .B(_abc_3576_new_n179_), .Y(_abc_3576_new_n180_));
AND2X2 AND2X2_150 ( .A(_abc_3576_new_n480_), .B(_abc_3576_new_n478_), .Y(_abc_3576_new_n481_));
AND2X2 AND2X2_151 ( .A(_abc_3576_new_n474_), .B(_abc_3576_new_n282_), .Y(_abc_3576_new_n482_));
AND2X2 AND2X2_152 ( .A(_abc_3576_new_n288_), .B(RLAST_REG_5_), .Y(_abc_3576_new_n483_));
AND2X2 AND2X2_153 ( .A(_abc_3576_new_n286_), .B(REG4_REG_5_), .Y(_abc_3576_new_n484_));
AND2X2 AND2X2_154 ( .A(_abc_3576_new_n290_), .B(DATA_OUT_REG_5_), .Y(_abc_3576_new_n485_));
AND2X2 AND2X2_155 ( .A(_abc_3576_new_n286_), .B(REG4_REG_6_), .Y(_abc_3576_new_n491_));
AND2X2 AND2X2_156 ( .A(_abc_3576_new_n288_), .B(RLAST_REG_6_), .Y(_abc_3576_new_n492_));
AND2X2 AND2X2_157 ( .A(_abc_3576_new_n290_), .B(DATA_OUT_REG_6_), .Y(_abc_3576_new_n493_));
AND2X2 AND2X2_158 ( .A(_abc_3576_new_n474_), .B(_abc_3576_new_n432_), .Y(_abc_3576_new_n497_));
AND2X2 AND2X2_159 ( .A(_abc_3576_new_n497_), .B(_abc_3576_new_n275_), .Y(_abc_3576_new_n498_));
AND2X2 AND2X2_16 ( .A(_abc_3576_new_n154_), .B(_abc_3576_new_n181_), .Y(_abc_3576_new_n182_));
AND2X2 AND2X2_160 ( .A(_abc_3576_new_n437_), .B(_abc_3576_new_n498_), .Y(_abc_3576_new_n499_));
AND2X2 AND2X2_161 ( .A(_abc_3576_new_n286_), .B(REG4_REG_7_), .Y(_abc_3576_new_n501_));
AND2X2 AND2X2_162 ( .A(_abc_3576_new_n288_), .B(RLAST_REG_7_), .Y(_abc_3576_new_n502_));
AND2X2 AND2X2_163 ( .A(_abc_3576_new_n290_), .B(DATA_OUT_REG_7_), .Y(_abc_3576_new_n503_));
AND2X2 AND2X2_164 ( .A(_abc_3576_new_n290_), .B(REG4_REG_0_), .Y(_abc_3576_new_n507_));
AND2X2 AND2X2_165 ( .A(_abc_3576_new_n147_), .B(REG3_REG_0_), .Y(_abc_3576_new_n508_));
AND2X2 AND2X2_166 ( .A(_abc_3576_new_n290_), .B(REG4_REG_1_), .Y(_abc_3576_new_n511_));
AND2X2 AND2X2_167 ( .A(_abc_3576_new_n147_), .B(REG3_REG_1_), .Y(_abc_3576_new_n512_));
AND2X2 AND2X2_168 ( .A(_abc_3576_new_n290_), .B(REG4_REG_2_), .Y(_abc_3576_new_n515_));
AND2X2 AND2X2_169 ( .A(_abc_3576_new_n147_), .B(REG3_REG_2_), .Y(_abc_3576_new_n516_));
AND2X2 AND2X2_17 ( .A(_abc_3576_new_n183_), .B(RESTART), .Y(_abc_3576_new_n184_));
AND2X2 AND2X2_170 ( .A(_abc_3576_new_n290_), .B(REG4_REG_3_), .Y(_abc_3576_new_n519_));
AND2X2 AND2X2_171 ( .A(_abc_3576_new_n147_), .B(REG3_REG_3_), .Y(_abc_3576_new_n520_));
AND2X2 AND2X2_172 ( .A(_abc_3576_new_n290_), .B(REG4_REG_4_), .Y(_abc_3576_new_n523_));
AND2X2 AND2X2_173 ( .A(_abc_3576_new_n147_), .B(REG3_REG_4_), .Y(_abc_3576_new_n524_));
AND2X2 AND2X2_174 ( .A(_abc_3576_new_n290_), .B(REG4_REG_5_), .Y(_abc_3576_new_n527_));
AND2X2 AND2X2_175 ( .A(_abc_3576_new_n147_), .B(REG3_REG_5_), .Y(_abc_3576_new_n528_));
AND2X2 AND2X2_176 ( .A(_abc_3576_new_n290_), .B(REG4_REG_6_), .Y(_abc_3576_new_n531_));
AND2X2 AND2X2_177 ( .A(_abc_3576_new_n147_), .B(REG3_REG_6_), .Y(_abc_3576_new_n532_));
AND2X2 AND2X2_178 ( .A(_abc_3576_new_n290_), .B(REG4_REG_7_), .Y(_abc_3576_new_n535_));
AND2X2 AND2X2_179 ( .A(_abc_3576_new_n147_), .B(REG3_REG_7_), .Y(_abc_3576_new_n536_));
AND2X2 AND2X2_18 ( .A(_abc_3576_new_n187_), .B(_abc_3576_new_n188_), .Y(_abc_3576_new_n189_));
AND2X2 AND2X2_180 ( .A(_abc_3576_new_n290_), .B(REG3_REG_0_), .Y(_abc_3576_new_n539_));
AND2X2 AND2X2_181 ( .A(_abc_3576_new_n147_), .B(REG2_REG_0_), .Y(_abc_3576_new_n540_));
AND2X2 AND2X2_182 ( .A(_abc_3576_new_n290_), .B(REG3_REG_1_), .Y(_abc_3576_new_n543_));
AND2X2 AND2X2_183 ( .A(_abc_3576_new_n147_), .B(REG2_REG_1_), .Y(_abc_3576_new_n544_));
AND2X2 AND2X2_184 ( .A(_abc_3576_new_n290_), .B(REG3_REG_2_), .Y(_abc_3576_new_n547_));
AND2X2 AND2X2_185 ( .A(_abc_3576_new_n147_), .B(REG2_REG_2_), .Y(_abc_3576_new_n548_));
AND2X2 AND2X2_186 ( .A(_abc_3576_new_n290_), .B(REG3_REG_3_), .Y(_abc_3576_new_n551_));
AND2X2 AND2X2_187 ( .A(_abc_3576_new_n147_), .B(REG2_REG_3_), .Y(_abc_3576_new_n552_));
AND2X2 AND2X2_188 ( .A(_abc_3576_new_n290_), .B(REG3_REG_4_), .Y(_abc_3576_new_n555_));
AND2X2 AND2X2_189 ( .A(_abc_3576_new_n147_), .B(REG2_REG_4_), .Y(_abc_3576_new_n556_));
AND2X2 AND2X2_19 ( .A(_abc_3576_new_n185_), .B(_abc_3576_new_n189_), .Y(_abc_3576_new_n190_));
AND2X2 AND2X2_190 ( .A(_abc_3576_new_n290_), .B(REG3_REG_5_), .Y(_abc_3576_new_n559_));
AND2X2 AND2X2_191 ( .A(_abc_3576_new_n147_), .B(REG2_REG_5_), .Y(_abc_3576_new_n560_));
AND2X2 AND2X2_192 ( .A(_abc_3576_new_n290_), .B(REG3_REG_6_), .Y(_abc_3576_new_n563_));
AND2X2 AND2X2_193 ( .A(_abc_3576_new_n147_), .B(REG2_REG_6_), .Y(_abc_3576_new_n564_));
AND2X2 AND2X2_194 ( .A(_abc_3576_new_n290_), .B(REG3_REG_7_), .Y(_abc_3576_new_n567_));
AND2X2 AND2X2_195 ( .A(_abc_3576_new_n147_), .B(REG2_REG_7_), .Y(_abc_3576_new_n568_));
AND2X2 AND2X2_196 ( .A(_abc_3576_new_n290_), .B(REG2_REG_0_), .Y(_abc_3576_new_n571_));
AND2X2 AND2X2_197 ( .A(_abc_3576_new_n147_), .B(REG1_REG_0_), .Y(_abc_3576_new_n572_));
AND2X2 AND2X2_198 ( .A(_abc_3576_new_n290_), .B(REG2_REG_1_), .Y(_abc_3576_new_n575_));
AND2X2 AND2X2_199 ( .A(_abc_3576_new_n147_), .B(REG1_REG_1_), .Y(_abc_3576_new_n576_));
AND2X2 AND2X2_2 ( .A(_abc_3576_new_n149_), .B(STATO_REG_0_), .Y(_abc_3576_new_n150_));
AND2X2 AND2X2_20 ( .A(_abc_3576_new_n192_), .B(_abc_3576_new_n173_), .Y(_abc_3576_new_n193_));
AND2X2 AND2X2_200 ( .A(_abc_3576_new_n290_), .B(REG2_REG_2_), .Y(_abc_3576_new_n579_));
AND2X2 AND2X2_201 ( .A(_abc_3576_new_n147_), .B(REG1_REG_2_), .Y(_abc_3576_new_n580_));
AND2X2 AND2X2_202 ( .A(_abc_3576_new_n290_), .B(REG2_REG_3_), .Y(_abc_3576_new_n583_));
AND2X2 AND2X2_203 ( .A(_abc_3576_new_n147_), .B(REG1_REG_3_), .Y(_abc_3576_new_n584_));
AND2X2 AND2X2_204 ( .A(_abc_3576_new_n290_), .B(REG2_REG_4_), .Y(_abc_3576_new_n587_));
AND2X2 AND2X2_205 ( .A(_abc_3576_new_n147_), .B(REG1_REG_4_), .Y(_abc_3576_new_n588_));
AND2X2 AND2X2_206 ( .A(_abc_3576_new_n290_), .B(REG2_REG_5_), .Y(_abc_3576_new_n591_));
AND2X2 AND2X2_207 ( .A(_abc_3576_new_n147_), .B(REG1_REG_5_), .Y(_abc_3576_new_n592_));
AND2X2 AND2X2_208 ( .A(_abc_3576_new_n290_), .B(REG2_REG_6_), .Y(_abc_3576_new_n595_));
AND2X2 AND2X2_209 ( .A(_abc_3576_new_n147_), .B(REG1_REG_6_), .Y(_abc_3576_new_n596_));
AND2X2 AND2X2_21 ( .A(_abc_3576_new_n196_), .B(_abc_3576_new_n198_), .Y(_abc_3576_new_n199_));
AND2X2 AND2X2_210 ( .A(_abc_3576_new_n290_), .B(REG2_REG_7_), .Y(_abc_3576_new_n599_));
AND2X2 AND2X2_211 ( .A(_abc_3576_new_n147_), .B(REG1_REG_7_), .Y(_abc_3576_new_n600_));
AND2X2 AND2X2_212 ( .A(_abc_3576_new_n290_), .B(REG1_REG_0_), .Y(_abc_3576_new_n603_));
AND2X2 AND2X2_213 ( .A(_abc_3576_new_n147_), .B(DATA_IN_0_), .Y(_abc_3576_new_n604_));
AND2X2 AND2X2_214 ( .A(_abc_3576_new_n290_), .B(REG1_REG_1_), .Y(_abc_3576_new_n607_));
AND2X2 AND2X2_215 ( .A(_abc_3576_new_n147_), .B(DATA_IN_1_), .Y(_abc_3576_new_n608_));
AND2X2 AND2X2_216 ( .A(_abc_3576_new_n290_), .B(REG1_REG_2_), .Y(_abc_3576_new_n611_));
AND2X2 AND2X2_217 ( .A(_abc_3576_new_n147_), .B(DATA_IN_2_), .Y(_abc_3576_new_n612_));
AND2X2 AND2X2_218 ( .A(_abc_3576_new_n290_), .B(REG1_REG_3_), .Y(_abc_3576_new_n615_));
AND2X2 AND2X2_219 ( .A(_abc_3576_new_n147_), .B(DATA_IN_3_), .Y(_abc_3576_new_n616_));
AND2X2 AND2X2_22 ( .A(_abc_3576_new_n199_), .B(_abc_3576_new_n191_), .Y(_abc_3576_new_n200_));
AND2X2 AND2X2_220 ( .A(_abc_3576_new_n290_), .B(REG1_REG_4_), .Y(_abc_3576_new_n619_));
AND2X2 AND2X2_221 ( .A(_abc_3576_new_n147_), .B(DATA_IN_4_), .Y(_abc_3576_new_n620_));
AND2X2 AND2X2_222 ( .A(_abc_3576_new_n290_), .B(REG1_REG_5_), .Y(_abc_3576_new_n623_));
AND2X2 AND2X2_223 ( .A(_abc_3576_new_n147_), .B(DATA_IN_5_), .Y(_abc_3576_new_n624_));
AND2X2 AND2X2_224 ( .A(_abc_3576_new_n290_), .B(REG1_REG_6_), .Y(_abc_3576_new_n627_));
AND2X2 AND2X2_225 ( .A(_abc_3576_new_n147_), .B(DATA_IN_6_), .Y(_abc_3576_new_n628_));
AND2X2 AND2X2_226 ( .A(_abc_3576_new_n290_), .B(REG1_REG_7_), .Y(_abc_3576_new_n631_));
AND2X2 AND2X2_227 ( .A(_abc_3576_new_n147_), .B(DATA_IN_7_), .Y(_abc_3576_new_n632_));
AND2X2 AND2X2_228 ( .A(_abc_3576_new_n146_), .B(_abc_3576_new_n269_), .Y(_abc_3576_new_n635_));
AND2X2 AND2X2_229 ( .A(_abc_3576_new_n636_), .B(STATO_REG_1_), .Y(_abc_3576_new_n637_));
AND2X2 AND2X2_23 ( .A(_abc_3576_new_n201_), .B(_abc_3576_new_n194_), .Y(_abc_3576_new_n202_));
AND2X2 AND2X2_230 ( .A(_abc_3576_new_n637_), .B(DATA_IN_0_), .Y(_abc_3576_new_n638_));
AND2X2 AND2X2_231 ( .A(_abc_3576_new_n149_), .B(_abc_3576_new_n146_), .Y(_abc_3576_new_n639_));
AND2X2 AND2X2_232 ( .A(_abc_3576_new_n640_), .B(RLAST_REG_0_), .Y(_abc_3576_new_n641_));
AND2X2 AND2X2_233 ( .A(_abc_3576_new_n637_), .B(DATA_IN_1_), .Y(_abc_3576_new_n644_));
AND2X2 AND2X2_234 ( .A(_abc_3576_new_n640_), .B(RLAST_REG_1_), .Y(_abc_3576_new_n645_));
AND2X2 AND2X2_235 ( .A(_abc_3576_new_n637_), .B(DATA_IN_2_), .Y(_abc_3576_new_n648_));
AND2X2 AND2X2_236 ( .A(_abc_3576_new_n640_), .B(RLAST_REG_2_), .Y(_abc_3576_new_n649_));
AND2X2 AND2X2_237 ( .A(_abc_3576_new_n637_), .B(DATA_IN_3_), .Y(_abc_3576_new_n652_));
AND2X2 AND2X2_238 ( .A(_abc_3576_new_n640_), .B(RLAST_REG_3_), .Y(_abc_3576_new_n653_));
AND2X2 AND2X2_239 ( .A(_abc_3576_new_n637_), .B(DATA_IN_4_), .Y(_abc_3576_new_n656_));
AND2X2 AND2X2_24 ( .A(n356), .B(STATO_REG_1_), .Y(_abc_3576_new_n203_));
AND2X2 AND2X2_240 ( .A(_abc_3576_new_n640_), .B(RLAST_REG_4_), .Y(_abc_3576_new_n657_));
AND2X2 AND2X2_241 ( .A(_abc_3576_new_n637_), .B(DATA_IN_5_), .Y(_abc_3576_new_n660_));
AND2X2 AND2X2_242 ( .A(_abc_3576_new_n640_), .B(RLAST_REG_5_), .Y(_abc_3576_new_n661_));
AND2X2 AND2X2_243 ( .A(_abc_3576_new_n637_), .B(DATA_IN_6_), .Y(_abc_3576_new_n664_));
AND2X2 AND2X2_244 ( .A(_abc_3576_new_n640_), .B(RLAST_REG_6_), .Y(_abc_3576_new_n665_));
AND2X2 AND2X2_245 ( .A(_abc_3576_new_n637_), .B(DATA_IN_7_), .Y(_abc_3576_new_n668_));
AND2X2 AND2X2_246 ( .A(_abc_3576_new_n640_), .B(RLAST_REG_7_), .Y(_abc_3576_new_n669_));
AND2X2 AND2X2_247 ( .A(_abc_3576_new_n262_), .B(RMAX_REG_7_), .Y(_abc_3576_new_n672_));
AND2X2 AND2X2_248 ( .A(_abc_3576_new_n168_), .B(RMAX_REG_1_), .Y(_abc_3576_new_n674_));
AND2X2 AND2X2_249 ( .A(_abc_3576_new_n183_), .B(DATA_IN_0_), .Y(_abc_3576_new_n676_));
AND2X2 AND2X2_25 ( .A(RMIN_REG_7_), .B(RMAX_REG_7_), .Y(_abc_3576_new_n204_));
AND2X2 AND2X2_250 ( .A(_abc_3576_new_n675_), .B(_abc_3576_new_n676_), .Y(_abc_3576_new_n677_));
AND2X2 AND2X2_251 ( .A(_abc_3576_new_n304_), .B(DATA_IN_2_), .Y(_abc_3576_new_n679_));
AND2X2 AND2X2_252 ( .A(_abc_3576_new_n680_), .B(_abc_3576_new_n681_), .Y(_abc_3576_new_n682_));
AND2X2 AND2X2_253 ( .A(_abc_3576_new_n678_), .B(_abc_3576_new_n682_), .Y(_abc_3576_new_n683_));
AND2X2 AND2X2_254 ( .A(_abc_3576_new_n684_), .B(RMAX_REG_3_), .Y(_abc_3576_new_n685_));
AND2X2 AND2X2_255 ( .A(_abc_3576_new_n302_), .B(RMAX_REG_2_), .Y(_abc_3576_new_n686_));
AND2X2 AND2X2_256 ( .A(_abc_3576_new_n689_), .B(DATA_IN_4_), .Y(_abc_3576_new_n690_));
AND2X2 AND2X2_257 ( .A(_abc_3576_new_n691_), .B(_abc_3576_new_n692_), .Y(_abc_3576_new_n693_));
AND2X2 AND2X2_258 ( .A(_abc_3576_new_n688_), .B(_abc_3576_new_n693_), .Y(_abc_3576_new_n694_));
AND2X2 AND2X2_259 ( .A(_abc_3576_new_n695_), .B(RMAX_REG_5_), .Y(_abc_3576_new_n696_));
AND2X2 AND2X2_26 ( .A(RMAX_REG_6_), .B(RMIN_REG_6_), .Y(_abc_3576_new_n206_));
AND2X2 AND2X2_260 ( .A(_abc_3576_new_n697_), .B(RMAX_REG_4_), .Y(_abc_3576_new_n698_));
AND2X2 AND2X2_261 ( .A(_abc_3576_new_n701_), .B(DATA_IN_6_), .Y(_abc_3576_new_n702_));
AND2X2 AND2X2_262 ( .A(_abc_3576_new_n703_), .B(_abc_3576_new_n704_), .Y(_abc_3576_new_n705_));
AND2X2 AND2X2_263 ( .A(_abc_3576_new_n700_), .B(_abc_3576_new_n705_), .Y(_abc_3576_new_n706_));
AND2X2 AND2X2_264 ( .A(_abc_3576_new_n233_), .B(DATA_IN_7_), .Y(_abc_3576_new_n707_));
AND2X2 AND2X2_265 ( .A(_abc_3576_new_n708_), .B(RMAX_REG_6_), .Y(_abc_3576_new_n709_));
AND2X2 AND2X2_266 ( .A(_abc_3576_new_n711_), .B(_abc_3576_new_n673_), .Y(_abc_3576_new_n712_));
AND2X2 AND2X2_267 ( .A(_abc_3576_new_n232_), .B(DATA_IN_7_), .Y(_abc_3576_new_n713_));
AND2X2 AND2X2_268 ( .A(_abc_3576_new_n714_), .B(DATA_IN_6_), .Y(_abc_3576_new_n715_));
AND2X2 AND2X2_269 ( .A(_abc_3576_new_n164_), .B(DATA_IN_1_), .Y(_abc_3576_new_n717_));
AND2X2 AND2X2_27 ( .A(RMIN_REG_1_), .B(RMAX_REG_1_), .Y(_abc_3576_new_n207_));
AND2X2 AND2X2_270 ( .A(_abc_3576_new_n181_), .B(RMIN_REG_0_), .Y(_abc_3576_new_n719_));
AND2X2 AND2X2_271 ( .A(_abc_3576_new_n718_), .B(_abc_3576_new_n719_), .Y(_abc_3576_new_n720_));
AND2X2 AND2X2_272 ( .A(_abc_3576_new_n302_), .B(RMIN_REG_2_), .Y(_abc_3576_new_n721_));
AND2X2 AND2X2_273 ( .A(_abc_3576_new_n168_), .B(RMIN_REG_1_), .Y(_abc_3576_new_n722_));
AND2X2 AND2X2_274 ( .A(_abc_3576_new_n725_), .B(DATA_IN_3_), .Y(_abc_3576_new_n726_));
AND2X2 AND2X2_275 ( .A(_abc_3576_new_n298_), .B(DATA_IN_2_), .Y(_abc_3576_new_n727_));
AND2X2 AND2X2_276 ( .A(_abc_3576_new_n724_), .B(_abc_3576_new_n729_), .Y(_abc_3576_new_n730_));
AND2X2 AND2X2_277 ( .A(_abc_3576_new_n697_), .B(RMIN_REG_4_), .Y(_abc_3576_new_n731_));
AND2X2 AND2X2_278 ( .A(_abc_3576_new_n684_), .B(RMIN_REG_3_), .Y(_abc_3576_new_n732_));
AND2X2 AND2X2_279 ( .A(_abc_3576_new_n735_), .B(_abc_3576_new_n736_), .Y(_abc_3576_new_n737_));
AND2X2 AND2X2_28 ( .A(RMIN_REG_0_), .B(RMAX_REG_0_), .Y(_abc_3576_new_n208_));
AND2X2 AND2X2_280 ( .A(_abc_3576_new_n734_), .B(_abc_3576_new_n737_), .Y(_abc_3576_new_n738_));
AND2X2 AND2X2_281 ( .A(_abc_3576_new_n695_), .B(RMIN_REG_5_), .Y(_abc_3576_new_n739_));
AND2X2 AND2X2_282 ( .A(_abc_3576_new_n708_), .B(RMIN_REG_6_), .Y(_abc_3576_new_n740_));
AND2X2 AND2X2_283 ( .A(_abc_3576_new_n742_), .B(_abc_3576_new_n716_), .Y(_abc_3576_new_n743_));
AND2X2 AND2X2_284 ( .A(_abc_3576_new_n262_), .B(RMIN_REG_7_), .Y(_abc_3576_new_n745_));
AND2X2 AND2X2_285 ( .A(_abc_3576_new_n746_), .B(STATO_REG_1_), .Y(_abc_3576_new_n747_));
AND2X2 AND2X2_286 ( .A(_abc_3576_new_n744_), .B(_abc_3576_new_n747_), .Y(_abc_3576_new_n748_));
AND2X2 AND2X2_287 ( .A(_abc_3576_new_n748_), .B(_abc_3576_new_n712_), .Y(_abc_3576_new_n749_));
AND2X2 AND2X2_288 ( .A(_abc_3576_new_n751_), .B(RMIN_REG_0_), .Y(_abc_3576_new_n752_));
AND2X2 AND2X2_289 ( .A(_abc_3576_new_n750_), .B(DATA_IN_0_), .Y(_abc_3576_new_n753_));
AND2X2 AND2X2_29 ( .A(_abc_3576_new_n210_), .B(_abc_3576_new_n211_), .Y(_abc_3576_new_n212_));
AND2X2 AND2X2_290 ( .A(_abc_3576_new_n751_), .B(RMIN_REG_1_), .Y(_abc_3576_new_n756_));
AND2X2 AND2X2_291 ( .A(_abc_3576_new_n750_), .B(DATA_IN_1_), .Y(_abc_3576_new_n757_));
AND2X2 AND2X2_292 ( .A(_abc_3576_new_n751_), .B(RMIN_REG_2_), .Y(_abc_3576_new_n760_));
AND2X2 AND2X2_293 ( .A(_abc_3576_new_n750_), .B(DATA_IN_2_), .Y(_abc_3576_new_n761_));
AND2X2 AND2X2_294 ( .A(_abc_3576_new_n751_), .B(RMIN_REG_3_), .Y(_abc_3576_new_n764_));
AND2X2 AND2X2_295 ( .A(_abc_3576_new_n750_), .B(DATA_IN_3_), .Y(_abc_3576_new_n765_));
AND2X2 AND2X2_296 ( .A(_abc_3576_new_n751_), .B(RMIN_REG_4_), .Y(_abc_3576_new_n768_));
AND2X2 AND2X2_297 ( .A(_abc_3576_new_n750_), .B(DATA_IN_4_), .Y(_abc_3576_new_n769_));
AND2X2 AND2X2_298 ( .A(_abc_3576_new_n751_), .B(RMIN_REG_5_), .Y(_abc_3576_new_n772_));
AND2X2 AND2X2_299 ( .A(_abc_3576_new_n750_), .B(DATA_IN_5_), .Y(_abc_3576_new_n773_));
AND2X2 AND2X2_3 ( .A(_abc_3576_new_n155_), .B(_abc_3576_new_n153_), .Y(_abc_3576_new_n156_));
AND2X2 AND2X2_30 ( .A(_abc_3576_new_n209_), .B(_abc_3576_new_n212_), .Y(_abc_3576_new_n213_));
AND2X2 AND2X2_300 ( .A(_abc_3576_new_n751_), .B(RMIN_REG_6_), .Y(_abc_3576_new_n776_));
AND2X2 AND2X2_301 ( .A(_abc_3576_new_n750_), .B(DATA_IN_6_), .Y(_abc_3576_new_n777_));
AND2X2 AND2X2_302 ( .A(_abc_3576_new_n751_), .B(RMIN_REG_7_), .Y(_abc_3576_new_n780_));
AND2X2 AND2X2_303 ( .A(_abc_3576_new_n750_), .B(DATA_IN_7_), .Y(_abc_3576_new_n781_));
AND2X2 AND2X2_304 ( .A(_abc_3576_new_n784_), .B(_abc_3576_new_n146_), .Y(_abc_3576_new_n785_));
AND2X2 AND2X2_305 ( .A(_abc_3576_new_n786_), .B(DATA_IN_0_), .Y(_abc_3576_new_n787_));
AND2X2 AND2X2_306 ( .A(_abc_3576_new_n785_), .B(RMAX_REG_0_), .Y(_abc_3576_new_n788_));
AND2X2 AND2X2_307 ( .A(_abc_3576_new_n786_), .B(DATA_IN_1_), .Y(_abc_3576_new_n791_));
AND2X2 AND2X2_308 ( .A(_abc_3576_new_n785_), .B(RMAX_REG_1_), .Y(_abc_3576_new_n792_));
AND2X2 AND2X2_309 ( .A(_abc_3576_new_n786_), .B(DATA_IN_2_), .Y(_abc_3576_new_n795_));
AND2X2 AND2X2_31 ( .A(RMIN_REG_2_), .B(RMAX_REG_2_), .Y(_abc_3576_new_n214_));
AND2X2 AND2X2_310 ( .A(_abc_3576_new_n785_), .B(RMAX_REG_2_), .Y(_abc_3576_new_n796_));
AND2X2 AND2X2_311 ( .A(_abc_3576_new_n786_), .B(DATA_IN_3_), .Y(_abc_3576_new_n799_));
AND2X2 AND2X2_312 ( .A(_abc_3576_new_n785_), .B(RMAX_REG_3_), .Y(_abc_3576_new_n800_));
AND2X2 AND2X2_313 ( .A(_abc_3576_new_n786_), .B(DATA_IN_4_), .Y(_abc_3576_new_n803_));
AND2X2 AND2X2_314 ( .A(_abc_3576_new_n785_), .B(RMAX_REG_4_), .Y(_abc_3576_new_n804_));
AND2X2 AND2X2_315 ( .A(_abc_3576_new_n786_), .B(DATA_IN_5_), .Y(_abc_3576_new_n807_));
AND2X2 AND2X2_316 ( .A(_abc_3576_new_n785_), .B(RMAX_REG_5_), .Y(_abc_3576_new_n808_));
AND2X2 AND2X2_317 ( .A(_abc_3576_new_n786_), .B(DATA_IN_6_), .Y(_abc_3576_new_n811_));
AND2X2 AND2X2_318 ( .A(_abc_3576_new_n785_), .B(RMAX_REG_6_), .Y(_abc_3576_new_n812_));
AND2X2 AND2X2_319 ( .A(_abc_3576_new_n786_), .B(DATA_IN_7_), .Y(_abc_3576_new_n815_));
AND2X2 AND2X2_32 ( .A(RMIN_REG_3_), .B(RMAX_REG_3_), .Y(_abc_3576_new_n215_));
AND2X2 AND2X2_320 ( .A(_abc_3576_new_n785_), .B(RMAX_REG_7_), .Y(_abc_3576_new_n816_));
AND2X2 AND2X2_321 ( .A(_abc_3576_new_n639_), .B(_abc_3576_new_n819_), .Y(n361));
AND2X2 AND2X2_33 ( .A(_abc_3576_new_n218_), .B(_abc_3576_new_n219_), .Y(_abc_3576_new_n220_));
AND2X2 AND2X2_34 ( .A(_abc_3576_new_n217_), .B(_abc_3576_new_n220_), .Y(_abc_3576_new_n221_));
AND2X2 AND2X2_35 ( .A(RMIN_REG_5_), .B(RMAX_REG_5_), .Y(_abc_3576_new_n222_));
AND2X2 AND2X2_36 ( .A(RMIN_REG_4_), .B(RMAX_REG_4_), .Y(_abc_3576_new_n223_));
AND2X2 AND2X2_37 ( .A(_abc_3576_new_n226_), .B(_abc_3576_new_n227_), .Y(_abc_3576_new_n228_));
AND2X2 AND2X2_38 ( .A(_abc_3576_new_n225_), .B(_abc_3576_new_n228_), .Y(_abc_3576_new_n229_));
AND2X2 AND2X2_39 ( .A(_abc_3576_new_n230_), .B(_abc_3576_new_n205_), .Y(_abc_3576_new_n231_));
AND2X2 AND2X2_4 ( .A(RESTART), .B(RMAX_REG_1_), .Y(_abc_3576_new_n157_));
AND2X2 AND2X2_40 ( .A(_abc_3576_new_n232_), .B(_abc_3576_new_n233_), .Y(_abc_3576_new_n234_));
AND2X2 AND2X2_41 ( .A(DATA_IN_7_), .B(REG4_REG_7_), .Y(_abc_3576_new_n237_));
AND2X2 AND2X2_42 ( .A(REG4_REG_1_), .B(DATA_IN_1_), .Y(_abc_3576_new_n239_));
AND2X2 AND2X2_43 ( .A(REG4_REG_0_), .B(DATA_IN_0_), .Y(_abc_3576_new_n240_));
AND2X2 AND2X2_44 ( .A(_abc_3576_new_n242_), .B(_abc_3576_new_n243_), .Y(_abc_3576_new_n244_));
AND2X2 AND2X2_45 ( .A(_abc_3576_new_n241_), .B(_abc_3576_new_n244_), .Y(_abc_3576_new_n245_));
AND2X2 AND2X2_46 ( .A(REG4_REG_2_), .B(DATA_IN_2_), .Y(_abc_3576_new_n246_));
AND2X2 AND2X2_47 ( .A(DATA_IN_3_), .B(REG4_REG_3_), .Y(_abc_3576_new_n247_));
AND2X2 AND2X2_48 ( .A(_abc_3576_new_n250_), .B(_abc_3576_new_n251_), .Y(_abc_3576_new_n252_));
AND2X2 AND2X2_49 ( .A(_abc_3576_new_n249_), .B(_abc_3576_new_n252_), .Y(_abc_3576_new_n253_));
AND2X2 AND2X2_5 ( .A(_abc_3576_new_n154_), .B(DATA_IN_1_), .Y(_abc_3576_new_n158_));
AND2X2 AND2X2_50 ( .A(REG4_REG_5_), .B(DATA_IN_5_), .Y(_abc_3576_new_n254_));
AND2X2 AND2X2_51 ( .A(REG4_REG_4_), .B(DATA_IN_4_), .Y(_abc_3576_new_n255_));
AND2X2 AND2X2_52 ( .A(_abc_3576_new_n258_), .B(_abc_3576_new_n259_), .Y(_abc_3576_new_n260_));
AND2X2 AND2X2_53 ( .A(_abc_3576_new_n257_), .B(_abc_3576_new_n260_), .Y(_abc_3576_new_n261_));
AND2X2 AND2X2_54 ( .A(_abc_3576_new_n262_), .B(_abc_3576_new_n263_), .Y(_abc_3576_new_n264_));
AND2X2 AND2X2_55 ( .A(DATA_IN_6_), .B(REG4_REG_6_), .Y(_abc_3576_new_n265_));
AND2X2 AND2X2_56 ( .A(_abc_3576_new_n267_), .B(_abc_3576_new_n238_), .Y(_abc_3576_new_n268_));
AND2X2 AND2X2_57 ( .A(_abc_3576_new_n272_), .B(_abc_3576_new_n236_), .Y(_abc_3576_new_n273_));
AND2X2 AND2X2_58 ( .A(_abc_3576_new_n274_), .B(_abc_3576_new_n203_), .Y(_abc_3576_new_n275_));
AND2X2 AND2X2_59 ( .A(_abc_3576_new_n275_), .B(_abc_3576_new_n202_), .Y(_abc_3576_new_n276_));
AND2X2 AND2X2_6 ( .A(_abc_3576_new_n156_), .B(_abc_3576_new_n159_), .Y(_abc_3576_new_n160_));
AND2X2 AND2X2_60 ( .A(_abc_3576_new_n268_), .B(_abc_3576_new_n278_), .Y(_abc_3576_new_n279_));
AND2X2 AND2X2_61 ( .A(_abc_3576_new_n236_), .B(_abc_3576_new_n203_), .Y(_abc_3576_new_n281_));
AND2X2 AND2X2_62 ( .A(_abc_3576_new_n280_), .B(_abc_3576_new_n281_), .Y(_abc_3576_new_n282_));
AND2X2 AND2X2_63 ( .A(_abc_3576_new_n282_), .B(_abc_3576_new_n277_), .Y(_abc_3576_new_n283_));
AND2X2 AND2X2_64 ( .A(_abc_3576_new_n203_), .B(_abc_3576_new_n154_), .Y(_abc_3576_new_n284_));
AND2X2 AND2X2_65 ( .A(AVERAGE), .B(ENABLE), .Y(_abc_3576_new_n285_));
AND2X2 AND2X2_66 ( .A(_abc_3576_new_n284_), .B(_abc_3576_new_n285_), .Y(_abc_3576_new_n286_));
AND2X2 AND2X2_67 ( .A(_abc_3576_new_n286_), .B(REG4_REG_0_), .Y(_abc_3576_new_n287_));
AND2X2 AND2X2_68 ( .A(_abc_3576_new_n284_), .B(_abc_3576_new_n269_), .Y(_abc_3576_new_n288_));
AND2X2 AND2X2_69 ( .A(_abc_3576_new_n288_), .B(RLAST_REG_0_), .Y(_abc_3576_new_n289_));
AND2X2 AND2X2_7 ( .A(_abc_3576_new_n154_), .B(_abc_3576_new_n162_), .Y(_abc_3576_new_n163_));
AND2X2 AND2X2_70 ( .A(_abc_3576_new_n290_), .B(DATA_OUT_REG_0_), .Y(_abc_3576_new_n291_));
AND2X2 AND2X2_71 ( .A(_abc_3576_new_n298_), .B(RESTART), .Y(_abc_3576_new_n299_));
AND2X2 AND2X2_72 ( .A(_abc_3576_new_n300_), .B(_abc_3576_new_n297_), .Y(_abc_3576_new_n301_));
AND2X2 AND2X2_73 ( .A(_abc_3576_new_n154_), .B(_abc_3576_new_n302_), .Y(_abc_3576_new_n303_));
AND2X2 AND2X2_74 ( .A(_abc_3576_new_n304_), .B(RESTART), .Y(_abc_3576_new_n305_));
AND2X2 AND2X2_75 ( .A(_abc_3576_new_n307_), .B(_abc_3576_new_n301_), .Y(_abc_3576_new_n309_));
AND2X2 AND2X2_76 ( .A(_abc_3576_new_n310_), .B(_abc_3576_new_n308_), .Y(_abc_3576_new_n311_));
AND2X2 AND2X2_77 ( .A(_abc_3576_new_n312_), .B(_abc_3576_new_n161_), .Y(_abc_3576_new_n313_));
AND2X2 AND2X2_78 ( .A(_abc_3576_new_n313_), .B(_abc_3576_new_n311_), .Y(_abc_3576_new_n314_));
AND2X2 AND2X2_79 ( .A(_abc_3576_new_n315_), .B(_abc_3576_new_n316_), .Y(_abc_3576_new_n317_));
AND2X2 AND2X2_8 ( .A(_abc_3576_new_n164_), .B(RESTART), .Y(_abc_3576_new_n165_));
AND2X2 AND2X2_80 ( .A(_abc_3576_new_n318_), .B(_abc_3576_new_n193_), .Y(_abc_3576_new_n319_));
AND2X2 AND2X2_81 ( .A(_abc_3576_new_n320_), .B(_abc_3576_new_n321_), .Y(_abc_3576_new_n322_));
AND2X2 AND2X2_82 ( .A(_abc_3576_new_n275_), .B(_abc_3576_new_n322_), .Y(_abc_3576_new_n323_));
AND2X2 AND2X2_83 ( .A(_abc_3576_new_n282_), .B(_abc_3576_new_n318_), .Y(_abc_3576_new_n324_));
AND2X2 AND2X2_84 ( .A(_abc_3576_new_n286_), .B(REG4_REG_1_), .Y(_abc_3576_new_n325_));
AND2X2 AND2X2_85 ( .A(_abc_3576_new_n288_), .B(RLAST_REG_1_), .Y(_abc_3576_new_n326_));
AND2X2 AND2X2_86 ( .A(_abc_3576_new_n290_), .B(DATA_OUT_REG_1_), .Y(_abc_3576_new_n327_));
AND2X2 AND2X2_87 ( .A(_abc_3576_new_n334_), .B(_abc_3576_new_n333_), .Y(_abc_3576_new_n335_));
AND2X2 AND2X2_88 ( .A(_abc_3576_new_n338_), .B(_abc_3576_new_n337_), .Y(_abc_3576_new_n339_));
AND2X2 AND2X2_89 ( .A(_abc_3576_new_n336_), .B(_abc_3576_new_n340_), .Y(_abc_3576_new_n341_));
AND2X2 AND2X2_9 ( .A(_abc_3576_new_n169_), .B(_abc_3576_new_n167_), .Y(_abc_3576_new_n170_));
AND2X2 AND2X2_90 ( .A(_abc_3576_new_n335_), .B(_abc_3576_new_n339_), .Y(_abc_3576_new_n343_));
AND2X2 AND2X2_91 ( .A(_abc_3576_new_n342_), .B(_abc_3576_new_n344_), .Y(_abc_3576_new_n345_));
AND2X2 AND2X2_92 ( .A(_abc_3576_new_n347_), .B(_abc_3576_new_n310_), .Y(_abc_3576_new_n348_));
AND2X2 AND2X2_93 ( .A(_abc_3576_new_n348_), .B(_abc_3576_new_n345_), .Y(_abc_3576_new_n349_));
AND2X2 AND2X2_94 ( .A(_abc_3576_new_n282_), .B(_abc_3576_new_n352_), .Y(_abc_3576_new_n353_));
AND2X2 AND2X2_95 ( .A(_abc_3576_new_n352_), .B(_abc_3576_new_n320_), .Y(_abc_3576_new_n354_));
AND2X2 AND2X2_96 ( .A(_abc_3576_new_n355_), .B(_abc_3576_new_n319_), .Y(_abc_3576_new_n356_));
AND2X2 AND2X2_97 ( .A(_abc_3576_new_n357_), .B(_abc_3576_new_n275_), .Y(_abc_3576_new_n358_));
AND2X2 AND2X2_98 ( .A(_abc_3576_new_n286_), .B(REG4_REG_2_), .Y(_abc_3576_new_n359_));
AND2X2 AND2X2_99 ( .A(_abc_3576_new_n288_), .B(RLAST_REG_2_), .Y(_abc_3576_new_n360_));
DFFPOSX1 DFFPOSX1_1 ( .CLK(clock), .D(n324), .Q(DATA_OUT_REG_7_));
DFFPOSX1 DFFPOSX1_10 ( .CLK(clock), .D(n49), .Q(RMAX_REG_6_));
DFFPOSX1 DFFPOSX1_11 ( .CLK(clock), .D(n54), .Q(RMAX_REG_5_));
DFFPOSX1 DFFPOSX1_12 ( .CLK(clock), .D(n59), .Q(RMAX_REG_4_));
DFFPOSX1 DFFPOSX1_13 ( .CLK(clock), .D(n64), .Q(RMAX_REG_3_));
DFFPOSX1 DFFPOSX1_14 ( .CLK(clock), .D(n69), .Q(RMAX_REG_2_));
DFFPOSX1 DFFPOSX1_15 ( .CLK(clock), .D(n74), .Q(RMAX_REG_1_));
DFFPOSX1 DFFPOSX1_16 ( .CLK(clock), .D(n79), .Q(RMAX_REG_0_));
DFFPOSX1 DFFPOSX1_17 ( .CLK(clock), .D(n84), .Q(RMIN_REG_7_));
DFFPOSX1 DFFPOSX1_18 ( .CLK(clock), .D(n89), .Q(RMIN_REG_6_));
DFFPOSX1 DFFPOSX1_19 ( .CLK(clock), .D(n94), .Q(RMIN_REG_5_));
DFFPOSX1 DFFPOSX1_2 ( .CLK(clock), .D(n332), .Q(DATA_OUT_REG_5_));
DFFPOSX1 DFFPOSX1_20 ( .CLK(clock), .D(n99), .Q(RMIN_REG_4_));
DFFPOSX1 DFFPOSX1_21 ( .CLK(clock), .D(n104), .Q(RMIN_REG_3_));
DFFPOSX1 DFFPOSX1_22 ( .CLK(clock), .D(n109), .Q(RMIN_REG_2_));
DFFPOSX1 DFFPOSX1_23 ( .CLK(clock), .D(n114), .Q(RMIN_REG_1_));
DFFPOSX1 DFFPOSX1_24 ( .CLK(clock), .D(n119), .Q(RMIN_REG_0_));
DFFPOSX1 DFFPOSX1_25 ( .CLK(clock), .D(n124), .Q(RLAST_REG_7_));
DFFPOSX1 DFFPOSX1_26 ( .CLK(clock), .D(n129), .Q(RLAST_REG_6_));
DFFPOSX1 DFFPOSX1_27 ( .CLK(clock), .D(n134), .Q(RLAST_REG_5_));
DFFPOSX1 DFFPOSX1_28 ( .CLK(clock), .D(n139), .Q(RLAST_REG_4_));
DFFPOSX1 DFFPOSX1_29 ( .CLK(clock), .D(n144), .Q(RLAST_REG_3_));
DFFPOSX1 DFFPOSX1_3 ( .CLK(clock), .D(n344), .Q(DATA_OUT_REG_2_));
DFFPOSX1 DFFPOSX1_30 ( .CLK(clock), .D(n149), .Q(RLAST_REG_2_));
DFFPOSX1 DFFPOSX1_31 ( .CLK(clock), .D(n154), .Q(RLAST_REG_1_));
DFFPOSX1 DFFPOSX1_32 ( .CLK(clock), .D(n159), .Q(RLAST_REG_0_));
DFFPOSX1 DFFPOSX1_33 ( .CLK(clock), .D(n164), .Q(REG1_REG_7_));
DFFPOSX1 DFFPOSX1_34 ( .CLK(clock), .D(n169), .Q(REG1_REG_6_));
DFFPOSX1 DFFPOSX1_35 ( .CLK(clock), .D(n174), .Q(REG1_REG_5_));
DFFPOSX1 DFFPOSX1_36 ( .CLK(clock), .D(n179), .Q(REG1_REG_4_));
DFFPOSX1 DFFPOSX1_37 ( .CLK(clock), .D(n184), .Q(REG1_REG_3_));
DFFPOSX1 DFFPOSX1_38 ( .CLK(clock), .D(n189), .Q(REG1_REG_2_));
DFFPOSX1 DFFPOSX1_39 ( .CLK(clock), .D(n194), .Q(REG1_REG_1_));
DFFPOSX1 DFFPOSX1_4 ( .CLK(clock), .D(n336), .Q(DATA_OUT_REG_4_));
DFFPOSX1 DFFPOSX1_40 ( .CLK(clock), .D(n199), .Q(REG1_REG_0_));
DFFPOSX1 DFFPOSX1_41 ( .CLK(clock), .D(n204), .Q(REG2_REG_7_));
DFFPOSX1 DFFPOSX1_42 ( .CLK(clock), .D(n209), .Q(REG2_REG_6_));
DFFPOSX1 DFFPOSX1_43 ( .CLK(clock), .D(n214), .Q(REG2_REG_5_));
DFFPOSX1 DFFPOSX1_44 ( .CLK(clock), .D(n219), .Q(REG2_REG_4_));
DFFPOSX1 DFFPOSX1_45 ( .CLK(clock), .D(n224), .Q(REG2_REG_3_));
DFFPOSX1 DFFPOSX1_46 ( .CLK(clock), .D(n229), .Q(REG2_REG_2_));
DFFPOSX1 DFFPOSX1_47 ( .CLK(clock), .D(n234), .Q(REG2_REG_1_));
DFFPOSX1 DFFPOSX1_48 ( .CLK(clock), .D(n239), .Q(REG2_REG_0_));
DFFPOSX1 DFFPOSX1_49 ( .CLK(clock), .D(n244), .Q(REG3_REG_7_));
DFFPOSX1 DFFPOSX1_5 ( .CLK(clock), .D(n340), .Q(DATA_OUT_REG_3_));
DFFPOSX1 DFFPOSX1_50 ( .CLK(clock), .D(n249), .Q(REG3_REG_6_));
DFFPOSX1 DFFPOSX1_51 ( .CLK(clock), .D(n254), .Q(REG3_REG_5_));
DFFPOSX1 DFFPOSX1_52 ( .CLK(clock), .D(n259), .Q(REG3_REG_4_));
DFFPOSX1 DFFPOSX1_53 ( .CLK(clock), .D(n264), .Q(REG3_REG_3_));
DFFPOSX1 DFFPOSX1_54 ( .CLK(clock), .D(n269), .Q(REG3_REG_2_));
DFFPOSX1 DFFPOSX1_55 ( .CLK(clock), .D(n274), .Q(REG3_REG_1_));
DFFPOSX1 DFFPOSX1_56 ( .CLK(clock), .D(n279), .Q(REG3_REG_0_));
DFFPOSX1 DFFPOSX1_57 ( .CLK(clock), .D(n284), .Q(REG4_REG_7_));
DFFPOSX1 DFFPOSX1_58 ( .CLK(clock), .D(n289), .Q(REG4_REG_6_));
DFFPOSX1 DFFPOSX1_59 ( .CLK(clock), .D(n294), .Q(REG4_REG_5_));
DFFPOSX1 DFFPOSX1_6 ( .CLK(clock), .D(n328), .Q(DATA_OUT_REG_6_));
DFFPOSX1 DFFPOSX1_60 ( .CLK(clock), .D(n299), .Q(REG4_REG_4_));
DFFPOSX1 DFFPOSX1_61 ( .CLK(clock), .D(n304), .Q(REG4_REG_3_));
DFFPOSX1 DFFPOSX1_62 ( .CLK(clock), .D(n309), .Q(REG4_REG_2_));
DFFPOSX1 DFFPOSX1_63 ( .CLK(clock), .D(n314), .Q(REG4_REG_1_));
DFFPOSX1 DFFPOSX1_64 ( .CLK(clock), .D(n319), .Q(REG4_REG_0_));
DFFPOSX1 DFFPOSX1_65 ( .CLK(clock), .D(n356), .Q(STATO_REG_1_));
DFFPOSX1 DFFPOSX1_66 ( .CLK(clock), .D(n361), .Q(STATO_REG_0_));
DFFPOSX1 DFFPOSX1_7 ( .CLK(clock), .D(n348), .Q(DATA_OUT_REG_1_));
DFFPOSX1 DFFPOSX1_8 ( .CLK(clock), .D(n352), .Q(DATA_OUT_REG_0_));
DFFPOSX1 DFFPOSX1_9 ( .CLK(clock), .D(n44), .Q(RMAX_REG_7_));
INVX1 INVX1_1 ( .A(STATO_REG_0_), .Y(_abc_3576_new_n146_));
INVX1 INVX1_10 ( .A(_abc_3576_new_n171_), .Y(_abc_3576_new_n172_));
INVX1 INVX1_11 ( .A(DATA_IN_0_), .Y(_abc_3576_new_n181_));
INVX1 INVX1_12 ( .A(RMAX_REG_0_), .Y(_abc_3576_new_n183_));
INVX1 INVX1_13 ( .A(REG4_REG_0_), .Y(_abc_3576_new_n186_));
INVX1 INVX1_14 ( .A(_abc_3576_new_n178_), .Y(_abc_3576_new_n188_));
INVX1 INVX1_15 ( .A(_abc_3576_new_n191_), .Y(_abc_3576_new_n192_));
INVX1 INVX1_16 ( .A(_abc_3576_new_n193_), .Y(_abc_3576_new_n194_));
INVX1 INVX1_17 ( .A(_abc_3576_new_n173_), .Y(_abc_3576_new_n195_));
INVX1 INVX1_18 ( .A(_abc_3576_new_n200_), .Y(_abc_3576_new_n201_));
INVX1 INVX1_19 ( .A(_abc_3576_new_n204_), .Y(_abc_3576_new_n205_));
INVX1 INVX1_2 ( .A(nRESET_G), .Y(_abc_3576_new_n148_));
INVX1 INVX1_20 ( .A(RMIN_REG_7_), .Y(_abc_3576_new_n232_));
INVX1 INVX1_21 ( .A(RMAX_REG_7_), .Y(_abc_3576_new_n233_));
INVX1 INVX1_22 ( .A(_abc_3576_new_n237_), .Y(_abc_3576_new_n238_));
INVX1 INVX1_23 ( .A(DATA_IN_7_), .Y(_abc_3576_new_n262_));
INVX1 INVX1_24 ( .A(REG4_REG_7_), .Y(_abc_3576_new_n263_));
INVX1 INVX1_25 ( .A(ENABLE), .Y(_abc_3576_new_n269_));
INVX1 INVX1_26 ( .A(_abc_3576_new_n273_), .Y(_abc_3576_new_n274_));
INVX1 INVX1_27 ( .A(_abc_3576_new_n199_), .Y(_abc_3576_new_n277_));
INVX1 INVX1_28 ( .A(_abc_3576_new_n270_), .Y(_abc_3576_new_n278_));
INVX1 INVX1_29 ( .A(n356), .Y(_abc_3576_new_n290_));
INVX1 INVX1_3 ( .A(STATO_REG_1_), .Y(_abc_3576_new_n149_));
INVX1 INVX1_30 ( .A(RMIN_REG_2_), .Y(_abc_3576_new_n298_));
INVX1 INVX1_31 ( .A(_abc_3576_new_n299_), .Y(_abc_3576_new_n300_));
INVX1 INVX1_32 ( .A(DATA_IN_2_), .Y(_abc_3576_new_n302_));
INVX1 INVX1_33 ( .A(RMAX_REG_2_), .Y(_abc_3576_new_n304_));
INVX1 INVX1_34 ( .A(_abc_3576_new_n306_), .Y(_abc_3576_new_n307_));
INVX1 INVX1_35 ( .A(_abc_3576_new_n309_), .Y(_abc_3576_new_n310_));
INVX1 INVX1_36 ( .A(_abc_3576_new_n314_), .Y(_abc_3576_new_n315_));
INVX1 INVX1_37 ( .A(_abc_3576_new_n317_), .Y(_abc_3576_new_n318_));
INVX1 INVX1_38 ( .A(_abc_3576_new_n319_), .Y(_abc_3576_new_n320_));
INVX1 INVX1_39 ( .A(_abc_3576_new_n335_), .Y(_abc_3576_new_n336_));
INVX1 INVX1_4 ( .A(RESTART), .Y(_abc_3576_new_n154_));
INVX1 INVX1_40 ( .A(_abc_3576_new_n339_), .Y(_abc_3576_new_n340_));
INVX1 INVX1_41 ( .A(_abc_3576_new_n341_), .Y(_abc_3576_new_n342_));
INVX1 INVX1_42 ( .A(_abc_3576_new_n343_), .Y(_abc_3576_new_n344_));
INVX1 INVX1_43 ( .A(_abc_3576_new_n308_), .Y(_abc_3576_new_n346_));
INVX1 INVX1_44 ( .A(_abc_3576_new_n350_), .Y(_abc_3576_new_n351_));
INVX1 INVX1_45 ( .A(_abc_3576_new_n352_), .Y(_abc_3576_new_n355_));
INVX1 INVX1_46 ( .A(_abc_3576_new_n379_), .Y(_abc_3576_new_n380_));
INVX1 INVX1_47 ( .A(_abc_3576_new_n382_), .Y(_abc_3576_new_n383_));
INVX1 INVX1_48 ( .A(_abc_3576_new_n392_), .Y(_abc_3576_new_n393_));
INVX1 INVX1_49 ( .A(_abc_3576_new_n368_), .Y(_abc_3576_new_n396_));
INVX1 INVX1_5 ( .A(_abc_3576_new_n160_), .Y(_abc_3576_new_n161_));
INVX1 INVX1_50 ( .A(_abc_3576_new_n399_), .Y(_abc_3576_new_n400_));
INVX1 INVX1_51 ( .A(_abc_3576_new_n418_), .Y(_abc_3576_new_n419_));
INVX1 INVX1_52 ( .A(_abc_3576_new_n421_), .Y(_abc_3576_new_n422_));
INVX1 INVX1_53 ( .A(_abc_3576_new_n381_), .Y(_abc_3576_new_n423_));
INVX1 INVX1_54 ( .A(_abc_3576_new_n431_), .Y(_abc_3576_new_n432_));
INVX1 INVX1_55 ( .A(_abc_3576_new_n434_), .Y(_abc_3576_new_n435_));
INVX1 INVX1_56 ( .A(_abc_3576_new_n437_), .Y(_abc_3576_new_n438_));
INVX1 INVX1_57 ( .A(_abc_3576_new_n430_), .Y(_abc_3576_new_n441_));
INVX1 INVX1_58 ( .A(_abc_3576_new_n420_), .Y(_abc_3576_new_n451_));
INVX1 INVX1_59 ( .A(_abc_3576_new_n456_), .Y(_abc_3576_new_n457_));
INVX1 INVX1_6 ( .A(REG4_REG_1_), .Y(_abc_3576_new_n162_));
INVX1 INVX1_60 ( .A(_abc_3576_new_n462_), .Y(_abc_3576_new_n463_));
INVX1 INVX1_61 ( .A(_abc_3576_new_n464_), .Y(_abc_3576_new_n465_));
INVX1 INVX1_62 ( .A(_abc_3576_new_n476_), .Y(_abc_3576_new_n477_));
INVX1 INVX1_63 ( .A(_abc_3576_new_n635_), .Y(_abc_3576_new_n636_));
INVX1 INVX1_64 ( .A(_abc_3576_new_n672_), .Y(_abc_3576_new_n673_));
INVX1 INVX1_65 ( .A(_abc_3576_new_n674_), .Y(_abc_3576_new_n675_));
INVX1 INVX1_66 ( .A(_abc_3576_new_n677_), .Y(_abc_3576_new_n678_));
INVX1 INVX1_67 ( .A(_abc_3576_new_n679_), .Y(_abc_3576_new_n680_));
INVX1 INVX1_68 ( .A(DATA_IN_3_), .Y(_abc_3576_new_n684_));
INVX1 INVX1_69 ( .A(RMAX_REG_4_), .Y(_abc_3576_new_n689_));
INVX1 INVX1_7 ( .A(RMIN_REG_1_), .Y(_abc_3576_new_n164_));
INVX1 INVX1_70 ( .A(_abc_3576_new_n690_), .Y(_abc_3576_new_n691_));
INVX1 INVX1_71 ( .A(DATA_IN_5_), .Y(_abc_3576_new_n695_));
INVX1 INVX1_72 ( .A(DATA_IN_4_), .Y(_abc_3576_new_n697_));
INVX1 INVX1_73 ( .A(RMAX_REG_6_), .Y(_abc_3576_new_n701_));
INVX1 INVX1_74 ( .A(_abc_3576_new_n702_), .Y(_abc_3576_new_n703_));
INVX1 INVX1_75 ( .A(DATA_IN_6_), .Y(_abc_3576_new_n708_));
INVX1 INVX1_76 ( .A(RMIN_REG_6_), .Y(_abc_3576_new_n714_));
INVX1 INVX1_77 ( .A(_abc_3576_new_n715_), .Y(_abc_3576_new_n716_));
INVX1 INVX1_78 ( .A(_abc_3576_new_n717_), .Y(_abc_3576_new_n718_));
INVX1 INVX1_79 ( .A(RMIN_REG_3_), .Y(_abc_3576_new_n725_));
INVX1 INVX1_8 ( .A(_abc_3576_new_n157_), .Y(_abc_3576_new_n167_));
INVX1 INVX1_80 ( .A(_abc_3576_new_n728_), .Y(_abc_3576_new_n729_));
INVX1 INVX1_81 ( .A(_abc_3576_new_n745_), .Y(_abc_3576_new_n746_));
INVX1 INVX1_82 ( .A(_abc_3576_new_n750_), .Y(_abc_3576_new_n751_));
INVX1 INVX1_83 ( .A(_abc_3576_new_n785_), .Y(_abc_3576_new_n786_));
INVX1 INVX1_84 ( .A(RESET_G), .Y(_abc_3576_new_n819_));
INVX1 INVX1_9 ( .A(DATA_IN_1_), .Y(_abc_3576_new_n168_));
OR2X2 OR2X2_1 ( .A(_abc_3576_new_n150_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n151_));
OR2X2 OR2X2_10 ( .A(_abc_3576_new_n177_), .B(_abc_3576_new_n178_), .Y(_abc_3576_new_n179_));
OR2X2 OR2X2_100 ( .A(_abc_3576_new_n372_), .B(_abc_3576_new_n423_), .Y(_abc_3576_new_n424_));
OR2X2 OR2X2_101 ( .A(_abc_3576_new_n427_), .B(_abc_3576_new_n379_), .Y(_abc_3576_new_n428_));
OR2X2 OR2X2_102 ( .A(_abc_3576_new_n426_), .B(_abc_3576_new_n429_), .Y(_abc_3576_new_n430_));
OR2X2 OR2X2_103 ( .A(_abc_3576_new_n430_), .B(_abc_3576_new_n395_), .Y(_abc_3576_new_n433_));
OR2X2 OR2X2_104 ( .A(_abc_3576_new_n435_), .B(_abc_3576_new_n399_), .Y(_abc_3576_new_n436_));
OR2X2 OR2X2_105 ( .A(_abc_3576_new_n445_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n446_));
OR2X2 OR2X2_106 ( .A(_abc_3576_new_n444_), .B(_abc_3576_new_n446_), .Y(_abc_3576_new_n447_));
OR2X2 OR2X2_107 ( .A(_abc_3576_new_n447_), .B(_abc_3576_new_n443_), .Y(_abc_3576_new_n448_));
OR2X2 OR2X2_108 ( .A(_abc_3576_new_n442_), .B(_abc_3576_new_n448_), .Y(_abc_3576_new_n449_));
OR2X2 OR2X2_109 ( .A(_abc_3576_new_n440_), .B(_abc_3576_new_n449_), .Y(n336));
OR2X2 OR2X2_11 ( .A(_abc_3576_new_n182_), .B(_abc_3576_new_n184_), .Y(_abc_3576_new_n185_));
OR2X2 OR2X2_110 ( .A(_abc_3576_new_n425_), .B(_abc_3576_new_n451_), .Y(_abc_3576_new_n452_));
OR2X2 OR2X2_111 ( .A(RESTART), .B(REG4_REG_6_), .Y(_abc_3576_new_n454_));
OR2X2 OR2X2_112 ( .A(_abc_3576_new_n154_), .B(RMIN_REG_6_), .Y(_abc_3576_new_n455_));
OR2X2 OR2X2_113 ( .A(RESTART), .B(DATA_IN_6_), .Y(_abc_3576_new_n458_));
OR2X2 OR2X2_114 ( .A(_abc_3576_new_n154_), .B(RMAX_REG_6_), .Y(_abc_3576_new_n459_));
OR2X2 OR2X2_115 ( .A(_abc_3576_new_n457_), .B(_abc_3576_new_n460_), .Y(_abc_3576_new_n462_));
OR2X2 OR2X2_116 ( .A(_abc_3576_new_n463_), .B(_abc_3576_new_n461_), .Y(_abc_3576_new_n464_));
OR2X2 OR2X2_117 ( .A(_abc_3576_new_n467_), .B(_abc_3576_new_n418_), .Y(_abc_3576_new_n468_));
OR2X2 OR2X2_118 ( .A(_abc_3576_new_n466_), .B(_abc_3576_new_n469_), .Y(_abc_3576_new_n470_));
OR2X2 OR2X2_119 ( .A(_abc_3576_new_n470_), .B(_abc_3576_new_n432_), .Y(_abc_3576_new_n471_));
OR2X2 OR2X2_12 ( .A(_abc_3576_new_n186_), .B(RESTART), .Y(_abc_3576_new_n187_));
OR2X2 OR2X2_120 ( .A(_abc_3576_new_n468_), .B(_abc_3576_new_n464_), .Y(_abc_3576_new_n472_));
OR2X2 OR2X2_121 ( .A(_abc_3576_new_n453_), .B(_abc_3576_new_n465_), .Y(_abc_3576_new_n473_));
OR2X2 OR2X2_122 ( .A(_abc_3576_new_n474_), .B(_abc_3576_new_n431_), .Y(_abc_3576_new_n475_));
OR2X2 OR2X2_123 ( .A(_abc_3576_new_n477_), .B(_abc_3576_new_n438_), .Y(_abc_3576_new_n478_));
OR2X2 OR2X2_124 ( .A(_abc_3576_new_n476_), .B(_abc_3576_new_n437_), .Y(_abc_3576_new_n479_));
OR2X2 OR2X2_125 ( .A(_abc_3576_new_n485_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n486_));
OR2X2 OR2X2_126 ( .A(_abc_3576_new_n484_), .B(_abc_3576_new_n486_), .Y(_abc_3576_new_n487_));
OR2X2 OR2X2_127 ( .A(_abc_3576_new_n487_), .B(_abc_3576_new_n483_), .Y(_abc_3576_new_n488_));
OR2X2 OR2X2_128 ( .A(_abc_3576_new_n482_), .B(_abc_3576_new_n488_), .Y(_abc_3576_new_n489_));
OR2X2 OR2X2_129 ( .A(_abc_3576_new_n481_), .B(_abc_3576_new_n489_), .Y(n332));
OR2X2 OR2X2_13 ( .A(_abc_3576_new_n190_), .B(_abc_3576_new_n180_), .Y(_abc_3576_new_n191_));
OR2X2 OR2X2_130 ( .A(_abc_3576_new_n493_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n494_));
OR2X2 OR2X2_131 ( .A(_abc_3576_new_n492_), .B(_abc_3576_new_n494_), .Y(_abc_3576_new_n495_));
OR2X2 OR2X2_132 ( .A(_abc_3576_new_n495_), .B(_abc_3576_new_n491_), .Y(_abc_3576_new_n496_));
OR2X2 OR2X2_133 ( .A(_abc_3576_new_n499_), .B(_abc_3576_new_n496_), .Y(n328));
OR2X2 OR2X2_134 ( .A(_abc_3576_new_n503_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n504_));
OR2X2 OR2X2_135 ( .A(_abc_3576_new_n502_), .B(_abc_3576_new_n504_), .Y(_abc_3576_new_n505_));
OR2X2 OR2X2_136 ( .A(_abc_3576_new_n505_), .B(_abc_3576_new_n501_), .Y(n324));
OR2X2 OR2X2_137 ( .A(_abc_3576_new_n508_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n509_));
OR2X2 OR2X2_138 ( .A(_abc_3576_new_n507_), .B(_abc_3576_new_n509_), .Y(n319));
OR2X2 OR2X2_139 ( .A(_abc_3576_new_n512_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n513_));
OR2X2 OR2X2_14 ( .A(_abc_3576_new_n195_), .B(_abc_3576_new_n180_), .Y(_abc_3576_new_n196_));
OR2X2 OR2X2_140 ( .A(_abc_3576_new_n511_), .B(_abc_3576_new_n513_), .Y(n314));
OR2X2 OR2X2_141 ( .A(_abc_3576_new_n516_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n517_));
OR2X2 OR2X2_142 ( .A(_abc_3576_new_n515_), .B(_abc_3576_new_n517_), .Y(n309));
OR2X2 OR2X2_143 ( .A(_abc_3576_new_n520_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n521_));
OR2X2 OR2X2_144 ( .A(_abc_3576_new_n519_), .B(_abc_3576_new_n521_), .Y(n304));
OR2X2 OR2X2_145 ( .A(_abc_3576_new_n524_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n525_));
OR2X2 OR2X2_146 ( .A(_abc_3576_new_n523_), .B(_abc_3576_new_n525_), .Y(n299));
OR2X2 OR2X2_147 ( .A(_abc_3576_new_n528_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n529_));
OR2X2 OR2X2_148 ( .A(_abc_3576_new_n527_), .B(_abc_3576_new_n529_), .Y(n294));
OR2X2 OR2X2_149 ( .A(_abc_3576_new_n532_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n533_));
OR2X2 OR2X2_15 ( .A(_abc_3576_new_n185_), .B(_abc_3576_new_n189_), .Y(_abc_3576_new_n197_));
OR2X2 OR2X2_150 ( .A(_abc_3576_new_n531_), .B(_abc_3576_new_n533_), .Y(n289));
OR2X2 OR2X2_151 ( .A(_abc_3576_new_n536_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n537_));
OR2X2 OR2X2_152 ( .A(_abc_3576_new_n535_), .B(_abc_3576_new_n537_), .Y(n284));
OR2X2 OR2X2_153 ( .A(_abc_3576_new_n540_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n541_));
OR2X2 OR2X2_154 ( .A(_abc_3576_new_n539_), .B(_abc_3576_new_n541_), .Y(n279));
OR2X2 OR2X2_155 ( .A(_abc_3576_new_n544_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n545_));
OR2X2 OR2X2_156 ( .A(_abc_3576_new_n543_), .B(_abc_3576_new_n545_), .Y(n274));
OR2X2 OR2X2_157 ( .A(_abc_3576_new_n548_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n549_));
OR2X2 OR2X2_158 ( .A(_abc_3576_new_n547_), .B(_abc_3576_new_n549_), .Y(n269));
OR2X2 OR2X2_159 ( .A(_abc_3576_new_n552_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n553_));
OR2X2 OR2X2_16 ( .A(_abc_3576_new_n173_), .B(_abc_3576_new_n197_), .Y(_abc_3576_new_n198_));
OR2X2 OR2X2_160 ( .A(_abc_3576_new_n551_), .B(_abc_3576_new_n553_), .Y(n264));
OR2X2 OR2X2_161 ( .A(_abc_3576_new_n556_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n557_));
OR2X2 OR2X2_162 ( .A(_abc_3576_new_n555_), .B(_abc_3576_new_n557_), .Y(n259));
OR2X2 OR2X2_163 ( .A(_abc_3576_new_n560_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n561_));
OR2X2 OR2X2_164 ( .A(_abc_3576_new_n559_), .B(_abc_3576_new_n561_), .Y(n254));
OR2X2 OR2X2_165 ( .A(_abc_3576_new_n564_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n565_));
OR2X2 OR2X2_166 ( .A(_abc_3576_new_n563_), .B(_abc_3576_new_n565_), .Y(n249));
OR2X2 OR2X2_167 ( .A(_abc_3576_new_n568_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n569_));
OR2X2 OR2X2_168 ( .A(_abc_3576_new_n567_), .B(_abc_3576_new_n569_), .Y(n244));
OR2X2 OR2X2_169 ( .A(_abc_3576_new_n572_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n573_));
OR2X2 OR2X2_17 ( .A(_abc_3576_new_n207_), .B(_abc_3576_new_n208_), .Y(_abc_3576_new_n209_));
OR2X2 OR2X2_170 ( .A(_abc_3576_new_n571_), .B(_abc_3576_new_n573_), .Y(n239));
OR2X2 OR2X2_171 ( .A(_abc_3576_new_n576_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n577_));
OR2X2 OR2X2_172 ( .A(_abc_3576_new_n575_), .B(_abc_3576_new_n577_), .Y(n234));
OR2X2 OR2X2_173 ( .A(_abc_3576_new_n580_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n581_));
OR2X2 OR2X2_174 ( .A(_abc_3576_new_n579_), .B(_abc_3576_new_n581_), .Y(n229));
OR2X2 OR2X2_175 ( .A(_abc_3576_new_n584_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n585_));
OR2X2 OR2X2_176 ( .A(_abc_3576_new_n583_), .B(_abc_3576_new_n585_), .Y(n224));
OR2X2 OR2X2_177 ( .A(_abc_3576_new_n588_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n589_));
OR2X2 OR2X2_178 ( .A(_abc_3576_new_n587_), .B(_abc_3576_new_n589_), .Y(n219));
OR2X2 OR2X2_179 ( .A(_abc_3576_new_n592_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n593_));
OR2X2 OR2X2_18 ( .A(RMIN_REG_2_), .B(RMAX_REG_2_), .Y(_abc_3576_new_n210_));
OR2X2 OR2X2_180 ( .A(_abc_3576_new_n591_), .B(_abc_3576_new_n593_), .Y(n214));
OR2X2 OR2X2_181 ( .A(_abc_3576_new_n596_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n597_));
OR2X2 OR2X2_182 ( .A(_abc_3576_new_n595_), .B(_abc_3576_new_n597_), .Y(n209));
OR2X2 OR2X2_183 ( .A(_abc_3576_new_n600_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n601_));
OR2X2 OR2X2_184 ( .A(_abc_3576_new_n599_), .B(_abc_3576_new_n601_), .Y(n204));
OR2X2 OR2X2_185 ( .A(_abc_3576_new_n604_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n605_));
OR2X2 OR2X2_186 ( .A(_abc_3576_new_n603_), .B(_abc_3576_new_n605_), .Y(n199));
OR2X2 OR2X2_187 ( .A(_abc_3576_new_n608_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n609_));
OR2X2 OR2X2_188 ( .A(_abc_3576_new_n607_), .B(_abc_3576_new_n609_), .Y(n194));
OR2X2 OR2X2_189 ( .A(_abc_3576_new_n612_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n613_));
OR2X2 OR2X2_19 ( .A(RMIN_REG_1_), .B(RMAX_REG_1_), .Y(_abc_3576_new_n211_));
OR2X2 OR2X2_190 ( .A(_abc_3576_new_n611_), .B(_abc_3576_new_n613_), .Y(n189));
OR2X2 OR2X2_191 ( .A(_abc_3576_new_n616_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n617_));
OR2X2 OR2X2_192 ( .A(_abc_3576_new_n615_), .B(_abc_3576_new_n617_), .Y(n184));
OR2X2 OR2X2_193 ( .A(_abc_3576_new_n620_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n621_));
OR2X2 OR2X2_194 ( .A(_abc_3576_new_n619_), .B(_abc_3576_new_n621_), .Y(n179));
OR2X2 OR2X2_195 ( .A(_abc_3576_new_n624_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n625_));
OR2X2 OR2X2_196 ( .A(_abc_3576_new_n623_), .B(_abc_3576_new_n625_), .Y(n174));
OR2X2 OR2X2_197 ( .A(_abc_3576_new_n628_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n629_));
OR2X2 OR2X2_198 ( .A(_abc_3576_new_n627_), .B(_abc_3576_new_n629_), .Y(n169));
OR2X2 OR2X2_199 ( .A(_abc_3576_new_n632_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n633_));
OR2X2 OR2X2_2 ( .A(_abc_3576_new_n151_), .B(_abc_3576_new_n147_), .Y(n356));
OR2X2 OR2X2_20 ( .A(_abc_3576_new_n214_), .B(_abc_3576_new_n215_), .Y(_abc_3576_new_n216_));
OR2X2 OR2X2_200 ( .A(_abc_3576_new_n631_), .B(_abc_3576_new_n633_), .Y(n164));
OR2X2 OR2X2_201 ( .A(_abc_3576_new_n635_), .B(_abc_3576_new_n639_), .Y(_abc_3576_new_n640_));
OR2X2 OR2X2_202 ( .A(_abc_3576_new_n641_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n642_));
OR2X2 OR2X2_203 ( .A(_abc_3576_new_n642_), .B(_abc_3576_new_n638_), .Y(n159));
OR2X2 OR2X2_204 ( .A(_abc_3576_new_n645_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n646_));
OR2X2 OR2X2_205 ( .A(_abc_3576_new_n646_), .B(_abc_3576_new_n644_), .Y(n154));
OR2X2 OR2X2_206 ( .A(_abc_3576_new_n649_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n650_));
OR2X2 OR2X2_207 ( .A(_abc_3576_new_n650_), .B(_abc_3576_new_n648_), .Y(n149));
OR2X2 OR2X2_208 ( .A(_abc_3576_new_n653_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n654_));
OR2X2 OR2X2_209 ( .A(_abc_3576_new_n654_), .B(_abc_3576_new_n652_), .Y(n144));
OR2X2 OR2X2_21 ( .A(_abc_3576_new_n213_), .B(_abc_3576_new_n216_), .Y(_abc_3576_new_n217_));
OR2X2 OR2X2_210 ( .A(_abc_3576_new_n657_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n658_));
OR2X2 OR2X2_211 ( .A(_abc_3576_new_n658_), .B(_abc_3576_new_n656_), .Y(n139));
OR2X2 OR2X2_212 ( .A(_abc_3576_new_n661_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n662_));
OR2X2 OR2X2_213 ( .A(_abc_3576_new_n662_), .B(_abc_3576_new_n660_), .Y(n134));
OR2X2 OR2X2_214 ( .A(_abc_3576_new_n665_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n666_));
OR2X2 OR2X2_215 ( .A(_abc_3576_new_n666_), .B(_abc_3576_new_n664_), .Y(n129));
OR2X2 OR2X2_216 ( .A(_abc_3576_new_n669_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n670_));
OR2X2 OR2X2_217 ( .A(_abc_3576_new_n670_), .B(_abc_3576_new_n668_), .Y(n124));
OR2X2 OR2X2_218 ( .A(_abc_3576_new_n168_), .B(RMAX_REG_1_), .Y(_abc_3576_new_n681_));
OR2X2 OR2X2_219 ( .A(_abc_3576_new_n685_), .B(_abc_3576_new_n686_), .Y(_abc_3576_new_n687_));
OR2X2 OR2X2_22 ( .A(RMIN_REG_4_), .B(RMAX_REG_4_), .Y(_abc_3576_new_n218_));
OR2X2 OR2X2_220 ( .A(_abc_3576_new_n683_), .B(_abc_3576_new_n687_), .Y(_abc_3576_new_n688_));
OR2X2 OR2X2_221 ( .A(_abc_3576_new_n684_), .B(RMAX_REG_3_), .Y(_abc_3576_new_n692_));
OR2X2 OR2X2_222 ( .A(_abc_3576_new_n696_), .B(_abc_3576_new_n698_), .Y(_abc_3576_new_n699_));
OR2X2 OR2X2_223 ( .A(_abc_3576_new_n694_), .B(_abc_3576_new_n699_), .Y(_abc_3576_new_n700_));
OR2X2 OR2X2_224 ( .A(_abc_3576_new_n695_), .B(RMAX_REG_5_), .Y(_abc_3576_new_n704_));
OR2X2 OR2X2_225 ( .A(_abc_3576_new_n707_), .B(_abc_3576_new_n709_), .Y(_abc_3576_new_n710_));
OR2X2 OR2X2_226 ( .A(_abc_3576_new_n706_), .B(_abc_3576_new_n710_), .Y(_abc_3576_new_n711_));
OR2X2 OR2X2_227 ( .A(_abc_3576_new_n721_), .B(_abc_3576_new_n722_), .Y(_abc_3576_new_n723_));
OR2X2 OR2X2_228 ( .A(_abc_3576_new_n720_), .B(_abc_3576_new_n723_), .Y(_abc_3576_new_n724_));
OR2X2 OR2X2_229 ( .A(_abc_3576_new_n726_), .B(_abc_3576_new_n727_), .Y(_abc_3576_new_n728_));
OR2X2 OR2X2_23 ( .A(RMIN_REG_3_), .B(RMAX_REG_3_), .Y(_abc_3576_new_n219_));
OR2X2 OR2X2_230 ( .A(_abc_3576_new_n731_), .B(_abc_3576_new_n732_), .Y(_abc_3576_new_n733_));
OR2X2 OR2X2_231 ( .A(_abc_3576_new_n730_), .B(_abc_3576_new_n733_), .Y(_abc_3576_new_n734_));
OR2X2 OR2X2_232 ( .A(_abc_3576_new_n695_), .B(RMIN_REG_5_), .Y(_abc_3576_new_n735_));
OR2X2 OR2X2_233 ( .A(_abc_3576_new_n697_), .B(RMIN_REG_4_), .Y(_abc_3576_new_n736_));
OR2X2 OR2X2_234 ( .A(_abc_3576_new_n739_), .B(_abc_3576_new_n740_), .Y(_abc_3576_new_n741_));
OR2X2 OR2X2_235 ( .A(_abc_3576_new_n738_), .B(_abc_3576_new_n741_), .Y(_abc_3576_new_n742_));
OR2X2 OR2X2_236 ( .A(_abc_3576_new_n743_), .B(_abc_3576_new_n713_), .Y(_abc_3576_new_n744_));
OR2X2 OR2X2_237 ( .A(_abc_3576_new_n749_), .B(STATO_REG_0_), .Y(_abc_3576_new_n750_));
OR2X2 OR2X2_238 ( .A(_abc_3576_new_n753_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n754_));
OR2X2 OR2X2_239 ( .A(_abc_3576_new_n754_), .B(_abc_3576_new_n752_), .Y(n119));
OR2X2 OR2X2_24 ( .A(_abc_3576_new_n222_), .B(_abc_3576_new_n223_), .Y(_abc_3576_new_n224_));
OR2X2 OR2X2_240 ( .A(_abc_3576_new_n757_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n758_));
OR2X2 OR2X2_241 ( .A(_abc_3576_new_n758_), .B(_abc_3576_new_n756_), .Y(n114));
OR2X2 OR2X2_242 ( .A(_abc_3576_new_n761_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n762_));
OR2X2 OR2X2_243 ( .A(_abc_3576_new_n762_), .B(_abc_3576_new_n760_), .Y(n109));
OR2X2 OR2X2_244 ( .A(_abc_3576_new_n765_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n766_));
OR2X2 OR2X2_245 ( .A(_abc_3576_new_n766_), .B(_abc_3576_new_n764_), .Y(n104));
OR2X2 OR2X2_246 ( .A(_abc_3576_new_n769_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n770_));
OR2X2 OR2X2_247 ( .A(_abc_3576_new_n770_), .B(_abc_3576_new_n768_), .Y(n99));
OR2X2 OR2X2_248 ( .A(_abc_3576_new_n773_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n774_));
OR2X2 OR2X2_249 ( .A(_abc_3576_new_n774_), .B(_abc_3576_new_n772_), .Y(n94));
OR2X2 OR2X2_25 ( .A(_abc_3576_new_n221_), .B(_abc_3576_new_n224_), .Y(_abc_3576_new_n225_));
OR2X2 OR2X2_250 ( .A(_abc_3576_new_n777_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n778_));
OR2X2 OR2X2_251 ( .A(_abc_3576_new_n778_), .B(_abc_3576_new_n776_), .Y(n89));
OR2X2 OR2X2_252 ( .A(_abc_3576_new_n781_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n782_));
OR2X2 OR2X2_253 ( .A(_abc_3576_new_n782_), .B(_abc_3576_new_n780_), .Y(n84));
OR2X2 OR2X2_254 ( .A(_abc_3576_new_n712_), .B(_abc_3576_new_n149_), .Y(_abc_3576_new_n784_));
OR2X2 OR2X2_255 ( .A(_abc_3576_new_n788_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n789_));
OR2X2 OR2X2_256 ( .A(_abc_3576_new_n789_), .B(_abc_3576_new_n787_), .Y(n79));
OR2X2 OR2X2_257 ( .A(_abc_3576_new_n792_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n793_));
OR2X2 OR2X2_258 ( .A(_abc_3576_new_n793_), .B(_abc_3576_new_n791_), .Y(n74));
OR2X2 OR2X2_259 ( .A(_abc_3576_new_n796_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n797_));
OR2X2 OR2X2_26 ( .A(RMIN_REG_5_), .B(RMAX_REG_5_), .Y(_abc_3576_new_n226_));
OR2X2 OR2X2_260 ( .A(_abc_3576_new_n797_), .B(_abc_3576_new_n795_), .Y(n69));
OR2X2 OR2X2_261 ( .A(_abc_3576_new_n800_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n801_));
OR2X2 OR2X2_262 ( .A(_abc_3576_new_n801_), .B(_abc_3576_new_n799_), .Y(n64));
OR2X2 OR2X2_263 ( .A(_abc_3576_new_n804_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n805_));
OR2X2 OR2X2_264 ( .A(_abc_3576_new_n805_), .B(_abc_3576_new_n803_), .Y(n59));
OR2X2 OR2X2_265 ( .A(_abc_3576_new_n808_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n809_));
OR2X2 OR2X2_266 ( .A(_abc_3576_new_n809_), .B(_abc_3576_new_n807_), .Y(n54));
OR2X2 OR2X2_267 ( .A(_abc_3576_new_n812_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n813_));
OR2X2 OR2X2_268 ( .A(_abc_3576_new_n813_), .B(_abc_3576_new_n811_), .Y(n49));
OR2X2 OR2X2_269 ( .A(_abc_3576_new_n816_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n817_));
OR2X2 OR2X2_27 ( .A(RMAX_REG_6_), .B(RMIN_REG_6_), .Y(_abc_3576_new_n227_));
OR2X2 OR2X2_270 ( .A(_abc_3576_new_n817_), .B(_abc_3576_new_n815_), .Y(n44));
OR2X2 OR2X2_28 ( .A(_abc_3576_new_n229_), .B(_abc_3576_new_n206_), .Y(_abc_3576_new_n230_));
OR2X2 OR2X2_29 ( .A(_abc_3576_new_n234_), .B(_abc_3576_new_n154_), .Y(_abc_3576_new_n235_));
OR2X2 OR2X2_3 ( .A(RESTART), .B(REG4_REG_1_), .Y(_abc_3576_new_n153_));
OR2X2 OR2X2_30 ( .A(_abc_3576_new_n231_), .B(_abc_3576_new_n235_), .Y(_abc_3576_new_n236_));
OR2X2 OR2X2_31 ( .A(_abc_3576_new_n239_), .B(_abc_3576_new_n240_), .Y(_abc_3576_new_n241_));
OR2X2 OR2X2_32 ( .A(REG4_REG_2_), .B(DATA_IN_2_), .Y(_abc_3576_new_n242_));
OR2X2 OR2X2_33 ( .A(REG4_REG_1_), .B(DATA_IN_1_), .Y(_abc_3576_new_n243_));
OR2X2 OR2X2_34 ( .A(_abc_3576_new_n246_), .B(_abc_3576_new_n247_), .Y(_abc_3576_new_n248_));
OR2X2 OR2X2_35 ( .A(_abc_3576_new_n245_), .B(_abc_3576_new_n248_), .Y(_abc_3576_new_n249_));
OR2X2 OR2X2_36 ( .A(REG4_REG_4_), .B(DATA_IN_4_), .Y(_abc_3576_new_n250_));
OR2X2 OR2X2_37 ( .A(DATA_IN_3_), .B(REG4_REG_3_), .Y(_abc_3576_new_n251_));
OR2X2 OR2X2_38 ( .A(_abc_3576_new_n254_), .B(_abc_3576_new_n255_), .Y(_abc_3576_new_n256_));
OR2X2 OR2X2_39 ( .A(_abc_3576_new_n253_), .B(_abc_3576_new_n256_), .Y(_abc_3576_new_n257_));
OR2X2 OR2X2_4 ( .A(_abc_3576_new_n154_), .B(RMIN_REG_1_), .Y(_abc_3576_new_n155_));
OR2X2 OR2X2_40 ( .A(REG4_REG_5_), .B(DATA_IN_5_), .Y(_abc_3576_new_n258_));
OR2X2 OR2X2_41 ( .A(DATA_IN_6_), .B(REG4_REG_6_), .Y(_abc_3576_new_n259_));
OR2X2 OR2X2_42 ( .A(_abc_3576_new_n264_), .B(_abc_3576_new_n265_), .Y(_abc_3576_new_n266_));
OR2X2 OR2X2_43 ( .A(_abc_3576_new_n261_), .B(_abc_3576_new_n266_), .Y(_abc_3576_new_n267_));
OR2X2 OR2X2_44 ( .A(_abc_3576_new_n269_), .B(AVERAGE), .Y(_abc_3576_new_n270_));
OR2X2 OR2X2_45 ( .A(_abc_3576_new_n270_), .B(RESTART), .Y(_abc_3576_new_n271_));
OR2X2 OR2X2_46 ( .A(_abc_3576_new_n268_), .B(_abc_3576_new_n271_), .Y(_abc_3576_new_n272_));
OR2X2 OR2X2_47 ( .A(_abc_3576_new_n279_), .B(RESTART), .Y(_abc_3576_new_n280_));
OR2X2 OR2X2_48 ( .A(_abc_3576_new_n291_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n292_));
OR2X2 OR2X2_49 ( .A(_abc_3576_new_n289_), .B(_abc_3576_new_n292_), .Y(_abc_3576_new_n293_));
OR2X2 OR2X2_5 ( .A(_abc_3576_new_n158_), .B(_abc_3576_new_n157_), .Y(_abc_3576_new_n159_));
OR2X2 OR2X2_50 ( .A(_abc_3576_new_n293_), .B(_abc_3576_new_n287_), .Y(_abc_3576_new_n294_));
OR2X2 OR2X2_51 ( .A(_abc_3576_new_n283_), .B(_abc_3576_new_n294_), .Y(_abc_3576_new_n295_));
OR2X2 OR2X2_52 ( .A(_abc_3576_new_n295_), .B(_abc_3576_new_n276_), .Y(n352));
OR2X2 OR2X2_53 ( .A(RESTART), .B(REG4_REG_2_), .Y(_abc_3576_new_n297_));
OR2X2 OR2X2_54 ( .A(_abc_3576_new_n303_), .B(_abc_3576_new_n305_), .Y(_abc_3576_new_n306_));
OR2X2 OR2X2_55 ( .A(_abc_3576_new_n307_), .B(_abc_3576_new_n301_), .Y(_abc_3576_new_n308_));
OR2X2 OR2X2_56 ( .A(_abc_3576_new_n197_), .B(_abc_3576_new_n171_), .Y(_abc_3576_new_n312_));
OR2X2 OR2X2_57 ( .A(_abc_3576_new_n313_), .B(_abc_3576_new_n311_), .Y(_abc_3576_new_n316_));
OR2X2 OR2X2_58 ( .A(_abc_3576_new_n318_), .B(_abc_3576_new_n193_), .Y(_abc_3576_new_n321_));
OR2X2 OR2X2_59 ( .A(_abc_3576_new_n327_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n328_));
OR2X2 OR2X2_6 ( .A(_abc_3576_new_n163_), .B(_abc_3576_new_n165_), .Y(_abc_3576_new_n166_));
OR2X2 OR2X2_60 ( .A(_abc_3576_new_n326_), .B(_abc_3576_new_n328_), .Y(_abc_3576_new_n329_));
OR2X2 OR2X2_61 ( .A(_abc_3576_new_n329_), .B(_abc_3576_new_n325_), .Y(_abc_3576_new_n330_));
OR2X2 OR2X2_62 ( .A(_abc_3576_new_n324_), .B(_abc_3576_new_n330_), .Y(_abc_3576_new_n331_));
OR2X2 OR2X2_63 ( .A(_abc_3576_new_n331_), .B(_abc_3576_new_n323_), .Y(n348));
OR2X2 OR2X2_64 ( .A(RESTART), .B(REG4_REG_3_), .Y(_abc_3576_new_n333_));
OR2X2 OR2X2_65 ( .A(_abc_3576_new_n154_), .B(RMIN_REG_3_), .Y(_abc_3576_new_n334_));
OR2X2 OR2X2_66 ( .A(RESTART), .B(DATA_IN_3_), .Y(_abc_3576_new_n337_));
OR2X2 OR2X2_67 ( .A(_abc_3576_new_n154_), .B(RMAX_REG_3_), .Y(_abc_3576_new_n338_));
OR2X2 OR2X2_68 ( .A(_abc_3576_new_n313_), .B(_abc_3576_new_n346_), .Y(_abc_3576_new_n347_));
OR2X2 OR2X2_69 ( .A(_abc_3576_new_n348_), .B(_abc_3576_new_n345_), .Y(_abc_3576_new_n350_));
OR2X2 OR2X2_7 ( .A(_abc_3576_new_n168_), .B(RESTART), .Y(_abc_3576_new_n169_));
OR2X2 OR2X2_70 ( .A(_abc_3576_new_n351_), .B(_abc_3576_new_n349_), .Y(_abc_3576_new_n352_));
OR2X2 OR2X2_71 ( .A(_abc_3576_new_n356_), .B(_abc_3576_new_n354_), .Y(_abc_3576_new_n357_));
OR2X2 OR2X2_72 ( .A(_abc_3576_new_n361_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n362_));
OR2X2 OR2X2_73 ( .A(_abc_3576_new_n360_), .B(_abc_3576_new_n362_), .Y(_abc_3576_new_n363_));
OR2X2 OR2X2_74 ( .A(_abc_3576_new_n363_), .B(_abc_3576_new_n359_), .Y(_abc_3576_new_n364_));
OR2X2 OR2X2_75 ( .A(_abc_3576_new_n358_), .B(_abc_3576_new_n364_), .Y(_abc_3576_new_n365_));
OR2X2 OR2X2_76 ( .A(_abc_3576_new_n365_), .B(_abc_3576_new_n353_), .Y(n344));
OR2X2 OR2X2_77 ( .A(_abc_3576_new_n368_), .B(_abc_3576_new_n369_), .Y(_abc_3576_new_n370_));
OR2X2 OR2X2_78 ( .A(_abc_3576_new_n348_), .B(_abc_3576_new_n341_), .Y(_abc_3576_new_n371_));
OR2X2 OR2X2_79 ( .A(RESTART), .B(REG4_REG_4_), .Y(_abc_3576_new_n373_));
OR2X2 OR2X2_8 ( .A(RESTART), .B(DATA_IN_0_), .Y(_abc_3576_new_n174_));
OR2X2 OR2X2_80 ( .A(_abc_3576_new_n154_), .B(RMIN_REG_4_), .Y(_abc_3576_new_n374_));
OR2X2 OR2X2_81 ( .A(RESTART), .B(DATA_IN_4_), .Y(_abc_3576_new_n376_));
OR2X2 OR2X2_82 ( .A(_abc_3576_new_n154_), .B(RMAX_REG_4_), .Y(_abc_3576_new_n377_));
OR2X2 OR2X2_83 ( .A(_abc_3576_new_n375_), .B(_abc_3576_new_n378_), .Y(_abc_3576_new_n381_));
OR2X2 OR2X2_84 ( .A(_abc_3576_new_n180_), .B(_abc_3576_new_n160_), .Y(_abc_3576_new_n385_));
OR2X2 OR2X2_85 ( .A(_abc_3576_new_n387_), .B(_abc_3576_new_n309_), .Y(_abc_3576_new_n388_));
OR2X2 OR2X2_86 ( .A(_abc_3576_new_n389_), .B(_abc_3576_new_n343_), .Y(_abc_3576_new_n390_));
OR2X2 OR2X2_87 ( .A(_abc_3576_new_n384_), .B(_abc_3576_new_n391_), .Y(_abc_3576_new_n392_));
OR2X2 OR2X2_88 ( .A(_abc_3576_new_n370_), .B(_abc_3576_new_n393_), .Y(_abc_3576_new_n394_));
OR2X2 OR2X2_89 ( .A(_abc_3576_new_n397_), .B(_abc_3576_new_n395_), .Y(_abc_3576_new_n398_));
OR2X2 OR2X2_9 ( .A(_abc_3576_new_n154_), .B(RMAX_REG_0_), .Y(_abc_3576_new_n175_));
OR2X2 OR2X2_90 ( .A(_abc_3576_new_n405_), .B(_abc_3576_new_n148_), .Y(_abc_3576_new_n406_));
OR2X2 OR2X2_91 ( .A(_abc_3576_new_n404_), .B(_abc_3576_new_n406_), .Y(_abc_3576_new_n407_));
OR2X2 OR2X2_92 ( .A(_abc_3576_new_n407_), .B(_abc_3576_new_n403_), .Y(_abc_3576_new_n408_));
OR2X2 OR2X2_93 ( .A(_abc_3576_new_n409_), .B(_abc_3576_new_n408_), .Y(_abc_3576_new_n410_));
OR2X2 OR2X2_94 ( .A(_abc_3576_new_n402_), .B(_abc_3576_new_n410_), .Y(n340));
OR2X2 OR2X2_95 ( .A(RESTART), .B(DATA_IN_5_), .Y(_abc_3576_new_n412_));
OR2X2 OR2X2_96 ( .A(_abc_3576_new_n154_), .B(RMAX_REG_5_), .Y(_abc_3576_new_n413_));
OR2X2 OR2X2_97 ( .A(RESTART), .B(REG4_REG_5_), .Y(_abc_3576_new_n415_));
OR2X2 OR2X2_98 ( .A(_abc_3576_new_n154_), .B(RMIN_REG_5_), .Y(_abc_3576_new_n416_));
OR2X2 OR2X2_99 ( .A(_abc_3576_new_n414_), .B(_abc_3576_new_n417_), .Y(_abc_3576_new_n420_));


endmodule