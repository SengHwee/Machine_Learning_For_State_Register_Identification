
module sdrc_top(\cfg_sdr_width[0] , \cfg_sdr_width[1] , \cfg_colbits[0] , \cfg_colbits[1] , wb_rst_i, wb_clk_i, wb_stb_i, \wb_addr_i[0] , \wb_addr_i[1] , \wb_addr_i[2] , \wb_addr_i[3] , \wb_addr_i[4] , \wb_addr_i[5] , \wb_addr_i[6] , \wb_addr_i[7] , \wb_addr_i[8] , \wb_addr_i[9] , \wb_addr_i[10] , \wb_addr_i[11] , \wb_addr_i[12] , \wb_addr_i[13] , \wb_addr_i[14] , \wb_addr_i[15] , \wb_addr_i[16] , \wb_addr_i[17] , \wb_addr_i[18] , \wb_addr_i[19] , \wb_addr_i[20] , \wb_addr_i[21] , \wb_addr_i[22] , \wb_addr_i[23] , \wb_addr_i[24] , \wb_addr_i[25] , wb_we_i, \wb_dat_i[0] , \wb_dat_i[1] , \wb_dat_i[2] , \wb_dat_i[3] , \wb_dat_i[4] , \wb_dat_i[5] , \wb_dat_i[6] , \wb_dat_i[7] , \wb_dat_i[8] , \wb_dat_i[9] , \wb_dat_i[10] , \wb_dat_i[11] , \wb_dat_i[12] , \wb_dat_i[13] , \wb_dat_i[14] , \wb_dat_i[15] , \wb_dat_i[16] , \wb_dat_i[17] , \wb_dat_i[18] , \wb_dat_i[19] , \wb_dat_i[20] , \wb_dat_i[21] , \wb_dat_i[22] , \wb_dat_i[23] , \wb_dat_i[24] , \wb_dat_i[25] , \wb_dat_i[26] , \wb_dat_i[27] , \wb_dat_i[28] , \wb_dat_i[29] , \wb_dat_i[30] , \wb_dat_i[31] , \wb_sel_i[0] , \wb_sel_i[1] , \wb_sel_i[2] , \wb_sel_i[3] , wb_cyc_i, \wb_cti_i[0] , \wb_cti_i[1] , \wb_cti_i[2] , sdram_clk, sdram_resetn, \sdr_dq[0] , \sdr_dq[1] , \sdr_dq[2] , \sdr_dq[3] , \sdr_dq[4] , \sdr_dq[5] , \sdr_dq[6] , \sdr_dq[7] , \sdr_dq[8] , \sdr_dq[9] , \sdr_dq[10] , \sdr_dq[11] , \sdr_dq[12] , \sdr_dq[13] , \sdr_dq[14] , \sdr_dq[15] , \cfg_req_depth[0] , \cfg_req_depth[1] , cfg_sdr_en, \cfg_sdr_mode_reg[0] , \cfg_sdr_mode_reg[1] , \cfg_sdr_mode_reg[2] , \cfg_sdr_mode_reg[3] , \cfg_sdr_mode_reg[4] , \cfg_sdr_mode_reg[5] , \cfg_sdr_mode_reg[6] , \cfg_sdr_mode_reg[7] , \cfg_sdr_mode_reg[8] , \cfg_sdr_mode_reg[9] , \cfg_sdr_mode_reg[10] , \cfg_sdr_mode_reg[11] , \cfg_sdr_mode_reg[12] , \cfg_sdr_tras_d[0] , \cfg_sdr_tras_d[1] , \cfg_sdr_tras_d[2] , \cfg_sdr_tras_d[3] , \cfg_sdr_trp_d[0] , \cfg_sdr_trp_d[1] , \cfg_sdr_trp_d[2] , \cfg_sdr_trp_d[3] , \cfg_sdr_trcd_d[0] , \cfg_sdr_trcd_d[1] , \cfg_sdr_trcd_d[2] , \cfg_sdr_trcd_d[3] , \cfg_sdr_cas[0] , \cfg_sdr_cas[1] , \cfg_sdr_cas[2] , \cfg_sdr_trcar_d[0] , \cfg_sdr_trcar_d[1] , \cfg_sdr_trcar_d[2] , \cfg_sdr_trcar_d[3] , \cfg_sdr_twr_d[0] , \cfg_sdr_twr_d[1] , \cfg_sdr_twr_d[2] , \cfg_sdr_twr_d[3] , \cfg_sdr_rfsh[0] , \cfg_sdr_rfsh[1] , \cfg_sdr_rfsh[2] , \cfg_sdr_rfsh[3] , \cfg_sdr_rfsh[4] , \cfg_sdr_rfsh[5] , \cfg_sdr_rfsh[6] , \cfg_sdr_rfsh[7] , \cfg_sdr_rfsh[8] , \cfg_sdr_rfsh[9] , \cfg_sdr_rfsh[10] , \cfg_sdr_rfsh[11] , \cfg_sdr_rfmax[0] , \cfg_sdr_rfmax[1] , \cfg_sdr_rfmax[2] , wb_ack_o, \wb_dat_o[0] , \wb_dat_o[1] , \wb_dat_o[2] , \wb_dat_o[3] , \wb_dat_o[4] , \wb_dat_o[5] , \wb_dat_o[6] , \wb_dat_o[7] , \wb_dat_o[8] , \wb_dat_o[9] , \wb_dat_o[10] , \wb_dat_o[11] , \wb_dat_o[12] , \wb_dat_o[13] , \wb_dat_o[14] , \wb_dat_o[15] , \wb_dat_o[16] , \wb_dat_o[17] , \wb_dat_o[18] , \wb_dat_o[19] , \wb_dat_o[20] , \wb_dat_o[21] , \wb_dat_o[22] , \wb_dat_o[23] , \wb_dat_o[24] , \wb_dat_o[25] , \wb_dat_o[26] , \wb_dat_o[27] , \wb_dat_o[28] , \wb_dat_o[29] , \wb_dat_o[30] , \wb_dat_o[31] , sdr_cs_n, sdr_cke, sdr_ras_n, sdr_cas_n, sdr_we_n, \sdr_dqm[0] , \sdr_dqm[1] , \sdr_ba[0] , \sdr_ba[1] , \sdr_addr[0] , \sdr_addr[1] , \sdr_addr[2] , \sdr_addr[3] , \sdr_addr[4] , \sdr_addr[5] , \sdr_addr[6] , \sdr_addr[7] , \sdr_addr[8] , \sdr_addr[9] , \sdr_addr[10] , \sdr_addr[11] , \sdr_addr[12] , sdr_init_done);
  wire _auto_iopadmap_cc_313_execute_24675_0_;
  wire _auto_iopadmap_cc_313_execute_24675_10_;
  wire _auto_iopadmap_cc_313_execute_24675_11_;
  wire _auto_iopadmap_cc_313_execute_24675_12_;
  wire _auto_iopadmap_cc_313_execute_24675_1_;
  wire _auto_iopadmap_cc_313_execute_24675_2_;
  wire _auto_iopadmap_cc_313_execute_24675_3_;
  wire _auto_iopadmap_cc_313_execute_24675_4_;
  wire _auto_iopadmap_cc_313_execute_24675_5_;
  wire _auto_iopadmap_cc_313_execute_24675_6_;
  wire _auto_iopadmap_cc_313_execute_24675_7_;
  wire _auto_iopadmap_cc_313_execute_24675_8_;
  wire _auto_iopadmap_cc_313_execute_24675_9_;
  wire _auto_iopadmap_cc_313_execute_24689_0_;
  wire _auto_iopadmap_cc_313_execute_24689_1_;
  wire _auto_iopadmap_cc_313_execute_24692;
  wire _auto_iopadmap_cc_313_execute_24694;
  wire _auto_iopadmap_cc_313_execute_24696;
  wire _auto_iopadmap_cc_313_execute_24698_0_;
  wire _auto_iopadmap_cc_313_execute_24698_1_;
  wire _auto_iopadmap_cc_313_execute_24701;
  wire _auto_iopadmap_cc_313_execute_24703;
  wire _auto_iopadmap_cc_313_execute_24705;
  wire _auto_iopadmap_cc_313_execute_24707;
  wire _auto_iopadmap_cc_313_execute_24709_0_;
  wire _auto_iopadmap_cc_313_execute_24709_10_;
  wire _auto_iopadmap_cc_313_execute_24709_11_;
  wire _auto_iopadmap_cc_313_execute_24709_12_;
  wire _auto_iopadmap_cc_313_execute_24709_13_;
  wire _auto_iopadmap_cc_313_execute_24709_14_;
  wire _auto_iopadmap_cc_313_execute_24709_15_;
  wire _auto_iopadmap_cc_313_execute_24709_16_;
  wire _auto_iopadmap_cc_313_execute_24709_17_;
  wire _auto_iopadmap_cc_313_execute_24709_18_;
  wire _auto_iopadmap_cc_313_execute_24709_19_;
  wire _auto_iopadmap_cc_313_execute_24709_1_;
  wire _auto_iopadmap_cc_313_execute_24709_20_;
  wire _auto_iopadmap_cc_313_execute_24709_21_;
  wire _auto_iopadmap_cc_313_execute_24709_22_;
  wire _auto_iopadmap_cc_313_execute_24709_23_;
  wire _auto_iopadmap_cc_313_execute_24709_24_;
  wire _auto_iopadmap_cc_313_execute_24709_25_;
  wire _auto_iopadmap_cc_313_execute_24709_26_;
  wire _auto_iopadmap_cc_313_execute_24709_27_;
  wire _auto_iopadmap_cc_313_execute_24709_28_;
  wire _auto_iopadmap_cc_313_execute_24709_29_;
  wire _auto_iopadmap_cc_313_execute_24709_2_;
  wire _auto_iopadmap_cc_313_execute_24709_30_;
  wire _auto_iopadmap_cc_313_execute_24709_31_;
  wire _auto_iopadmap_cc_313_execute_24709_3_;
  wire _auto_iopadmap_cc_313_execute_24709_4_;
  wire _auto_iopadmap_cc_313_execute_24709_5_;
  wire _auto_iopadmap_cc_313_execute_24709_6_;
  wire _auto_iopadmap_cc_313_execute_24709_7_;
  wire _auto_iopadmap_cc_313_execute_24709_8_;
  wire _auto_iopadmap_cc_313_execute_24709_9_;
  wire app_last_rd;
  wire app_last_wr;
  wire app_rd_data_0_;
  wire app_rd_data_10_;
  wire app_rd_data_11_;
  wire app_rd_data_12_;
  wire app_rd_data_13_;
  wire app_rd_data_14_;
  wire app_rd_data_15_;
  wire app_rd_data_16_;
  wire app_rd_data_17_;
  wire app_rd_data_18_;
  wire app_rd_data_19_;
  wire app_rd_data_1_;
  wire app_rd_data_20_;
  wire app_rd_data_21_;
  wire app_rd_data_22_;
  wire app_rd_data_23_;
  wire app_rd_data_24_;
  wire app_rd_data_25_;
  wire app_rd_data_26_;
  wire app_rd_data_27_;
  wire app_rd_data_28_;
  wire app_rd_data_29_;
  wire app_rd_data_2_;
  wire app_rd_data_30_;
  wire app_rd_data_31_;
  wire app_rd_data_3_;
  wire app_rd_data_4_;
  wire app_rd_data_5_;
  wire app_rd_data_6_;
  wire app_rd_data_7_;
  wire app_rd_data_8_;
  wire app_rd_data_9_;
  wire app_rd_valid;
  wire app_req;
  wire app_req_ack;
  wire app_req_ack_bF_buf0;
  wire app_req_ack_bF_buf1;
  wire app_req_ack_bF_buf2;
  wire app_req_ack_bF_buf3;
  wire app_req_ack_bF_buf4;
  wire app_req_ack_bF_buf5;
  wire app_req_ack_bF_buf6;
  wire app_req_addr_0_;
  wire app_req_addr_10_;
  wire app_req_addr_11_;
  wire app_req_addr_12_;
  wire app_req_addr_13_;
  wire app_req_addr_14_;
  wire app_req_addr_15_;
  wire app_req_addr_16_;
  wire app_req_addr_17_;
  wire app_req_addr_18_;
  wire app_req_addr_19_;
  wire app_req_addr_1_;
  wire app_req_addr_20_;
  wire app_req_addr_21_;
  wire app_req_addr_22_;
  wire app_req_addr_23_;
  wire app_req_addr_24_;
  wire app_req_addr_25_;
  wire app_req_addr_2_;
  wire app_req_addr_3_;
  wire app_req_addr_4_;
  wire app_req_addr_5_;
  wire app_req_addr_6_;
  wire app_req_addr_7_;
  wire app_req_addr_8_;
  wire app_req_addr_9_;
  wire app_req_len_0_;
  wire app_req_len_1_;
  wire app_req_len_2_;
  wire app_req_len_3_;
  wire app_req_len_4_;
  wire app_req_len_5_;
  wire app_req_len_6_;
  wire app_req_len_7_;
  wire app_req_len_8_;
  wire app_req_wr_n;
  wire app_wr_data_0_;
  wire app_wr_data_10_;
  wire app_wr_data_11_;
  wire app_wr_data_12_;
  wire app_wr_data_13_;
  wire app_wr_data_14_;
  wire app_wr_data_15_;
  wire app_wr_data_16_;
  wire app_wr_data_17_;
  wire app_wr_data_18_;
  wire app_wr_data_19_;
  wire app_wr_data_1_;
  wire app_wr_data_20_;
  wire app_wr_data_21_;
  wire app_wr_data_22_;
  wire app_wr_data_23_;
  wire app_wr_data_24_;
  wire app_wr_data_25_;
  wire app_wr_data_26_;
  wire app_wr_data_27_;
  wire app_wr_data_28_;
  wire app_wr_data_29_;
  wire app_wr_data_2_;
  wire app_wr_data_30_;
  wire app_wr_data_31_;
  wire app_wr_data_3_;
  wire app_wr_data_4_;
  wire app_wr_data_5_;
  wire app_wr_data_6_;
  wire app_wr_data_7_;
  wire app_wr_data_8_;
  wire app_wr_data_9_;
  wire app_wr_en_n_0_;
  wire app_wr_en_n_1_;
  wire app_wr_en_n_2_;
  wire app_wr_en_n_3_;
  wire app_wr_next_req;
  input \cfg_colbits[0] ;
  input \cfg_colbits[1] ;
  input \cfg_req_depth[0] ;
  input \cfg_req_depth[1] ;
  input \cfg_sdr_cas[0] ;
  input \cfg_sdr_cas[1] ;
  input \cfg_sdr_cas[2] ;
  input cfg_sdr_en;
  input \cfg_sdr_mode_reg[0] ;
  input \cfg_sdr_mode_reg[10] ;
  input \cfg_sdr_mode_reg[11] ;
  input \cfg_sdr_mode_reg[12] ;
  input \cfg_sdr_mode_reg[1] ;
  input \cfg_sdr_mode_reg[2] ;
  input \cfg_sdr_mode_reg[3] ;
  input \cfg_sdr_mode_reg[4] ;
  input \cfg_sdr_mode_reg[5] ;
  input \cfg_sdr_mode_reg[6] ;
  input \cfg_sdr_mode_reg[7] ;
  input \cfg_sdr_mode_reg[8] ;
  input \cfg_sdr_mode_reg[9] ;
  input \cfg_sdr_rfmax[0] ;
  input \cfg_sdr_rfmax[1] ;
  input \cfg_sdr_rfmax[2] ;
  input \cfg_sdr_rfsh[0] ;
  input \cfg_sdr_rfsh[10] ;
  input \cfg_sdr_rfsh[11] ;
  input \cfg_sdr_rfsh[1] ;
  input \cfg_sdr_rfsh[2] ;
  input \cfg_sdr_rfsh[3] ;
  input \cfg_sdr_rfsh[4] ;
  input \cfg_sdr_rfsh[5] ;
  input \cfg_sdr_rfsh[6] ;
  input \cfg_sdr_rfsh[7] ;
  input \cfg_sdr_rfsh[8] ;
  input \cfg_sdr_rfsh[9] ;
  input \cfg_sdr_tras_d[0] ;
  input \cfg_sdr_tras_d[1] ;
  input \cfg_sdr_tras_d[2] ;
  input \cfg_sdr_tras_d[3] ;
  input \cfg_sdr_trcar_d[0] ;
  input \cfg_sdr_trcar_d[1] ;
  input \cfg_sdr_trcar_d[2] ;
  input \cfg_sdr_trcar_d[3] ;
  input \cfg_sdr_trcd_d[0] ;
  input \cfg_sdr_trcd_d[1] ;
  input \cfg_sdr_trcd_d[2] ;
  input \cfg_sdr_trcd_d[3] ;
  input \cfg_sdr_trp_d[0] ;
  input \cfg_sdr_trp_d[1] ;
  input \cfg_sdr_trp_d[2] ;
  input \cfg_sdr_trp_d[3] ;
  input \cfg_sdr_twr_d[0] ;
  input \cfg_sdr_twr_d[1] ;
  input \cfg_sdr_twr_d[2] ;
  input \cfg_sdr_twr_d[3] ;
  input \cfg_sdr_width[0] ;
  input \cfg_sdr_width[1] ;
  wire cfg_sdr_width_1_bF_buf0;
  wire cfg_sdr_width_1_bF_buf1;
  wire cfg_sdr_width_1_bF_buf2;
  wire cfg_sdr_width_1_bF_buf3;
  wire cfg_sdr_width_1_bF_buf4;
  wire cfg_sdr_width_1_bF_buf5;
  output \sdr_addr[0] ;
  output \sdr_addr[10] ;
  output \sdr_addr[11] ;
  output \sdr_addr[12] ;
  output \sdr_addr[1] ;
  output \sdr_addr[2] ;
  output \sdr_addr[3] ;
  output \sdr_addr[4] ;
  output \sdr_addr[5] ;
  output \sdr_addr[6] ;
  output \sdr_addr[7] ;
  output \sdr_addr[8] ;
  output \sdr_addr[9] ;
  output \sdr_ba[0] ;
  output \sdr_ba[1] ;
  output sdr_cas_n;
  output sdr_cke;
  output sdr_cs_n;
  input \sdr_dq[0] ;
  input \sdr_dq[10] ;
  input \sdr_dq[11] ;
  input \sdr_dq[12] ;
  input \sdr_dq[13] ;
  input \sdr_dq[14] ;
  input \sdr_dq[15] ;
  input \sdr_dq[1] ;
  input \sdr_dq[2] ;
  input \sdr_dq[3] ;
  input \sdr_dq[4] ;
  input \sdr_dq[5] ;
  input \sdr_dq[6] ;
  input \sdr_dq[7] ;
  input \sdr_dq[8] ;
  input \sdr_dq[9] ;
  output \sdr_dqm[0] ;
  output \sdr_dqm[1] ;
  output sdr_init_done;
  output sdr_ras_n;
  output sdr_we_n;
  input sdram_clk;
  wire sdram_clk_bF_buf0;
  wire sdram_clk_bF_buf1;
  wire sdram_clk_bF_buf10;
  wire sdram_clk_bF_buf11;
  wire sdram_clk_bF_buf12;
  wire sdram_clk_bF_buf13;
  wire sdram_clk_bF_buf14;
  wire sdram_clk_bF_buf15;
  wire sdram_clk_bF_buf16;
  wire sdram_clk_bF_buf17;
  wire sdram_clk_bF_buf18;
  wire sdram_clk_bF_buf19;
  wire sdram_clk_bF_buf2;
  wire sdram_clk_bF_buf20;
  wire sdram_clk_bF_buf21;
  wire sdram_clk_bF_buf22;
  wire sdram_clk_bF_buf23;
  wire sdram_clk_bF_buf24;
  wire sdram_clk_bF_buf25;
  wire sdram_clk_bF_buf26;
  wire sdram_clk_bF_buf27;
  wire sdram_clk_bF_buf28;
  wire sdram_clk_bF_buf29;
  wire sdram_clk_bF_buf3;
  wire sdram_clk_bF_buf30;
  wire sdram_clk_bF_buf31;
  wire sdram_clk_bF_buf32;
  wire sdram_clk_bF_buf33;
  wire sdram_clk_bF_buf34;
  wire sdram_clk_bF_buf35;
  wire sdram_clk_bF_buf36;
  wire sdram_clk_bF_buf37;
  wire sdram_clk_bF_buf38;
  wire sdram_clk_bF_buf39;
  wire sdram_clk_bF_buf4;
  wire sdram_clk_bF_buf40;
  wire sdram_clk_bF_buf41;
  wire sdram_clk_bF_buf42;
  wire sdram_clk_bF_buf43;
  wire sdram_clk_bF_buf44;
  wire sdram_clk_bF_buf45;
  wire sdram_clk_bF_buf46;
  wire sdram_clk_bF_buf47;
  wire sdram_clk_bF_buf48;
  wire sdram_clk_bF_buf49;
  wire sdram_clk_bF_buf5;
  wire sdram_clk_bF_buf50;
  wire sdram_clk_bF_buf51;
  wire sdram_clk_bF_buf52;
  wire sdram_clk_bF_buf53;
  wire sdram_clk_bF_buf54;
  wire sdram_clk_bF_buf55;
  wire sdram_clk_bF_buf56;
  wire sdram_clk_bF_buf57;
  wire sdram_clk_bF_buf58;
  wire sdram_clk_bF_buf59;
  wire sdram_clk_bF_buf6;
  wire sdram_clk_bF_buf60;
  wire sdram_clk_bF_buf61;
  wire sdram_clk_bF_buf62;
  wire sdram_clk_bF_buf63;
  wire sdram_clk_bF_buf64;
  wire sdram_clk_bF_buf65;
  wire sdram_clk_bF_buf66;
  wire sdram_clk_bF_buf67;
  wire sdram_clk_bF_buf68;
  wire sdram_clk_bF_buf69;
  wire sdram_clk_bF_buf7;
  wire sdram_clk_bF_buf70;
  wire sdram_clk_bF_buf71;
  wire sdram_clk_bF_buf72;
  wire sdram_clk_bF_buf73;
  wire sdram_clk_bF_buf74;
  wire sdram_clk_bF_buf75;
  wire sdram_clk_bF_buf76;
  wire sdram_clk_bF_buf77;
  wire sdram_clk_bF_buf78;
  wire sdram_clk_bF_buf79;
  wire sdram_clk_bF_buf8;
  wire sdram_clk_bF_buf80;
  wire sdram_clk_bF_buf9;
  wire sdram_clk_hier0_bF_buf0;
  wire sdram_clk_hier0_bF_buf1;
  wire sdram_clk_hier0_bF_buf2;
  wire sdram_clk_hier0_bF_buf3;
  wire sdram_clk_hier0_bF_buf4;
  wire sdram_clk_hier0_bF_buf5;
  wire sdram_clk_hier0_bF_buf6;
  wire sdram_clk_hier0_bF_buf7;
  wire sdram_clk_hier0_bF_buf8;
  input sdram_resetn;
  wire sdram_resetn_bF_buf0;
  wire sdram_resetn_bF_buf1;
  wire sdram_resetn_bF_buf10;
  wire sdram_resetn_bF_buf11;
  wire sdram_resetn_bF_buf12;
  wire sdram_resetn_bF_buf13;
  wire sdram_resetn_bF_buf14;
  wire sdram_resetn_bF_buf15;
  wire sdram_resetn_bF_buf16;
  wire sdram_resetn_bF_buf17;
  wire sdram_resetn_bF_buf18;
  wire sdram_resetn_bF_buf19;
  wire sdram_resetn_bF_buf2;
  wire sdram_resetn_bF_buf20;
  wire sdram_resetn_bF_buf21;
  wire sdram_resetn_bF_buf22;
  wire sdram_resetn_bF_buf23;
  wire sdram_resetn_bF_buf24;
  wire sdram_resetn_bF_buf25;
  wire sdram_resetn_bF_buf26;
  wire sdram_resetn_bF_buf27;
  wire sdram_resetn_bF_buf28;
  wire sdram_resetn_bF_buf29;
  wire sdram_resetn_bF_buf3;
  wire sdram_resetn_bF_buf30;
  wire sdram_resetn_bF_buf31;
  wire sdram_resetn_bF_buf32;
  wire sdram_resetn_bF_buf33;
  wire sdram_resetn_bF_buf34;
  wire sdram_resetn_bF_buf35;
  wire sdram_resetn_bF_buf36;
  wire sdram_resetn_bF_buf37;
  wire sdram_resetn_bF_buf38;
  wire sdram_resetn_bF_buf39;
  wire sdram_resetn_bF_buf4;
  wire sdram_resetn_bF_buf40;
  wire sdram_resetn_bF_buf41;
  wire sdram_resetn_bF_buf42;
  wire sdram_resetn_bF_buf43;
  wire sdram_resetn_bF_buf44;
  wire sdram_resetn_bF_buf45;
  wire sdram_resetn_bF_buf46;
  wire sdram_resetn_bF_buf47;
  wire sdram_resetn_bF_buf48;
  wire sdram_resetn_bF_buf49;
  wire sdram_resetn_bF_buf5;
  wire sdram_resetn_bF_buf6;
  wire sdram_resetn_bF_buf7;
  wire sdram_resetn_bF_buf8;
  wire sdram_resetn_bF_buf9;
  wire sdram_resetn_hier0_bF_buf0;
  wire sdram_resetn_hier0_bF_buf1;
  wire sdram_resetn_hier0_bF_buf2;
  wire sdram_resetn_hier0_bF_buf3;
  wire sdram_resetn_hier0_bF_buf4;
  wire sdram_resetn_hier0_bF_buf5;
  wire sdram_resetn_hier0_bF_buf6;
  wire u_sdrc_core_a2x_wrdt_0_;
  wire u_sdrc_core_a2x_wrdt_10_;
  wire u_sdrc_core_a2x_wrdt_11_;
  wire u_sdrc_core_a2x_wrdt_12_;
  wire u_sdrc_core_a2x_wrdt_13_;
  wire u_sdrc_core_a2x_wrdt_14_;
  wire u_sdrc_core_a2x_wrdt_15_;
  wire u_sdrc_core_a2x_wrdt_1_;
  wire u_sdrc_core_a2x_wrdt_2_;
  wire u_sdrc_core_a2x_wrdt_3_;
  wire u_sdrc_core_a2x_wrdt_4_;
  wire u_sdrc_core_a2x_wrdt_5_;
  wire u_sdrc_core_a2x_wrdt_6_;
  wire u_sdrc_core_a2x_wrdt_7_;
  wire u_sdrc_core_a2x_wrdt_8_;
  wire u_sdrc_core_a2x_wrdt_9_;
  wire u_sdrc_core_a2x_wren_n_0_;
  wire u_sdrc_core_a2x_wren_n_1_;
  wire u_sdrc_core_b2r_ack;
  wire u_sdrc_core_b2r_arb_ok;
  wire u_sdrc_core_b2x_addr_0_;
  wire u_sdrc_core_b2x_addr_10_;
  wire u_sdrc_core_b2x_addr_11_;
  wire u_sdrc_core_b2x_addr_12_;
  wire u_sdrc_core_b2x_addr_1_;
  wire u_sdrc_core_b2x_addr_2_;
  wire u_sdrc_core_b2x_addr_3_;
  wire u_sdrc_core_b2x_addr_4_;
  wire u_sdrc_core_b2x_addr_5_;
  wire u_sdrc_core_b2x_addr_6_;
  wire u_sdrc_core_b2x_addr_7_;
  wire u_sdrc_core_b2x_addr_8_;
  wire u_sdrc_core_b2x_addr_9_;
  wire u_sdrc_core_b2x_ba_0_;
  wire u_sdrc_core_b2x_ba_1_;
  wire u_sdrc_core_b2x_cmd_0_;
  wire u_sdrc_core_b2x_cmd_1_;
  wire u_sdrc_core_b2x_idle;
  wire u_sdrc_core_b2x_last;
  wire u_sdrc_core_b2x_len_0_;
  wire u_sdrc_core_b2x_len_1_;
  wire u_sdrc_core_b2x_len_2_;
  wire u_sdrc_core_b2x_len_3_;
  wire u_sdrc_core_b2x_len_4_;
  wire u_sdrc_core_b2x_len_5_;
  wire u_sdrc_core_b2x_len_6_;
  wire u_sdrc_core_b2x_req;
  wire u_sdrc_core_b2x_tras_ok;
  wire u_sdrc_core_b2x_wrap;
  wire u_sdrc_core_pad_sdr_din1_0_;
  wire u_sdrc_core_pad_sdr_din1_10_;
  wire u_sdrc_core_pad_sdr_din1_11_;
  wire u_sdrc_core_pad_sdr_din1_12_;
  wire u_sdrc_core_pad_sdr_din1_13_;
  wire u_sdrc_core_pad_sdr_din1_14_;
  wire u_sdrc_core_pad_sdr_din1_15_;
  wire u_sdrc_core_pad_sdr_din1_1_;
  wire u_sdrc_core_pad_sdr_din1_2_;
  wire u_sdrc_core_pad_sdr_din1_3_;
  wire u_sdrc_core_pad_sdr_din1_4_;
  wire u_sdrc_core_pad_sdr_din1_5_;
  wire u_sdrc_core_pad_sdr_din1_6_;
  wire u_sdrc_core_pad_sdr_din1_7_;
  wire u_sdrc_core_pad_sdr_din1_8_;
  wire u_sdrc_core_pad_sdr_din1_9_;
  wire u_sdrc_core_pad_sdr_din2_0_;
  wire u_sdrc_core_pad_sdr_din2_10_;
  wire u_sdrc_core_pad_sdr_din2_11_;
  wire u_sdrc_core_pad_sdr_din2_12_;
  wire u_sdrc_core_pad_sdr_din2_13_;
  wire u_sdrc_core_pad_sdr_din2_14_;
  wire u_sdrc_core_pad_sdr_din2_15_;
  wire u_sdrc_core_pad_sdr_din2_1_;
  wire u_sdrc_core_pad_sdr_din2_2_;
  wire u_sdrc_core_pad_sdr_din2_3_;
  wire u_sdrc_core_pad_sdr_din2_4_;
  wire u_sdrc_core_pad_sdr_din2_5_;
  wire u_sdrc_core_pad_sdr_din2_6_;
  wire u_sdrc_core_pad_sdr_din2_7_;
  wire u_sdrc_core_pad_sdr_din2_8_;
  wire u_sdrc_core_pad_sdr_din2_9_;
  wire u_sdrc_core_r2b_ba_0_;
  wire u_sdrc_core_r2b_ba_1_;
  wire u_sdrc_core_r2b_caddr_0_;
  wire u_sdrc_core_r2b_caddr_10_;
  wire u_sdrc_core_r2b_caddr_1_;
  wire u_sdrc_core_r2b_caddr_2_;
  wire u_sdrc_core_r2b_caddr_3_;
  wire u_sdrc_core_r2b_caddr_4_;
  wire u_sdrc_core_r2b_caddr_5_;
  wire u_sdrc_core_r2b_caddr_6_;
  wire u_sdrc_core_r2b_caddr_7_;
  wire u_sdrc_core_r2b_caddr_8_;
  wire u_sdrc_core_r2b_caddr_9_;
  wire u_sdrc_core_r2b_last;
  wire u_sdrc_core_r2b_len_0_;
  wire u_sdrc_core_r2b_len_1_;
  wire u_sdrc_core_r2b_len_2_;
  wire u_sdrc_core_r2b_len_3_;
  wire u_sdrc_core_r2b_len_4_;
  wire u_sdrc_core_r2b_len_5_;
  wire u_sdrc_core_r2b_len_6_;
  wire u_sdrc_core_r2b_raddr_0_;
  wire u_sdrc_core_r2b_raddr_10_;
  wire u_sdrc_core_r2b_raddr_11_;
  wire u_sdrc_core_r2b_raddr_12_;
  wire u_sdrc_core_r2b_raddr_1_;
  wire u_sdrc_core_r2b_raddr_2_;
  wire u_sdrc_core_r2b_raddr_3_;
  wire u_sdrc_core_r2b_raddr_4_;
  wire u_sdrc_core_r2b_raddr_5_;
  wire u_sdrc_core_r2b_raddr_6_;
  wire u_sdrc_core_r2b_raddr_7_;
  wire u_sdrc_core_r2b_raddr_8_;
  wire u_sdrc_core_r2b_raddr_9_;
  wire u_sdrc_core_r2b_req;
  wire u_sdrc_core_r2b_start;
  wire u_sdrc_core_r2b_wrap;
  wire u_sdrc_core_r2b_write;
  wire u_sdrc_core_r2x_idle;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n204_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n205_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n207_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n208;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n211_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n213;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n216_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n217_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n218_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n219_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n221_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n222;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n223_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n223_1_bF_buf0;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n223_1_bF_buf1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n223_1_bF_buf2;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n223_1_bF_buf3;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n224_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n225_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n226_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n227;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n227_bF_buf0;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n227_bF_buf1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n227_bF_buf2;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n227_bF_buf3;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n228_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n229;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n230_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n232_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n233_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n234;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n235_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n236;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n237_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n239_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n240_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n241;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n242_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n243;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n244_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n245_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n246_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n247_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n248;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n249_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n251_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n252_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n253_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n254_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n255;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n256_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n257;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n258_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n259_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n260_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n261_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n262;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n264;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n265_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n266_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n267_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n268_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n269;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n270_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n271;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n272_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n273_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n274_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n275_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n276;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n278;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n279_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n280_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n281_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n282_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n283;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n283_bF_buf0;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n283_bF_buf1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n283_bF_buf2;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n283_bF_buf3;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n284_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n285;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n286_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n287_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n288_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n289_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n290;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n291_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n292_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n293;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n294_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n295_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n296_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n297;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n298_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n299_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n300;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n301_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n302_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n303_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n304;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n305_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n306_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n308_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n309_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n310;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n311_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n312;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n313_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n315;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n316;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n317_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n318;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n319;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n320_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n321;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n322_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n323;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n324_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n325_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n326_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n328_1;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n329;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n330;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n331;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n332;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n333;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n335;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n336;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n337;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n338;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n339;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n340;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n341;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n342;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n343;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n344;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n345;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n347;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n348;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n349;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n350;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n351;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n352;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n354;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n355;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n356;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n357;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n358;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n359;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n360;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n361;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n362;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n363;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n365;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n366;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n367;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n368;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n370;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n371;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n372;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n373;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n374;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n375;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n376;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n377;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n379;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n380;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n381;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n382;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n383;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n384;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n385;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n386;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n388;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n389;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n390;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n391;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n392;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n393;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n394;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n395;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n397;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n398;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n399;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n400;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n401;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n402;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n403;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n404;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n406;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n407;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n408;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n409;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n410;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n411;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n412;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n413;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n415;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n416;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n417;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n418;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n419;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n420;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n421;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n422;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n424;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n425;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n426;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n427;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n428;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n429;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n430;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n431;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n433;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n434;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n435;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n436;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n437;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n438;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n439;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n440;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n442;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n443;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n444;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n445;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n446;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n447;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n448;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n449;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n451;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n452;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n453;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n454;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n455;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n456;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n457;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n458;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n460;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n461;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n462;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n463;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n464;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n465;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n466;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n467;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n469;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n470;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n471;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n472;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n473;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n474;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n475;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n476;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n478;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n479;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n480;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n481;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n482;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n483;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n484;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n485;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n487;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n488;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n489;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n490;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n491;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n492;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n493;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n494;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n496;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n497;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n498;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n499;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n500;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n501;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n502;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n503;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n505;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n506;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n507;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n508;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n509;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n510;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n511;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n512;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n514;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n515;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n516;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n517;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n518;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n519;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n520;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n521;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n523;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n524;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n525;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n526;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n527;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n528;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n529;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n530;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n532;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n533;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n534;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n535;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n536;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n537;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n538;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n539;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n541;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n542;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n543;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n544;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n545;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n546;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n547;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n548;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n550;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n551;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n552;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n553;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n554;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n555;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n556;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n557;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n594;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n595;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n596;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n597;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n598;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n599;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n608;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n609;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n610;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n611;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n612;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n613;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n615;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n616;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n617;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n618;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n619;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n620;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n621;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n622;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n623;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n625;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n626;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n627;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n628;
  wire u_sdrc_core_u_bank_ctl__abc_21249_n631;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_17422_n55;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_17422_n61;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_17422_n66;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_17422_n82;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_17422_n90;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n249_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n250_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n251;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n253_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n254;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n255_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n256_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n257;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n258_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n259_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n260;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n261_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n262_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n263;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n264_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n265_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n266;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n267_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n268_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n269;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n270_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n271_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n272;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n273_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n274_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n275;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n276_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n277_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n278;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n279_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n280_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n281;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n282_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n283_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n284_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n285;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n286_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n287_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n288_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n289;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n290_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n291_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n292_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n293;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n294_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n295_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n296_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n297;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n298_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n299_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n300_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n301;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n302_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n303_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n304_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n305;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n306_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n307_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n308_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n309;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n310_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n311_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n312_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n313;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n314_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n315_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n316_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n317;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n318_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n319_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n320_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n321;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n322_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n323_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n324_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n325;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n326_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n327_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n328_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n329;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n330_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n331_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n332_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n333;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n335;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n336;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n337;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n338_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n339_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n340;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n342;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n343_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n344_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n345;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n346;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n348_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n349_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n350;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n351;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n353_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n354_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n355;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n356;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n357;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n358_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n359_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n360;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n361;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n362;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n364_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n365;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n366;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n367;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n368_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n369_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n370;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n371;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n372;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n373_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n374_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n376;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n377;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n379_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n380;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n381;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n382;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n383_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n384_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n385;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n386_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n387_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n388;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n389;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n390;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n392_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n393;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n394_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n395_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n396_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n397_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n399_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n400_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n401_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n402_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n403_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n404_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n406_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n407_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n408_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n409_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n411_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n412_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n413_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n414_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n415_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n416;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n417_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n418;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n419_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n420_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n421;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n422;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n424;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n425;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n426;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n427_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n428_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n429;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n430;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n431_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n432;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n433;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n434_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n435_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n437_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n438_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n439_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n440_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n441;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n442;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n443;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n444_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n445_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n446_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n448_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n449_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n450;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n451;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n452;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n453_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n454;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf0;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf2;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf3;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf4;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf5;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n473;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n474;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n475;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n477;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n478;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n479;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n481;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n482;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n483;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n485;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n486;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n487;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n489;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n490;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n491;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n493;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n494;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n495;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n497;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n498;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n499;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n501;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n502;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n503;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n505;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n506;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n507;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n509;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n510;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n511;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n513;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n514;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n515;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n517;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n518;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n519;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n521;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n522;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n523;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n525;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n526;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n527;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n529;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n530;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n531;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n533;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n534;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n535;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n537;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n538;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n539;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n541;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n542;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n543;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n545;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n546;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n547;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n549;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n550;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n551;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n553;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n554;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n555;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n557;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n558;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n559;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n561;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n562;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n563;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n565;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n566;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n567;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n569;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n570;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n571;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n573;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n574;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n575;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n577;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n578;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n579;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n581;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n582;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n583;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n585;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n586;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n587;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n589;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n590;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n591;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n593;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n594;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n595;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n597;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n598;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n599;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n601;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n602;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n603;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n605;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n606;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n607;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n609;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n610;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n612;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n613;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n615;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n616;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n618;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n619;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n621;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n622;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n624;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n625;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n627;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n628;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n630;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n631;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n633;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n634;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n636;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n637;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n639;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n640;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n642;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n643;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n645;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n646;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n648;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n649;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n651;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n652;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n654;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n655;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n657;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n658;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n660;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n661;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n663;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n664;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n666;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n667;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n669;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n670;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n672;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n673;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n675;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n676;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n678;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n679;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n681;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n682;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n685;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n688;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n689;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n703;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n704;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n706;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n707;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n709;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n710;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n712;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n713;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n715;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n716;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n718;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n719;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n721;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n722;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n724;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n725;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n727;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n728;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n729;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n730;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n731;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n732;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n733;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n734;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n735;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n736;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n737;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n742;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n743;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n745;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n749;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n750;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n756;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n757;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n758;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n760;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n761;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n762;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n764;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n765;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n766;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n768;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n769;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n770;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf0;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf2;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf3;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf4;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_0_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_10_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_11_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_12_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_1_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_2_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_3_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_4_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_5_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_6_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_7_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_8_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_9_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_cmd_0_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_cmd_1_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_cmd_r_0__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_cmd_r_1__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_last;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_len_0_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_len_1_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_len_2_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_len_3_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_len_4_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_len_5_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_len_6_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_req;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_wrap;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_prech_page_closed;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_0_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_0__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_10_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_10__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_11_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_11__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_12_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_12__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_1_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_1__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_2_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_2__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_3_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_3__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_4_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_4__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_5_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_5__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_6_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_6__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_7_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_7__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_8_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_8__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_9_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_9__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_0_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_2_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_2_bF_buf0;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_2_bF_buf1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_2_bF_buf2;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_2_bF_buf3;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_3_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_4_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_4_bF_buf0;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_4_bF_buf1;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_4_bF_buf2;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_4_bF_buf3;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_valid;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_bank_valid_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_0_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_0__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_10_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_10__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_11_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_11__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_12_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_12__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_1_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_1__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_2_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_2__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_3_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_3__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_4_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_4__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_5_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_5__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_6_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_6__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_7_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_7__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_8_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_8__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_9_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_9__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_last;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_last_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_0_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_0__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_1_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_1__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_2_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_2__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_3_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_3__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_4_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_4__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_5_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_5__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_6_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_6__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_0_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_0__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_10_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_10__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_11_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_11__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_12_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_12__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_1_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_1__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_2_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_2__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_3_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_3__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_4_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_4__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_5_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_5__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_6_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_6__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_7_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_7__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_8_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_8__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_9_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_9__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_sdr_dma_last;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_sdr_dma_last_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_wrap;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_wrap_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_write;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_l_write_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_r2b_req;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_timer0_0_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_timer0_0__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_timer0_1_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_timer0_1__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_timer0_2_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_timer0_2__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_timer0_3_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_timer0_3__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_timer0_tc;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_timer0_tc_r_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_tras_cntr_0_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_tras_cntr_0__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_tras_cntr_1_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_tras_cntr_1__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_tras_cntr_2_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_tras_cntr_2__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_tras_cntr_3_;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_tras_cntr_3__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_tras_ok;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_tras_ok_r_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_ack;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_act_ok;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_act_ok_r_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_act_ok_t;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_pre_ok;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_pre_ok_r_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_pre_ok_t;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_rdok;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_rdok_r;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_rdok_r_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_refresh;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_wrok;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_wrok_r;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_wrok_r_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_xfr_ok;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_xfr_ok_r;
  wire u_sdrc_core_u_bank_ctl_bank0_fsm_xfr_ok_r_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_17422_n55;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_17422_n61;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_17422_n66;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_17422_n82;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_17422_n90;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n249_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n250_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n251;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n253_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n254;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n255_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n256_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n257;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n258_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n259_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n260;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n261_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n262_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n263;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n264_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n265_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n266;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n267_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n268_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n269;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n270_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n271_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n272;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n273_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n274_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n275;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n276_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n277_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n278;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n279_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n280_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n281;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n282_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n283_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n284_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n285;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n286_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n287_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n288_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n289;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n290_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n291_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n292_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n293;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n294_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n295_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n296_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n297;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n298_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n299_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n300_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n301;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n302_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n303_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n304_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n305;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n306_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n307_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n308_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n309;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n310_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n311_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n312_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n313;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n314_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n315_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n316_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n317;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n318_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n319_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n320_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n321;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n322_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n323_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n324_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n325;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n326_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n327_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n328_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n329;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n330_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n331_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n332_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n333;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n335;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n336;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n337;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n338_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n339_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n340;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n342;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n343_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n344_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n345;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n346;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n348_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n349_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n350;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n351;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n353_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n354_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n355;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n356;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n357;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n358_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n359_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n360;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n361;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n362;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n364_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n365;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n366;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n367;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n368_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n369_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n370;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n371;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n372;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n373_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n374_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n376;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n377;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n379_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n380;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n381;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n382;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n383_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n384_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n385;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n386_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n387_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n388;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n389;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n390;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n392_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n393;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n394_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n395_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n396_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n397_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n399_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n400_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n401_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n402_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n403_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n404_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n406_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n407_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n408_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n409_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n411_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n412_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n413_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n414_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n415_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n416;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n417_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n418;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n419_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n420_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n421;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n422;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n424;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n425;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n426;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n427_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n428_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n429;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n430;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n431_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n432;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n433;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n434_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n435_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n437_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n438_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n439_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n440_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n441;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n442;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n443;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n444_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n445_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n446_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n448_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n449_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n450;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n451;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n452;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n453_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n454;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf0;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf2;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf3;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf4;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf5;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n473;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n474;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n475;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n477;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n478;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n479;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n481;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n482;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n483;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n485;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n486;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n487;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n489;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n490;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n491;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n493;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n494;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n495;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n497;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n498;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n499;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n501;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n502;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n503;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n505;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n506;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n507;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n509;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n510;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n511;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n513;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n514;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n515;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n517;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n518;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n519;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n521;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n522;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n523;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n525;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n526;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n527;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n529;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n530;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n531;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n533;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n534;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n535;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n537;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n538;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n539;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n541;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n542;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n543;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n545;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n546;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n547;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n549;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n550;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n551;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n553;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n554;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n555;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n557;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n558;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n559;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n561;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n562;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n563;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n565;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n566;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n567;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n569;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n570;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n571;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n573;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n574;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n575;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n577;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n578;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n579;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n581;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n582;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n583;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n585;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n586;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n587;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n589;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n590;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n591;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n593;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n594;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n595;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n597;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n598;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n599;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n601;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n602;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n603;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n605;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n606;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n607;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n609;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n610;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n612;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n613;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n615;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n616;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n618;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n619;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n621;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n622;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n624;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n625;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n627;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n628;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n630;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n631;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n633;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n634;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n636;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n637;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n639;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n640;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n642;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n643;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n645;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n646;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n648;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n649;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n651;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n652;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n654;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n655;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n657;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n658;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n660;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n661;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n663;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n664;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n666;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n667;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n669;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n670;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n672;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n673;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n675;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n676;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n678;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n679;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n681;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n682;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n685;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n688;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n689;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n703;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n704;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n706;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n707;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n709;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n710;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n712;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n713;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n715;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n716;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n718;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n719;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n721;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n722;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n724;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n725;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n727;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n728;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n729;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n730;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n731;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n732;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n733;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n734;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n735;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n736;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n737;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n742;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n743;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n745;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n749;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n750;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n756;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n757;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n758;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n760;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n761;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n762;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n764;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n765;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n766;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n768;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n769;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n770;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf0;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf2;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf3;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf4;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_0_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_10_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_11_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_12_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_1_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_2_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_3_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_4_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_5_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_6_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_7_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_8_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_9_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_cmd_0_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_cmd_1_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_cmd_r_0__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_cmd_r_1__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_last;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_len_0_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_len_1_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_len_2_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_len_3_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_len_4_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_len_5_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_len_6_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_req;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_wrap;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_prech_page_closed;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_0_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_0__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_10_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_10__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_11_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_11__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_12_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_12__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_1_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_1__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_2_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_2__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_3_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_3__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_4_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_4__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_5_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_5__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_6_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_6__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_7_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_7__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_8_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_8__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_9_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_9__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_0_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_2_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_2_bF_buf0;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_2_bF_buf1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_2_bF_buf2;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_2_bF_buf3;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_3_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_4_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_4_bF_buf0;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_4_bF_buf1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_4_bF_buf2;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_4_bF_buf3;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_valid;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_bank_valid_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_0_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_0__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_10_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_10__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_11_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_11__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_12_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_12__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_1_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_1__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_2_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_2__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_3_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_3__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_4_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_4__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_5_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_5__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_6_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_6__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_7_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_7__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_8_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_8__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_9_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_9__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_last;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_last_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_0_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_0__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_1_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_1__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_2_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_2__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_3_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_3__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_4_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_4__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_5_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_5__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_6_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_6__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_0_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_0__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_10_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_10__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_11_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_11__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_12_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_12__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_1_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_1__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_2_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_2__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_3_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_3__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_4_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_4__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_5_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_5__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_6_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_6__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_7_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_7__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_8_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_8__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_9_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_9__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_sdr_dma_last;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_sdr_dma_last_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_wrap;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_wrap_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_write;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_l_write_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_r2b_req;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_timer0_0_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_timer0_0__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_timer0_1_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_timer0_1__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_timer0_2_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_timer0_2__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_timer0_3_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_timer0_3__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_timer0_tc;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_timer0_tc_r_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_tras_cntr_0_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_tras_cntr_0__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_tras_cntr_1_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_tras_cntr_1__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_tras_cntr_2_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_tras_cntr_2__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_tras_cntr_3_;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_tras_cntr_3__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_tras_ok;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_tras_ok_r_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_x2b_ack;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_x2b_act_ok_r_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_x2b_act_ok_t;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_x2b_pre_ok_r_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_x2b_pre_ok_t;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_x2b_rdok_r;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_x2b_rdok_r_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_x2b_wrok_r;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_x2b_wrok_r_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf0;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf1;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf2;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf3;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf4;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_r;
  wire u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_r_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_17422_n55;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_17422_n61;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_17422_n66;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_17422_n82;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_17422_n90;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n249_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n250_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n251;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n253_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n254;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n255_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n256_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n257;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n258_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n259_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n260;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n261_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n262_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n263;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n264_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n265_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n266;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n267_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n268_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n269;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n270_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n271_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n272;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n273_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n274_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n275;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n276_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n277_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n278;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n279_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n280_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n281;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n282_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n283_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n284_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n285;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n286_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n287_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n288_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n289;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n290_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n291_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n292_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n293;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n294_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n295_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n296_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n297;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n298_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n299_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n300_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n301;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n302_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n303_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n304_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n305;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n306_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n307_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n308_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n309;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n310_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n311_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n312_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n313;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n314_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n315_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n316_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n317;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n318_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n319_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n320_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n321;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n322_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n323_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n324_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n325;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n326_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n327_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n328_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n329;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n330_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n331_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n332_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n333;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n335;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n336;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n337;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n338_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n339_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n340;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n342;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n343_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n344_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n345;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n346;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n348_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n349_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n350;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n351;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n353_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n354_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n355;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n356;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n357;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n358_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n359_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n360;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n361;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n362;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n364_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n365;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n366;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n367;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n368_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n369_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n370;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n371;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n372;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n373_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n374_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n376;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n377;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n379_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n380;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n381;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n382;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n383_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n384_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n385;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n386_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n387_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n388;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n389;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n390;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n392_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n393;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n394_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n395_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n396_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n397_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n399_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n400_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n401_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n402_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n403_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n404_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n406_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n407_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n408_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n409_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n411_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n412_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n413_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n414_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n415_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n416;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n417_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n418;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n419_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n420_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n421;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n422;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n424;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n425;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n426;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n427_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n428_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n429;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n430;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n431_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n432;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n433;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n434_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n435_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n437_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n438_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n439_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n440_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n441;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n442;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n443;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n444_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n445_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n446_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n448_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n449_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n450;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n451;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n452;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n453_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n454;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf0;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf2;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf3;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf4;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf5;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n473;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n474;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n475;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n477;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n478;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n479;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n481;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n482;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n483;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n485;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n486;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n487;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n489;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n490;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n491;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n493;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n494;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n495;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n497;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n498;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n499;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n501;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n502;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n503;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n505;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n506;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n507;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n509;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n510;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n511;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n513;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n514;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n515;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n517;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n518;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n519;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n521;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n522;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n523;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n525;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n526;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n527;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n529;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n530;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n531;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n533;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n534;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n535;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n537;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n538;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n539;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n541;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n542;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n543;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n545;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n546;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n547;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n549;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n550;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n551;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n553;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n554;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n555;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n557;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n558;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n559;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n561;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n562;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n563;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n565;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n566;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n567;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n569;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n570;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n571;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n573;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n574;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n575;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n577;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n578;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n579;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n581;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n582;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n583;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n585;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n586;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n587;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n589;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n590;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n591;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n593;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n594;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n595;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n597;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n598;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n599;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n601;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n602;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n603;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n605;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n606;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n607;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n609;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n610;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n612;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n613;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n615;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n616;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n618;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n619;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n621;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n622;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n624;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n625;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n627;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n628;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n630;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n631;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n633;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n634;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n636;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n637;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n639;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n640;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n642;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n643;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n645;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n646;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n648;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n649;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n651;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n652;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n654;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n655;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n657;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n658;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n660;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n661;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n663;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n664;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n666;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n667;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n669;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n670;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n672;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n673;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n675;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n676;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n678;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n679;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n681;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n682;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n685;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n688;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n689;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n703;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n704;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n706;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n707;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n709;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n710;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n712;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n713;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n715;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n716;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n718;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n719;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n721;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n722;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n724;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n725;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n727;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n728;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n729;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n730;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n731;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n732;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n733;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n734;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n735;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n736;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n737;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n742;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n743;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n745;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n749;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n750;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n756;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n757;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n758;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n760;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n761;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n762;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n764;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n765;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n766;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n768;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n769;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n770;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf0;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf2;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf3;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf4;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_0_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_10_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_11_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_12_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_1_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_2_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_3_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_4_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_5_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_6_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_7_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_8_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_9_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_cmd_0_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_cmd_1_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_cmd_r_0__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_cmd_r_1__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_last;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_len_0_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_len_1_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_len_2_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_len_3_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_len_4_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_len_5_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_len_6_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_req;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_wrap;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_prech_page_closed;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_0_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_0__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_10_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_10__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_11_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_11__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_12_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_12__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_1_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_1__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_2_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_2__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_3_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_3__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_4_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_4__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_5_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_5__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_6_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_6__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_7_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_7__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_8_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_8__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_9_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_9__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_0_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_2_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_2_bF_buf0;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_2_bF_buf1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_2_bF_buf2;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_2_bF_buf3;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_3_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_4_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_4_bF_buf0;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_4_bF_buf1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_4_bF_buf2;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_4_bF_buf3;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_valid;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_bank_valid_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_0_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_0__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_10_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_10__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_11_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_11__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_12_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_12__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_1_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_1__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_2_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_2__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_3_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_3__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_4_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_4__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_5_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_5__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_6_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_6__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_7_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_7__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_8_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_8__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_9_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_9__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_last;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_last_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_0_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_0__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_1_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_1__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_2_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_2__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_3_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_3__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_4_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_4__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_5_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_5__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_6_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_6__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_0_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_0__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_10_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_10__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_11_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_11__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_12_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_12__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_1_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_1__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_2_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_2__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_3_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_3__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_4_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_4__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_5_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_5__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_6_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_6__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_7_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_7__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_8_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_8__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_9_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_9__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_sdr_dma_last;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_sdr_dma_last_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_wrap;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_wrap_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_write;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_l_write_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_r2b_req;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_timer0_0_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_timer0_0__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_timer0_1_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_timer0_1__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_timer0_2_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_timer0_2__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_timer0_3_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_timer0_3__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_timer0_tc;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_timer0_tc_r_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_tras_cntr_0_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_tras_cntr_0__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_tras_cntr_1_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_tras_cntr_1__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_tras_cntr_2_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_tras_cntr_2__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_tras_cntr_3_;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_tras_cntr_3__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_tras_ok;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_tras_ok_r_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_x2b_ack;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_x2b_act_ok_r_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_x2b_act_ok_t;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_x2b_pre_ok_r_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_x2b_pre_ok_t;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_x2b_rdok_r;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_x2b_rdok_r_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_x2b_wrok_r;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_x2b_wrok_r_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf0;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf1;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf2;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf3;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf4;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_r;
  wire u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_r_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_17422_n55;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_17422_n61;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_17422_n66;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_17422_n82;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_17422_n90;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n249_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n250_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n251;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n253_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n254;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n255_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n256_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n257;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n258_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n259_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n260;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n261_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n262_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n263;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n264_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n265_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n266;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n267_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n268_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n269;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n270_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n271_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n272;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n273_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n274_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n275;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n276_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n277_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n278;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n279_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n280_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n281;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n282_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n283_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n284_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n285;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n286_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n287_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n288_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n289;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n290_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n291_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n292_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n293;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n294_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n295_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n296_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n297;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n298_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n299_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n300_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n301;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n302_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n303_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n304_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n305;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n306_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n307_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n308_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n309;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n310_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n311_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n312_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n313;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n314_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n315_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n316_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n317;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n318_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n319_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n320_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n321;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n322_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n323_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n324_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n325;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n326_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n327_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n328_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n329;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n330_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n331_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n332_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n333;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n335;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n336;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n337;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n338_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n339_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n340;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n342;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n343_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n344_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n345;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n346;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n348_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n349_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n350;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n351;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n353_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n354_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n355;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n356;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n357;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n358_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n359_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n360;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n361;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n362;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n364_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n365;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n366;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n367;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n368_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n369_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n370;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n371;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n372;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n373_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n374_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n376;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n377;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n379_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n380;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n381;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n382;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n383_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n384_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n385;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n386_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n387_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n388;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n389;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n390;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n392_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n393;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n394_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n395_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n396_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n397_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n399_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n400_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n401_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n402_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n403_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n404_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n406_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n407_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n408_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n409_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n411_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n412_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n413_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n414_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n415_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n416;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n417_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n418;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n419_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n420_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n421;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n422;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n424;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n425;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n426;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n427_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n428_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n429;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n430;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n431_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n432;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n433;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n434_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n435_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n437_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n438_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n439_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n440_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n441;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n442;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n443;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n444_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n445_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n446_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n448_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n449_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n450;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n451;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n452;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n453_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n454;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf0;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf2;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf3;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf4;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf5;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n473;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n474;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n475;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n477;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n478;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n479;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n481;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n482;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n483;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n485;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n486;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n487;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n489;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n490;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n491;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n493;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n494;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n495;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n497;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n498;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n499;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n501;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n502;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n503;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n505;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n506;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n507;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n509;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n510;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n511;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n513;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n514;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n515;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n517;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n518;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n519;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n521;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n522;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n523;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n525;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n526;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n527;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n529;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n530;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n531;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n533;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n534;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n535;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n537;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n538;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n539;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n541;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n542;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n543;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n545;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n546;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n547;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n549;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n550;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n551;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n553;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n554;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n555;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n557;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n558;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n559;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n561;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n562;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n563;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n565;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n566;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n567;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n569;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n570;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n571;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n573;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n574;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n575;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n577;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n578;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n579;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n581;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n582;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n583;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n585;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n586;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n587;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n589;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n590;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n591;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n593;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n594;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n595;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n597;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n598;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n599;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n601;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n602;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n603;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n605;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n606;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n607;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n609;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n610;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n612;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n613;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n615;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n616;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n618;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n619;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n621;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n622;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n624;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n625;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n627;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n628;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n630;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n631;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n633;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n634;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n636;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n637;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n639;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n640;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n642;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n643;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n645;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n646;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n648;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n649;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n651;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n652;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n654;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n655;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n657;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n658;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n660;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n661;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n663;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n664;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n666;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n667;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n669;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n670;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n672;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n673;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n675;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n676;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n678;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n679;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n681;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n682;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n685;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n688;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n689;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n703;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n704;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n706;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n707;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n709;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n710;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n712;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n713;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n715;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n716;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n718;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n719;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n721;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n722;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n724;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n725;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n727;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n728;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n729;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n730;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n731;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n732;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n733;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n734;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n735;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n736;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n737;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n742;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n743;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n745;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n749;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n750;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n756;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n757;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n758;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n760;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n761;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n762;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n764;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n765;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n766;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n768;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n769;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n770;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf0;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf2;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf3;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf4;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_0_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_10_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_11_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_12_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_1_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_2_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_3_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_4_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_5_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_6_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_7_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_8_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_9_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_cmd_0_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_cmd_1_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_cmd_r_0__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_cmd_r_1__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_last;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_len_0_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_len_1_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_len_2_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_len_3_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_len_4_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_len_5_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_len_6_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_req;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_wrap;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_prech_page_closed;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_0_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_0__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_10_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_10__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_11_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_11__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_12_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_12__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_1_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_1__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_2_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_2__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_3_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_3__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_4_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_4__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_5_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_5__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_6_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_6__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_7_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_7__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_8_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_8__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_9_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_9__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_0_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_2_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_2_bF_buf0;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_2_bF_buf1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_2_bF_buf2;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_2_bF_buf3;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_3_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_4_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_4_bF_buf0;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_4_bF_buf1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_4_bF_buf2;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_4_bF_buf3;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_valid;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_bank_valid_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_0_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_0__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_10_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_10__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_11_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_11__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_12_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_12__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_1_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_1__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_2_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_2__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_3_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_3__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_4_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_4__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_5_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_5__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_6_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_6__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_7_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_7__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_8_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_8__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_9_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_9__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_last;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_last_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_0_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_0__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_1_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_1__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_2_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_2__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_3_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_3__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_4_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_4__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_5_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_5__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_6_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_6__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_0_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_0__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_10_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_10__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_11_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_11__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_12_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_12__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_1_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_1__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_2_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_2__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_3_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_3__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_4_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_4__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_5_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_5__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_6_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_6__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_7_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_7__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_8_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_8__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_9_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_9__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_sdr_dma_last;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_sdr_dma_last_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_wrap;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_wrap_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_write;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_l_write_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_r2b_req;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_timer0_0_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_timer0_0__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_timer0_1_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_timer0_1__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_timer0_2_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_timer0_2__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_timer0_3_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_timer0_3__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_timer0_tc;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_timer0_tc_r_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_tras_cntr_0_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_tras_cntr_0__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_tras_cntr_1_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_tras_cntr_1__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_tras_cntr_2_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_tras_cntr_2__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_tras_cntr_3_;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_tras_cntr_3__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_tras_ok;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_tras_ok_r_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_x2b_ack;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_x2b_act_ok_r_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_x2b_act_ok_t;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_x2b_pre_ok_r_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_x2b_pre_ok_t;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_x2b_rdok_r;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_x2b_rdok_r_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_x2b_wrok_r;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_x2b_wrok_r_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf0;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf1;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf2;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf3;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf4;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_r;
  wire u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_r_FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_rank_ba_0__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_rank_ba_1__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_rank_ba_2_;
  wire u_sdrc_core_u_bank_ctl_rank_ba_2__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_rank_ba_3_;
  wire u_sdrc_core_u_bank_ctl_rank_ba_3__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_rank_ba_4_;
  wire u_sdrc_core_u_bank_ctl_rank_ba_4__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_rank_ba_5_;
  wire u_sdrc_core_u_bank_ctl_rank_ba_5__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_rank_ba_6_;
  wire u_sdrc_core_u_bank_ctl_rank_ba_6__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_rank_ba_7_;
  wire u_sdrc_core_u_bank_ctl_rank_ba_7__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_rank_cnt_0_;
  wire u_sdrc_core_u_bank_ctl_rank_cnt_0__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_rank_cnt_1_;
  wire u_sdrc_core_u_bank_ctl_rank_cnt_1__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_rank_cnt_2_;
  wire u_sdrc_core_u_bank_ctl_rank_cnt_2__FF_INPUT;
  wire u_sdrc_core_u_bank_ctl_x2b_ack;
  wire u_sdrc_core_u_bank_ctl_x2b_ack_bF_buf0;
  wire u_sdrc_core_u_bank_ctl_x2b_ack_bF_buf1;
  wire u_sdrc_core_u_bank_ctl_x2b_ack_bF_buf2;
  wire u_sdrc_core_u_bank_ctl_x2b_ack_bF_buf3;
  wire u_sdrc_core_u_bank_ctl_xfr_bank_sel_0_;
  wire u_sdrc_core_u_bank_ctl_xfr_bank_sel_1_;
  wire u_sdrc_core_u_bs_convert__abc_21684_n168_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n169_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n170_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n170_1_bF_buf0;
  wire u_sdrc_core_u_bs_convert__abc_21684_n170_1_bF_buf1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n170_1_bF_buf2;
  wire u_sdrc_core_u_bs_convert__abc_21684_n170_1_bF_buf3;
  wire u_sdrc_core_u_bs_convert__abc_21684_n171_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n171_1_bF_buf0;
  wire u_sdrc_core_u_bs_convert__abc_21684_n171_1_bF_buf1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n171_1_bF_buf2;
  wire u_sdrc_core_u_bs_convert__abc_21684_n171_1_bF_buf3;
  wire u_sdrc_core_u_bs_convert__abc_21684_n172_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n173_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n174_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n175_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n176_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n177_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n178_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n179_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n180_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n181_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n182_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n183_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n184_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf0;
  wire u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf2;
  wire u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf3;
  wire u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf4;
  wire u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf5;
  wire u_sdrc_core_u_bs_convert__abc_21684_n185_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n186_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n187_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n188_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n189_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n190_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n191_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n192_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n193_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n194_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n195_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n196;
  wire u_sdrc_core_u_bs_convert__abc_21684_n197_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n199;
  wire u_sdrc_core_u_bs_convert__abc_21684_n200_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n201_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n202;
  wire u_sdrc_core_u_bs_convert__abc_21684_n203_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n204_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n205;
  wire u_sdrc_core_u_bs_convert__abc_21684_n206_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n207_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n208;
  wire u_sdrc_core_u_bs_convert__abc_21684_n209_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n210_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n211;
  wire u_sdrc_core_u_bs_convert__abc_21684_n212_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n213_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n214;
  wire u_sdrc_core_u_bs_convert__abc_21684_n215_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n217;
  wire u_sdrc_core_u_bs_convert__abc_21684_n218_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n219;
  wire u_sdrc_core_u_bs_convert__abc_21684_n220_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n221;
  wire u_sdrc_core_u_bs_convert__abc_21684_n222_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n223;
  wire u_sdrc_core_u_bs_convert__abc_21684_n224_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n225;
  wire u_sdrc_core_u_bs_convert__abc_21684_n226_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n227;
  wire u_sdrc_core_u_bs_convert__abc_21684_n228_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n229;
  wire u_sdrc_core_u_bs_convert__abc_21684_n230_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n231;
  wire u_sdrc_core_u_bs_convert__abc_21684_n233;
  wire u_sdrc_core_u_bs_convert__abc_21684_n234_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n235_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n236_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n237;
  wire u_sdrc_core_u_bs_convert__abc_21684_n238_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n239;
  wire u_sdrc_core_u_bs_convert__abc_21684_n240;
  wire u_sdrc_core_u_bs_convert__abc_21684_n241;
  wire u_sdrc_core_u_bs_convert__abc_21684_n242_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n243;
  wire u_sdrc_core_u_bs_convert__abc_21684_n244_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n245;
  wire u_sdrc_core_u_bs_convert__abc_21684_n246_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n247;
  wire u_sdrc_core_u_bs_convert__abc_21684_n249;
  wire u_sdrc_core_u_bs_convert__abc_21684_n250;
  wire u_sdrc_core_u_bs_convert__abc_21684_n251_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n252;
  wire u_sdrc_core_u_bs_convert__abc_21684_n253_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n254;
  wire u_sdrc_core_u_bs_convert__abc_21684_n255_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n256;
  wire u_sdrc_core_u_bs_convert__abc_21684_n257;
  wire u_sdrc_core_u_bs_convert__abc_21684_n258_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n259;
  wire u_sdrc_core_u_bs_convert__abc_21684_n260;
  wire u_sdrc_core_u_bs_convert__abc_21684_n261;
  wire u_sdrc_core_u_bs_convert__abc_21684_n262;
  wire u_sdrc_core_u_bs_convert__abc_21684_n263;
  wire u_sdrc_core_u_bs_convert__abc_21684_n264;
  wire u_sdrc_core_u_bs_convert__abc_21684_n265;
  wire u_sdrc_core_u_bs_convert__abc_21684_n266;
  wire u_sdrc_core_u_bs_convert__abc_21684_n268;
  wire u_sdrc_core_u_bs_convert__abc_21684_n269;
  wire u_sdrc_core_u_bs_convert__abc_21684_n270_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n271;
  wire u_sdrc_core_u_bs_convert__abc_21684_n272;
  wire u_sdrc_core_u_bs_convert__abc_21684_n273;
  wire u_sdrc_core_u_bs_convert__abc_21684_n274;
  wire u_sdrc_core_u_bs_convert__abc_21684_n275;
  wire u_sdrc_core_u_bs_convert__abc_21684_n276;
  wire u_sdrc_core_u_bs_convert__abc_21684_n277;
  wire u_sdrc_core_u_bs_convert__abc_21684_n278;
  wire u_sdrc_core_u_bs_convert__abc_21684_n279_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n280;
  wire u_sdrc_core_u_bs_convert__abc_21684_n281;
  wire u_sdrc_core_u_bs_convert__abc_21684_n282;
  wire u_sdrc_core_u_bs_convert__abc_21684_n283;
  wire u_sdrc_core_u_bs_convert__abc_21684_n284;
  wire u_sdrc_core_u_bs_convert__abc_21684_n285;
  wire u_sdrc_core_u_bs_convert__abc_21684_n287;
  wire u_sdrc_core_u_bs_convert__abc_21684_n288_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n289;
  wire u_sdrc_core_u_bs_convert__abc_21684_n290;
  wire u_sdrc_core_u_bs_convert__abc_21684_n291;
  wire u_sdrc_core_u_bs_convert__abc_21684_n292;
  wire u_sdrc_core_u_bs_convert__abc_21684_n293;
  wire u_sdrc_core_u_bs_convert__abc_21684_n294;
  wire u_sdrc_core_u_bs_convert__abc_21684_n295;
  wire u_sdrc_core_u_bs_convert__abc_21684_n296;
  wire u_sdrc_core_u_bs_convert__abc_21684_n297_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n298;
  wire u_sdrc_core_u_bs_convert__abc_21684_n299;
  wire u_sdrc_core_u_bs_convert__abc_21684_n300;
  wire u_sdrc_core_u_bs_convert__abc_21684_n301;
  wire u_sdrc_core_u_bs_convert__abc_21684_n303;
  wire u_sdrc_core_u_bs_convert__abc_21684_n304;
  wire u_sdrc_core_u_bs_convert__abc_21684_n305;
  wire u_sdrc_core_u_bs_convert__abc_21684_n306_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n307;
  wire u_sdrc_core_u_bs_convert__abc_21684_n308;
  wire u_sdrc_core_u_bs_convert__abc_21684_n309;
  wire u_sdrc_core_u_bs_convert__abc_21684_n310;
  wire u_sdrc_core_u_bs_convert__abc_21684_n311;
  wire u_sdrc_core_u_bs_convert__abc_21684_n312;
  wire u_sdrc_core_u_bs_convert__abc_21684_n313;
  wire u_sdrc_core_u_bs_convert__abc_21684_n314;
  wire u_sdrc_core_u_bs_convert__abc_21684_n315_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n316;
  wire u_sdrc_core_u_bs_convert__abc_21684_n317;
  wire u_sdrc_core_u_bs_convert__abc_21684_n318;
  wire u_sdrc_core_u_bs_convert__abc_21684_n319;
  wire u_sdrc_core_u_bs_convert__abc_21684_n320;
  wire u_sdrc_core_u_bs_convert__abc_21684_n322;
  wire u_sdrc_core_u_bs_convert__abc_21684_n323;
  wire u_sdrc_core_u_bs_convert__abc_21684_n324_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n326;
  wire u_sdrc_core_u_bs_convert__abc_21684_n327;
  wire u_sdrc_core_u_bs_convert__abc_21684_n328;
  wire u_sdrc_core_u_bs_convert__abc_21684_n330;
  wire u_sdrc_core_u_bs_convert__abc_21684_n331;
  wire u_sdrc_core_u_bs_convert__abc_21684_n332;
  wire u_sdrc_core_u_bs_convert__abc_21684_n334;
  wire u_sdrc_core_u_bs_convert__abc_21684_n335;
  wire u_sdrc_core_u_bs_convert__abc_21684_n336;
  wire u_sdrc_core_u_bs_convert__abc_21684_n338;
  wire u_sdrc_core_u_bs_convert__abc_21684_n339;
  wire u_sdrc_core_u_bs_convert__abc_21684_n340;
  wire u_sdrc_core_u_bs_convert__abc_21684_n342;
  wire u_sdrc_core_u_bs_convert__abc_21684_n343;
  wire u_sdrc_core_u_bs_convert__abc_21684_n344;
  wire u_sdrc_core_u_bs_convert__abc_21684_n346;
  wire u_sdrc_core_u_bs_convert__abc_21684_n347;
  wire u_sdrc_core_u_bs_convert__abc_21684_n348;
  wire u_sdrc_core_u_bs_convert__abc_21684_n350;
  wire u_sdrc_core_u_bs_convert__abc_21684_n351;
  wire u_sdrc_core_u_bs_convert__abc_21684_n352;
  wire u_sdrc_core_u_bs_convert__abc_21684_n354;
  wire u_sdrc_core_u_bs_convert__abc_21684_n355;
  wire u_sdrc_core_u_bs_convert__abc_21684_n356;
  wire u_sdrc_core_u_bs_convert__abc_21684_n357_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n358;
  wire u_sdrc_core_u_bs_convert__abc_21684_n359;
  wire u_sdrc_core_u_bs_convert__abc_21684_n360;
  wire u_sdrc_core_u_bs_convert__abc_21684_n361_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n362;
  wire u_sdrc_core_u_bs_convert__abc_21684_n363;
  wire u_sdrc_core_u_bs_convert__abc_21684_n364;
  wire u_sdrc_core_u_bs_convert__abc_21684_n365_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n366;
  wire u_sdrc_core_u_bs_convert__abc_21684_n367;
  wire u_sdrc_core_u_bs_convert__abc_21684_n368;
  wire u_sdrc_core_u_bs_convert__abc_21684_n369;
  wire u_sdrc_core_u_bs_convert__abc_21684_n370;
  wire u_sdrc_core_u_bs_convert__abc_21684_n371_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n373;
  wire u_sdrc_core_u_bs_convert__abc_21684_n374;
  wire u_sdrc_core_u_bs_convert__abc_21684_n375;
  wire u_sdrc_core_u_bs_convert__abc_21684_n377;
  wire u_sdrc_core_u_bs_convert__abc_21684_n378;
  wire u_sdrc_core_u_bs_convert__abc_21684_n379;
  wire u_sdrc_core_u_bs_convert__abc_21684_n381_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n382;
  wire u_sdrc_core_u_bs_convert__abc_21684_n384;
  wire u_sdrc_core_u_bs_convert__abc_21684_n385;
  wire u_sdrc_core_u_bs_convert__abc_21684_n387;
  wire u_sdrc_core_u_bs_convert__abc_21684_n388;
  wire u_sdrc_core_u_bs_convert__abc_21684_n390;
  wire u_sdrc_core_u_bs_convert__abc_21684_n391_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n393;
  wire u_sdrc_core_u_bs_convert__abc_21684_n394;
  wire u_sdrc_core_u_bs_convert__abc_21684_n396_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n397;
  wire u_sdrc_core_u_bs_convert__abc_21684_n399;
  wire u_sdrc_core_u_bs_convert__abc_21684_n400;
  wire u_sdrc_core_u_bs_convert__abc_21684_n402;
  wire u_sdrc_core_u_bs_convert__abc_21684_n403;
  wire u_sdrc_core_u_bs_convert__abc_21684_n405;
  wire u_sdrc_core_u_bs_convert__abc_21684_n406_1;
  wire u_sdrc_core_u_bs_convert__abc_21684_n408;
  wire u_sdrc_core_u_bs_convert__abc_21684_n409;
  wire u_sdrc_core_u_bs_convert__abc_21684_n411;
  wire u_sdrc_core_u_bs_convert__abc_21684_n412;
  wire u_sdrc_core_u_bs_convert__abc_21684_n414;
  wire u_sdrc_core_u_bs_convert__abc_21684_n415;
  wire u_sdrc_core_u_bs_convert__abc_21684_n417;
  wire u_sdrc_core_u_bs_convert__abc_21684_n418;
  wire u_sdrc_core_u_bs_convert__abc_21684_n420;
  wire u_sdrc_core_u_bs_convert__abc_21684_n421;
  wire u_sdrc_core_u_bs_convert__abc_21684_n423;
  wire u_sdrc_core_u_bs_convert__abc_21684_n424;
  wire u_sdrc_core_u_bs_convert__abc_21684_n426;
  wire u_sdrc_core_u_bs_convert__abc_21684_n427;
  wire u_sdrc_core_u_bs_convert__abc_21684_n429;
  wire u_sdrc_core_u_bs_convert__abc_21684_n430;
  wire u_sdrc_core_u_bs_convert__abc_21684_n432;
  wire u_sdrc_core_u_bs_convert__abc_21684_n433;
  wire u_sdrc_core_u_bs_convert__abc_21684_n435;
  wire u_sdrc_core_u_bs_convert__abc_21684_n436;
  wire u_sdrc_core_u_bs_convert__abc_21684_n438;
  wire u_sdrc_core_u_bs_convert__abc_21684_n439;
  wire u_sdrc_core_u_bs_convert__abc_21684_n441;
  wire u_sdrc_core_u_bs_convert__abc_21684_n442;
  wire u_sdrc_core_u_bs_convert__abc_21684_n444;
  wire u_sdrc_core_u_bs_convert__abc_21684_n445;
  wire u_sdrc_core_u_bs_convert__abc_21684_n447;
  wire u_sdrc_core_u_bs_convert__abc_21684_n448;
  wire u_sdrc_core_u_bs_convert__abc_21684_n450;
  wire u_sdrc_core_u_bs_convert__abc_21684_n451;
  wire u_sdrc_core_u_bs_convert__abc_21684_n453;
  wire u_sdrc_core_u_bs_convert__abc_21684_n454;
  wire u_sdrc_core_u_bs_convert__abc_21684_n456;
  wire u_sdrc_core_u_bs_convert__abc_21684_n457;
  wire u_sdrc_core_u_bs_convert__abc_21684_n459;
  wire u_sdrc_core_u_bs_convert__abc_21684_n460;
  wire u_sdrc_core_u_bs_convert__abc_21684_n462;
  wire u_sdrc_core_u_bs_convert__abc_21684_n463;
  wire u_sdrc_core_u_bs_convert__abc_21684_n465;
  wire u_sdrc_core_u_bs_convert__abc_21684_n466;
  wire u_sdrc_core_u_bs_convert__abc_21684_n468;
  wire u_sdrc_core_u_bs_convert__abc_21684_n469;
  wire u_sdrc_core_u_bs_convert__abc_21684_n471;
  wire u_sdrc_core_u_bs_convert__abc_21684_n472;
  wire u_sdrc_core_u_bs_convert__abc_21684_n474;
  wire u_sdrc_core_u_bs_convert__abc_21684_n475;
  wire u_sdrc_core_u_bs_convert__abc_21684_n477;
  wire u_sdrc_core_u_bs_convert__abc_21684_n478;
  wire u_sdrc_core_u_bs_convert__abc_21684_n479;
  wire u_sdrc_core_u_bs_convert__abc_21684_n481;
  wire u_sdrc_core_u_bs_convert__abc_21684_n482;
  wire u_sdrc_core_u_bs_convert__abc_21684_n483;
  wire u_sdrc_core_u_bs_convert__abc_21684_n484;
  wire u_sdrc_core_u_bs_convert__abc_21684_n485;
  wire u_sdrc_core_u_bs_convert__abc_21684_n486;
  wire u_sdrc_core_u_bs_convert__abc_21684_n488;
  wire u_sdrc_core_u_bs_convert__abc_21684_n489;
  wire u_sdrc_core_u_bs_convert__abc_21684_n490;
  wire u_sdrc_core_u_bs_convert__abc_21684_n491;
  wire u_sdrc_core_u_bs_convert__abc_21684_n493;
  wire u_sdrc_core_u_bs_convert__abc_21684_n494;
  wire u_sdrc_core_u_bs_convert__abc_21684_n495;
  wire u_sdrc_core_u_bs_convert__abc_21684_n496;
  wire u_sdrc_core_u_bs_convert__abc_21684_n497;
  wire u_sdrc_core_u_bs_convert__abc_21684_n498;
  wire u_sdrc_core_u_bs_convert__abc_21684_n500;
  wire u_sdrc_core_u_bs_convert__abc_21684_n501;
  wire u_sdrc_core_u_bs_convert__abc_21684_n502;
  wire u_sdrc_core_u_bs_convert__abc_21684_n503;
  wire u_sdrc_core_u_bs_convert__abc_21684_n505;
  wire u_sdrc_core_u_bs_convert__abc_21684_n506;
  wire u_sdrc_core_u_bs_convert__abc_21684_n507;
  wire u_sdrc_core_u_bs_convert__abc_21684_n508;
  wire u_sdrc_core_u_bs_convert__abc_21684_n509;
  wire u_sdrc_core_u_bs_convert__abc_21684_n510;
  wire u_sdrc_core_u_bs_convert__abc_21684_n511;
  wire u_sdrc_core_u_bs_convert__abc_21684_n512;
  wire u_sdrc_core_u_bs_convert__abc_21684_n514;
  wire u_sdrc_core_u_bs_convert__abc_21684_n515;
  wire u_sdrc_core_u_bs_convert__abc_21684_n516;
  wire u_sdrc_core_u_bs_convert__abc_21684_n518;
  wire u_sdrc_core_u_bs_convert__abc_21684_n519;
  wire u_sdrc_core_u_bs_convert__abc_21684_n520;
  wire u_sdrc_core_u_bs_convert__abc_21684_n522;
  wire u_sdrc_core_u_bs_convert__abc_21684_n523;
  wire u_sdrc_core_u_bs_convert__abc_21684_n524;
  wire u_sdrc_core_u_bs_convert__abc_21684_n526;
  wire u_sdrc_core_u_bs_convert__abc_21684_n527;
  wire u_sdrc_core_u_bs_convert__abc_21684_n528;
  wire u_sdrc_core_u_bs_convert__abc_21684_n530;
  wire u_sdrc_core_u_bs_convert__abc_21684_n531;
  wire u_sdrc_core_u_bs_convert__abc_21684_n532;
  wire u_sdrc_core_u_bs_convert__abc_21684_n534;
  wire u_sdrc_core_u_bs_convert__abc_21684_n535;
  wire u_sdrc_core_u_bs_convert__abc_21684_n536;
  wire u_sdrc_core_u_bs_convert__abc_21684_n538;
  wire u_sdrc_core_u_bs_convert__abc_21684_n539;
  wire u_sdrc_core_u_bs_convert__abc_21684_n540;
  wire u_sdrc_core_u_bs_convert__abc_21684_n542;
  wire u_sdrc_core_u_bs_convert__abc_21684_n543;
  wire u_sdrc_core_u_bs_convert__abc_21684_n544;
  wire u_sdrc_core_u_bs_convert__abc_21684_n545;
  wire u_sdrc_core_u_bs_convert__abc_21684_n546;
  wire u_sdrc_core_u_bs_convert__abc_21684_n547;
  wire u_sdrc_core_u_bs_convert__abc_21684_n548;
  wire u_sdrc_core_u_bs_convert__abc_21684_n549;
  wire u_sdrc_core_u_bs_convert__abc_21684_n551;
  wire u_sdrc_core_u_bs_convert__abc_21684_n552;
  wire u_sdrc_core_u_bs_convert__abc_21684_n553;
  wire u_sdrc_core_u_bs_convert__abc_21684_n555;
  wire u_sdrc_core_u_bs_convert__abc_21684_n556;
  wire u_sdrc_core_u_bs_convert__abc_21684_n557;
  wire u_sdrc_core_u_bs_convert__abc_21684_n559;
  wire u_sdrc_core_u_bs_convert__abc_21684_n560;
  wire u_sdrc_core_u_bs_convert__abc_21684_n561;
  wire u_sdrc_core_u_bs_convert__abc_21684_n563;
  wire u_sdrc_core_u_bs_convert__abc_21684_n564;
  wire u_sdrc_core_u_bs_convert__abc_21684_n565;
  wire u_sdrc_core_u_bs_convert__abc_21684_n567;
  wire u_sdrc_core_u_bs_convert__abc_21684_n568;
  wire u_sdrc_core_u_bs_convert__abc_21684_n569;
  wire u_sdrc_core_u_bs_convert__abc_21684_n571;
  wire u_sdrc_core_u_bs_convert__abc_21684_n572;
  wire u_sdrc_core_u_bs_convert__abc_21684_n573;
  wire u_sdrc_core_u_bs_convert__abc_21684_n575;
  wire u_sdrc_core_u_bs_convert__abc_21684_n576;
  wire u_sdrc_core_u_bs_convert__abc_21684_n577;
  wire u_sdrc_core_u_bs_convert__abc_21684_n579;
  wire u_sdrc_core_u_bs_convert__abc_21684_n580;
  wire u_sdrc_core_u_bs_convert__abc_21684_n581;
  wire u_sdrc_core_u_bs_convert__abc_21684_n582;
  wire u_sdrc_core_u_bs_convert__abc_21684_n583;
  wire u_sdrc_core_u_bs_convert__abc_21684_n584;
  wire u_sdrc_core_u_bs_convert__abc_21684_n585;
  wire u_sdrc_core_u_bs_convert__abc_21684_n586;
  wire u_sdrc_core_u_bs_convert__abc_21684_n587;
  wire u_sdrc_core_u_bs_convert__abc_21684_n588;
  wire u_sdrc_core_u_bs_convert__abc_21684_n590;
  wire u_sdrc_core_u_bs_convert__abc_21684_n591;
  wire u_sdrc_core_u_bs_convert__abc_21684_n592;
  wire u_sdrc_core_u_bs_convert__abc_21684_n593;
  wire u_sdrc_core_u_bs_convert__abc_21684_n594;
  wire u_sdrc_core_u_bs_convert__abc_21684_n595;
  wire u_sdrc_core_u_bs_convert__abc_21684_n596;
  wire u_sdrc_core_u_bs_convert__abc_21684_n597;
  wire u_sdrc_core_u_bs_convert__abc_21684_n599;
  wire u_sdrc_core_u_bs_convert__abc_21684_n600;
  wire u_sdrc_core_u_bs_convert__abc_21684_n601;
  wire u_sdrc_core_u_bs_convert__abc_21684_n602;
  wire u_sdrc_core_u_bs_convert__abc_21684_n603;
  wire u_sdrc_core_u_bs_convert__abc_21684_n604;
  wire u_sdrc_core_u_bs_convert__abc_21684_n605;
  wire u_sdrc_core_u_bs_convert__abc_21684_n606;
  wire u_sdrc_core_u_bs_convert__abc_21684_n608;
  wire u_sdrc_core_u_bs_convert__abc_21684_n609;
  wire u_sdrc_core_u_bs_convert__abc_21684_n610;
  wire u_sdrc_core_u_bs_convert__abc_21684_n611;
  wire u_sdrc_core_u_bs_convert__abc_21684_n612;
  wire u_sdrc_core_u_bs_convert__abc_21684_n613;
  wire u_sdrc_core_u_bs_convert__abc_21684_n614;
  wire u_sdrc_core_u_bs_convert__abc_21684_n615;
  wire u_sdrc_core_u_bs_convert__abc_21684_n617;
  wire u_sdrc_core_u_bs_convert__abc_21684_n618;
  wire u_sdrc_core_u_bs_convert__abc_21684_n619;
  wire u_sdrc_core_u_bs_convert__abc_21684_n620;
  wire u_sdrc_core_u_bs_convert__abc_21684_n621;
  wire u_sdrc_core_u_bs_convert__abc_21684_n622;
  wire u_sdrc_core_u_bs_convert__abc_21684_n623;
  wire u_sdrc_core_u_bs_convert__abc_21684_n624;
  wire u_sdrc_core_u_bs_convert__abc_21684_n626;
  wire u_sdrc_core_u_bs_convert__abc_21684_n627;
  wire u_sdrc_core_u_bs_convert__abc_21684_n628;
  wire u_sdrc_core_u_bs_convert__abc_21684_n629;
  wire u_sdrc_core_u_bs_convert__abc_21684_n630;
  wire u_sdrc_core_u_bs_convert__abc_21684_n631;
  wire u_sdrc_core_u_bs_convert__abc_21684_n632;
  wire u_sdrc_core_u_bs_convert__abc_21684_n633;
  wire u_sdrc_core_u_bs_convert__abc_21684_n635;
  wire u_sdrc_core_u_bs_convert__abc_21684_n636;
  wire u_sdrc_core_u_bs_convert__abc_21684_n637;
  wire u_sdrc_core_u_bs_convert__abc_21684_n638;
  wire u_sdrc_core_u_bs_convert__abc_21684_n639;
  wire u_sdrc_core_u_bs_convert__abc_21684_n640;
  wire u_sdrc_core_u_bs_convert__abc_21684_n641;
  wire u_sdrc_core_u_bs_convert__abc_21684_n642;
  wire u_sdrc_core_u_bs_convert__abc_21684_n644;
  wire u_sdrc_core_u_bs_convert__abc_21684_n645;
  wire u_sdrc_core_u_bs_convert__abc_21684_n646;
  wire u_sdrc_core_u_bs_convert__abc_21684_n647;
  wire u_sdrc_core_u_bs_convert__abc_21684_n648;
  wire u_sdrc_core_u_bs_convert__abc_21684_n649;
  wire u_sdrc_core_u_bs_convert__abc_21684_n650;
  wire u_sdrc_core_u_bs_convert__abc_21684_n651;
  wire u_sdrc_core_u_bs_convert_rd_xfr_count_0_;
  wire u_sdrc_core_u_bs_convert_rd_xfr_count_0__FF_INPUT;
  wire u_sdrc_core_u_bs_convert_rd_xfr_count_1_;
  wire u_sdrc_core_u_bs_convert_rd_xfr_count_1__FF_INPUT;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_0_;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_0__FF_INPUT;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_10_;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_10__FF_INPUT;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_11_;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_11__FF_INPUT;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_12_;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_12__FF_INPUT;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_13_;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_13__FF_INPUT;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_14_;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_14__FF_INPUT;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_15_;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_15__FF_INPUT;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_16_;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_16__FF_INPUT;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_17_;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_17__FF_INPUT;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_18_;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_18__FF_INPUT;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_19_;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_19__FF_INPUT;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_1_;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_1__FF_INPUT;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_20_;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_20__FF_INPUT;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_21_;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_21__FF_INPUT;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_22_;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_22__FF_INPUT;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_23_;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_23__FF_INPUT;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_2_;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_2__FF_INPUT;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_3_;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_3__FF_INPUT;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_4_;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_4__FF_INPUT;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_5_;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_5__FF_INPUT;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_6_;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_6__FF_INPUT;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_7_;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_7__FF_INPUT;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_8_;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_8__FF_INPUT;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_9_;
  wire u_sdrc_core_u_bs_convert_saved_rd_data_9__FF_INPUT;
  wire u_sdrc_core_u_bs_convert_wr_xfr_count_0_;
  wire u_sdrc_core_u_bs_convert_wr_xfr_count_0__FF_INPUT;
  wire u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf0;
  wire u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf1;
  wire u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf2;
  wire u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf3;
  wire u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf4;
  wire u_sdrc_core_u_bs_convert_wr_xfr_count_1_;
  wire u_sdrc_core_u_bs_convert_wr_xfr_count_1__FF_INPUT;
  wire u_sdrc_core_u_bs_convert_x2a_rdok;
  wire u_sdrc_core_u_bs_convert_x2a_wrnext;
  wire u_sdrc_core_u_bs_convert_x2a_wrnext_bF_buf0;
  wire u_sdrc_core_u_bs_convert_x2a_wrnext_bF_buf1;
  wire u_sdrc_core_u_bs_convert_x2a_wrnext_bF_buf2;
  wire u_sdrc_core_u_bs_convert_x2a_wrnext_bF_buf3;
  wire u_sdrc_core_u_req_gen__abc_16238_n30;
  wire u_sdrc_core_u_req_gen__abc_16238_n38;
  wire u_sdrc_core_u_req_gen__abc_16238_n57;
  wire u_sdrc_core_u_req_gen__abc_22171_n1000;
  wire u_sdrc_core_u_req_gen__abc_22171_n1001;
  wire u_sdrc_core_u_req_gen__abc_22171_n1002;
  wire u_sdrc_core_u_req_gen__abc_22171_n1003;
  wire u_sdrc_core_u_req_gen__abc_22171_n1005;
  wire u_sdrc_core_u_req_gen__abc_22171_n1007;
  wire u_sdrc_core_u_req_gen__abc_22171_n1009;
  wire u_sdrc_core_u_req_gen__abc_22171_n1010;
  wire u_sdrc_core_u_req_gen__abc_22171_n1011;
  wire u_sdrc_core_u_req_gen__abc_22171_n1012;
  wire u_sdrc_core_u_req_gen__abc_22171_n1013;
  wire u_sdrc_core_u_req_gen__abc_22171_n1014;
  wire u_sdrc_core_u_req_gen__abc_22171_n1015;
  wire u_sdrc_core_u_req_gen__abc_22171_n1016;
  wire u_sdrc_core_u_req_gen__abc_22171_n1017;
  wire u_sdrc_core_u_req_gen__abc_22171_n1018;
  wire u_sdrc_core_u_req_gen__abc_22171_n1019;
  wire u_sdrc_core_u_req_gen__abc_22171_n1020;
  wire u_sdrc_core_u_req_gen__abc_22171_n1021;
  wire u_sdrc_core_u_req_gen__abc_22171_n1022;
  wire u_sdrc_core_u_req_gen__abc_22171_n1023;
  wire u_sdrc_core_u_req_gen__abc_22171_n1024;
  wire u_sdrc_core_u_req_gen__abc_22171_n1025;
  wire u_sdrc_core_u_req_gen__abc_22171_n1026;
  wire u_sdrc_core_u_req_gen__abc_22171_n1027;
  wire u_sdrc_core_u_req_gen__abc_22171_n1028;
  wire u_sdrc_core_u_req_gen__abc_22171_n1029;
  wire u_sdrc_core_u_req_gen__abc_22171_n1030;
  wire u_sdrc_core_u_req_gen__abc_22171_n1031;
  wire u_sdrc_core_u_req_gen__abc_22171_n1032;
  wire u_sdrc_core_u_req_gen__abc_22171_n1033;
  wire u_sdrc_core_u_req_gen__abc_22171_n1034;
  wire u_sdrc_core_u_req_gen__abc_22171_n1035;
  wire u_sdrc_core_u_req_gen__abc_22171_n1036;
  wire u_sdrc_core_u_req_gen__abc_22171_n1037;
  wire u_sdrc_core_u_req_gen__abc_22171_n1038;
  wire u_sdrc_core_u_req_gen__abc_22171_n1039;
  wire u_sdrc_core_u_req_gen__abc_22171_n1040;
  wire u_sdrc_core_u_req_gen__abc_22171_n1041;
  wire u_sdrc_core_u_req_gen__abc_22171_n1042;
  wire u_sdrc_core_u_req_gen__abc_22171_n1043;
  wire u_sdrc_core_u_req_gen__abc_22171_n1044;
  wire u_sdrc_core_u_req_gen__abc_22171_n1045;
  wire u_sdrc_core_u_req_gen__abc_22171_n1046;
  wire u_sdrc_core_u_req_gen__abc_22171_n1047;
  wire u_sdrc_core_u_req_gen__abc_22171_n1048;
  wire u_sdrc_core_u_req_gen__abc_22171_n1049;
  wire u_sdrc_core_u_req_gen__abc_22171_n1050;
  wire u_sdrc_core_u_req_gen__abc_22171_n1051;
  wire u_sdrc_core_u_req_gen__abc_22171_n1052;
  wire u_sdrc_core_u_req_gen__abc_22171_n1053;
  wire u_sdrc_core_u_req_gen__abc_22171_n1054;
  wire u_sdrc_core_u_req_gen__abc_22171_n1055;
  wire u_sdrc_core_u_req_gen__abc_22171_n1056;
  wire u_sdrc_core_u_req_gen__abc_22171_n1057;
  wire u_sdrc_core_u_req_gen__abc_22171_n1058;
  wire u_sdrc_core_u_req_gen__abc_22171_n1059;
  wire u_sdrc_core_u_req_gen__abc_22171_n1060;
  wire u_sdrc_core_u_req_gen__abc_22171_n1061;
  wire u_sdrc_core_u_req_gen__abc_22171_n1062;
  wire u_sdrc_core_u_req_gen__abc_22171_n1063;
  wire u_sdrc_core_u_req_gen__abc_22171_n1064;
  wire u_sdrc_core_u_req_gen__abc_22171_n1065;
  wire u_sdrc_core_u_req_gen__abc_22171_n1066;
  wire u_sdrc_core_u_req_gen__abc_22171_n1067;
  wire u_sdrc_core_u_req_gen__abc_22171_n1068;
  wire u_sdrc_core_u_req_gen__abc_22171_n1069;
  wire u_sdrc_core_u_req_gen__abc_22171_n1070;
  wire u_sdrc_core_u_req_gen__abc_22171_n1071;
  wire u_sdrc_core_u_req_gen__abc_22171_n1072;
  wire u_sdrc_core_u_req_gen__abc_22171_n1073;
  wire u_sdrc_core_u_req_gen__abc_22171_n1074;
  wire u_sdrc_core_u_req_gen__abc_22171_n1075;
  wire u_sdrc_core_u_req_gen__abc_22171_n1076;
  wire u_sdrc_core_u_req_gen__abc_22171_n1077;
  wire u_sdrc_core_u_req_gen__abc_22171_n1078;
  wire u_sdrc_core_u_req_gen__abc_22171_n1079;
  wire u_sdrc_core_u_req_gen__abc_22171_n1080;
  wire u_sdrc_core_u_req_gen__abc_22171_n1081;
  wire u_sdrc_core_u_req_gen__abc_22171_n1082;
  wire u_sdrc_core_u_req_gen__abc_22171_n1083;
  wire u_sdrc_core_u_req_gen__abc_22171_n1084;
  wire u_sdrc_core_u_req_gen__abc_22171_n1085;
  wire u_sdrc_core_u_req_gen__abc_22171_n1086;
  wire u_sdrc_core_u_req_gen__abc_22171_n1087;
  wire u_sdrc_core_u_req_gen__abc_22171_n1088;
  wire u_sdrc_core_u_req_gen__abc_22171_n1089;
  wire u_sdrc_core_u_req_gen__abc_22171_n1090;
  wire u_sdrc_core_u_req_gen__abc_22171_n1091;
  wire u_sdrc_core_u_req_gen__abc_22171_n1092;
  wire u_sdrc_core_u_req_gen__abc_22171_n1093;
  wire u_sdrc_core_u_req_gen__abc_22171_n1094;
  wire u_sdrc_core_u_req_gen__abc_22171_n1095;
  wire u_sdrc_core_u_req_gen__abc_22171_n1096;
  wire u_sdrc_core_u_req_gen__abc_22171_n1097;
  wire u_sdrc_core_u_req_gen__abc_22171_n1098;
  wire u_sdrc_core_u_req_gen__abc_22171_n1099;
  wire u_sdrc_core_u_req_gen__abc_22171_n1100;
  wire u_sdrc_core_u_req_gen__abc_22171_n1101;
  wire u_sdrc_core_u_req_gen__abc_22171_n1102;
  wire u_sdrc_core_u_req_gen__abc_22171_n1103;
  wire u_sdrc_core_u_req_gen__abc_22171_n1105;
  wire u_sdrc_core_u_req_gen__abc_22171_n181;
  wire u_sdrc_core_u_req_gen__abc_22171_n182_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n183;
  wire u_sdrc_core_u_req_gen__abc_22171_n184;
  wire u_sdrc_core_u_req_gen__abc_22171_n185;
  wire u_sdrc_core_u_req_gen__abc_22171_n186;
  wire u_sdrc_core_u_req_gen__abc_22171_n188;
  wire u_sdrc_core_u_req_gen__abc_22171_n189;
  wire u_sdrc_core_u_req_gen__abc_22171_n190;
  wire u_sdrc_core_u_req_gen__abc_22171_n191;
  wire u_sdrc_core_u_req_gen__abc_22171_n193;
  wire u_sdrc_core_u_req_gen__abc_22171_n194;
  wire u_sdrc_core_u_req_gen__abc_22171_n195_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n196;
  wire u_sdrc_core_u_req_gen__abc_22171_n197;
  wire u_sdrc_core_u_req_gen__abc_22171_n198;
  wire u_sdrc_core_u_req_gen__abc_22171_n199;
  wire u_sdrc_core_u_req_gen__abc_22171_n200_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n202;
  wire u_sdrc_core_u_req_gen__abc_22171_n203;
  wire u_sdrc_core_u_req_gen__abc_22171_n204;
  wire u_sdrc_core_u_req_gen__abc_22171_n205;
  wire u_sdrc_core_u_req_gen__abc_22171_n207;
  wire u_sdrc_core_u_req_gen__abc_22171_n208;
  wire u_sdrc_core_u_req_gen__abc_22171_n209;
  wire u_sdrc_core_u_req_gen__abc_22171_n210_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n212;
  wire u_sdrc_core_u_req_gen__abc_22171_n213;
  wire u_sdrc_core_u_req_gen__abc_22171_n214;
  wire u_sdrc_core_u_req_gen__abc_22171_n215_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n216_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n218;
  wire u_sdrc_core_u_req_gen__abc_22171_n219_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n220;
  wire u_sdrc_core_u_req_gen__abc_22171_n221_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n222;
  wire u_sdrc_core_u_req_gen__abc_22171_n224;
  wire u_sdrc_core_u_req_gen__abc_22171_n225;
  wire u_sdrc_core_u_req_gen__abc_22171_n226_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n227;
  wire u_sdrc_core_u_req_gen__abc_22171_n229;
  wire u_sdrc_core_u_req_gen__abc_22171_n230;
  wire u_sdrc_core_u_req_gen__abc_22171_n231;
  wire u_sdrc_core_u_req_gen__abc_22171_n232;
  wire u_sdrc_core_u_req_gen__abc_22171_n234_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n235;
  wire u_sdrc_core_u_req_gen__abc_22171_n236_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n237;
  wire u_sdrc_core_u_req_gen__abc_22171_n240;
  wire u_sdrc_core_u_req_gen__abc_22171_n241;
  wire u_sdrc_core_u_req_gen__abc_22171_n242;
  wire u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf0;
  wire u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf1;
  wire u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf2;
  wire u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf3;
  wire u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf4;
  wire u_sdrc_core_u_req_gen__abc_22171_n243_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n245_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf0;
  wire u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf1;
  wire u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf2;
  wire u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf3;
  wire u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf4;
  wire u_sdrc_core_u_req_gen__abc_22171_n246;
  wire u_sdrc_core_u_req_gen__abc_22171_n247;
  wire u_sdrc_core_u_req_gen__abc_22171_n248;
  wire u_sdrc_core_u_req_gen__abc_22171_n249;
  wire u_sdrc_core_u_req_gen__abc_22171_n250;
  wire u_sdrc_core_u_req_gen__abc_22171_n251;
  wire u_sdrc_core_u_req_gen__abc_22171_n252;
  wire u_sdrc_core_u_req_gen__abc_22171_n253;
  wire u_sdrc_core_u_req_gen__abc_22171_n255;
  wire u_sdrc_core_u_req_gen__abc_22171_n256_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n257;
  wire u_sdrc_core_u_req_gen__abc_22171_n258;
  wire u_sdrc_core_u_req_gen__abc_22171_n259;
  wire u_sdrc_core_u_req_gen__abc_22171_n260;
  wire u_sdrc_core_u_req_gen__abc_22171_n261;
  wire u_sdrc_core_u_req_gen__abc_22171_n262_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n263_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n264;
  wire u_sdrc_core_u_req_gen__abc_22171_n265;
  wire u_sdrc_core_u_req_gen__abc_22171_n266;
  wire u_sdrc_core_u_req_gen__abc_22171_n267;
  wire u_sdrc_core_u_req_gen__abc_22171_n269;
  wire u_sdrc_core_u_req_gen__abc_22171_n270;
  wire u_sdrc_core_u_req_gen__abc_22171_n271;
  wire u_sdrc_core_u_req_gen__abc_22171_n272;
  wire u_sdrc_core_u_req_gen__abc_22171_n273_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n274;
  wire u_sdrc_core_u_req_gen__abc_22171_n275;
  wire u_sdrc_core_u_req_gen__abc_22171_n276;
  wire u_sdrc_core_u_req_gen__abc_22171_n277_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n278;
  wire u_sdrc_core_u_req_gen__abc_22171_n280;
  wire u_sdrc_core_u_req_gen__abc_22171_n281_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n282;
  wire u_sdrc_core_u_req_gen__abc_22171_n283_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n284;
  wire u_sdrc_core_u_req_gen__abc_22171_n285;
  wire u_sdrc_core_u_req_gen__abc_22171_n286;
  wire u_sdrc_core_u_req_gen__abc_22171_n287;
  wire u_sdrc_core_u_req_gen__abc_22171_n288;
  wire u_sdrc_core_u_req_gen__abc_22171_n289;
  wire u_sdrc_core_u_req_gen__abc_22171_n290_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n292;
  wire u_sdrc_core_u_req_gen__abc_22171_n293;
  wire u_sdrc_core_u_req_gen__abc_22171_n294_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n295;
  wire u_sdrc_core_u_req_gen__abc_22171_n296_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n297;
  wire u_sdrc_core_u_req_gen__abc_22171_n298_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n299;
  wire u_sdrc_core_u_req_gen__abc_22171_n300;
  wire u_sdrc_core_u_req_gen__abc_22171_n301;
  wire u_sdrc_core_u_req_gen__abc_22171_n303;
  wire u_sdrc_core_u_req_gen__abc_22171_n304_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n305;
  wire u_sdrc_core_u_req_gen__abc_22171_n306;
  wire u_sdrc_core_u_req_gen__abc_22171_n307_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n308;
  wire u_sdrc_core_u_req_gen__abc_22171_n309;
  wire u_sdrc_core_u_req_gen__abc_22171_n310_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n311;
  wire u_sdrc_core_u_req_gen__abc_22171_n312;
  wire u_sdrc_core_u_req_gen__abc_22171_n314;
  wire u_sdrc_core_u_req_gen__abc_22171_n315;
  wire u_sdrc_core_u_req_gen__abc_22171_n316;
  wire u_sdrc_core_u_req_gen__abc_22171_n318;
  wire u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf0;
  wire u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf1;
  wire u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf2;
  wire u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf3;
  wire u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf4;
  wire u_sdrc_core_u_req_gen__abc_22171_n331;
  wire u_sdrc_core_u_req_gen__abc_22171_n332;
  wire u_sdrc_core_u_req_gen__abc_22171_n335_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n335_1_bF_buf0;
  wire u_sdrc_core_u_req_gen__abc_22171_n335_1_bF_buf1;
  wire u_sdrc_core_u_req_gen__abc_22171_n335_1_bF_buf2;
  wire u_sdrc_core_u_req_gen__abc_22171_n335_1_bF_buf3;
  wire u_sdrc_core_u_req_gen__abc_22171_n336;
  wire u_sdrc_core_u_req_gen__abc_22171_n337_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n338;
  wire u_sdrc_core_u_req_gen__abc_22171_n339;
  wire u_sdrc_core_u_req_gen__abc_22171_n340;
  wire u_sdrc_core_u_req_gen__abc_22171_n341_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n342;
  wire u_sdrc_core_u_req_gen__abc_22171_n343_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n344;
  wire u_sdrc_core_u_req_gen__abc_22171_n346_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n347;
  wire u_sdrc_core_u_req_gen__abc_22171_n348;
  wire u_sdrc_core_u_req_gen__abc_22171_n349;
  wire u_sdrc_core_u_req_gen__abc_22171_n350_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n351;
  wire u_sdrc_core_u_req_gen__abc_22171_n352_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n353;
  wire u_sdrc_core_u_req_gen__abc_22171_n354_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n355;
  wire u_sdrc_core_u_req_gen__abc_22171_n356;
  wire u_sdrc_core_u_req_gen__abc_22171_n357;
  wire u_sdrc_core_u_req_gen__abc_22171_n358_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n359;
  wire u_sdrc_core_u_req_gen__abc_22171_n360_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n361;
  wire u_sdrc_core_u_req_gen__abc_22171_n362;
  wire u_sdrc_core_u_req_gen__abc_22171_n363;
  wire u_sdrc_core_u_req_gen__abc_22171_n364;
  wire u_sdrc_core_u_req_gen__abc_22171_n366;
  wire u_sdrc_core_u_req_gen__abc_22171_n367;
  wire u_sdrc_core_u_req_gen__abc_22171_n368;
  wire u_sdrc_core_u_req_gen__abc_22171_n369_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n370;
  wire u_sdrc_core_u_req_gen__abc_22171_n371_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n372;
  wire u_sdrc_core_u_req_gen__abc_22171_n373_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n374;
  wire u_sdrc_core_u_req_gen__abc_22171_n375;
  wire u_sdrc_core_u_req_gen__abc_22171_n376;
  wire u_sdrc_core_u_req_gen__abc_22171_n377_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n378;
  wire u_sdrc_core_u_req_gen__abc_22171_n379_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n380;
  wire u_sdrc_core_u_req_gen__abc_22171_n381;
  wire u_sdrc_core_u_req_gen__abc_22171_n382_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n383;
  wire u_sdrc_core_u_req_gen__abc_22171_n384;
  wire u_sdrc_core_u_req_gen__abc_22171_n385;
  wire u_sdrc_core_u_req_gen__abc_22171_n386_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n387;
  wire u_sdrc_core_u_req_gen__abc_22171_n388_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n389;
  wire u_sdrc_core_u_req_gen__abc_22171_n391;
  wire u_sdrc_core_u_req_gen__abc_22171_n392;
  wire u_sdrc_core_u_req_gen__abc_22171_n393;
  wire u_sdrc_core_u_req_gen__abc_22171_n394_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n395;
  wire u_sdrc_core_u_req_gen__abc_22171_n396_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n397;
  wire u_sdrc_core_u_req_gen__abc_22171_n398;
  wire u_sdrc_core_u_req_gen__abc_22171_n399;
  wire u_sdrc_core_u_req_gen__abc_22171_n400_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n401;
  wire u_sdrc_core_u_req_gen__abc_22171_n402;
  wire u_sdrc_core_u_req_gen__abc_22171_n403;
  wire u_sdrc_core_u_req_gen__abc_22171_n404_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n405;
  wire u_sdrc_core_u_req_gen__abc_22171_n406_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n407;
  wire u_sdrc_core_u_req_gen__abc_22171_n408_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n409;
  wire u_sdrc_core_u_req_gen__abc_22171_n410;
  wire u_sdrc_core_u_req_gen__abc_22171_n411;
  wire u_sdrc_core_u_req_gen__abc_22171_n412_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n414_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n415;
  wire u_sdrc_core_u_req_gen__abc_22171_n416;
  wire u_sdrc_core_u_req_gen__abc_22171_n417_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n418;
  wire u_sdrc_core_u_req_gen__abc_22171_n419;
  wire u_sdrc_core_u_req_gen__abc_22171_n420;
  wire u_sdrc_core_u_req_gen__abc_22171_n421_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n422;
  wire u_sdrc_core_u_req_gen__abc_22171_n423_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n424;
  wire u_sdrc_core_u_req_gen__abc_22171_n425_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n426;
  wire u_sdrc_core_u_req_gen__abc_22171_n427;
  wire u_sdrc_core_u_req_gen__abc_22171_n428;
  wire u_sdrc_core_u_req_gen__abc_22171_n429_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n430;
  wire u_sdrc_core_u_req_gen__abc_22171_n431_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n432;
  wire u_sdrc_core_u_req_gen__abc_22171_n433;
  wire u_sdrc_core_u_req_gen__abc_22171_n434;
  wire u_sdrc_core_u_req_gen__abc_22171_n435;
  wire u_sdrc_core_u_req_gen__abc_22171_n436_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n438;
  wire u_sdrc_core_u_req_gen__abc_22171_n439;
  wire u_sdrc_core_u_req_gen__abc_22171_n440_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n441;
  wire u_sdrc_core_u_req_gen__abc_22171_n442_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n443;
  wire u_sdrc_core_u_req_gen__abc_22171_n444_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n445;
  wire u_sdrc_core_u_req_gen__abc_22171_n446;
  wire u_sdrc_core_u_req_gen__abc_22171_n447;
  wire u_sdrc_core_u_req_gen__abc_22171_n448_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n449;
  wire u_sdrc_core_u_req_gen__abc_22171_n450_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n451_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n452_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n453;
  wire u_sdrc_core_u_req_gen__abc_22171_n454;
  wire u_sdrc_core_u_req_gen__abc_22171_n455;
  wire u_sdrc_core_u_req_gen__abc_22171_n456;
  wire u_sdrc_core_u_req_gen__abc_22171_n457;
  wire u_sdrc_core_u_req_gen__abc_22171_n458;
  wire u_sdrc_core_u_req_gen__abc_22171_n460;
  wire u_sdrc_core_u_req_gen__abc_22171_n461;
  wire u_sdrc_core_u_req_gen__abc_22171_n462_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n463;
  wire u_sdrc_core_u_req_gen__abc_22171_n464_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n465;
  wire u_sdrc_core_u_req_gen__abc_22171_n466_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n467;
  wire u_sdrc_core_u_req_gen__abc_22171_n468_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n469;
  wire u_sdrc_core_u_req_gen__abc_22171_n470;
  wire u_sdrc_core_u_req_gen__abc_22171_n471_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n472;
  wire u_sdrc_core_u_req_gen__abc_22171_n473;
  wire u_sdrc_core_u_req_gen__abc_22171_n474_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n475;
  wire u_sdrc_core_u_req_gen__abc_22171_n476;
  wire u_sdrc_core_u_req_gen__abc_22171_n477_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n479;
  wire u_sdrc_core_u_req_gen__abc_22171_n480_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n481;
  wire u_sdrc_core_u_req_gen__abc_22171_n482;
  wire u_sdrc_core_u_req_gen__abc_22171_n483_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n484;
  wire u_sdrc_core_u_req_gen__abc_22171_n486_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n487;
  wire u_sdrc_core_u_req_gen__abc_22171_n488;
  wire u_sdrc_core_u_req_gen__abc_22171_n489_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n490;
  wire u_sdrc_core_u_req_gen__abc_22171_n491;
  wire u_sdrc_core_u_req_gen__abc_22171_n492_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n493;
  wire u_sdrc_core_u_req_gen__abc_22171_n494;
  wire u_sdrc_core_u_req_gen__abc_22171_n495_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n496;
  wire u_sdrc_core_u_req_gen__abc_22171_n497;
  wire u_sdrc_core_u_req_gen__abc_22171_n498_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n499;
  wire u_sdrc_core_u_req_gen__abc_22171_n500;
  wire u_sdrc_core_u_req_gen__abc_22171_n502;
  wire u_sdrc_core_u_req_gen__abc_22171_n503;
  wire u_sdrc_core_u_req_gen__abc_22171_n504_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n505;
  wire u_sdrc_core_u_req_gen__abc_22171_n506;
  wire u_sdrc_core_u_req_gen__abc_22171_n507_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n508_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n509_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n510_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n511;
  wire u_sdrc_core_u_req_gen__abc_22171_n512;
  wire u_sdrc_core_u_req_gen__abc_22171_n513;
  wire u_sdrc_core_u_req_gen__abc_22171_n514;
  wire u_sdrc_core_u_req_gen__abc_22171_n515;
  wire u_sdrc_core_u_req_gen__abc_22171_n516;
  wire u_sdrc_core_u_req_gen__abc_22171_n518;
  wire u_sdrc_core_u_req_gen__abc_22171_n519;
  wire u_sdrc_core_u_req_gen__abc_22171_n520;
  wire u_sdrc_core_u_req_gen__abc_22171_n521;
  wire u_sdrc_core_u_req_gen__abc_22171_n522;
  wire u_sdrc_core_u_req_gen__abc_22171_n523;
  wire u_sdrc_core_u_req_gen__abc_22171_n524;
  wire u_sdrc_core_u_req_gen__abc_22171_n525;
  wire u_sdrc_core_u_req_gen__abc_22171_n526;
  wire u_sdrc_core_u_req_gen__abc_22171_n527_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n528;
  wire u_sdrc_core_u_req_gen__abc_22171_n529_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n530;
  wire u_sdrc_core_u_req_gen__abc_22171_n531;
  wire u_sdrc_core_u_req_gen__abc_22171_n532;
  wire u_sdrc_core_u_req_gen__abc_22171_n533;
  wire u_sdrc_core_u_req_gen__abc_22171_n534;
  wire u_sdrc_core_u_req_gen__abc_22171_n536;
  wire u_sdrc_core_u_req_gen__abc_22171_n537;
  wire u_sdrc_core_u_req_gen__abc_22171_n538;
  wire u_sdrc_core_u_req_gen__abc_22171_n539;
  wire u_sdrc_core_u_req_gen__abc_22171_n540;
  wire u_sdrc_core_u_req_gen__abc_22171_n541;
  wire u_sdrc_core_u_req_gen__abc_22171_n542;
  wire u_sdrc_core_u_req_gen__abc_22171_n543;
  wire u_sdrc_core_u_req_gen__abc_22171_n544;
  wire u_sdrc_core_u_req_gen__abc_22171_n545;
  wire u_sdrc_core_u_req_gen__abc_22171_n546;
  wire u_sdrc_core_u_req_gen__abc_22171_n547;
  wire u_sdrc_core_u_req_gen__abc_22171_n548;
  wire u_sdrc_core_u_req_gen__abc_22171_n549;
  wire u_sdrc_core_u_req_gen__abc_22171_n550;
  wire u_sdrc_core_u_req_gen__abc_22171_n551;
  wire u_sdrc_core_u_req_gen__abc_22171_n552;
  wire u_sdrc_core_u_req_gen__abc_22171_n553;
  wire u_sdrc_core_u_req_gen__abc_22171_n554;
  wire u_sdrc_core_u_req_gen__abc_22171_n556;
  wire u_sdrc_core_u_req_gen__abc_22171_n557;
  wire u_sdrc_core_u_req_gen__abc_22171_n558;
  wire u_sdrc_core_u_req_gen__abc_22171_n559;
  wire u_sdrc_core_u_req_gen__abc_22171_n560;
  wire u_sdrc_core_u_req_gen__abc_22171_n561;
  wire u_sdrc_core_u_req_gen__abc_22171_n562;
  wire u_sdrc_core_u_req_gen__abc_22171_n563;
  wire u_sdrc_core_u_req_gen__abc_22171_n564;
  wire u_sdrc_core_u_req_gen__abc_22171_n565;
  wire u_sdrc_core_u_req_gen__abc_22171_n566;
  wire u_sdrc_core_u_req_gen__abc_22171_n567;
  wire u_sdrc_core_u_req_gen__abc_22171_n568;
  wire u_sdrc_core_u_req_gen__abc_22171_n569;
  wire u_sdrc_core_u_req_gen__abc_22171_n570;
  wire u_sdrc_core_u_req_gen__abc_22171_n571;
  wire u_sdrc_core_u_req_gen__abc_22171_n573;
  wire u_sdrc_core_u_req_gen__abc_22171_n574;
  wire u_sdrc_core_u_req_gen__abc_22171_n575;
  wire u_sdrc_core_u_req_gen__abc_22171_n576;
  wire u_sdrc_core_u_req_gen__abc_22171_n577;
  wire u_sdrc_core_u_req_gen__abc_22171_n578;
  wire u_sdrc_core_u_req_gen__abc_22171_n579;
  wire u_sdrc_core_u_req_gen__abc_22171_n580;
  wire u_sdrc_core_u_req_gen__abc_22171_n581;
  wire u_sdrc_core_u_req_gen__abc_22171_n582;
  wire u_sdrc_core_u_req_gen__abc_22171_n583;
  wire u_sdrc_core_u_req_gen__abc_22171_n584;
  wire u_sdrc_core_u_req_gen__abc_22171_n585;
  wire u_sdrc_core_u_req_gen__abc_22171_n586;
  wire u_sdrc_core_u_req_gen__abc_22171_n587_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n588_1;
  wire u_sdrc_core_u_req_gen__abc_22171_n589;
  wire u_sdrc_core_u_req_gen__abc_22171_n590;
  wire u_sdrc_core_u_req_gen__abc_22171_n592;
  wire u_sdrc_core_u_req_gen__abc_22171_n593;
  wire u_sdrc_core_u_req_gen__abc_22171_n594;
  wire u_sdrc_core_u_req_gen__abc_22171_n595;
  wire u_sdrc_core_u_req_gen__abc_22171_n596;
  wire u_sdrc_core_u_req_gen__abc_22171_n597;
  wire u_sdrc_core_u_req_gen__abc_22171_n598;
  wire u_sdrc_core_u_req_gen__abc_22171_n599;
  wire u_sdrc_core_u_req_gen__abc_22171_n600;
  wire u_sdrc_core_u_req_gen__abc_22171_n601;
  wire u_sdrc_core_u_req_gen__abc_22171_n602;
  wire u_sdrc_core_u_req_gen__abc_22171_n603;
  wire u_sdrc_core_u_req_gen__abc_22171_n604;
  wire u_sdrc_core_u_req_gen__abc_22171_n605;
  wire u_sdrc_core_u_req_gen__abc_22171_n607;
  wire u_sdrc_core_u_req_gen__abc_22171_n608;
  wire u_sdrc_core_u_req_gen__abc_22171_n609;
  wire u_sdrc_core_u_req_gen__abc_22171_n610;
  wire u_sdrc_core_u_req_gen__abc_22171_n611;
  wire u_sdrc_core_u_req_gen__abc_22171_n612;
  wire u_sdrc_core_u_req_gen__abc_22171_n613;
  wire u_sdrc_core_u_req_gen__abc_22171_n614;
  wire u_sdrc_core_u_req_gen__abc_22171_n615;
  wire u_sdrc_core_u_req_gen__abc_22171_n616;
  wire u_sdrc_core_u_req_gen__abc_22171_n617;
  wire u_sdrc_core_u_req_gen__abc_22171_n618;
  wire u_sdrc_core_u_req_gen__abc_22171_n619;
  wire u_sdrc_core_u_req_gen__abc_22171_n620;
  wire u_sdrc_core_u_req_gen__abc_22171_n621;
  wire u_sdrc_core_u_req_gen__abc_22171_n622;
  wire u_sdrc_core_u_req_gen__abc_22171_n623;
  wire u_sdrc_core_u_req_gen__abc_22171_n624;
  wire u_sdrc_core_u_req_gen__abc_22171_n625;
  wire u_sdrc_core_u_req_gen__abc_22171_n627;
  wire u_sdrc_core_u_req_gen__abc_22171_n628;
  wire u_sdrc_core_u_req_gen__abc_22171_n629;
  wire u_sdrc_core_u_req_gen__abc_22171_n630;
  wire u_sdrc_core_u_req_gen__abc_22171_n631;
  wire u_sdrc_core_u_req_gen__abc_22171_n632;
  wire u_sdrc_core_u_req_gen__abc_22171_n633;
  wire u_sdrc_core_u_req_gen__abc_22171_n634;
  wire u_sdrc_core_u_req_gen__abc_22171_n635;
  wire u_sdrc_core_u_req_gen__abc_22171_n636;
  wire u_sdrc_core_u_req_gen__abc_22171_n637;
  wire u_sdrc_core_u_req_gen__abc_22171_n638;
  wire u_sdrc_core_u_req_gen__abc_22171_n640;
  wire u_sdrc_core_u_req_gen__abc_22171_n641;
  wire u_sdrc_core_u_req_gen__abc_22171_n642;
  wire u_sdrc_core_u_req_gen__abc_22171_n643;
  wire u_sdrc_core_u_req_gen__abc_22171_n644;
  wire u_sdrc_core_u_req_gen__abc_22171_n645;
  wire u_sdrc_core_u_req_gen__abc_22171_n646;
  wire u_sdrc_core_u_req_gen__abc_22171_n647;
  wire u_sdrc_core_u_req_gen__abc_22171_n648;
  wire u_sdrc_core_u_req_gen__abc_22171_n649;
  wire u_sdrc_core_u_req_gen__abc_22171_n650;
  wire u_sdrc_core_u_req_gen__abc_22171_n652;
  wire u_sdrc_core_u_req_gen__abc_22171_n653;
  wire u_sdrc_core_u_req_gen__abc_22171_n654;
  wire u_sdrc_core_u_req_gen__abc_22171_n655;
  wire u_sdrc_core_u_req_gen__abc_22171_n656;
  wire u_sdrc_core_u_req_gen__abc_22171_n657;
  wire u_sdrc_core_u_req_gen__abc_22171_n658;
  wire u_sdrc_core_u_req_gen__abc_22171_n659;
  wire u_sdrc_core_u_req_gen__abc_22171_n660;
  wire u_sdrc_core_u_req_gen__abc_22171_n661;
  wire u_sdrc_core_u_req_gen__abc_22171_n662;
  wire u_sdrc_core_u_req_gen__abc_22171_n663;
  wire u_sdrc_core_u_req_gen__abc_22171_n664;
  wire u_sdrc_core_u_req_gen__abc_22171_n666;
  wire u_sdrc_core_u_req_gen__abc_22171_n667;
  wire u_sdrc_core_u_req_gen__abc_22171_n668;
  wire u_sdrc_core_u_req_gen__abc_22171_n669;
  wire u_sdrc_core_u_req_gen__abc_22171_n670;
  wire u_sdrc_core_u_req_gen__abc_22171_n671;
  wire u_sdrc_core_u_req_gen__abc_22171_n672;
  wire u_sdrc_core_u_req_gen__abc_22171_n673;
  wire u_sdrc_core_u_req_gen__abc_22171_n674;
  wire u_sdrc_core_u_req_gen__abc_22171_n675;
  wire u_sdrc_core_u_req_gen__abc_22171_n676;
  wire u_sdrc_core_u_req_gen__abc_22171_n678;
  wire u_sdrc_core_u_req_gen__abc_22171_n679;
  wire u_sdrc_core_u_req_gen__abc_22171_n680;
  wire u_sdrc_core_u_req_gen__abc_22171_n681;
  wire u_sdrc_core_u_req_gen__abc_22171_n682;
  wire u_sdrc_core_u_req_gen__abc_22171_n683;
  wire u_sdrc_core_u_req_gen__abc_22171_n684;
  wire u_sdrc_core_u_req_gen__abc_22171_n685;
  wire u_sdrc_core_u_req_gen__abc_22171_n686;
  wire u_sdrc_core_u_req_gen__abc_22171_n687;
  wire u_sdrc_core_u_req_gen__abc_22171_n688;
  wire u_sdrc_core_u_req_gen__abc_22171_n689;
  wire u_sdrc_core_u_req_gen__abc_22171_n690;
  wire u_sdrc_core_u_req_gen__abc_22171_n692;
  wire u_sdrc_core_u_req_gen__abc_22171_n693;
  wire u_sdrc_core_u_req_gen__abc_22171_n694;
  wire u_sdrc_core_u_req_gen__abc_22171_n695;
  wire u_sdrc_core_u_req_gen__abc_22171_n696;
  wire u_sdrc_core_u_req_gen__abc_22171_n697;
  wire u_sdrc_core_u_req_gen__abc_22171_n698;
  wire u_sdrc_core_u_req_gen__abc_22171_n699;
  wire u_sdrc_core_u_req_gen__abc_22171_n700;
  wire u_sdrc_core_u_req_gen__abc_22171_n701;
  wire u_sdrc_core_u_req_gen__abc_22171_n702;
  wire u_sdrc_core_u_req_gen__abc_22171_n704;
  wire u_sdrc_core_u_req_gen__abc_22171_n705;
  wire u_sdrc_core_u_req_gen__abc_22171_n706;
  wire u_sdrc_core_u_req_gen__abc_22171_n707;
  wire u_sdrc_core_u_req_gen__abc_22171_n708;
  wire u_sdrc_core_u_req_gen__abc_22171_n709;
  wire u_sdrc_core_u_req_gen__abc_22171_n710;
  wire u_sdrc_core_u_req_gen__abc_22171_n711;
  wire u_sdrc_core_u_req_gen__abc_22171_n712;
  wire u_sdrc_core_u_req_gen__abc_22171_n713;
  wire u_sdrc_core_u_req_gen__abc_22171_n714;
  wire u_sdrc_core_u_req_gen__abc_22171_n715;
  wire u_sdrc_core_u_req_gen__abc_22171_n716;
  wire u_sdrc_core_u_req_gen__abc_22171_n717;
  wire u_sdrc_core_u_req_gen__abc_22171_n719;
  wire u_sdrc_core_u_req_gen__abc_22171_n720;
  wire u_sdrc_core_u_req_gen__abc_22171_n721;
  wire u_sdrc_core_u_req_gen__abc_22171_n722;
  wire u_sdrc_core_u_req_gen__abc_22171_n723;
  wire u_sdrc_core_u_req_gen__abc_22171_n724;
  wire u_sdrc_core_u_req_gen__abc_22171_n725;
  wire u_sdrc_core_u_req_gen__abc_22171_n726;
  wire u_sdrc_core_u_req_gen__abc_22171_n727;
  wire u_sdrc_core_u_req_gen__abc_22171_n728;
  wire u_sdrc_core_u_req_gen__abc_22171_n729;
  wire u_sdrc_core_u_req_gen__abc_22171_n731;
  wire u_sdrc_core_u_req_gen__abc_22171_n732;
  wire u_sdrc_core_u_req_gen__abc_22171_n733;
  wire u_sdrc_core_u_req_gen__abc_22171_n734;
  wire u_sdrc_core_u_req_gen__abc_22171_n735;
  wire u_sdrc_core_u_req_gen__abc_22171_n736;
  wire u_sdrc_core_u_req_gen__abc_22171_n737;
  wire u_sdrc_core_u_req_gen__abc_22171_n738;
  wire u_sdrc_core_u_req_gen__abc_22171_n739;
  wire u_sdrc_core_u_req_gen__abc_22171_n740;
  wire u_sdrc_core_u_req_gen__abc_22171_n741;
  wire u_sdrc_core_u_req_gen__abc_22171_n742;
  wire u_sdrc_core_u_req_gen__abc_22171_n744;
  wire u_sdrc_core_u_req_gen__abc_22171_n745;
  wire u_sdrc_core_u_req_gen__abc_22171_n746;
  wire u_sdrc_core_u_req_gen__abc_22171_n747;
  wire u_sdrc_core_u_req_gen__abc_22171_n748;
  wire u_sdrc_core_u_req_gen__abc_22171_n749;
  wire u_sdrc_core_u_req_gen__abc_22171_n750;
  wire u_sdrc_core_u_req_gen__abc_22171_n751;
  wire u_sdrc_core_u_req_gen__abc_22171_n752;
  wire u_sdrc_core_u_req_gen__abc_22171_n753;
  wire u_sdrc_core_u_req_gen__abc_22171_n754;
  wire u_sdrc_core_u_req_gen__abc_22171_n756;
  wire u_sdrc_core_u_req_gen__abc_22171_n757;
  wire u_sdrc_core_u_req_gen__abc_22171_n758;
  wire u_sdrc_core_u_req_gen__abc_22171_n759;
  wire u_sdrc_core_u_req_gen__abc_22171_n760;
  wire u_sdrc_core_u_req_gen__abc_22171_n761;
  wire u_sdrc_core_u_req_gen__abc_22171_n762;
  wire u_sdrc_core_u_req_gen__abc_22171_n763;
  wire u_sdrc_core_u_req_gen__abc_22171_n764;
  wire u_sdrc_core_u_req_gen__abc_22171_n765;
  wire u_sdrc_core_u_req_gen__abc_22171_n766;
  wire u_sdrc_core_u_req_gen__abc_22171_n767;
  wire u_sdrc_core_u_req_gen__abc_22171_n768;
  wire u_sdrc_core_u_req_gen__abc_22171_n769;
  wire u_sdrc_core_u_req_gen__abc_22171_n770;
  wire u_sdrc_core_u_req_gen__abc_22171_n772;
  wire u_sdrc_core_u_req_gen__abc_22171_n773;
  wire u_sdrc_core_u_req_gen__abc_22171_n774;
  wire u_sdrc_core_u_req_gen__abc_22171_n775;
  wire u_sdrc_core_u_req_gen__abc_22171_n776;
  wire u_sdrc_core_u_req_gen__abc_22171_n777;
  wire u_sdrc_core_u_req_gen__abc_22171_n778;
  wire u_sdrc_core_u_req_gen__abc_22171_n779;
  wire u_sdrc_core_u_req_gen__abc_22171_n780;
  wire u_sdrc_core_u_req_gen__abc_22171_n781;
  wire u_sdrc_core_u_req_gen__abc_22171_n782;
  wire u_sdrc_core_u_req_gen__abc_22171_n783;
  wire u_sdrc_core_u_req_gen__abc_22171_n785;
  wire u_sdrc_core_u_req_gen__abc_22171_n786;
  wire u_sdrc_core_u_req_gen__abc_22171_n787;
  wire u_sdrc_core_u_req_gen__abc_22171_n788;
  wire u_sdrc_core_u_req_gen__abc_22171_n789;
  wire u_sdrc_core_u_req_gen__abc_22171_n790;
  wire u_sdrc_core_u_req_gen__abc_22171_n791;
  wire u_sdrc_core_u_req_gen__abc_22171_n792;
  wire u_sdrc_core_u_req_gen__abc_22171_n793;
  wire u_sdrc_core_u_req_gen__abc_22171_n794;
  wire u_sdrc_core_u_req_gen__abc_22171_n795;
  wire u_sdrc_core_u_req_gen__abc_22171_n796;
  wire u_sdrc_core_u_req_gen__abc_22171_n797;
  wire u_sdrc_core_u_req_gen__abc_22171_n798;
  wire u_sdrc_core_u_req_gen__abc_22171_n800;
  wire u_sdrc_core_u_req_gen__abc_22171_n801;
  wire u_sdrc_core_u_req_gen__abc_22171_n802;
  wire u_sdrc_core_u_req_gen__abc_22171_n803;
  wire u_sdrc_core_u_req_gen__abc_22171_n804;
  wire u_sdrc_core_u_req_gen__abc_22171_n805;
  wire u_sdrc_core_u_req_gen__abc_22171_n806;
  wire u_sdrc_core_u_req_gen__abc_22171_n807;
  wire u_sdrc_core_u_req_gen__abc_22171_n808;
  wire u_sdrc_core_u_req_gen__abc_22171_n809;
  wire u_sdrc_core_u_req_gen__abc_22171_n810;
  wire u_sdrc_core_u_req_gen__abc_22171_n811;
  wire u_sdrc_core_u_req_gen__abc_22171_n812;
  wire u_sdrc_core_u_req_gen__abc_22171_n813;
  wire u_sdrc_core_u_req_gen__abc_22171_n815;
  wire u_sdrc_core_u_req_gen__abc_22171_n816;
  wire u_sdrc_core_u_req_gen__abc_22171_n817;
  wire u_sdrc_core_u_req_gen__abc_22171_n818;
  wire u_sdrc_core_u_req_gen__abc_22171_n819;
  wire u_sdrc_core_u_req_gen__abc_22171_n820;
  wire u_sdrc_core_u_req_gen__abc_22171_n821;
  wire u_sdrc_core_u_req_gen__abc_22171_n822;
  wire u_sdrc_core_u_req_gen__abc_22171_n823;
  wire u_sdrc_core_u_req_gen__abc_22171_n824;
  wire u_sdrc_core_u_req_gen__abc_22171_n825;
  wire u_sdrc_core_u_req_gen__abc_22171_n826;
  wire u_sdrc_core_u_req_gen__abc_22171_n827;
  wire u_sdrc_core_u_req_gen__abc_22171_n828;
  wire u_sdrc_core_u_req_gen__abc_22171_n829;
  wire u_sdrc_core_u_req_gen__abc_22171_n830;
  wire u_sdrc_core_u_req_gen__abc_22171_n831;
  wire u_sdrc_core_u_req_gen__abc_22171_n833;
  wire u_sdrc_core_u_req_gen__abc_22171_n834;
  wire u_sdrc_core_u_req_gen__abc_22171_n835;
  wire u_sdrc_core_u_req_gen__abc_22171_n836;
  wire u_sdrc_core_u_req_gen__abc_22171_n837;
  wire u_sdrc_core_u_req_gen__abc_22171_n838;
  wire u_sdrc_core_u_req_gen__abc_22171_n839;
  wire u_sdrc_core_u_req_gen__abc_22171_n840;
  wire u_sdrc_core_u_req_gen__abc_22171_n841;
  wire u_sdrc_core_u_req_gen__abc_22171_n842;
  wire u_sdrc_core_u_req_gen__abc_22171_n843;
  wire u_sdrc_core_u_req_gen__abc_22171_n844;
  wire u_sdrc_core_u_req_gen__abc_22171_n845;
  wire u_sdrc_core_u_req_gen__abc_22171_n846;
  wire u_sdrc_core_u_req_gen__abc_22171_n847;
  wire u_sdrc_core_u_req_gen__abc_22171_n848;
  wire u_sdrc_core_u_req_gen__abc_22171_n849;
  wire u_sdrc_core_u_req_gen__abc_22171_n850;
  wire u_sdrc_core_u_req_gen__abc_22171_n852;
  wire u_sdrc_core_u_req_gen__abc_22171_n853;
  wire u_sdrc_core_u_req_gen__abc_22171_n854;
  wire u_sdrc_core_u_req_gen__abc_22171_n855;
  wire u_sdrc_core_u_req_gen__abc_22171_n856;
  wire u_sdrc_core_u_req_gen__abc_22171_n857;
  wire u_sdrc_core_u_req_gen__abc_22171_n858;
  wire u_sdrc_core_u_req_gen__abc_22171_n859;
  wire u_sdrc_core_u_req_gen__abc_22171_n860;
  wire u_sdrc_core_u_req_gen__abc_22171_n861;
  wire u_sdrc_core_u_req_gen__abc_22171_n862;
  wire u_sdrc_core_u_req_gen__abc_22171_n863;
  wire u_sdrc_core_u_req_gen__abc_22171_n864;
  wire u_sdrc_core_u_req_gen__abc_22171_n865;
  wire u_sdrc_core_u_req_gen__abc_22171_n866;
  wire u_sdrc_core_u_req_gen__abc_22171_n867;
  wire u_sdrc_core_u_req_gen__abc_22171_n868;
  wire u_sdrc_core_u_req_gen__abc_22171_n869;
  wire u_sdrc_core_u_req_gen__abc_22171_n871;
  wire u_sdrc_core_u_req_gen__abc_22171_n872;
  wire u_sdrc_core_u_req_gen__abc_22171_n873;
  wire u_sdrc_core_u_req_gen__abc_22171_n874;
  wire u_sdrc_core_u_req_gen__abc_22171_n875;
  wire u_sdrc_core_u_req_gen__abc_22171_n876;
  wire u_sdrc_core_u_req_gen__abc_22171_n877;
  wire u_sdrc_core_u_req_gen__abc_22171_n878;
  wire u_sdrc_core_u_req_gen__abc_22171_n879;
  wire u_sdrc_core_u_req_gen__abc_22171_n880;
  wire u_sdrc_core_u_req_gen__abc_22171_n881;
  wire u_sdrc_core_u_req_gen__abc_22171_n882;
  wire u_sdrc_core_u_req_gen__abc_22171_n884;
  wire u_sdrc_core_u_req_gen__abc_22171_n885;
  wire u_sdrc_core_u_req_gen__abc_22171_n886;
  wire u_sdrc_core_u_req_gen__abc_22171_n887;
  wire u_sdrc_core_u_req_gen__abc_22171_n888;
  wire u_sdrc_core_u_req_gen__abc_22171_n889;
  wire u_sdrc_core_u_req_gen__abc_22171_n890;
  wire u_sdrc_core_u_req_gen__abc_22171_n891;
  wire u_sdrc_core_u_req_gen__abc_22171_n892;
  wire u_sdrc_core_u_req_gen__abc_22171_n893;
  wire u_sdrc_core_u_req_gen__abc_22171_n893_bF_buf0;
  wire u_sdrc_core_u_req_gen__abc_22171_n893_bF_buf1;
  wire u_sdrc_core_u_req_gen__abc_22171_n893_bF_buf2;
  wire u_sdrc_core_u_req_gen__abc_22171_n893_bF_buf3;
  wire u_sdrc_core_u_req_gen__abc_22171_n894;
  wire u_sdrc_core_u_req_gen__abc_22171_n899;
  wire u_sdrc_core_u_req_gen__abc_22171_n900;
  wire u_sdrc_core_u_req_gen__abc_22171_n901;
  wire u_sdrc_core_u_req_gen__abc_22171_n902;
  wire u_sdrc_core_u_req_gen__abc_22171_n903;
  wire u_sdrc_core_u_req_gen__abc_22171_n904;
  wire u_sdrc_core_u_req_gen__abc_22171_n905;
  wire u_sdrc_core_u_req_gen__abc_22171_n907;
  wire u_sdrc_core_u_req_gen__abc_22171_n908;
  wire u_sdrc_core_u_req_gen__abc_22171_n909;
  wire u_sdrc_core_u_req_gen__abc_22171_n910;
  wire u_sdrc_core_u_req_gen__abc_22171_n911;
  wire u_sdrc_core_u_req_gen__abc_22171_n912;
  wire u_sdrc_core_u_req_gen__abc_22171_n913;
  wire u_sdrc_core_u_req_gen__abc_22171_n915;
  wire u_sdrc_core_u_req_gen__abc_22171_n916;
  wire u_sdrc_core_u_req_gen__abc_22171_n917;
  wire u_sdrc_core_u_req_gen__abc_22171_n918;
  wire u_sdrc_core_u_req_gen__abc_22171_n919;
  wire u_sdrc_core_u_req_gen__abc_22171_n920;
  wire u_sdrc_core_u_req_gen__abc_22171_n921;
  wire u_sdrc_core_u_req_gen__abc_22171_n923;
  wire u_sdrc_core_u_req_gen__abc_22171_n924;
  wire u_sdrc_core_u_req_gen__abc_22171_n925;
  wire u_sdrc_core_u_req_gen__abc_22171_n926;
  wire u_sdrc_core_u_req_gen__abc_22171_n927;
  wire u_sdrc_core_u_req_gen__abc_22171_n928;
  wire u_sdrc_core_u_req_gen__abc_22171_n930;
  wire u_sdrc_core_u_req_gen__abc_22171_n931;
  wire u_sdrc_core_u_req_gen__abc_22171_n932;
  wire u_sdrc_core_u_req_gen__abc_22171_n933;
  wire u_sdrc_core_u_req_gen__abc_22171_n934;
  wire u_sdrc_core_u_req_gen__abc_22171_n935;
  wire u_sdrc_core_u_req_gen__abc_22171_n936;
  wire u_sdrc_core_u_req_gen__abc_22171_n938;
  wire u_sdrc_core_u_req_gen__abc_22171_n939;
  wire u_sdrc_core_u_req_gen__abc_22171_n940;
  wire u_sdrc_core_u_req_gen__abc_22171_n941;
  wire u_sdrc_core_u_req_gen__abc_22171_n942;
  wire u_sdrc_core_u_req_gen__abc_22171_n943;
  wire u_sdrc_core_u_req_gen__abc_22171_n944;
  wire u_sdrc_core_u_req_gen__abc_22171_n946;
  wire u_sdrc_core_u_req_gen__abc_22171_n947;
  wire u_sdrc_core_u_req_gen__abc_22171_n948;
  wire u_sdrc_core_u_req_gen__abc_22171_n949;
  wire u_sdrc_core_u_req_gen__abc_22171_n950;
  wire u_sdrc_core_u_req_gen__abc_22171_n951;
  wire u_sdrc_core_u_req_gen__abc_22171_n952;
  wire u_sdrc_core_u_req_gen__abc_22171_n954;
  wire u_sdrc_core_u_req_gen__abc_22171_n955;
  wire u_sdrc_core_u_req_gen__abc_22171_n956;
  wire u_sdrc_core_u_req_gen__abc_22171_n957;
  wire u_sdrc_core_u_req_gen__abc_22171_n958;
  wire u_sdrc_core_u_req_gen__abc_22171_n959;
  wire u_sdrc_core_u_req_gen__abc_22171_n960;
  wire u_sdrc_core_u_req_gen__abc_22171_n962;
  wire u_sdrc_core_u_req_gen__abc_22171_n963;
  wire u_sdrc_core_u_req_gen__abc_22171_n964;
  wire u_sdrc_core_u_req_gen__abc_22171_n965;
  wire u_sdrc_core_u_req_gen__abc_22171_n966;
  wire u_sdrc_core_u_req_gen__abc_22171_n967;
  wire u_sdrc_core_u_req_gen__abc_22171_n968;
  wire u_sdrc_core_u_req_gen__abc_22171_n970;
  wire u_sdrc_core_u_req_gen__abc_22171_n971;
  wire u_sdrc_core_u_req_gen__abc_22171_n972;
  wire u_sdrc_core_u_req_gen__abc_22171_n973;
  wire u_sdrc_core_u_req_gen__abc_22171_n974;
  wire u_sdrc_core_u_req_gen__abc_22171_n975;
  wire u_sdrc_core_u_req_gen__abc_22171_n977;
  wire u_sdrc_core_u_req_gen__abc_22171_n978;
  wire u_sdrc_core_u_req_gen__abc_22171_n979;
  wire u_sdrc_core_u_req_gen__abc_22171_n980;
  wire u_sdrc_core_u_req_gen__abc_22171_n981;
  wire u_sdrc_core_u_req_gen__abc_22171_n982;
  wire u_sdrc_core_u_req_gen__abc_22171_n983;
  wire u_sdrc_core_u_req_gen__abc_22171_n984;
  wire u_sdrc_core_u_req_gen__abc_22171_n985;
  wire u_sdrc_core_u_req_gen__abc_22171_n987;
  wire u_sdrc_core_u_req_gen__abc_22171_n988;
  wire u_sdrc_core_u_req_gen__abc_22171_n989;
  wire u_sdrc_core_u_req_gen__abc_22171_n990;
  wire u_sdrc_core_u_req_gen__abc_22171_n991;
  wire u_sdrc_core_u_req_gen__abc_22171_n992;
  wire u_sdrc_core_u_req_gen__abc_22171_n993;
  wire u_sdrc_core_u_req_gen__abc_22171_n994;
  wire u_sdrc_core_u_req_gen__abc_22171_n996;
  wire u_sdrc_core_u_req_gen__abc_22171_n997;
  wire u_sdrc_core_u_req_gen__abc_22171_n998;
  wire u_sdrc_core_u_req_gen__abc_22171_n999;
  wire u_sdrc_core_u_req_gen_curr_sdr_addr_10_;
  wire u_sdrc_core_u_req_gen_curr_sdr_addr_11_;
  wire u_sdrc_core_u_req_gen_curr_sdr_addr_12_;
  wire u_sdrc_core_u_req_gen_curr_sdr_addr_13_;
  wire u_sdrc_core_u_req_gen_curr_sdr_addr_14_;
  wire u_sdrc_core_u_req_gen_curr_sdr_addr_15_;
  wire u_sdrc_core_u_req_gen_curr_sdr_addr_16_;
  wire u_sdrc_core_u_req_gen_curr_sdr_addr_17_;
  wire u_sdrc_core_u_req_gen_curr_sdr_addr_18_;
  wire u_sdrc_core_u_req_gen_curr_sdr_addr_19_;
  wire u_sdrc_core_u_req_gen_curr_sdr_addr_20_;
  wire u_sdrc_core_u_req_gen_curr_sdr_addr_21_;
  wire u_sdrc_core_u_req_gen_curr_sdr_addr_22_;
  wire u_sdrc_core_u_req_gen_curr_sdr_addr_23_;
  wire u_sdrc_core_u_req_gen_curr_sdr_addr_24_;
  wire u_sdrc_core_u_req_gen_curr_sdr_addr_25_;
  wire u_sdrc_core_u_req_gen_curr_sdr_addr_8_;
  wire u_sdrc_core_u_req_gen_curr_sdr_addr_9_;
  wire u_sdrc_core_u_req_gen_lcl_req_len_0_;
  wire u_sdrc_core_u_req_gen_lcl_req_len_0__FF_INPUT;
  wire u_sdrc_core_u_req_gen_lcl_req_len_1_;
  wire u_sdrc_core_u_req_gen_lcl_req_len_1__FF_INPUT;
  wire u_sdrc_core_u_req_gen_lcl_req_len_2_;
  wire u_sdrc_core_u_req_gen_lcl_req_len_2__FF_INPUT;
  wire u_sdrc_core_u_req_gen_lcl_req_len_3_;
  wire u_sdrc_core_u_req_gen_lcl_req_len_3__FF_INPUT;
  wire u_sdrc_core_u_req_gen_lcl_req_len_4_;
  wire u_sdrc_core_u_req_gen_lcl_req_len_4__FF_INPUT;
  wire u_sdrc_core_u_req_gen_lcl_req_len_5_;
  wire u_sdrc_core_u_req_gen_lcl_req_len_5__FF_INPUT;
  wire u_sdrc_core_u_req_gen_lcl_req_len_6_;
  wire u_sdrc_core_u_req_gen_lcl_req_len_6__FF_INPUT;
  wire u_sdrc_core_u_req_gen_lcl_wrap_FF_INPUT;
  wire u_sdrc_core_u_req_gen_map_address_0_;
  wire u_sdrc_core_u_req_gen_map_address_10_;
  wire u_sdrc_core_u_req_gen_map_address_11_;
  wire u_sdrc_core_u_req_gen_map_address_12_;
  wire u_sdrc_core_u_req_gen_map_address_13_;
  wire u_sdrc_core_u_req_gen_map_address_14_;
  wire u_sdrc_core_u_req_gen_map_address_15_;
  wire u_sdrc_core_u_req_gen_map_address_16_;
  wire u_sdrc_core_u_req_gen_map_address_17_;
  wire u_sdrc_core_u_req_gen_map_address_18_;
  wire u_sdrc_core_u_req_gen_map_address_19_;
  wire u_sdrc_core_u_req_gen_map_address_1_;
  wire u_sdrc_core_u_req_gen_map_address_20_;
  wire u_sdrc_core_u_req_gen_map_address_21_;
  wire u_sdrc_core_u_req_gen_map_address_22_;
  wire u_sdrc_core_u_req_gen_map_address_23_;
  wire u_sdrc_core_u_req_gen_map_address_24_;
  wire u_sdrc_core_u_req_gen_map_address_25_;
  wire u_sdrc_core_u_req_gen_map_address_2_;
  wire u_sdrc_core_u_req_gen_map_address_3_;
  wire u_sdrc_core_u_req_gen_map_address_4_;
  wire u_sdrc_core_u_req_gen_map_address_5_;
  wire u_sdrc_core_u_req_gen_map_address_6_;
  wire u_sdrc_core_u_req_gen_map_address_7_;
  wire u_sdrc_core_u_req_gen_map_address_8_;
  wire u_sdrc_core_u_req_gen_map_address_9_;
  wire u_sdrc_core_u_req_gen_max_r2b_len_r_0_;
  wire u_sdrc_core_u_req_gen_max_r2b_len_r_0__FF_INPUT;
  wire u_sdrc_core_u_req_gen_max_r2b_len_r_1_;
  wire u_sdrc_core_u_req_gen_max_r2b_len_r_1__FF_INPUT;
  wire u_sdrc_core_u_req_gen_max_r2b_len_r_2_;
  wire u_sdrc_core_u_req_gen_max_r2b_len_r_2__FF_INPUT;
  wire u_sdrc_core_u_req_gen_max_r2b_len_r_3_;
  wire u_sdrc_core_u_req_gen_max_r2b_len_r_3__FF_INPUT;
  wire u_sdrc_core_u_req_gen_max_r2b_len_r_4_;
  wire u_sdrc_core_u_req_gen_max_r2b_len_r_4__FF_INPUT;
  wire u_sdrc_core_u_req_gen_max_r2b_len_r_5_;
  wire u_sdrc_core_u_req_gen_max_r2b_len_r_5__FF_INPUT;
  wire u_sdrc_core_u_req_gen_max_r2b_len_r_6_;
  wire u_sdrc_core_u_req_gen_max_r2b_len_r_6__FF_INPUT;
  wire u_sdrc_core_u_req_gen_page_ovflw_r;
  wire u_sdrc_core_u_req_gen_page_ovflw_r_FF_INPUT;
  wire u_sdrc_core_u_req_gen_r2b_ba_0__FF_INPUT;
  wire u_sdrc_core_u_req_gen_r2b_ba_1__FF_INPUT;
  wire u_sdrc_core_u_req_gen_r2b_caddr_10__FF_INPUT;
  wire u_sdrc_core_u_req_gen_r2b_caddr_8__FF_INPUT;
  wire u_sdrc_core_u_req_gen_r2b_caddr_9__FF_INPUT;
  wire u_sdrc_core_u_req_gen_r2b_raddr_0__FF_INPUT;
  wire u_sdrc_core_u_req_gen_r2b_raddr_10__FF_INPUT;
  wire u_sdrc_core_u_req_gen_r2b_raddr_11__FF_INPUT;
  wire u_sdrc_core_u_req_gen_r2b_raddr_12__FF_INPUT;
  wire u_sdrc_core_u_req_gen_r2b_raddr_1__FF_INPUT;
  wire u_sdrc_core_u_req_gen_r2b_raddr_2__FF_INPUT;
  wire u_sdrc_core_u_req_gen_r2b_raddr_3__FF_INPUT;
  wire u_sdrc_core_u_req_gen_r2b_raddr_4__FF_INPUT;
  wire u_sdrc_core_u_req_gen_r2b_raddr_5__FF_INPUT;
  wire u_sdrc_core_u_req_gen_r2b_raddr_6__FF_INPUT;
  wire u_sdrc_core_u_req_gen_r2b_raddr_7__FF_INPUT;
  wire u_sdrc_core_u_req_gen_r2b_raddr_8__FF_INPUT;
  wire u_sdrc_core_u_req_gen_r2b_raddr_9__FF_INPUT;
  wire u_sdrc_core_u_req_gen_r2b_start_FF_INPUT;
  wire u_sdrc_core_u_req_gen_r2b_write_FF_INPUT;
  wire u_sdrc_core_u_req_gen_req_st_0_;
  wire u_sdrc_core_u_req_gen_req_st_1_;
  wire u_sdrc_core_u_req_gen_req_st_2_;
  wire u_sdrc_core_u_xfr_ctl__abc_16728_n178;
  wire u_sdrc_core_u_xfr_ctl__abc_16728_n181;
  wire u_sdrc_core_u_xfr_ctl__abc_16728_n184;
  wire u_sdrc_core_u_xfr_ctl__abc_16728_n189;
  wire u_sdrc_core_u_xfr_ctl__abc_16728_n258;
  wire u_sdrc_core_u_xfr_ctl__abc_16728_n270;
  wire u_sdrc_core_u_xfr_ctl__abc_16728_n35;
  wire u_sdrc_core_u_xfr_ctl__abc_16728_n43;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1000;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1001;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1002;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1004;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1005;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1006;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1007;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1008;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1009;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1010;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1011;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1013;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1014;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1015;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1016;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1017;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1018;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1019;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1020;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1021;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1023;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1024;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1025;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1026;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1027;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1028;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1029;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1031;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1032;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1033;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1034;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1035;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1036;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1037;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1038;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1040;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1041;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1042;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1043;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1044;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1045;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1046;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1047;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1048;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1049;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1050;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1051;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1052;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1053;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1054;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1055;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1056;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1058;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1059;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1060;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1061;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1062;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1063;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1064;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1065;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1066;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1067;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1068;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1070;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1071;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1072;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1073;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1074;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1075;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1076;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1077;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1078;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1079;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1080;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1082;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1083;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1084;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1085;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1086;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1087;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1088;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1090;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1091;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1092;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1093;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1094;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1095;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1096;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1097;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1098;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1099;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1100;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1101;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1102;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1103;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1105;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1106;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1107;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1108;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1109;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1110;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1111;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1112;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1113;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1115;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1116;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1117;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1118;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1119;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1120;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1121;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1122;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1123;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1125;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1126;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1127;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1128;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1129;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1130;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1132;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1133;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1134;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1135;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1136;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1137;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1138;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1139;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1140;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1141;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1142;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1143;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1144;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1145;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1146;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1147;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1148;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1149;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1150;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1151;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1152;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1153;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1154;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1155;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1156;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1157;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1158;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1159;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1160;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1161;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1162;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1163;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1164;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1165;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1166;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1167;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1168;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1169;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1170;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1171;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1172;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1173;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1174;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1175;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1176;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1177;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1178;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1179;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1180;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1181;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1182;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1183;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1184;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1185;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1186;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1187;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1188;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1189;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1190;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1191;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1192;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1193;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1194;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1195;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1196;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1197;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1198;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1199;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1200;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1201;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1202;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1203;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1204;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1206;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1207;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1208;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1209;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1211;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1212;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1213;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1214;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1216;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1217;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1218;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1219;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1221;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1222;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1223;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1224;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1226;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1227;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1228;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1229;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1231;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1232;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1233;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1234;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1236;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1237;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1238;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1239;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1241;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1242;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1243;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1244;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1246;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1247;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1248;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1249;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1251;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1252;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1253;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1254;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1256;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1257;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1258;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1260;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1261;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1262;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1263;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1265;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1266;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1267;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1268;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1270;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1271;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1272;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1273;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1275;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1276;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1277;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1278;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1279;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1280;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1281;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1282;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1283;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1284;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1285;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1287;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1288;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1289;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1290;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1291;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1292;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1293;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1294;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1295;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1296;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1297;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1311;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1312;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1314;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1315;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1317;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1318;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1320;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1321;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1323;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1324;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1326;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1327;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1329;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1330;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1332;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1333;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1335;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1336;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1338;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1339;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1341;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1342;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1344;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1345;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1347;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1348;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1350;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1351;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1353;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1354;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1356;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1357;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1359;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1360;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1363;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1364;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1365;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1367;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1370;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1374;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n1375;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n351_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n352;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n353_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n354;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n355;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n356_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n357;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n358_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n359;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n360;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n361;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n362_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n363;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n364;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n365_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n366;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n367_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n368;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n369_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n370;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n371;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n372_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n373;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n374_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n375;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n376;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n377_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n378;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n379;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n380_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n381;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n382_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n383;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n385;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n386;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n387_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n388;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n389_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n390;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n392;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n393_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n394;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n395;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n396_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n397;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n398_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n399_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n400_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n401_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n402_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n403_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n404_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n405_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n405_1_bF_buf0;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n405_1_bF_buf1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n405_1_bF_buf2;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n405_1_bF_buf3;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n406_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n407_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n408_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n409_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n410_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n411_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n413_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n414_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n415;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n416_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n418_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n419;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n420_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n421;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n423;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n424;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n425_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n426;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n428_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n429;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n430;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n431;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n432_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n433;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n434_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n435;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n436_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n438_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n439;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n441;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n442_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n444_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n445;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n446_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n447;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n448_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n449_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n450_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n451_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n452_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n453_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n454_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n455_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n456_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n457;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n458;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n459_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n460_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n461_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n462_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n463_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n464_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n465_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n466_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n467_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n468_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n469_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n470_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n471_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n472;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n473;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n474;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n475;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n476;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n477;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n478;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n479;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n480;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n481;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n482;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n483;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n484_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n485_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n486;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n487;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n488_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n489_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n490_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n491_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n492_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n493_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n494_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n495_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n496_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n497_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n498_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n499_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n500_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n501_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n502;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n503;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n505_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n506_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n507;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n508;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n509;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n510;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n511_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n512_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n513_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n514;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n515;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n516_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n517_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n518_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n519;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n520_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n521_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n522;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n523_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n523_1_bF_buf0;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n523_1_bF_buf1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n523_1_bF_buf2;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n523_1_bF_buf3;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n524_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n525;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n526_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n527;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n528;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n529_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n530_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n531;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n532;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n533_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n534_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n535;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n536_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n537;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n538;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n539_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n540_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n541;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n542_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n543;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n544;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n546_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n547;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n548_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n549;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n550;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n551_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n552_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n553;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n554_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n555;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n556;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n557_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n558_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n559;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n560_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n561;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n562;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n563_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n564_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n565;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n566_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n567;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n568;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n569_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n570_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n571;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n572_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n573;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n574;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n575_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n576_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n577;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n578_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n579;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n580;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n581_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n582_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n583;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n584_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n585;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n587_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n588_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n589;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n590_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n591;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n592;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n593_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n594_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n595;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n597;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n598;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n599_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n600_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n601;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n602;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n602_bF_buf0;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n602_bF_buf1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n602_bF_buf2;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n602_bF_buf3;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n603_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n604_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n605;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n606_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n607;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n608;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n609_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf0;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf2;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf3;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf4;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n610_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n611;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n612;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n613;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n614;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n614_bF_buf0;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n614_bF_buf1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n614_bF_buf2;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n614_bF_buf3;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n615;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n616;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n618_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n619;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n620_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n621;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n622;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n623;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n624;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n625_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n626;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n628_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n629;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n630_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n631;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n632;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n633;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n634;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n635_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n636;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n637;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n639_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n640;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n641_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n642;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n643;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n644;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n645;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n646_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n647;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n648;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n650;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n651;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n652_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n653_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n654;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n655;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n656;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n657_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n658;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n659;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n661;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n662;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n663;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n664;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n665;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n666;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n667_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n668;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n669;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n670;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n672_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n673;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n674;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n675;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n676;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n677_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n678;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n679;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n680;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n681;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n683;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n684_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n685_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n686_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n687;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n688_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n689_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n690;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n691;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n692_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n694;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n695_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n696_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n697;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n698;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n699;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n700_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n701_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n702;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n703_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n705;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n706;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n707_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n708_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n709;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n710_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n711_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n712;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n713;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n714;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n716_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n717;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n718_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n719_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n720;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n721;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n722_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n723_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n724;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n725_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n727;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n728;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n729;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n730;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n731;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n732;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n733_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n734;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n735;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n736_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n738;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n739;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n740_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n741;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n742;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n743;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n744_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n745;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n746;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n747;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n765;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n766;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n767;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n769;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n770;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n771_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n773;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n774;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n775_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n776;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n777;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n779;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n780;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n781_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n782;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n783;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n784_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n786;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n787;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n788_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n789_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n790;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n791;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n792;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n794_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n795;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n796;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n797;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n798_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n799_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n800;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n802;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n803_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n804_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n805_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n806_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n807_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n808_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n810_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n811_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n812_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n813_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n814_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n815_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n816_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n818_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n819_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n820_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n821_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n822_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n823_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n824_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n826_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n843_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n844_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n845_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n846_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n847_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n848_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n849_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n850_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n851_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n852_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n853;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n854;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n855_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n856_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n857_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n858;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n859_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n860;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n869_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n871_1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n872;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n873;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n874;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n875;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n876;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n877;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n878;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n879;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n881;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n882;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n883;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n883_bF_buf0;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n883_bF_buf1;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n883_bF_buf2;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n883_bF_buf3;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n885;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n886;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n887;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n888;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n890;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n891;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n892;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n895;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n896;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n897;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n899;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n901;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n904;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n905;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n906;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n907;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n908;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n909;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n910;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n911;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n912;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n913;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n914;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n915;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n917;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n918;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n919;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n920;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n921;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n923;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n924;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n925;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n926;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n927;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n928;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n929;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n930;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n932;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n933;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n934;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n935;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n936;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n937;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n938;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n939;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n941;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n942;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n943;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n944;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n945;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n946;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n947;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n948;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n950;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n951;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n952;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n953;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n954;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n955;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n956;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n957;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n959;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n960;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n961;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n962;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n963;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n964;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n965;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n966;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n968;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n969;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n970;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n971;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n972;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n973;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n974;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n975;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n977;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n978;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n979;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n980;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n981;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n982;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n983;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n984;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n986;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n987;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n988;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n989;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n990;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n991;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n992;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n993;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n995;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n996;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n997;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n998;
  wire u_sdrc_core_u_xfr_ctl__abc_23098_n999;
  wire u_sdrc_core_u_xfr_ctl_act_cmd;
  wire u_sdrc_core_u_xfr_ctl_act_cmd_FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_cntr1_0_;
  wire u_sdrc_core_u_xfr_ctl_cntr1_0__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_cntr1_1_;
  wire u_sdrc_core_u_xfr_ctl_cntr1_1__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_cntr1_2_;
  wire u_sdrc_core_u_xfr_ctl_cntr1_2__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_cntr1_3_;
  wire u_sdrc_core_u_xfr_ctl_cntr1_3__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_d_act_cmd;
  wire u_sdrc_core_u_xfr_ctl_d_act_cmd_FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_l_ba_0__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_l_ba_1__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_l_last;
  wire u_sdrc_core_u_xfr_ctl_l_last_FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_l_len_0_;
  wire u_sdrc_core_u_xfr_ctl_l_len_0__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_l_len_1_;
  wire u_sdrc_core_u_xfr_ctl_l_len_1__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_l_len_2_;
  wire u_sdrc_core_u_xfr_ctl_l_len_2__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_l_len_3_;
  wire u_sdrc_core_u_xfr_ctl_l_len_3__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_l_len_4_;
  wire u_sdrc_core_u_xfr_ctl_l_len_4__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_l_len_5_;
  wire u_sdrc_core_u_xfr_ctl_l_len_5__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_l_len_6_;
  wire u_sdrc_core_u_xfr_ctl_l_len_6__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_l_rd_last_0_;
  wire u_sdrc_core_u_xfr_ctl_l_rd_last_0__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_l_rd_last_1_;
  wire u_sdrc_core_u_xfr_ctl_l_rd_last_1__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_l_rd_last_2_;
  wire u_sdrc_core_u_xfr_ctl_l_rd_last_2__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_l_rd_last_3_;
  wire u_sdrc_core_u_xfr_ctl_l_rd_last_3__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_l_rd_last_4_;
  wire u_sdrc_core_u_xfr_ctl_l_rd_last_4__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_l_rd_last_5_;
  wire u_sdrc_core_u_xfr_ctl_l_rd_last_5__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_l_rd_last_6_;
  wire u_sdrc_core_u_xfr_ctl_l_rd_last_6__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_l_rd_next_0_;
  wire u_sdrc_core_u_xfr_ctl_l_rd_next_0__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_l_rd_next_1_;
  wire u_sdrc_core_u_xfr_ctl_l_rd_next_1__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_l_rd_next_2_;
  wire u_sdrc_core_u_xfr_ctl_l_rd_next_2__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_l_rd_next_3_;
  wire u_sdrc_core_u_xfr_ctl_l_rd_next_3__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_l_rd_next_4_;
  wire u_sdrc_core_u_xfr_ctl_l_rd_next_4__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_l_rd_next_5_;
  wire u_sdrc_core_u_xfr_ctl_l_rd_next_5__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_l_rd_next_6_;
  wire u_sdrc_core_u_xfr_ctl_l_rd_next_6__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_l_wrap;
  wire u_sdrc_core_u_xfr_ctl_l_wrap_FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_mgmt_st_0_;
  wire u_sdrc_core_u_xfr_ctl_mgmt_st_1_;
  wire u_sdrc_core_u_xfr_ctl_mgmt_st_2_;
  wire u_sdrc_core_u_xfr_ctl_mgmt_st_3_;
  wire u_sdrc_core_u_xfr_ctl_mgmt_st_4_;
  wire u_sdrc_core_u_xfr_ctl_mgmt_st_5_;
  wire u_sdrc_core_u_xfr_ctl_mgmt_st_6_;
  wire u_sdrc_core_u_xfr_ctl_mgmt_st_7_;
  wire u_sdrc_core_u_xfr_ctl_rfsh_row_cnt_0_;
  wire u_sdrc_core_u_xfr_ctl_rfsh_row_cnt_0__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_rfsh_row_cnt_1_;
  wire u_sdrc_core_u_xfr_ctl_rfsh_row_cnt_1__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_rfsh_row_cnt_2_;
  wire u_sdrc_core_u_xfr_ctl_rfsh_row_cnt_2__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_rfsh_timer_0_;
  wire u_sdrc_core_u_xfr_ctl_rfsh_timer_0__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_rfsh_timer_10_;
  wire u_sdrc_core_u_xfr_ctl_rfsh_timer_10__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_rfsh_timer_11_;
  wire u_sdrc_core_u_xfr_ctl_rfsh_timer_11__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_rfsh_timer_1_;
  wire u_sdrc_core_u_xfr_ctl_rfsh_timer_1__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_rfsh_timer_2_;
  wire u_sdrc_core_u_xfr_ctl_rfsh_timer_2__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_rfsh_timer_3_;
  wire u_sdrc_core_u_xfr_ctl_rfsh_timer_3__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_rfsh_timer_4_;
  wire u_sdrc_core_u_xfr_ctl_rfsh_timer_4__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_rfsh_timer_5_;
  wire u_sdrc_core_u_xfr_ctl_rfsh_timer_5__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_rfsh_timer_6_;
  wire u_sdrc_core_u_xfr_ctl_rfsh_timer_6__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_rfsh_timer_7_;
  wire u_sdrc_core_u_xfr_ctl_rfsh_timer_7__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_rfsh_timer_8_;
  wire u_sdrc_core_u_xfr_ctl_rfsh_timer_8__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_rfsh_timer_9_;
  wire u_sdrc_core_u_xfr_ctl_rfsh_timer_9__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_addr_0__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_addr_10__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_addr_11__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_addr_12__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_addr_1__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_addr_2__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_addr_3__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_addr_4__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_addr_5__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_addr_6__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_addr_7__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_addr_8__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_addr_9__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_ba_0__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_ba_1__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_cas_n_FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_cke_FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_cs_n_FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_dout_0__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_dout_10__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_dout_11__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_dout_12__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_dout_13__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_dout_14__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_dout_15__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_dout_1__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_dout_2__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_dout_3__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_dout_4__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_dout_5__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_dout_6__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_dout_7__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_dout_8__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_dout_9__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_dqm_0__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_dqm_1__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_init_done_FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_ras_n_FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_sdr_we_n_FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_tmr0_0_;
  wire u_sdrc_core_u_xfr_ctl_tmr0_0__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_tmr0_1_;
  wire u_sdrc_core_u_xfr_ctl_tmr0_1__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_tmr0_2_;
  wire u_sdrc_core_u_xfr_ctl_tmr0_2__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_tmr0_3_;
  wire u_sdrc_core_u_xfr_ctl_tmr0_3__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_xfr_caddr_0_;
  wire u_sdrc_core_u_xfr_ctl_xfr_caddr_0__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_xfr_caddr_10_;
  wire u_sdrc_core_u_xfr_ctl_xfr_caddr_10__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_xfr_caddr_11_;
  wire u_sdrc_core_u_xfr_ctl_xfr_caddr_11__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_xfr_caddr_12_;
  wire u_sdrc_core_u_xfr_ctl_xfr_caddr_12__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_xfr_caddr_1_;
  wire u_sdrc_core_u_xfr_ctl_xfr_caddr_1__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_xfr_caddr_2_;
  wire u_sdrc_core_u_xfr_ctl_xfr_caddr_2__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_xfr_caddr_3_;
  wire u_sdrc_core_u_xfr_ctl_xfr_caddr_3__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_xfr_caddr_4_;
  wire u_sdrc_core_u_xfr_ctl_xfr_caddr_4__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_xfr_caddr_5_;
  wire u_sdrc_core_u_xfr_ctl_xfr_caddr_5__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_xfr_caddr_6_;
  wire u_sdrc_core_u_xfr_ctl_xfr_caddr_6__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_xfr_caddr_7_;
  wire u_sdrc_core_u_xfr_ctl_xfr_caddr_7__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_xfr_caddr_8_;
  wire u_sdrc_core_u_xfr_ctl_xfr_caddr_8__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_xfr_caddr_9_;
  wire u_sdrc_core_u_xfr_ctl_xfr_caddr_9__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_xfr_st_0_;
  wire u_sdrc_core_u_xfr_ctl_xfr_st_0__FF_INPUT;
  wire u_sdrc_core_u_xfr_ctl_xfr_st_1_;
  wire u_sdrc_core_u_xfr_ctl_xfr_st_1__FF_INPUT;
  wire u_wb2sdrc__abc_24125_n28_1;
  wire u_wb2sdrc__abc_24125_n29_1;
  wire u_wb2sdrc__abc_24125_n30;
  wire u_wb2sdrc__abc_24125_n31;
  wire u_wb2sdrc__abc_24125_n32;
  wire u_wb2sdrc__abc_24125_n34;
  wire u_wb2sdrc__abc_24125_n35_1;
  wire u_wb2sdrc__abc_24125_n36_1;
  wire u_wb2sdrc__abc_24125_n39_1;
  wire u_wb2sdrc__abc_24125_n40;
  wire u_wb2sdrc__abc_24125_n41;
  wire u_wb2sdrc__abc_24125_n47;
  wire u_wb2sdrc_cmdfifo_empty;
  wire u_wb2sdrc_cmdfifo_full;
  wire u_wb2sdrc_cmdfifo_wr;
  wire u_wb2sdrc_pending_read;
  wire u_wb2sdrc_pending_read_FF_INPUT;
  wire u_wb2sdrc_rddatafifo_empty;
  wire u_wb2sdrc_rddatafifo_rd;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n102;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n105;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n108;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n111;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n114;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n117;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n120;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n123;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n126;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n129;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n132;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n135;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n138;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n141;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n144;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n147;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n150;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n153;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n156;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n159;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n162;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n165;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n168;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n171;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n174;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n177;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n180;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n183;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n186;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n189;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n192;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n195;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n198;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n201;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n204;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n349;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n351;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n353;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n355;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n357;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n359;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n361;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n363;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n365;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n367;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n369;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n371;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n373;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n375;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n377;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n379;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n381;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n383;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n385;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n387;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n389;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n391;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n393;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n395;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n397;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n399;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n401;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n403;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n405;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n407;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n409;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n411;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n413;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n415;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n417;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n419;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n422;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n424;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n426;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n428;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n430;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n432;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n434;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n436;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n438;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n440;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n442;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n444;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n446;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n448;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n450;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n452;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n454;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n456;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n458;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n460;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n462;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n464;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n466;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n468;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n470;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n472;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n474;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n476;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n478;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n480;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n482;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n484;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n486;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n488;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n490;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n492;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n494;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n495;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n496;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n497;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n498;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n499;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n500;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n501;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n502;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n503;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n504;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n505;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n506;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n507;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n508;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n509;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n510;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n511;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n512;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n513;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n514;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n515;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n516;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n517;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n518;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n519;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n520;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n521;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n522;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n523;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n524;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n525;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n526;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n527;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n528;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n529;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n532;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n534;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n536;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n538;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n540;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n542;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n544;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n546;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n548;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n550;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n552;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n554;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n556;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n558;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n560;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n562;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n564;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n566;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n568;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n570;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n572;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n574;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n576;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n578;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n580;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n582;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n584;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n586;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n588;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n590;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n592;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n594;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n596;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n598;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n600;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n602;
  wire u_wb2sdrc_u_cmdfifo__abc_14585_n99;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1001;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1002;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1004;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1005;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1007;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1008;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1010;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1011;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1013;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1014;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1016;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1017;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1019;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1020;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1022;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1023;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1025;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1026;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1028;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1029;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1031;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1032;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1034;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1035;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1037;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1038;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1040;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1041;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1043;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1044;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1046;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1047;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1049;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1050;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1052;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1053;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1055;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1056;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1058;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1059;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1061;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1062;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1064;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1065;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1067;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1068;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1070;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1071;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1073;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1074;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1076;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1077;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1079;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1080;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1082;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1083;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1085;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1086;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1088;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1089;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1091;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1092;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf0;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf2;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf3;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf4;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf5;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1093;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1095;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1096;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1098;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1099;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1101;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1102;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1104;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1105;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1107;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1108;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1110;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1111;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1113;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1114;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1116;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1117;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1119;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1120;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1122;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1123;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1125;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1126;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1128;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1129;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1131;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1132;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1134;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1135;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1137;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1138;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1140;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1141;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1143;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1144;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1146;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1147;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1149;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1150;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1152;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1153;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1155;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1156;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1158;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1159;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1161;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1162;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1164;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1165;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1167;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1168;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1170;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1171;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1173;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1174;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1176;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1177;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1179;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1180;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1182;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1183;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1185;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1186;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1188;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1189;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1191;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1192;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1194;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1195;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1197;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1198;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1200;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1201;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf0;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf2;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf3;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf4;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf5;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1202;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1204;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1205;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1207;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1208;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1210;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1211;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1213;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1214;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1216;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1217;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1219;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1220;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1222;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1223;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1225;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1226;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1228;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1229;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1231;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1232;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1234;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1235;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1237;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1238;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1240;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1241;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1243;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1244;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1246;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1247;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1249;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1250;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1252;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1253;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1255;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1256;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1258;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1259;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1261;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1262;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1264;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1265;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1267;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1268;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1270;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1271;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1273;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1274;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1276;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1277;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1279;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1280;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1282;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1283;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1285;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1286;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1288;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1289;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1291;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1292;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1294;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1295;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1297;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1298;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1300;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1301;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1303;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1304;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1306;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n1307;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n399;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n400_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n401_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n402;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n403_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n404_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n405;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n406_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n407_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n408;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n409_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n410_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n411;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n412_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n413_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n414;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n415_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n416_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n417;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n418_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n419_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n420;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n421_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n422_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n423;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n424_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n425_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n426;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n427_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n428_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n429;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n430_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n431_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n432;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n433_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n434_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n436_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf0;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf2;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf3;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf4;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf5;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n437_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n438;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n439_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n440_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n441;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n442_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf0;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf2;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf3;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf4;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf5;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf6;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf7;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n443_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n444;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n445_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n446_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n447;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n448_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n449_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n450;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n451_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n452_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n453;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n454_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n455;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n456_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n457_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n458_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n459_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n460_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n461_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n462_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n463_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n464_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n465_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n466_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n467_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n468_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n469_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n470_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n471_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n472_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n473_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n474_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n475_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n476_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n478_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n479_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf0;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf2;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf3;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf4;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf5;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n480_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n481_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf0;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf2;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf3;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf4;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf5;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n482_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n484_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n485_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n487_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n488_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n490_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n491_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n493_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n494_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n496_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n497_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n499_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n500_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n502_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n503_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n505_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n506_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n508_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n509_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n511_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n512_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n514_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n515_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n517_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n518_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n520_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n521_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n523_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n524_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n526_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n527_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n529;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n530_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n532_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n533_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n535_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n536_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n538_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n539_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n541_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n542_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n544_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n545_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n547_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n548_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n550_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n551_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n553_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n554_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n556_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n557_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n559_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n560_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n562_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n563_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n565_1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n566;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n568;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n569;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n571;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n572;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n574;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n575;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n577;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n578;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n580;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n581;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n583;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n584;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n586;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n587;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n589;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n590;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n591;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n593;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n594;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n595;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n596;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n597;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n598;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n599;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n600;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n601;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n602;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n603;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n604;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n605;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n606;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n608;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n610;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n611;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n613;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n615;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n617;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n618;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n619;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n620;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n621;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n622;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n624;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n625;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n627;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf0;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf2;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf3;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf4;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf5;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n628;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n629;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n630;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf0;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf2;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf3;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf4;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf5;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n631;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n633;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n634;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n635;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n636;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n637;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n638;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n639;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n641;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n643;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n644;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n645;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n646;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n647;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n648;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n649;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n651;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n653;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n654;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n655;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n657;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n658;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n659;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n660;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n661;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n662;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n663;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n664;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n666;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n667;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n668;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n669;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n670;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n671;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n672;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n673;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n675;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n676;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n677;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n678;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n679;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n680;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n681;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n682;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n684;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n685;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n686;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n687;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n688;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n689;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n690;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n691;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n693;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n694;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n695;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n696;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n697;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n698;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n699;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n700;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n702;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n703;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n704;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n705;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n706;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n707;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n708;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n709;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n711;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n712;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n713;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n714;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n715;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n716;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n717;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n718;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n720;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n721;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n722;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n723;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n724;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n725;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n726;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n727;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n729;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n730;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n731;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n732;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n733;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n734;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n735;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n736;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n738;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n739;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n740;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n741;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n742;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n743;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n744;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n745;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n747;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n748;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n749;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n750;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n751;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n752;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n753;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n754;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n756;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n757;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n758;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n759;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n760;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n761;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n762;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n763;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n765;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n766;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n767;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n768;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n769;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n770;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n771;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n772;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n774;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n775;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n776;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n777;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n778;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n779;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n780;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n781;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n783;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n784;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n785;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n786;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n787;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n788;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n789;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n790;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n792;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n793;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n794;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n795;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n796;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n797;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n798;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n799;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n801;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n802;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n803;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n804;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n805;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n806;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n807;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n808;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n810;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n811;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n812;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n813;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n814;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n815;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n816;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n817;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n819;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n820;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n821;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n822;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n823;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n824;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n825;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n826;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n828;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n829;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n830;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n831;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n832;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n833;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n834;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n835;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n837;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n838;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n839;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n840;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n841;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n842;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n843;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n844;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n846;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n847;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n848;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n849;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n850;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n851;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n852;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n853;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n855;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n856;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n857;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n858;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n859;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n860;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n861;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n862;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n864;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n865;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n866;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n867;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n868;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n869;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n870;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n871;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n873;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n874;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n875;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n876;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n877;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n878;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n879;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n880;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n882;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n883;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n884;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n885;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n886;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n887;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n888;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n889;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n891;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n892;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n893;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n894;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n895;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n896;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n897;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n898;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n900;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n901;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n902;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n903;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n904;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n905;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n906;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n907;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n909;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n910;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n911;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n912;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n913;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n914;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n915;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n916;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n918;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n919;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n920;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n921;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n922;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n923;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n924;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n925;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n927;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n928;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n929;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n930;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n931;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n932;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n933;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n934;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n936;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n937;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n938;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n939;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n940;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n941;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n942;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n943;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n945;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n946;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n947;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n948;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n949;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n950;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n951;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n952;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n954;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n955;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n956;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n957;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n958;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n959;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n960;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n961;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n963;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n964;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n965;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n966;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n967;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n968;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n969;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n970;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n972;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n973;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n974;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n975;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n976;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n977;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n978;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n979;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n981;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf0;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf2;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf3;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf4;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf5;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n982;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf0;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf1;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf2;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf3;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf4;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf5;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n983;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n984;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n986;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n987;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n989;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n990;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n992;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n993;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n995;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n996;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n998;
  wire u_wb2sdrc_u_cmdfifo__abc_18561_n999;
  wire u_wb2sdrc_u_cmdfifo_aempty;
  wire u_wb2sdrc_u_cmdfifo_afull;
  wire u_wb2sdrc_u_cmdfifo_empty_q_FF_INPUT;
  wire u_wb2sdrc_u_cmdfifo_full_q_FF_INPUT;
  wire u_wb2sdrc_u_cmdfifo_grey_rd_ptr_0_;
  wire u_wb2sdrc_u_cmdfifo_grey_rd_ptr_0__FF_INPUT;
  wire u_wb2sdrc_u_cmdfifo_grey_rd_ptr_1_;
  wire u_wb2sdrc_u_cmdfifo_grey_rd_ptr_1__FF_INPUT;
  wire u_wb2sdrc_u_cmdfifo_grey_rd_ptr_2_;
  wire u_wb2sdrc_u_cmdfifo_grey_rd_ptr_2__FF_INPUT;
  wire u_wb2sdrc_u_cmdfifo_grey_wr_ptr_0_;
  wire u_wb2sdrc_u_cmdfifo_grey_wr_ptr_0__FF_INPUT;
  wire u_wb2sdrc_u_cmdfifo_grey_wr_ptr_1_;
  wire u_wb2sdrc_u_cmdfifo_grey_wr_ptr_1__FF_INPUT;
  wire u_wb2sdrc_u_cmdfifo_grey_wr_ptr_2_;
  wire u_wb2sdrc_u_cmdfifo_grey_wr_ptr_2__FF_INPUT;
  wire u_wb2sdrc_u_cmdfifo_mem_0__0_;
  wire u_wb2sdrc_u_cmdfifo_mem_0__10_;
  wire u_wb2sdrc_u_cmdfifo_mem_0__11_;
  wire u_wb2sdrc_u_cmdfifo_mem_0__12_;
  wire u_wb2sdrc_u_cmdfifo_mem_0__13_;
  wire u_wb2sdrc_u_cmdfifo_mem_0__14_;
  wire u_wb2sdrc_u_cmdfifo_mem_0__15_;
  wire u_wb2sdrc_u_cmdfifo_mem_0__16_;
  wire u_wb2sdrc_u_cmdfifo_mem_0__17_;
  wire u_wb2sdrc_u_cmdfifo_mem_0__18_;
  wire u_wb2sdrc_u_cmdfifo_mem_0__19_;
  wire u_wb2sdrc_u_cmdfifo_mem_0__1_;
  wire u_wb2sdrc_u_cmdfifo_mem_0__20_;
  wire u_wb2sdrc_u_cmdfifo_mem_0__21_;
  wire u_wb2sdrc_u_cmdfifo_mem_0__22_;
  wire u_wb2sdrc_u_cmdfifo_mem_0__23_;
  wire u_wb2sdrc_u_cmdfifo_mem_0__24_;
  wire u_wb2sdrc_u_cmdfifo_mem_0__25_;
  wire u_wb2sdrc_u_cmdfifo_mem_0__26_;
  wire u_wb2sdrc_u_cmdfifo_mem_0__27_;
  wire u_wb2sdrc_u_cmdfifo_mem_0__28_;
  wire u_wb2sdrc_u_cmdfifo_mem_0__29_;
  wire u_wb2sdrc_u_cmdfifo_mem_0__2_;
  wire u_wb2sdrc_u_cmdfifo_mem_0__30_;
  wire u_wb2sdrc_u_cmdfifo_mem_0__31_;
  wire u_wb2sdrc_u_cmdfifo_mem_0__32_;
  wire u_wb2sdrc_u_cmdfifo_mem_0__33_;
  wire u_wb2sdrc_u_cmdfifo_mem_0__34_;
  wire u_wb2sdrc_u_cmdfifo_mem_0__35_;
  wire u_wb2sdrc_u_cmdfifo_mem_0__3_;
  wire u_wb2sdrc_u_cmdfifo_mem_0__4_;
  wire u_wb2sdrc_u_cmdfifo_mem_0__5_;
  wire u_wb2sdrc_u_cmdfifo_mem_0__6_;
  wire u_wb2sdrc_u_cmdfifo_mem_0__7_;
  wire u_wb2sdrc_u_cmdfifo_mem_0__8_;
  wire u_wb2sdrc_u_cmdfifo_mem_0__9_;
  wire u_wb2sdrc_u_cmdfifo_mem_1__0_;
  wire u_wb2sdrc_u_cmdfifo_mem_1__10_;
  wire u_wb2sdrc_u_cmdfifo_mem_1__11_;
  wire u_wb2sdrc_u_cmdfifo_mem_1__12_;
  wire u_wb2sdrc_u_cmdfifo_mem_1__13_;
  wire u_wb2sdrc_u_cmdfifo_mem_1__14_;
  wire u_wb2sdrc_u_cmdfifo_mem_1__15_;
  wire u_wb2sdrc_u_cmdfifo_mem_1__16_;
  wire u_wb2sdrc_u_cmdfifo_mem_1__17_;
  wire u_wb2sdrc_u_cmdfifo_mem_1__18_;
  wire u_wb2sdrc_u_cmdfifo_mem_1__19_;
  wire u_wb2sdrc_u_cmdfifo_mem_1__1_;
  wire u_wb2sdrc_u_cmdfifo_mem_1__20_;
  wire u_wb2sdrc_u_cmdfifo_mem_1__21_;
  wire u_wb2sdrc_u_cmdfifo_mem_1__22_;
  wire u_wb2sdrc_u_cmdfifo_mem_1__23_;
  wire u_wb2sdrc_u_cmdfifo_mem_1__24_;
  wire u_wb2sdrc_u_cmdfifo_mem_1__25_;
  wire u_wb2sdrc_u_cmdfifo_mem_1__26_;
  wire u_wb2sdrc_u_cmdfifo_mem_1__27_;
  wire u_wb2sdrc_u_cmdfifo_mem_1__28_;
  wire u_wb2sdrc_u_cmdfifo_mem_1__29_;
  wire u_wb2sdrc_u_cmdfifo_mem_1__2_;
  wire u_wb2sdrc_u_cmdfifo_mem_1__30_;
  wire u_wb2sdrc_u_cmdfifo_mem_1__31_;
  wire u_wb2sdrc_u_cmdfifo_mem_1__32_;
  wire u_wb2sdrc_u_cmdfifo_mem_1__33_;
  wire u_wb2sdrc_u_cmdfifo_mem_1__34_;
  wire u_wb2sdrc_u_cmdfifo_mem_1__35_;
  wire u_wb2sdrc_u_cmdfifo_mem_1__3_;
  wire u_wb2sdrc_u_cmdfifo_mem_1__4_;
  wire u_wb2sdrc_u_cmdfifo_mem_1__5_;
  wire u_wb2sdrc_u_cmdfifo_mem_1__6_;
  wire u_wb2sdrc_u_cmdfifo_mem_1__7_;
  wire u_wb2sdrc_u_cmdfifo_mem_1__8_;
  wire u_wb2sdrc_u_cmdfifo_mem_1__9_;
  wire u_wb2sdrc_u_cmdfifo_mem_2__0_;
  wire u_wb2sdrc_u_cmdfifo_mem_2__10_;
  wire u_wb2sdrc_u_cmdfifo_mem_2__11_;
  wire u_wb2sdrc_u_cmdfifo_mem_2__12_;
  wire u_wb2sdrc_u_cmdfifo_mem_2__13_;
  wire u_wb2sdrc_u_cmdfifo_mem_2__14_;
  wire u_wb2sdrc_u_cmdfifo_mem_2__15_;
  wire u_wb2sdrc_u_cmdfifo_mem_2__16_;
  wire u_wb2sdrc_u_cmdfifo_mem_2__17_;
  wire u_wb2sdrc_u_cmdfifo_mem_2__18_;
  wire u_wb2sdrc_u_cmdfifo_mem_2__19_;
  wire u_wb2sdrc_u_cmdfifo_mem_2__1_;
  wire u_wb2sdrc_u_cmdfifo_mem_2__20_;
  wire u_wb2sdrc_u_cmdfifo_mem_2__21_;
  wire u_wb2sdrc_u_cmdfifo_mem_2__22_;
  wire u_wb2sdrc_u_cmdfifo_mem_2__23_;
  wire u_wb2sdrc_u_cmdfifo_mem_2__24_;
  wire u_wb2sdrc_u_cmdfifo_mem_2__25_;
  wire u_wb2sdrc_u_cmdfifo_mem_2__26_;
  wire u_wb2sdrc_u_cmdfifo_mem_2__27_;
  wire u_wb2sdrc_u_cmdfifo_mem_2__28_;
  wire u_wb2sdrc_u_cmdfifo_mem_2__29_;
  wire u_wb2sdrc_u_cmdfifo_mem_2__2_;
  wire u_wb2sdrc_u_cmdfifo_mem_2__30_;
  wire u_wb2sdrc_u_cmdfifo_mem_2__31_;
  wire u_wb2sdrc_u_cmdfifo_mem_2__32_;
  wire u_wb2sdrc_u_cmdfifo_mem_2__33_;
  wire u_wb2sdrc_u_cmdfifo_mem_2__34_;
  wire u_wb2sdrc_u_cmdfifo_mem_2__35_;
  wire u_wb2sdrc_u_cmdfifo_mem_2__3_;
  wire u_wb2sdrc_u_cmdfifo_mem_2__4_;
  wire u_wb2sdrc_u_cmdfifo_mem_2__5_;
  wire u_wb2sdrc_u_cmdfifo_mem_2__6_;
  wire u_wb2sdrc_u_cmdfifo_mem_2__7_;
  wire u_wb2sdrc_u_cmdfifo_mem_2__8_;
  wire u_wb2sdrc_u_cmdfifo_mem_2__9_;
  wire u_wb2sdrc_u_cmdfifo_mem_3__0_;
  wire u_wb2sdrc_u_cmdfifo_mem_3__10_;
  wire u_wb2sdrc_u_cmdfifo_mem_3__11_;
  wire u_wb2sdrc_u_cmdfifo_mem_3__12_;
  wire u_wb2sdrc_u_cmdfifo_mem_3__13_;
  wire u_wb2sdrc_u_cmdfifo_mem_3__14_;
  wire u_wb2sdrc_u_cmdfifo_mem_3__15_;
  wire u_wb2sdrc_u_cmdfifo_mem_3__16_;
  wire u_wb2sdrc_u_cmdfifo_mem_3__17_;
  wire u_wb2sdrc_u_cmdfifo_mem_3__18_;
  wire u_wb2sdrc_u_cmdfifo_mem_3__19_;
  wire u_wb2sdrc_u_cmdfifo_mem_3__1_;
  wire u_wb2sdrc_u_cmdfifo_mem_3__20_;
  wire u_wb2sdrc_u_cmdfifo_mem_3__21_;
  wire u_wb2sdrc_u_cmdfifo_mem_3__22_;
  wire u_wb2sdrc_u_cmdfifo_mem_3__23_;
  wire u_wb2sdrc_u_cmdfifo_mem_3__24_;
  wire u_wb2sdrc_u_cmdfifo_mem_3__25_;
  wire u_wb2sdrc_u_cmdfifo_mem_3__26_;
  wire u_wb2sdrc_u_cmdfifo_mem_3__27_;
  wire u_wb2sdrc_u_cmdfifo_mem_3__28_;
  wire u_wb2sdrc_u_cmdfifo_mem_3__29_;
  wire u_wb2sdrc_u_cmdfifo_mem_3__2_;
  wire u_wb2sdrc_u_cmdfifo_mem_3__30_;
  wire u_wb2sdrc_u_cmdfifo_mem_3__31_;
  wire u_wb2sdrc_u_cmdfifo_mem_3__32_;
  wire u_wb2sdrc_u_cmdfifo_mem_3__33_;
  wire u_wb2sdrc_u_cmdfifo_mem_3__34_;
  wire u_wb2sdrc_u_cmdfifo_mem_3__35_;
  wire u_wb2sdrc_u_cmdfifo_mem_3__3_;
  wire u_wb2sdrc_u_cmdfifo_mem_3__4_;
  wire u_wb2sdrc_u_cmdfifo_mem_3__5_;
  wire u_wb2sdrc_u_cmdfifo_mem_3__6_;
  wire u_wb2sdrc_u_cmdfifo_mem_3__7_;
  wire u_wb2sdrc_u_cmdfifo_mem_3__8_;
  wire u_wb2sdrc_u_cmdfifo_mem_3__9_;
  wire u_wb2sdrc_u_cmdfifo_rd_ptr_0_;
  wire u_wb2sdrc_u_cmdfifo_rd_ptr_0__FF_INPUT;
  wire u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf0;
  wire u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf1;
  wire u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf2;
  wire u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf3;
  wire u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf4;
  wire u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf5;
  wire u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf6;
  wire u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf7;
  wire u_wb2sdrc_u_cmdfifo_rd_ptr_1_;
  wire u_wb2sdrc_u_cmdfifo_rd_ptr_1__FF_INPUT;
  wire u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf0;
  wire u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf1;
  wire u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf2;
  wire u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf3;
  wire u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf4;
  wire u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf5;
  wire u_wb2sdrc_u_cmdfifo_rd_ptr_2_;
  wire u_wb2sdrc_u_cmdfifo_rd_ptr_2__FF_INPUT;
  wire u_wb2sdrc_u_cmdfifo_sync_rd_ptr_0_0_;
  wire u_wb2sdrc_u_cmdfifo_sync_rd_ptr_0_1_;
  wire u_wb2sdrc_u_cmdfifo_sync_rd_ptr_0_2_;
  wire u_wb2sdrc_u_cmdfifo_sync_rd_ptr_1_0_;
  wire u_wb2sdrc_u_cmdfifo_sync_rd_ptr_1_1_;
  wire u_wb2sdrc_u_cmdfifo_sync_rd_ptr_2_;
  wire u_wb2sdrc_u_cmdfifo_sync_wr_ptr_0_0_;
  wire u_wb2sdrc_u_cmdfifo_sync_wr_ptr_0_1_;
  wire u_wb2sdrc_u_cmdfifo_sync_wr_ptr_0_2_;
  wire u_wb2sdrc_u_cmdfifo_sync_wr_ptr_1_0_;
  wire u_wb2sdrc_u_cmdfifo_sync_wr_ptr_1_1_;
  wire u_wb2sdrc_u_cmdfifo_sync_wr_ptr_2_;
  wire u_wb2sdrc_u_cmdfifo_wr_data_26_;
  wire u_wb2sdrc_u_cmdfifo_wr_ptr_0_;
  wire u_wb2sdrc_u_cmdfifo_wr_ptr_0__FF_INPUT;
  wire u_wb2sdrc_u_cmdfifo_wr_ptr_1_;
  wire u_wb2sdrc_u_cmdfifo_wr_ptr_1__FF_INPUT;
  wire u_wb2sdrc_u_cmdfifo_wr_ptr_2_;
  wire u_wb2sdrc_u_cmdfifo_wr_ptr_2__FF_INPUT;
  wire u_wb2sdrc_u_cmdfifo_wr_reset_n;
  wire u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf0;
  wire u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf1;
  wire u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf2;
  wire u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf3;
  wire u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf4;
  wire u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf5;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n101;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n104;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n107;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n110;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n113;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n116;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n119;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n122;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n125;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n128;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n131;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n134;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n137;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n140;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n143;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n146;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n149;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n152;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n155;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n158;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n161;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n164;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n167;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n170;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n173;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n176;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n179;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n182;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n185;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n188;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n191;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n197;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n199;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n201;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n203;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n205;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n207;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n209;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n211;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n213;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n215;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n217;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n219;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n221;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n223;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n225;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n227;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n229;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n231;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n233;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n235;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n237;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n239;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n241;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n243;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n245;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n247;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n249;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n251;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n253;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n255;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n257;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n259;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n264;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n266;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n268;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n270;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n272;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n274;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n276;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n278;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n280;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n282;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n284;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n286;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n288;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n290;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n292;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n294;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n296;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n298;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n300;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n302;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n304;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n306;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n308;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n310;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n312;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n314;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n316;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n318;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n320;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n322;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n324;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n326;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n464;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n465;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n466;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n467;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n468;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n469;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n470;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n471;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n472;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n473;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n474;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n475;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n476;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n477;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n478;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n479;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n480;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n481;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n482;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n483;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n484;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n485;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n486;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n487;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n488;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n489;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n490;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n491;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n492;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n493;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n494;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n495;
  wire u_wb2sdrc_u_rddatafifo__abc_14216_n98;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1001;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1002;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1003;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1004;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1005;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1006;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1007;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1017;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1018;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf0;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf2;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf3;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf4;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1019;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1020;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf0;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf2;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf3;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf4;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1021;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1023;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1024;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1026;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1027;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1029;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1030;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1032;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1033;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1035;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1036;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1038;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1039;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1041;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1042;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1044;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1045;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1047;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1048;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1050;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1051;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1053;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1054;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1056;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1057;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1059;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1060;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1062;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1063;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1065;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1066;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1068;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1069;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1071;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1072;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1074;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1075;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1077;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1078;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1080;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1081;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1083;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1084;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1086;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1087;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1089;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1090;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1092;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1093;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1095;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1096;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1098;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1099;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1101;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1102;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1104;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1105;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1107;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1108;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1110;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1111;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1113;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1114;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1119;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1120;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1121;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1123;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1124;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1125;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1126;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1128;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1129;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1130;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1131;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1132;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1133;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1151;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1152;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1154;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1155;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1156;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1157;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1158;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1159;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1160;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1161;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1162;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1163;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1164;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1165;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1166;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1168;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1170;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1172;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n1174;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n375_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n384_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n389;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n409;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf0;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf2;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf3;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf4;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n410;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n411_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n412_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n413;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n414;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n415_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n416_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n417;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n418;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n419_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf0;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf2;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf3;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf4;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf5;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n420_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n421;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n422;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n423_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n424_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n425;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n426;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n427_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n428_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n429;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n430;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n431_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n432_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n433;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n446;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n447_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf0;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf2;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf3;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf4;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n448;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n449;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf0;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf2;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf3;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf4;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n450_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n452_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n453_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n455_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n456_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n458_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n459_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n461_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n462_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n464_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n465_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n467_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n468_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n470_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n471_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n473_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n474_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n476_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n477_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n479_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n480_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n482_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n483_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n485;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n486_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n488;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n489_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n491;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n492;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n494;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n495_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n497;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n498;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n500_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n501_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n503_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n504;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n506;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n507;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n509_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n510_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n512;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n513;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n515;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n516;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n518;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n519;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n521_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n522_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n524_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n525;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n527_1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n528;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n530;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n531;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n533;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n534;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n536;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n537;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n539;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n540;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n542;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n543;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n548;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n549;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf0;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf2;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf3;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf4;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n550;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n551;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf0;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf2;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf3;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf4;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n552;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n554;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n555;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n557;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n558;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n560;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n561;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n563;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n564;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n566;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n567;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n569;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n570;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n572;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n573;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n575;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n576;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n578;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n579;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n581;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n582;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n584;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n585;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n587;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n588;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n590;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n591;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n593;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n594;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n596;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n597;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n599;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n600;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n602;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n603;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n605;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n606;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n608;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n609;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n611;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n612;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n614;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n615;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n617;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n618;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n620;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n621;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n623;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n624;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n626;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n627;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n629;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n630;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n632;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n633;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n635;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n636;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n638;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n639;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n641;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n642;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n644;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n645;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n650;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf0;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf2;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf3;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf4;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n651;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n652;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf0;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf2;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf3;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf4;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n653;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n655;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n656;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n658;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n659;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n661;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n662;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n664;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n665;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n667;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n668;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n670;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n671;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n673;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n674;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n676;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n677;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n679;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n680;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n682;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n683;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n685;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n686;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n688;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n689;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n691;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n692;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n694;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n695;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n697;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n698;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n700;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n701;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n703;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n704;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n706;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n707;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n709;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n710;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n712;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n713;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n715;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n716;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n718;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n719;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n721;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n722;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n724;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n725;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n727;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n728;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n730;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n731;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n733;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n734;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n736;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n737;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n739;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n740;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n742;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n743;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n745;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n746;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n751;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n752;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n753;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n754;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n755;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf0;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf2;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf3;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf4;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n756;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n757;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf0;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf1;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf2;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf3;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf4;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n758;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n759;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n761;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n762;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n763;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n764;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n765;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n766;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n767;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n769;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n770;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n771;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n772;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n773;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n774;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n775;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n777;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n778;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n779;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n780;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n781;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n782;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n783;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n785;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n786;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n787;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n788;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n789;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n790;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n791;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n793;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n794;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n795;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n796;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n797;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n798;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n799;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n801;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n802;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n803;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n804;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n805;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n806;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n807;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n809;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n810;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n811;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n812;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n813;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n814;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n815;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n817;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n818;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n819;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n820;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n821;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n822;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n823;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n825;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n826;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n827;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n828;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n829;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n830;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n831;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n833;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n834;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n835;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n836;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n837;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n838;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n839;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n841;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n842;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n843;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n844;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n845;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n846;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n847;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n849;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n850;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n851;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n852;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n853;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n854;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n855;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n857;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n858;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n859;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n860;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n861;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n862;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n863;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n865;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n866;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n867;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n868;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n869;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n870;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n871;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n873;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n874;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n875;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n876;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n877;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n878;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n879;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n881;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n882;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n883;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n884;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n885;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n886;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n887;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n889;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n890;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n891;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n892;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n893;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n894;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n895;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n897;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n898;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n899;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n900;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n901;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n902;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n903;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n905;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n906;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n907;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n908;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n909;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n910;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n911;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n913;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n914;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n915;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n916;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n917;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n918;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n919;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n921;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n922;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n923;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n924;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n925;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n926;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n927;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n929;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n930;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n931;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n932;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n933;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n934;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n935;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n937;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n938;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n939;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n940;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n941;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n942;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n943;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n945;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n946;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n947;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n948;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n949;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n950;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n951;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n953;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n954;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n955;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n956;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n957;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n958;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n959;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n961;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n962;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n963;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n964;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n965;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n966;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n967;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n969;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n970;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n971;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n972;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n973;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n974;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n975;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n977;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n978;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n979;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n980;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n981;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n982;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n983;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n985;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n986;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n987;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n988;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n989;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n990;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n991;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n993;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n994;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n995;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n996;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n997;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n998;
  wire u_wb2sdrc_u_rddatafifo__abc_17752_n999;
  wire u_wb2sdrc_u_rddatafifo_grey_wr_ptr_0_;
  wire u_wb2sdrc_u_rddatafifo_grey_wr_ptr_0__FF_INPUT;
  wire u_wb2sdrc_u_rddatafifo_grey_wr_ptr_1_;
  wire u_wb2sdrc_u_rddatafifo_grey_wr_ptr_1__FF_INPUT;
  wire u_wb2sdrc_u_rddatafifo_grey_wr_ptr_2_;
  wire u_wb2sdrc_u_rddatafifo_grey_wr_ptr_2__FF_INPUT;
  wire u_wb2sdrc_u_rddatafifo_mem_0__0_;
  wire u_wb2sdrc_u_rddatafifo_mem_0__10_;
  wire u_wb2sdrc_u_rddatafifo_mem_0__11_;
  wire u_wb2sdrc_u_rddatafifo_mem_0__12_;
  wire u_wb2sdrc_u_rddatafifo_mem_0__13_;
  wire u_wb2sdrc_u_rddatafifo_mem_0__14_;
  wire u_wb2sdrc_u_rddatafifo_mem_0__15_;
  wire u_wb2sdrc_u_rddatafifo_mem_0__16_;
  wire u_wb2sdrc_u_rddatafifo_mem_0__17_;
  wire u_wb2sdrc_u_rddatafifo_mem_0__18_;
  wire u_wb2sdrc_u_rddatafifo_mem_0__19_;
  wire u_wb2sdrc_u_rddatafifo_mem_0__1_;
  wire u_wb2sdrc_u_rddatafifo_mem_0__20_;
  wire u_wb2sdrc_u_rddatafifo_mem_0__21_;
  wire u_wb2sdrc_u_rddatafifo_mem_0__22_;
  wire u_wb2sdrc_u_rddatafifo_mem_0__23_;
  wire u_wb2sdrc_u_rddatafifo_mem_0__24_;
  wire u_wb2sdrc_u_rddatafifo_mem_0__25_;
  wire u_wb2sdrc_u_rddatafifo_mem_0__26_;
  wire u_wb2sdrc_u_rddatafifo_mem_0__27_;
  wire u_wb2sdrc_u_rddatafifo_mem_0__28_;
  wire u_wb2sdrc_u_rddatafifo_mem_0__29_;
  wire u_wb2sdrc_u_rddatafifo_mem_0__2_;
  wire u_wb2sdrc_u_rddatafifo_mem_0__30_;
  wire u_wb2sdrc_u_rddatafifo_mem_0__31_;
  wire u_wb2sdrc_u_rddatafifo_mem_0__3_;
  wire u_wb2sdrc_u_rddatafifo_mem_0__4_;
  wire u_wb2sdrc_u_rddatafifo_mem_0__5_;
  wire u_wb2sdrc_u_rddatafifo_mem_0__6_;
  wire u_wb2sdrc_u_rddatafifo_mem_0__7_;
  wire u_wb2sdrc_u_rddatafifo_mem_0__8_;
  wire u_wb2sdrc_u_rddatafifo_mem_0__9_;
  wire u_wb2sdrc_u_rddatafifo_mem_1__0_;
  wire u_wb2sdrc_u_rddatafifo_mem_1__10_;
  wire u_wb2sdrc_u_rddatafifo_mem_1__11_;
  wire u_wb2sdrc_u_rddatafifo_mem_1__12_;
  wire u_wb2sdrc_u_rddatafifo_mem_1__13_;
  wire u_wb2sdrc_u_rddatafifo_mem_1__14_;
  wire u_wb2sdrc_u_rddatafifo_mem_1__15_;
  wire u_wb2sdrc_u_rddatafifo_mem_1__16_;
  wire u_wb2sdrc_u_rddatafifo_mem_1__17_;
  wire u_wb2sdrc_u_rddatafifo_mem_1__18_;
  wire u_wb2sdrc_u_rddatafifo_mem_1__19_;
  wire u_wb2sdrc_u_rddatafifo_mem_1__1_;
  wire u_wb2sdrc_u_rddatafifo_mem_1__20_;
  wire u_wb2sdrc_u_rddatafifo_mem_1__21_;
  wire u_wb2sdrc_u_rddatafifo_mem_1__22_;
  wire u_wb2sdrc_u_rddatafifo_mem_1__23_;
  wire u_wb2sdrc_u_rddatafifo_mem_1__24_;
  wire u_wb2sdrc_u_rddatafifo_mem_1__25_;
  wire u_wb2sdrc_u_rddatafifo_mem_1__26_;
  wire u_wb2sdrc_u_rddatafifo_mem_1__27_;
  wire u_wb2sdrc_u_rddatafifo_mem_1__28_;
  wire u_wb2sdrc_u_rddatafifo_mem_1__29_;
  wire u_wb2sdrc_u_rddatafifo_mem_1__2_;
  wire u_wb2sdrc_u_rddatafifo_mem_1__30_;
  wire u_wb2sdrc_u_rddatafifo_mem_1__31_;
  wire u_wb2sdrc_u_rddatafifo_mem_1__3_;
  wire u_wb2sdrc_u_rddatafifo_mem_1__4_;
  wire u_wb2sdrc_u_rddatafifo_mem_1__5_;
  wire u_wb2sdrc_u_rddatafifo_mem_1__6_;
  wire u_wb2sdrc_u_rddatafifo_mem_1__7_;
  wire u_wb2sdrc_u_rddatafifo_mem_1__8_;
  wire u_wb2sdrc_u_rddatafifo_mem_1__9_;
  wire u_wb2sdrc_u_rddatafifo_mem_2__0_;
  wire u_wb2sdrc_u_rddatafifo_mem_2__10_;
  wire u_wb2sdrc_u_rddatafifo_mem_2__11_;
  wire u_wb2sdrc_u_rddatafifo_mem_2__12_;
  wire u_wb2sdrc_u_rddatafifo_mem_2__13_;
  wire u_wb2sdrc_u_rddatafifo_mem_2__14_;
  wire u_wb2sdrc_u_rddatafifo_mem_2__15_;
  wire u_wb2sdrc_u_rddatafifo_mem_2__16_;
  wire u_wb2sdrc_u_rddatafifo_mem_2__17_;
  wire u_wb2sdrc_u_rddatafifo_mem_2__18_;
  wire u_wb2sdrc_u_rddatafifo_mem_2__19_;
  wire u_wb2sdrc_u_rddatafifo_mem_2__1_;
  wire u_wb2sdrc_u_rddatafifo_mem_2__20_;
  wire u_wb2sdrc_u_rddatafifo_mem_2__21_;
  wire u_wb2sdrc_u_rddatafifo_mem_2__22_;
  wire u_wb2sdrc_u_rddatafifo_mem_2__23_;
  wire u_wb2sdrc_u_rddatafifo_mem_2__24_;
  wire u_wb2sdrc_u_rddatafifo_mem_2__25_;
  wire u_wb2sdrc_u_rddatafifo_mem_2__26_;
  wire u_wb2sdrc_u_rddatafifo_mem_2__27_;
  wire u_wb2sdrc_u_rddatafifo_mem_2__28_;
  wire u_wb2sdrc_u_rddatafifo_mem_2__29_;
  wire u_wb2sdrc_u_rddatafifo_mem_2__2_;
  wire u_wb2sdrc_u_rddatafifo_mem_2__30_;
  wire u_wb2sdrc_u_rddatafifo_mem_2__31_;
  wire u_wb2sdrc_u_rddatafifo_mem_2__3_;
  wire u_wb2sdrc_u_rddatafifo_mem_2__4_;
  wire u_wb2sdrc_u_rddatafifo_mem_2__5_;
  wire u_wb2sdrc_u_rddatafifo_mem_2__6_;
  wire u_wb2sdrc_u_rddatafifo_mem_2__7_;
  wire u_wb2sdrc_u_rddatafifo_mem_2__8_;
  wire u_wb2sdrc_u_rddatafifo_mem_2__9_;
  wire u_wb2sdrc_u_rddatafifo_mem_3__0_;
  wire u_wb2sdrc_u_rddatafifo_mem_3__10_;
  wire u_wb2sdrc_u_rddatafifo_mem_3__11_;
  wire u_wb2sdrc_u_rddatafifo_mem_3__12_;
  wire u_wb2sdrc_u_rddatafifo_mem_3__13_;
  wire u_wb2sdrc_u_rddatafifo_mem_3__14_;
  wire u_wb2sdrc_u_rddatafifo_mem_3__15_;
  wire u_wb2sdrc_u_rddatafifo_mem_3__16_;
  wire u_wb2sdrc_u_rddatafifo_mem_3__17_;
  wire u_wb2sdrc_u_rddatafifo_mem_3__18_;
  wire u_wb2sdrc_u_rddatafifo_mem_3__19_;
  wire u_wb2sdrc_u_rddatafifo_mem_3__1_;
  wire u_wb2sdrc_u_rddatafifo_mem_3__20_;
  wire u_wb2sdrc_u_rddatafifo_mem_3__21_;
  wire u_wb2sdrc_u_rddatafifo_mem_3__22_;
  wire u_wb2sdrc_u_rddatafifo_mem_3__23_;
  wire u_wb2sdrc_u_rddatafifo_mem_3__24_;
  wire u_wb2sdrc_u_rddatafifo_mem_3__25_;
  wire u_wb2sdrc_u_rddatafifo_mem_3__26_;
  wire u_wb2sdrc_u_rddatafifo_mem_3__27_;
  wire u_wb2sdrc_u_rddatafifo_mem_3__28_;
  wire u_wb2sdrc_u_rddatafifo_mem_3__29_;
  wire u_wb2sdrc_u_rddatafifo_mem_3__2_;
  wire u_wb2sdrc_u_rddatafifo_mem_3__30_;
  wire u_wb2sdrc_u_rddatafifo_mem_3__31_;
  wire u_wb2sdrc_u_rddatafifo_mem_3__3_;
  wire u_wb2sdrc_u_rddatafifo_mem_3__4_;
  wire u_wb2sdrc_u_rddatafifo_mem_3__5_;
  wire u_wb2sdrc_u_rddatafifo_mem_3__6_;
  wire u_wb2sdrc_u_rddatafifo_mem_3__7_;
  wire u_wb2sdrc_u_rddatafifo_mem_3__8_;
  wire u_wb2sdrc_u_rddatafifo_mem_3__9_;
  wire u_wb2sdrc_u_rddatafifo_rd_ptr_0_;
  wire u_wb2sdrc_u_rddatafifo_rd_ptr_0__FF_INPUT;
  wire u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf0;
  wire u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf1;
  wire u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf2;
  wire u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf3;
  wire u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf4;
  wire u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf5;
  wire u_wb2sdrc_u_rddatafifo_rd_ptr_1_;
  wire u_wb2sdrc_u_rddatafifo_rd_ptr_1__FF_INPUT;
  wire u_wb2sdrc_u_rddatafifo_rd_ptr_2_;
  wire u_wb2sdrc_u_rddatafifo_rd_ptr_2__FF_INPUT;
  wire u_wb2sdrc_u_rddatafifo_sync_wr_ptr_0_0_;
  wire u_wb2sdrc_u_rddatafifo_sync_wr_ptr_0_1_;
  wire u_wb2sdrc_u_rddatafifo_sync_wr_ptr_0_2_;
  wire u_wb2sdrc_u_rddatafifo_sync_wr_ptr_1_0_;
  wire u_wb2sdrc_u_rddatafifo_sync_wr_ptr_1_1_;
  wire u_wb2sdrc_u_rddatafifo_sync_wr_ptr_2_;
  wire u_wb2sdrc_u_rddatafifo_wr_ptr_0_;
  wire u_wb2sdrc_u_rddatafifo_wr_ptr_0__FF_INPUT;
  wire u_wb2sdrc_u_rddatafifo_wr_ptr_1_;
  wire u_wb2sdrc_u_rddatafifo_wr_ptr_1__FF_INPUT;
  wire u_wb2sdrc_u_rddatafifo_wr_ptr_2_;
  wire u_wb2sdrc_u_rddatafifo_wr_ptr_2__FF_INPUT;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1000;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1001;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1002;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1003;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1004;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1005;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1006;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1007;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1008;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1009;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1010;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1011;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1012;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1013;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1014;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1015;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1016;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1017;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1018;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1019;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1020;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1021;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1070;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1071;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1072;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1073;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1074;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1075;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1076;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1077;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1078;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1079;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1080;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1081;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1082;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1083;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1084;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1085;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1086;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1087;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1088;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1089;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1090;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1091;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1092;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1093;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1094;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1095;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1096;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1097;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1098;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1099;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1100;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1101;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1102;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1103;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1104;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n1105;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n154;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n157;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n160;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n163;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n166;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n169;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n172;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n175;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n178;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n181;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n184;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n187;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n190;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n193;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n196;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n199;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n202;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n205;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n208;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n211;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n214;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n217;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n220;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n223;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n226;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n229;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n232;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n235;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n238;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n241;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n244;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n247;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n250;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n253;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n256;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n259;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n513;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n515;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n517;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n519;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n521;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n523;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n525;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n527;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n529;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n531;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n533;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n535;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n537;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n539;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n541;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n543;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n545;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n547;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n549;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n551;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n553;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n555;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n557;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n559;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n561;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n563;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n565;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n567;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n569;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n571;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n573;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n575;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n577;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n579;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n581;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n583;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n586;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n588;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n590;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n592;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n594;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n596;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n598;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n600;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n602;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n604;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n606;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n608;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n610;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n612;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n614;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n616;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n618;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n620;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n622;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n624;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n626;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n628;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n630;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n632;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n634;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n636;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n638;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n640;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n642;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n644;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n646;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n648;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n650;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n652;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n654;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n656;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n767;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n768;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n769;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n770;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n771;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n772;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n773;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n774;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n775;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n776;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n777;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n778;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n779;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n780;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n781;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n782;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n783;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n784;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n785;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n786;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n787;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n788;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n789;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n790;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n791;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n792;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n793;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n794;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n795;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n796;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n797;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n798;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n799;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n800;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n801;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n802;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n876;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n877;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n878;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n879;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n880;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n881;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n882;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n883;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n884;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n885;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n886;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n887;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n888;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n889;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n890;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n891;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n892;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n893;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n894;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n895;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n896;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n897;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n898;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n899;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n900;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n901;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n902;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n903;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n904;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n905;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n906;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n907;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n908;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n909;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n910;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n911;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n914;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n916;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n918;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n920;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n922;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n924;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n926;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n928;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n930;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n932;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n934;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n936;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n938;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n940;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n942;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n944;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n946;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n948;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n950;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n952;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n954;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n956;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n958;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n960;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n962;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n964;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n966;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n968;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n970;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n972;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n974;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n976;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n978;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n980;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n982;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n984;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n986;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n987;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n988;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n989;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n990;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n991;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n992;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n993;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n994;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n995;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n996;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n997;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n998;
  wire u_wb2sdrc_u_wrdatafifo__abc_14975_n999;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1001;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1002;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1004;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1005_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1007;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1008;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1010;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1011_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1013_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1014;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1016;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1017;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1019;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1020;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1022_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1023_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1025;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1026;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1028_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1029;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1031_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1032;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1034;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1035_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1037_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1038_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1040_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1041_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf0;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf2;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf3;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf4;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf5;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1043_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf0;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf2;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf3;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf4;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf5;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1045_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1047_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1048_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1050_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1051_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1053_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1054_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1056_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1057_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1059_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1060_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1062_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1063_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1065_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1066_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1068_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1069_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1071;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1072;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1074;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1075;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1077;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1078;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1080;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1081;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1083;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1084;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1086;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1087;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1089;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1090;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1092;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1093;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1095;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1096;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1098;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1099;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1101;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1102;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1104;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1105;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1107;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1108;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1110;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1111;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1113;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1114;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1116;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1117;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1119;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1120;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1122;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1123;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1125;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1126;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1128;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1129;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1131;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1132;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1134;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1135;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1137;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1138;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1140;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1141;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1143;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1144;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1146;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1147;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1149;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1150;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1152;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1153;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1154;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1155;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1156;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf0;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf2;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf3;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf4;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf5;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf6;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf7;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1157;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1158;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf0;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf2;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf3;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf4;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf5;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf6;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf7;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1159;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1160;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1161;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1162;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1163;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1164;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1165;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1166;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1167;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1168;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1169;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1170;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1171;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1173;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1174;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1175;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1176;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1177;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1178;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1179;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1180;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1181;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1182;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1183;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1184;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1185;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1186;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1187;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1188;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1189;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1190;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1192;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1193;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1194;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1195;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1196;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1197;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1198;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1199;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1200;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1201;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1202;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1203;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1204;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1205;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1206;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1207;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1208;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1209;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1211;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1212;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1213;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1214;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1215;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1216;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1217;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1218;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1219;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1220;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1221;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1222;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1223;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1224;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1225;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1226;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1227;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1228;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1230;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1231;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1232;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1233;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1234;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1235;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1236;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1237;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1238;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1239;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1240;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1241;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1242;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1243;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1244;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1245;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1246;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1247;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1249;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1250;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1251;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1252;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1253;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1254;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1255;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1256;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1257;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1258;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1259;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1260;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1261;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1262;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1263;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1264;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1265;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1266;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1268;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1269;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1270;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1271;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1272;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1273;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1274;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1275;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1276;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1277;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1278;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1279;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1280;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1281;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1282;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1283;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1284;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1285;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1287;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1288;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1289;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1290;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1291;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1292;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1293;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1294;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1295;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1296;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1297;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1298;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1299;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1300;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1301;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1302;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1303;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1304;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1306;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1307;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1308;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1309;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1310;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1311;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1312;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1313;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1314;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1315;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1316;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1317;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1318;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1319;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1320;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1321;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1322;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1323;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1325;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1326;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1327;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1328;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1329;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1330;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1331;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1332;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1333;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1334;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1335;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1336;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1337;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1338;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1339;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1340;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1341;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1342;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1344;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1345;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1346;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1347;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1348;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1349;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1350;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1351;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1352;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1353;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1354;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1355;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1356;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1357;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1358;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1359;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1360;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1361;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1363;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1364;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1365;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1366;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1367;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1368;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1369;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1370;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1371;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1372;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1373;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1374;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1375;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1376;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1377;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1378;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1379;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1380;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1382;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1383;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1384;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1385;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1386;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1387;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1388;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1389;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1390;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1391;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1392;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1393;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1394;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1395;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1396;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1397;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1398;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1399;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1401;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1402;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1403;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1404;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1405;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1406;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1407;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1408;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1409;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1410;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1411;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1412;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1413;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1414;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1415;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1416;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1417;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1418;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1420;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1421;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1422;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1423;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1424;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1425;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1426;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1427;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1428;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1429;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1430;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1431;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1432;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1433;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1434;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1435;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1436;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1437;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1439;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1440;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1441;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1442;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1443;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1444;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1445;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1446;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1447;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1448;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1449;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1450;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1451;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1452;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1453;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1454;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1455;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1456;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1458;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1459;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1460;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1461;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1462;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1463;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1464;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1465;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1466;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1467;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1468;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1469;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1470;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1471;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1472;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1473;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1474;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1475;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1477;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1478;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1479;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1480;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1481;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1482;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1483;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1484;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1485;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1486;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1487;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1488;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1489;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1490;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1491;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1492;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1493;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1494;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1496;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1497;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1498;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1499;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1500;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1501;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1502;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1503;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1504;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1505;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1506;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1507;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1508;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1509;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1510;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1511;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1512;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1513;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1515;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1516;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1517;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1518;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1519;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1520;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1521;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1522;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1523;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1524;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1525;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1526;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1527;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1528;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1529;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1530;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1531;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1532;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1534;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1535;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1536;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1537;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1538;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1539;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1540;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1541;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1542;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1543;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1544;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1545;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1546;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1547;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1548;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1549;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1550;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1551;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1553;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1554;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1555;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1556;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1557;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1558;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1559;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1560;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1561;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1562;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1563;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1564;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1565;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1566;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1567;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1568;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1569;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1570;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1572;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1573;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1574;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1575;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1576;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1577;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1578;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1579;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1580;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1581;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1582;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1583;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1584;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1585;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1586;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1587;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1588;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1589;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1591;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1592;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1593;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1594;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1595;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1596;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1597;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1598;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1599;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1600;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1601;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1602;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1603;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1604;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1605;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1606;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1607;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1608;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1610;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1611;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1612;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1613;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1614;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1615;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1616;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1617;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1618;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1619;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1620;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1621;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1622;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1623;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1624;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1625;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1626;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1627;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1629;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1630;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1631;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1632;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1633;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1634;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1635;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1636;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1637;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1638;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1639;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1640;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1641;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1642;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1643;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1644;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1645;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1646;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1648;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1649;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1650;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1651;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1652;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1653;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1654;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1655;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1656;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1657;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1658;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1659;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1660;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1661;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1662;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1663;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1664;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1665;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1667;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1668;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1669;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1670;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1671;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1672;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1673;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1674;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1675;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1676;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1677;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1678;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1679;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1680;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1681;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1682;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1683;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1684;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1686;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1687;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1688;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1689;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1690;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1691;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1692;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1693;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1694;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1695;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1696;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1697;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1698;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1699;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1700;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1701;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1702;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1703;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1705;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1706;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1707;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1708;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1709;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1710;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1711;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1712;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1713;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1714;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1715;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1716;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1717;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1718;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1719;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1720;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1721;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1722;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1724;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1725;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1726;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1727;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1728;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1729;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1730;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1731;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1732;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1733;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1734;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1735;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1736;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1737;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1738;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1739;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1740;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1741;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1743;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1744;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1745;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1746;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1747;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1748;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1749;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1750;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1751;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1752;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1753;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1754;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1755;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1756;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1757;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1758;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1759;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1760;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1762;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1763;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1764;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1765;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1766;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1767;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1768;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1769;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1770;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1771;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1772;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1773;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1774;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1775;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1776;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1777;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1778;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1779;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1781;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1782;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1783;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1784;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1785;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1786;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1787;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1788;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1789;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1790;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1791;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1792;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1793;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1794;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1795;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1796;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1797;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1798;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1800;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1801;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1802;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1803;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1804;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1805;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1806;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1807;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1808;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1809;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1810;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1811;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1812;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1813;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1814;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1815;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1816;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1817;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1819;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1820;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1821;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1822;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1823;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1824;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1825;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1826;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1827;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1828;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1829;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1830;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1831;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1832;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1833;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1834;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1835;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1836;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1838;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1839;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf0;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf2;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf3;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf4;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf5;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1840;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1841;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf0;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf2;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf3;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf4;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf5;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1842;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1844;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1845;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1847;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1848;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1850;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1851;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1853;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1854;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1856;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1857;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1859;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1860;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1862;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1863;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1865;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1866;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1868;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1869;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1871;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1872;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1874;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1875;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1877;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1878;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1880;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1881;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1883;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1884;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1886;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1887;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1889;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1890;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1892;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1893;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1895;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1896;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1898;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1899;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1901;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1902;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1904;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1905;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1907;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1908;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1910;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1911;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1913;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1914;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1916;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1917;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1919;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1920;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1922;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1923;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1925;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1926;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1928;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1929;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1931;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1932;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1934;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1935;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1937;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1938;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1940;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1941;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1943;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1944;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1946;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1947;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1949;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf0;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf2;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf3;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf4;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf5;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1950;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1951;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf0;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf2;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf3;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf4;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf5;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1952;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1954;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1955;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1957;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1958;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1960;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1961;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1963;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1964;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1966;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1967;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1969;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1970;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1972;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1973;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1975;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1976;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1978;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1979;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1981;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1982;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1984;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1985;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1987;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1988;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1990;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1991;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1993;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1994;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1996;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1997;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n1999;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2000;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2002;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2003;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2005;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2006;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2008;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2009;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2011;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2012;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2014;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2015;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2017;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2018;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2020;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2021;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2023;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2024;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2026;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2027;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2029;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2030;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2032;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2033;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2035;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2036;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2038;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2039;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2041;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2042;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2044;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2045;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2047;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2048;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2050;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2051;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2053;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2054;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2056;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2057;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2059;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf0;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf2;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf3;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf4;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf5;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2060;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2061;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf0;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf2;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf3;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf4;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf5;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2062;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2064;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2065;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2067;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2068;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2070;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2071;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2073;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2074;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2076;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2077;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2079;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2080;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2082;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2083;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2085;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2086;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2088;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2089;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2091;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2092;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2094;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2095;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2097;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2098;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2100;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2101;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2103;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2104;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2106;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2107;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2109;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2110;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2112;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2113;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2115;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2116;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2118;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2119;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2121;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2122;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2124;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2125;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2127;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2128;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2130;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2131;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2133;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2134;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2136;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2137;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2139;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2140;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2142;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2143;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2145;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2146;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2148;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2149;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2151;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2152;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2154;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2155;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2157;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2158;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2160;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2161;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2163;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2164;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2166;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2167;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2169;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf0;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf2;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf3;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf4;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf5;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2170;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2171;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf0;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf2;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf3;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf4;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf5;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2172;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2174;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2175;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2177;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2178;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2180;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2181;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2183;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2184;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2186;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2187;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2189;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2190;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2192;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2193;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2195;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2196;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2198;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2199;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2201;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2202;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2204;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2205;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2207;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2208;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2210;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2211;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2213;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2214;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2216;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2217;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2219;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2220;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2222;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2223;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2225;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2226;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2228;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2229;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2231;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2232;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2234;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2235;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2237;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2238;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2240;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2241;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2243;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2244;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2246;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2247;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2249;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2250;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2252;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2253;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2255;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2256;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2258;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2259;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2261;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2262;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2264;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2265;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2267;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2268;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2270;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2271;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2273;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2274;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2276;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2277;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2279;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2280;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2281;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2283;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2284;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2285;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2286;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2287;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2289;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2290;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2291;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2292;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2293;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2294;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2296;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2297;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2298;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2299;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2300;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2302;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2303;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2305;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2306;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2307;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2308;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2310;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2311;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2312;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2313;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2314;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2316;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2318;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2319;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2320;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2323;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2326;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2327;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2328;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2329;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2330;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2331;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2332;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2333;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2334;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2335;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2342;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2343;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2344;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2345;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2346;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2354;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2356;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2358;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2360;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2362;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf0;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf2;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf3;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf4;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf5;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2363;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf0;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf2;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf3;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf4;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf5;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2364;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2365;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2367;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2368;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2370;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2371;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2373;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2374;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2376;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2377;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2379;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2380;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2382;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2383;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2385;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2386;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2388;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2389;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2391;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2392;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2394;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2395;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2397;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2398;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2400;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2401;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2403;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2404;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2406;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2407;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2409;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2410;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2412;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2413;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2415;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2416;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2418;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2419;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2421;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2422;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2424;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2425;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2427;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2428;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2430;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2431;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2433;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2434;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2436;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2437;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2439;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2440;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2442;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2443;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2445;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2446;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2448;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2449;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2451;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2452;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2454;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2455;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2457;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2458;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2460;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2461;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2463;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2464;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2466;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2467;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2469;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n2470;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n696_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n697_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n698;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n699_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n700;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n701;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n702_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n703;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n704_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n705_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n706;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n707;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n708_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n709_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n710;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n711_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n712;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n713;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n714_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n715;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n716_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n717_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n718;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n719;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n720_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n721_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n722;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n723_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n724;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n725;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n726_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n727;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n728_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n729_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n730;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n731;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n732_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n733_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n734;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n735_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n736;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n737;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n738_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n739;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n740_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n741_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n742;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n743;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n744_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n745_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n746;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n747_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n748;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n749;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n750_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n751;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n752_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n753_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n754;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n755;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n756_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n757_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n758;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n759_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n760;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n761;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n762_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf0;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf2;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf3;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf4;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf5;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf6;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf7;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n782;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf0;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf2;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf3;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf4;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf5;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf6;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf7;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n792_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf0;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf2;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf3;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf4;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf5;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n817_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n818_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf0;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf2;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf3;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf4;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf5;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n820_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf0;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf2;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf3;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf4;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf5;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n822_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n824_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n825_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n827_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n828_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n830_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n831_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n833_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n834_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n836_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n837_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n839_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n840_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n842_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n843;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n845_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n846_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n848_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n849_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n851_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n852_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n854_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n855_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n857_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n858_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n860_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n861_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n863_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n864_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n866_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n867_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n869_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n870_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n872_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n873_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n875_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n876_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n878_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n879_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n881_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n882_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n884_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n885_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n887_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n888_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n890_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n891_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n893_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n894_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n896_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n897_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n899_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n900_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n902_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n903_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n905_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n906_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n908_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n909_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n911_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n912_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n914_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n915_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n917;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n918_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n920_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n921_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n923_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n924_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n926_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n927_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n929_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf0;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf2;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf3;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf4;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf5;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n931_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf0;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf2;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf3;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf4;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf5;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n933_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n935_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n936_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n938_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n939_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n941_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n942_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n944_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n945_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n947_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n948_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n950_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n951_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n953_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n954_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n956;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n957_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n959;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n960;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n962;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n963;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n965_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n966_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n968;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n969;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n971_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n972;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n974;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n975;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n977_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n978_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n980;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n981;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n983;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n984_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n986;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n987;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n989_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n990;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n992;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n993_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n995;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n996;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n998_1;
  wire u_wb2sdrc_u_wrdatafifo__abc_19472_n999_1;
  wire u_wb2sdrc_u_wrdatafifo_afull;
  wire u_wb2sdrc_u_wrdatafifo_full;
  wire u_wb2sdrc_u_wrdatafifo_full_q_FF_INPUT;
  wire u_wb2sdrc_u_wrdatafifo_grey_rd_ptr_0_;
  wire u_wb2sdrc_u_wrdatafifo_grey_rd_ptr_0__FF_INPUT;
  wire u_wb2sdrc_u_wrdatafifo_grey_rd_ptr_1_;
  wire u_wb2sdrc_u_wrdatafifo_grey_rd_ptr_1__FF_INPUT;
  wire u_wb2sdrc_u_wrdatafifo_grey_rd_ptr_2_;
  wire u_wb2sdrc_u_wrdatafifo_grey_rd_ptr_2__FF_INPUT;
  wire u_wb2sdrc_u_wrdatafifo_grey_rd_ptr_3_;
  wire u_wb2sdrc_u_wrdatafifo_grey_rd_ptr_3__FF_INPUT;
  wire u_wb2sdrc_u_wrdatafifo_mem_0__0_;
  wire u_wb2sdrc_u_wrdatafifo_mem_0__10_;
  wire u_wb2sdrc_u_wrdatafifo_mem_0__11_;
  wire u_wb2sdrc_u_wrdatafifo_mem_0__12_;
  wire u_wb2sdrc_u_wrdatafifo_mem_0__13_;
  wire u_wb2sdrc_u_wrdatafifo_mem_0__14_;
  wire u_wb2sdrc_u_wrdatafifo_mem_0__15_;
  wire u_wb2sdrc_u_wrdatafifo_mem_0__16_;
  wire u_wb2sdrc_u_wrdatafifo_mem_0__17_;
  wire u_wb2sdrc_u_wrdatafifo_mem_0__18_;
  wire u_wb2sdrc_u_wrdatafifo_mem_0__19_;
  wire u_wb2sdrc_u_wrdatafifo_mem_0__1_;
  wire u_wb2sdrc_u_wrdatafifo_mem_0__20_;
  wire u_wb2sdrc_u_wrdatafifo_mem_0__21_;
  wire u_wb2sdrc_u_wrdatafifo_mem_0__22_;
  wire u_wb2sdrc_u_wrdatafifo_mem_0__23_;
  wire u_wb2sdrc_u_wrdatafifo_mem_0__24_;
  wire u_wb2sdrc_u_wrdatafifo_mem_0__25_;
  wire u_wb2sdrc_u_wrdatafifo_mem_0__26_;
  wire u_wb2sdrc_u_wrdatafifo_mem_0__27_;
  wire u_wb2sdrc_u_wrdatafifo_mem_0__28_;
  wire u_wb2sdrc_u_wrdatafifo_mem_0__29_;
  wire u_wb2sdrc_u_wrdatafifo_mem_0__2_;
  wire u_wb2sdrc_u_wrdatafifo_mem_0__30_;
  wire u_wb2sdrc_u_wrdatafifo_mem_0__31_;
  wire u_wb2sdrc_u_wrdatafifo_mem_0__32_;
  wire u_wb2sdrc_u_wrdatafifo_mem_0__33_;
  wire u_wb2sdrc_u_wrdatafifo_mem_0__34_;
  wire u_wb2sdrc_u_wrdatafifo_mem_0__35_;
  wire u_wb2sdrc_u_wrdatafifo_mem_0__3_;
  wire u_wb2sdrc_u_wrdatafifo_mem_0__4_;
  wire u_wb2sdrc_u_wrdatafifo_mem_0__5_;
  wire u_wb2sdrc_u_wrdatafifo_mem_0__6_;
  wire u_wb2sdrc_u_wrdatafifo_mem_0__7_;
  wire u_wb2sdrc_u_wrdatafifo_mem_0__8_;
  wire u_wb2sdrc_u_wrdatafifo_mem_0__9_;
  wire u_wb2sdrc_u_wrdatafifo_mem_1__0_;
  wire u_wb2sdrc_u_wrdatafifo_mem_1__10_;
  wire u_wb2sdrc_u_wrdatafifo_mem_1__11_;
  wire u_wb2sdrc_u_wrdatafifo_mem_1__12_;
  wire u_wb2sdrc_u_wrdatafifo_mem_1__13_;
  wire u_wb2sdrc_u_wrdatafifo_mem_1__14_;
  wire u_wb2sdrc_u_wrdatafifo_mem_1__15_;
  wire u_wb2sdrc_u_wrdatafifo_mem_1__16_;
  wire u_wb2sdrc_u_wrdatafifo_mem_1__17_;
  wire u_wb2sdrc_u_wrdatafifo_mem_1__18_;
  wire u_wb2sdrc_u_wrdatafifo_mem_1__19_;
  wire u_wb2sdrc_u_wrdatafifo_mem_1__1_;
  wire u_wb2sdrc_u_wrdatafifo_mem_1__20_;
  wire u_wb2sdrc_u_wrdatafifo_mem_1__21_;
  wire u_wb2sdrc_u_wrdatafifo_mem_1__22_;
  wire u_wb2sdrc_u_wrdatafifo_mem_1__23_;
  wire u_wb2sdrc_u_wrdatafifo_mem_1__24_;
  wire u_wb2sdrc_u_wrdatafifo_mem_1__25_;
  wire u_wb2sdrc_u_wrdatafifo_mem_1__26_;
  wire u_wb2sdrc_u_wrdatafifo_mem_1__27_;
  wire u_wb2sdrc_u_wrdatafifo_mem_1__28_;
  wire u_wb2sdrc_u_wrdatafifo_mem_1__29_;
  wire u_wb2sdrc_u_wrdatafifo_mem_1__2_;
  wire u_wb2sdrc_u_wrdatafifo_mem_1__30_;
  wire u_wb2sdrc_u_wrdatafifo_mem_1__31_;
  wire u_wb2sdrc_u_wrdatafifo_mem_1__32_;
  wire u_wb2sdrc_u_wrdatafifo_mem_1__33_;
  wire u_wb2sdrc_u_wrdatafifo_mem_1__34_;
  wire u_wb2sdrc_u_wrdatafifo_mem_1__35_;
  wire u_wb2sdrc_u_wrdatafifo_mem_1__3_;
  wire u_wb2sdrc_u_wrdatafifo_mem_1__4_;
  wire u_wb2sdrc_u_wrdatafifo_mem_1__5_;
  wire u_wb2sdrc_u_wrdatafifo_mem_1__6_;
  wire u_wb2sdrc_u_wrdatafifo_mem_1__7_;
  wire u_wb2sdrc_u_wrdatafifo_mem_1__8_;
  wire u_wb2sdrc_u_wrdatafifo_mem_1__9_;
  wire u_wb2sdrc_u_wrdatafifo_mem_2__0_;
  wire u_wb2sdrc_u_wrdatafifo_mem_2__10_;
  wire u_wb2sdrc_u_wrdatafifo_mem_2__11_;
  wire u_wb2sdrc_u_wrdatafifo_mem_2__12_;
  wire u_wb2sdrc_u_wrdatafifo_mem_2__13_;
  wire u_wb2sdrc_u_wrdatafifo_mem_2__14_;
  wire u_wb2sdrc_u_wrdatafifo_mem_2__15_;
  wire u_wb2sdrc_u_wrdatafifo_mem_2__16_;
  wire u_wb2sdrc_u_wrdatafifo_mem_2__17_;
  wire u_wb2sdrc_u_wrdatafifo_mem_2__18_;
  wire u_wb2sdrc_u_wrdatafifo_mem_2__19_;
  wire u_wb2sdrc_u_wrdatafifo_mem_2__1_;
  wire u_wb2sdrc_u_wrdatafifo_mem_2__20_;
  wire u_wb2sdrc_u_wrdatafifo_mem_2__21_;
  wire u_wb2sdrc_u_wrdatafifo_mem_2__22_;
  wire u_wb2sdrc_u_wrdatafifo_mem_2__23_;
  wire u_wb2sdrc_u_wrdatafifo_mem_2__24_;
  wire u_wb2sdrc_u_wrdatafifo_mem_2__25_;
  wire u_wb2sdrc_u_wrdatafifo_mem_2__26_;
  wire u_wb2sdrc_u_wrdatafifo_mem_2__27_;
  wire u_wb2sdrc_u_wrdatafifo_mem_2__28_;
  wire u_wb2sdrc_u_wrdatafifo_mem_2__29_;
  wire u_wb2sdrc_u_wrdatafifo_mem_2__2_;
  wire u_wb2sdrc_u_wrdatafifo_mem_2__30_;
  wire u_wb2sdrc_u_wrdatafifo_mem_2__31_;
  wire u_wb2sdrc_u_wrdatafifo_mem_2__32_;
  wire u_wb2sdrc_u_wrdatafifo_mem_2__33_;
  wire u_wb2sdrc_u_wrdatafifo_mem_2__34_;
  wire u_wb2sdrc_u_wrdatafifo_mem_2__35_;
  wire u_wb2sdrc_u_wrdatafifo_mem_2__3_;
  wire u_wb2sdrc_u_wrdatafifo_mem_2__4_;
  wire u_wb2sdrc_u_wrdatafifo_mem_2__5_;
  wire u_wb2sdrc_u_wrdatafifo_mem_2__6_;
  wire u_wb2sdrc_u_wrdatafifo_mem_2__7_;
  wire u_wb2sdrc_u_wrdatafifo_mem_2__8_;
  wire u_wb2sdrc_u_wrdatafifo_mem_2__9_;
  wire u_wb2sdrc_u_wrdatafifo_mem_3__0_;
  wire u_wb2sdrc_u_wrdatafifo_mem_3__10_;
  wire u_wb2sdrc_u_wrdatafifo_mem_3__11_;
  wire u_wb2sdrc_u_wrdatafifo_mem_3__12_;
  wire u_wb2sdrc_u_wrdatafifo_mem_3__13_;
  wire u_wb2sdrc_u_wrdatafifo_mem_3__14_;
  wire u_wb2sdrc_u_wrdatafifo_mem_3__15_;
  wire u_wb2sdrc_u_wrdatafifo_mem_3__16_;
  wire u_wb2sdrc_u_wrdatafifo_mem_3__17_;
  wire u_wb2sdrc_u_wrdatafifo_mem_3__18_;
  wire u_wb2sdrc_u_wrdatafifo_mem_3__19_;
  wire u_wb2sdrc_u_wrdatafifo_mem_3__1_;
  wire u_wb2sdrc_u_wrdatafifo_mem_3__20_;
  wire u_wb2sdrc_u_wrdatafifo_mem_3__21_;
  wire u_wb2sdrc_u_wrdatafifo_mem_3__22_;
  wire u_wb2sdrc_u_wrdatafifo_mem_3__23_;
  wire u_wb2sdrc_u_wrdatafifo_mem_3__24_;
  wire u_wb2sdrc_u_wrdatafifo_mem_3__25_;
  wire u_wb2sdrc_u_wrdatafifo_mem_3__26_;
  wire u_wb2sdrc_u_wrdatafifo_mem_3__27_;
  wire u_wb2sdrc_u_wrdatafifo_mem_3__28_;
  wire u_wb2sdrc_u_wrdatafifo_mem_3__29_;
  wire u_wb2sdrc_u_wrdatafifo_mem_3__2_;
  wire u_wb2sdrc_u_wrdatafifo_mem_3__30_;
  wire u_wb2sdrc_u_wrdatafifo_mem_3__31_;
  wire u_wb2sdrc_u_wrdatafifo_mem_3__32_;
  wire u_wb2sdrc_u_wrdatafifo_mem_3__33_;
  wire u_wb2sdrc_u_wrdatafifo_mem_3__34_;
  wire u_wb2sdrc_u_wrdatafifo_mem_3__35_;
  wire u_wb2sdrc_u_wrdatafifo_mem_3__3_;
  wire u_wb2sdrc_u_wrdatafifo_mem_3__4_;
  wire u_wb2sdrc_u_wrdatafifo_mem_3__5_;
  wire u_wb2sdrc_u_wrdatafifo_mem_3__6_;
  wire u_wb2sdrc_u_wrdatafifo_mem_3__7_;
  wire u_wb2sdrc_u_wrdatafifo_mem_3__8_;
  wire u_wb2sdrc_u_wrdatafifo_mem_3__9_;
  wire u_wb2sdrc_u_wrdatafifo_mem_4__0_;
  wire u_wb2sdrc_u_wrdatafifo_mem_4__10_;
  wire u_wb2sdrc_u_wrdatafifo_mem_4__11_;
  wire u_wb2sdrc_u_wrdatafifo_mem_4__12_;
  wire u_wb2sdrc_u_wrdatafifo_mem_4__13_;
  wire u_wb2sdrc_u_wrdatafifo_mem_4__14_;
  wire u_wb2sdrc_u_wrdatafifo_mem_4__15_;
  wire u_wb2sdrc_u_wrdatafifo_mem_4__16_;
  wire u_wb2sdrc_u_wrdatafifo_mem_4__17_;
  wire u_wb2sdrc_u_wrdatafifo_mem_4__18_;
  wire u_wb2sdrc_u_wrdatafifo_mem_4__19_;
  wire u_wb2sdrc_u_wrdatafifo_mem_4__1_;
  wire u_wb2sdrc_u_wrdatafifo_mem_4__20_;
  wire u_wb2sdrc_u_wrdatafifo_mem_4__21_;
  wire u_wb2sdrc_u_wrdatafifo_mem_4__22_;
  wire u_wb2sdrc_u_wrdatafifo_mem_4__23_;
  wire u_wb2sdrc_u_wrdatafifo_mem_4__24_;
  wire u_wb2sdrc_u_wrdatafifo_mem_4__25_;
  wire u_wb2sdrc_u_wrdatafifo_mem_4__26_;
  wire u_wb2sdrc_u_wrdatafifo_mem_4__27_;
  wire u_wb2sdrc_u_wrdatafifo_mem_4__28_;
  wire u_wb2sdrc_u_wrdatafifo_mem_4__29_;
  wire u_wb2sdrc_u_wrdatafifo_mem_4__2_;
  wire u_wb2sdrc_u_wrdatafifo_mem_4__30_;
  wire u_wb2sdrc_u_wrdatafifo_mem_4__31_;
  wire u_wb2sdrc_u_wrdatafifo_mem_4__32_;
  wire u_wb2sdrc_u_wrdatafifo_mem_4__33_;
  wire u_wb2sdrc_u_wrdatafifo_mem_4__34_;
  wire u_wb2sdrc_u_wrdatafifo_mem_4__35_;
  wire u_wb2sdrc_u_wrdatafifo_mem_4__3_;
  wire u_wb2sdrc_u_wrdatafifo_mem_4__4_;
  wire u_wb2sdrc_u_wrdatafifo_mem_4__5_;
  wire u_wb2sdrc_u_wrdatafifo_mem_4__6_;
  wire u_wb2sdrc_u_wrdatafifo_mem_4__7_;
  wire u_wb2sdrc_u_wrdatafifo_mem_4__8_;
  wire u_wb2sdrc_u_wrdatafifo_mem_4__9_;
  wire u_wb2sdrc_u_wrdatafifo_mem_5__0_;
  wire u_wb2sdrc_u_wrdatafifo_mem_5__10_;
  wire u_wb2sdrc_u_wrdatafifo_mem_5__11_;
  wire u_wb2sdrc_u_wrdatafifo_mem_5__12_;
  wire u_wb2sdrc_u_wrdatafifo_mem_5__13_;
  wire u_wb2sdrc_u_wrdatafifo_mem_5__14_;
  wire u_wb2sdrc_u_wrdatafifo_mem_5__15_;
  wire u_wb2sdrc_u_wrdatafifo_mem_5__16_;
  wire u_wb2sdrc_u_wrdatafifo_mem_5__17_;
  wire u_wb2sdrc_u_wrdatafifo_mem_5__18_;
  wire u_wb2sdrc_u_wrdatafifo_mem_5__19_;
  wire u_wb2sdrc_u_wrdatafifo_mem_5__1_;
  wire u_wb2sdrc_u_wrdatafifo_mem_5__20_;
  wire u_wb2sdrc_u_wrdatafifo_mem_5__21_;
  wire u_wb2sdrc_u_wrdatafifo_mem_5__22_;
  wire u_wb2sdrc_u_wrdatafifo_mem_5__23_;
  wire u_wb2sdrc_u_wrdatafifo_mem_5__24_;
  wire u_wb2sdrc_u_wrdatafifo_mem_5__25_;
  wire u_wb2sdrc_u_wrdatafifo_mem_5__26_;
  wire u_wb2sdrc_u_wrdatafifo_mem_5__27_;
  wire u_wb2sdrc_u_wrdatafifo_mem_5__28_;
  wire u_wb2sdrc_u_wrdatafifo_mem_5__29_;
  wire u_wb2sdrc_u_wrdatafifo_mem_5__2_;
  wire u_wb2sdrc_u_wrdatafifo_mem_5__30_;
  wire u_wb2sdrc_u_wrdatafifo_mem_5__31_;
  wire u_wb2sdrc_u_wrdatafifo_mem_5__32_;
  wire u_wb2sdrc_u_wrdatafifo_mem_5__33_;
  wire u_wb2sdrc_u_wrdatafifo_mem_5__34_;
  wire u_wb2sdrc_u_wrdatafifo_mem_5__35_;
  wire u_wb2sdrc_u_wrdatafifo_mem_5__3_;
  wire u_wb2sdrc_u_wrdatafifo_mem_5__4_;
  wire u_wb2sdrc_u_wrdatafifo_mem_5__5_;
  wire u_wb2sdrc_u_wrdatafifo_mem_5__6_;
  wire u_wb2sdrc_u_wrdatafifo_mem_5__7_;
  wire u_wb2sdrc_u_wrdatafifo_mem_5__8_;
  wire u_wb2sdrc_u_wrdatafifo_mem_5__9_;
  wire u_wb2sdrc_u_wrdatafifo_mem_6__0_;
  wire u_wb2sdrc_u_wrdatafifo_mem_6__10_;
  wire u_wb2sdrc_u_wrdatafifo_mem_6__11_;
  wire u_wb2sdrc_u_wrdatafifo_mem_6__12_;
  wire u_wb2sdrc_u_wrdatafifo_mem_6__13_;
  wire u_wb2sdrc_u_wrdatafifo_mem_6__14_;
  wire u_wb2sdrc_u_wrdatafifo_mem_6__15_;
  wire u_wb2sdrc_u_wrdatafifo_mem_6__16_;
  wire u_wb2sdrc_u_wrdatafifo_mem_6__17_;
  wire u_wb2sdrc_u_wrdatafifo_mem_6__18_;
  wire u_wb2sdrc_u_wrdatafifo_mem_6__19_;
  wire u_wb2sdrc_u_wrdatafifo_mem_6__1_;
  wire u_wb2sdrc_u_wrdatafifo_mem_6__20_;
  wire u_wb2sdrc_u_wrdatafifo_mem_6__21_;
  wire u_wb2sdrc_u_wrdatafifo_mem_6__22_;
  wire u_wb2sdrc_u_wrdatafifo_mem_6__23_;
  wire u_wb2sdrc_u_wrdatafifo_mem_6__24_;
  wire u_wb2sdrc_u_wrdatafifo_mem_6__25_;
  wire u_wb2sdrc_u_wrdatafifo_mem_6__26_;
  wire u_wb2sdrc_u_wrdatafifo_mem_6__27_;
  wire u_wb2sdrc_u_wrdatafifo_mem_6__28_;
  wire u_wb2sdrc_u_wrdatafifo_mem_6__29_;
  wire u_wb2sdrc_u_wrdatafifo_mem_6__2_;
  wire u_wb2sdrc_u_wrdatafifo_mem_6__30_;
  wire u_wb2sdrc_u_wrdatafifo_mem_6__31_;
  wire u_wb2sdrc_u_wrdatafifo_mem_6__32_;
  wire u_wb2sdrc_u_wrdatafifo_mem_6__33_;
  wire u_wb2sdrc_u_wrdatafifo_mem_6__34_;
  wire u_wb2sdrc_u_wrdatafifo_mem_6__35_;
  wire u_wb2sdrc_u_wrdatafifo_mem_6__3_;
  wire u_wb2sdrc_u_wrdatafifo_mem_6__4_;
  wire u_wb2sdrc_u_wrdatafifo_mem_6__5_;
  wire u_wb2sdrc_u_wrdatafifo_mem_6__6_;
  wire u_wb2sdrc_u_wrdatafifo_mem_6__7_;
  wire u_wb2sdrc_u_wrdatafifo_mem_6__8_;
  wire u_wb2sdrc_u_wrdatafifo_mem_6__9_;
  wire u_wb2sdrc_u_wrdatafifo_mem_7__0_;
  wire u_wb2sdrc_u_wrdatafifo_mem_7__10_;
  wire u_wb2sdrc_u_wrdatafifo_mem_7__11_;
  wire u_wb2sdrc_u_wrdatafifo_mem_7__12_;
  wire u_wb2sdrc_u_wrdatafifo_mem_7__13_;
  wire u_wb2sdrc_u_wrdatafifo_mem_7__14_;
  wire u_wb2sdrc_u_wrdatafifo_mem_7__15_;
  wire u_wb2sdrc_u_wrdatafifo_mem_7__16_;
  wire u_wb2sdrc_u_wrdatafifo_mem_7__17_;
  wire u_wb2sdrc_u_wrdatafifo_mem_7__18_;
  wire u_wb2sdrc_u_wrdatafifo_mem_7__19_;
  wire u_wb2sdrc_u_wrdatafifo_mem_7__1_;
  wire u_wb2sdrc_u_wrdatafifo_mem_7__20_;
  wire u_wb2sdrc_u_wrdatafifo_mem_7__21_;
  wire u_wb2sdrc_u_wrdatafifo_mem_7__22_;
  wire u_wb2sdrc_u_wrdatafifo_mem_7__23_;
  wire u_wb2sdrc_u_wrdatafifo_mem_7__24_;
  wire u_wb2sdrc_u_wrdatafifo_mem_7__25_;
  wire u_wb2sdrc_u_wrdatafifo_mem_7__26_;
  wire u_wb2sdrc_u_wrdatafifo_mem_7__27_;
  wire u_wb2sdrc_u_wrdatafifo_mem_7__28_;
  wire u_wb2sdrc_u_wrdatafifo_mem_7__29_;
  wire u_wb2sdrc_u_wrdatafifo_mem_7__2_;
  wire u_wb2sdrc_u_wrdatafifo_mem_7__30_;
  wire u_wb2sdrc_u_wrdatafifo_mem_7__31_;
  wire u_wb2sdrc_u_wrdatafifo_mem_7__32_;
  wire u_wb2sdrc_u_wrdatafifo_mem_7__33_;
  wire u_wb2sdrc_u_wrdatafifo_mem_7__34_;
  wire u_wb2sdrc_u_wrdatafifo_mem_7__35_;
  wire u_wb2sdrc_u_wrdatafifo_mem_7__3_;
  wire u_wb2sdrc_u_wrdatafifo_mem_7__4_;
  wire u_wb2sdrc_u_wrdatafifo_mem_7__5_;
  wire u_wb2sdrc_u_wrdatafifo_mem_7__6_;
  wire u_wb2sdrc_u_wrdatafifo_mem_7__7_;
  wire u_wb2sdrc_u_wrdatafifo_mem_7__8_;
  wire u_wb2sdrc_u_wrdatafifo_mem_7__9_;
  wire u_wb2sdrc_u_wrdatafifo_rd_ptr_0_;
  wire u_wb2sdrc_u_wrdatafifo_rd_ptr_0__FF_INPUT;
  wire u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf0;
  wire u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf1;
  wire u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf2;
  wire u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf3;
  wire u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf4;
  wire u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf5;
  wire u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf6;
  wire u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf7;
  wire u_wb2sdrc_u_wrdatafifo_rd_ptr_1_;
  wire u_wb2sdrc_u_wrdatafifo_rd_ptr_1__FF_INPUT;
  wire u_wb2sdrc_u_wrdatafifo_rd_ptr_2_;
  wire u_wb2sdrc_u_wrdatafifo_rd_ptr_2__FF_INPUT;
  wire u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf0;
  wire u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf1;
  wire u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf2;
  wire u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf3;
  wire u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf4;
  wire u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf5;
  wire u_wb2sdrc_u_wrdatafifo_rd_ptr_3_;
  wire u_wb2sdrc_u_wrdatafifo_rd_ptr_3__FF_INPUT;
  wire u_wb2sdrc_u_wrdatafifo_sync_rd_ptr_0_0_;
  wire u_wb2sdrc_u_wrdatafifo_sync_rd_ptr_0_1_;
  wire u_wb2sdrc_u_wrdatafifo_sync_rd_ptr_0_2_;
  wire u_wb2sdrc_u_wrdatafifo_sync_rd_ptr_0_3_;
  wire u_wb2sdrc_u_wrdatafifo_sync_rd_ptr_1_0_;
  wire u_wb2sdrc_u_wrdatafifo_sync_rd_ptr_1_1_;
  wire u_wb2sdrc_u_wrdatafifo_sync_rd_ptr_1_2_;
  wire u_wb2sdrc_u_wrdatafifo_sync_rd_ptr_1_3_;
  wire u_wb2sdrc_u_wrdatafifo_wr_data_32_;
  wire u_wb2sdrc_u_wrdatafifo_wr_data_33_;
  wire u_wb2sdrc_u_wrdatafifo_wr_data_34_;
  wire u_wb2sdrc_u_wrdatafifo_wr_data_35_;
  wire u_wb2sdrc_u_wrdatafifo_wr_en;
  wire u_wb2sdrc_u_wrdatafifo_wr_ptr_0_;
  wire u_wb2sdrc_u_wrdatafifo_wr_ptr_0__FF_INPUT;
  wire u_wb2sdrc_u_wrdatafifo_wr_ptr_1_;
  wire u_wb2sdrc_u_wrdatafifo_wr_ptr_1__FF_INPUT;
  wire u_wb2sdrc_u_wrdatafifo_wr_ptr_2_;
  wire u_wb2sdrc_u_wrdatafifo_wr_ptr_2__FF_INPUT;
  wire u_wb2sdrc_u_wrdatafifo_wr_ptr_3_;
  wire u_wb2sdrc_u_wrdatafifo_wr_ptr_3__FF_INPUT;
  output wb_ack_o;
  input \wb_addr_i[0] ;
  input \wb_addr_i[10] ;
  input \wb_addr_i[11] ;
  input \wb_addr_i[12] ;
  input \wb_addr_i[13] ;
  input \wb_addr_i[14] ;
  input \wb_addr_i[15] ;
  input \wb_addr_i[16] ;
  input \wb_addr_i[17] ;
  input \wb_addr_i[18] ;
  input \wb_addr_i[19] ;
  input \wb_addr_i[1] ;
  input \wb_addr_i[20] ;
  input \wb_addr_i[21] ;
  input \wb_addr_i[22] ;
  input \wb_addr_i[23] ;
  input \wb_addr_i[24] ;
  input \wb_addr_i[25] ;
  input \wb_addr_i[2] ;
  input \wb_addr_i[3] ;
  input \wb_addr_i[4] ;
  input \wb_addr_i[5] ;
  input \wb_addr_i[6] ;
  input \wb_addr_i[7] ;
  input \wb_addr_i[8] ;
  input \wb_addr_i[9] ;
  input wb_clk_i;
  wire wb_clk_i_bF_buf0;
  wire wb_clk_i_bF_buf1;
  wire wb_clk_i_bF_buf10;
  wire wb_clk_i_bF_buf11;
  wire wb_clk_i_bF_buf12;
  wire wb_clk_i_bF_buf13;
  wire wb_clk_i_bF_buf14;
  wire wb_clk_i_bF_buf15;
  wire wb_clk_i_bF_buf16;
  wire wb_clk_i_bF_buf17;
  wire wb_clk_i_bF_buf18;
  wire wb_clk_i_bF_buf19;
  wire wb_clk_i_bF_buf2;
  wire wb_clk_i_bF_buf20;
  wire wb_clk_i_bF_buf21;
  wire wb_clk_i_bF_buf22;
  wire wb_clk_i_bF_buf23;
  wire wb_clk_i_bF_buf24;
  wire wb_clk_i_bF_buf25;
  wire wb_clk_i_bF_buf26;
  wire wb_clk_i_bF_buf27;
  wire wb_clk_i_bF_buf28;
  wire wb_clk_i_bF_buf29;
  wire wb_clk_i_bF_buf3;
  wire wb_clk_i_bF_buf30;
  wire wb_clk_i_bF_buf31;
  wire wb_clk_i_bF_buf32;
  wire wb_clk_i_bF_buf33;
  wire wb_clk_i_bF_buf34;
  wire wb_clk_i_bF_buf35;
  wire wb_clk_i_bF_buf36;
  wire wb_clk_i_bF_buf37;
  wire wb_clk_i_bF_buf38;
  wire wb_clk_i_bF_buf39;
  wire wb_clk_i_bF_buf4;
  wire wb_clk_i_bF_buf40;
  wire wb_clk_i_bF_buf41;
  wire wb_clk_i_bF_buf42;
  wire wb_clk_i_bF_buf43;
  wire wb_clk_i_bF_buf44;
  wire wb_clk_i_bF_buf45;
  wire wb_clk_i_bF_buf46;
  wire wb_clk_i_bF_buf47;
  wire wb_clk_i_bF_buf48;
  wire wb_clk_i_bF_buf49;
  wire wb_clk_i_bF_buf5;
  wire wb_clk_i_bF_buf50;
  wire wb_clk_i_bF_buf51;
  wire wb_clk_i_bF_buf52;
  wire wb_clk_i_bF_buf53;
  wire wb_clk_i_bF_buf54;
  wire wb_clk_i_bF_buf55;
  wire wb_clk_i_bF_buf56;
  wire wb_clk_i_bF_buf57;
  wire wb_clk_i_bF_buf58;
  wire wb_clk_i_bF_buf59;
  wire wb_clk_i_bF_buf6;
  wire wb_clk_i_bF_buf7;
  wire wb_clk_i_bF_buf8;
  wire wb_clk_i_bF_buf9;
  wire wb_clk_i_hier0_bF_buf0;
  wire wb_clk_i_hier0_bF_buf1;
  wire wb_clk_i_hier0_bF_buf2;
  wire wb_clk_i_hier0_bF_buf3;
  wire wb_clk_i_hier0_bF_buf4;
  wire wb_clk_i_hier0_bF_buf5;
  wire wb_clk_i_hier0_bF_buf6;
  input \wb_cti_i[0] ;
  input \wb_cti_i[1] ;
  input \wb_cti_i[2] ;
  input wb_cyc_i;
  input \wb_dat_i[0] ;
  input \wb_dat_i[10] ;
  input \wb_dat_i[11] ;
  input \wb_dat_i[12] ;
  input \wb_dat_i[13] ;
  input \wb_dat_i[14] ;
  input \wb_dat_i[15] ;
  input \wb_dat_i[16] ;
  input \wb_dat_i[17] ;
  input \wb_dat_i[18] ;
  input \wb_dat_i[19] ;
  input \wb_dat_i[1] ;
  input \wb_dat_i[20] ;
  input \wb_dat_i[21] ;
  input \wb_dat_i[22] ;
  input \wb_dat_i[23] ;
  input \wb_dat_i[24] ;
  input \wb_dat_i[25] ;
  input \wb_dat_i[26] ;
  input \wb_dat_i[27] ;
  input \wb_dat_i[28] ;
  input \wb_dat_i[29] ;
  input \wb_dat_i[2] ;
  input \wb_dat_i[30] ;
  input \wb_dat_i[31] ;
  input \wb_dat_i[3] ;
  input \wb_dat_i[4] ;
  input \wb_dat_i[5] ;
  input \wb_dat_i[6] ;
  input \wb_dat_i[7] ;
  input \wb_dat_i[8] ;
  input \wb_dat_i[9] ;
  output \wb_dat_o[0] ;
  output \wb_dat_o[10] ;
  output \wb_dat_o[11] ;
  output \wb_dat_o[12] ;
  output \wb_dat_o[13] ;
  output \wb_dat_o[14] ;
  output \wb_dat_o[15] ;
  output \wb_dat_o[16] ;
  output \wb_dat_o[17] ;
  output \wb_dat_o[18] ;
  output \wb_dat_o[19] ;
  output \wb_dat_o[1] ;
  output \wb_dat_o[20] ;
  output \wb_dat_o[21] ;
  output \wb_dat_o[22] ;
  output \wb_dat_o[23] ;
  output \wb_dat_o[24] ;
  output \wb_dat_o[25] ;
  output \wb_dat_o[26] ;
  output \wb_dat_o[27] ;
  output \wb_dat_o[28] ;
  output \wb_dat_o[29] ;
  output \wb_dat_o[2] ;
  output \wb_dat_o[30] ;
  output \wb_dat_o[31] ;
  output \wb_dat_o[3] ;
  output \wb_dat_o[4] ;
  output \wb_dat_o[5] ;
  output \wb_dat_o[6] ;
  output \wb_dat_o[7] ;
  output \wb_dat_o[8] ;
  output \wb_dat_o[9] ;
  input wb_rst_i;
  input \wb_sel_i[0] ;
  input \wb_sel_i[1] ;
  input \wb_sel_i[2] ;
  input \wb_sel_i[3] ;
  input wb_stb_i;
  input wb_we_i;
  AND2X2 AND2X2_1 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_tras_ok), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_tras_ok), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n204_1) );
  AND2X2 AND2X2_10 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_cmd_1_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n221_1) );
  AND2X2 AND2X2_100 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_4_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n406) );
  AND2X2 AND2X2_1000 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n257), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n259_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n260) );
  AND2X2 AND2X2_1001 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n260), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n255_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n261_1) );
  AND2X2 AND2X2_1002 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n263), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n265_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n266) );
  AND2X2 AND2X2_1003 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n268_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n270_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n271_1) );
  AND2X2 AND2X2_1004 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n266), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n271_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n272) );
  AND2X2 AND2X2_1005 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n272), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n261_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n273_1) );
  AND2X2 AND2X2_1006 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n275), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n277_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n278) );
  AND2X2 AND2X2_1007 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n280_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n282_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n283_1) );
  AND2X2 AND2X2_1008 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n278), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n283_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n284_1) );
  AND2X2 AND2X2_1009 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n286_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n288_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n289) );
  AND2X2 AND2X2_101 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n408), .B(u_sdrc_core_u_bank_ctl__abc_21249_n407), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n409) );
  AND2X2 AND2X2_1010 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n291_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n293), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n294_1) );
  AND2X2 AND2X2_1011 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n289), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n294_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n295_1) );
  AND2X2 AND2X2_1012 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n284_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n295_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n296_1) );
  AND2X2 AND2X2_1013 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n296_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n273_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n297) );
  AND2X2 AND2X2_1014 ( .A(u_sdrc_core_r2b_raddr_10_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_10_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n298_1) );
  AND2X2 AND2X2_1015 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n299_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n300_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n301) );
  AND2X2 AND2X2_1016 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_8_), .B(u_sdrc_core_r2b_raddr_8_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n303_1) );
  AND2X2 AND2X2_1017 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n304_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n305), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n306_1) );
  AND2X2 AND2X2_1018 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n302_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n307_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n308_1) );
  AND2X2 AND2X2_1019 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n310_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n312_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n313) );
  AND2X2 AND2X2_102 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n410), .B(u_sdrc_core_u_bank_ctl__abc_21249_n411), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n412) );
  AND2X2 AND2X2_1020 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n315_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n317), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n318_1) );
  AND2X2 AND2X2_1021 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n313), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n318_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n319_1) );
  AND2X2 AND2X2_1022 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n321), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n323_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n324_1) );
  AND2X2 AND2X2_1023 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n326_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_valid), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n327_1) );
  AND2X2 AND2X2_1024 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n324_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n327_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n328_1) );
  AND2X2 AND2X2_1025 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n319_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n328_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n329) );
  AND2X2 AND2X2_1026 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n329), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n308_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n330_1) );
  AND2X2 AND2X2_1027 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n297), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n330_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n331_1) );
  AND2X2 AND2X2_1028 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n332_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n253_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n333) );
  AND2X2 AND2X2_1029 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n250_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_prech_page_closed), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n335) );
  AND2X2 AND2X2_103 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n412), .B(u_sdrc_core_u_bank_ctl__abc_21249_n227_bF_buf2), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n413) );
  AND2X2 AND2X2_1030 ( .A(sdram_resetn_bF_buf9), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_4_bF_buf3), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n337) );
  AND2X2 AND2X2_1031 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n337), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n336), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n338_1) );
  AND2X2 AND2X2_1032 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n338_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_x2b_ack), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n339_1) );
  AND2X2 AND2X2_1033 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n339_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_sdr_dma_last), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n340) );
  AND2X2 AND2X2_1034 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n250_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_2_bF_buf3), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n342) );
  AND2X2 AND2X2_1035 ( .A(sdram_resetn_bF_buf8), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_x2b_ack), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n343_1) );
  AND2X2 AND2X2_1036 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n343_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_3_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n344_1) );
  AND2X2 AND2X2_1037 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n337), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_refresh), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n345) );
  AND2X2 AND2X2_1038 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n343_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_2_bF_buf2), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n348_1) );
  AND2X2 AND2X2_1039 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n338_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n249_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n349_1) );
  AND2X2 AND2X2_104 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_5_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n415) );
  AND2X2 AND2X2_1040 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n331_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n253_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n351) );
  AND2X2 AND2X2_1041 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n339_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n353_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n354_1) );
  AND2X2 AND2X2_1042 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n356), .B(sdram_resetn_bF_buf7), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n357) );
  AND2X2 AND2X2_1043 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n355), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n358_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n359_1) );
  AND2X2 AND2X2_1044 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n360), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_0_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n361) );
  AND2X2 AND2X2_1045 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_4_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_write), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n364_1) );
  AND2X2 AND2X2_1046 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n369_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n367), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n370) );
  AND2X2 AND2X2_1047 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n370), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n371) );
  AND2X2 AND2X2_1048 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n371), .B(u_sdrc_core_r2b_write), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n372) );
  AND2X2 AND2X2_1049 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n331_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n372), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n373_1) );
  AND2X2 AND2X2_105 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n417), .B(u_sdrc_core_u_bank_ctl__abc_21249_n416), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n418) );
  AND2X2 AND2X2_1050 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n374_1), .B(sdram_resetn_bF_buf6), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_cmd_r_0__FF_INPUT) );
  AND2X2 AND2X2_1051 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n371), .B(sdram_resetn_bF_buf5), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n376) );
  AND2X2 AND2X2_1052 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n331_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n376), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n377) );
  AND2X2 AND2X2_1053 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n381), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_cmd_0_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n382) );
  AND2X2 AND2X2_1054 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n383_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n386_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n387_1) );
  AND2X2 AND2X2_1055 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n387_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n379_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n388) );
  AND2X2 AND2X2_1056 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n382), .B(\cfg_sdr_tras_d[0] ), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n389) );
  AND2X2 AND2X2_1057 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n390), .B(sdram_resetn_bF_buf4), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_tras_cntr_0__FF_INPUT) );
  AND2X2 AND2X2_1058 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n382), .B(\cfg_sdr_tras_d[1] ), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n392_1) );
  AND2X2 AND2X2_1059 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_tras_cntr_0_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_tras_cntr_1_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n394_1) );
  AND2X2 AND2X2_106 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n419), .B(u_sdrc_core_u_bank_ctl__abc_21249_n420), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n421) );
  AND2X2 AND2X2_1060 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n387_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n395_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n396_1) );
  AND2X2 AND2X2_1061 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n397_1), .B(sdram_resetn_bF_buf3), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_tras_cntr_1__FF_INPUT) );
  AND2X2 AND2X2_1062 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n382), .B(\cfg_sdr_tras_d[2] ), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n399_1) );
  AND2X2 AND2X2_1063 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n384_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_tras_cntr_2_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n401_1) );
  AND2X2 AND2X2_1064 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n387_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n402_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n403_1) );
  AND2X2 AND2X2_1065 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n404_1), .B(sdram_resetn_bF_buf2), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_tras_cntr_2__FF_INPUT) );
  AND2X2 AND2X2_1066 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n385), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_tras_cntr_3_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n406_1) );
  AND2X2 AND2X2_1067 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n408_1), .B(sdram_resetn_bF_buf1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n409_1) );
  AND2X2 AND2X2_1068 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n409_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n407_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_tras_cntr_3__FF_INPUT) );
  AND2X2 AND2X2_1069 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n415_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n413_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n416) );
  AND2X2 AND2X2_107 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n421), .B(u_sdrc_core_u_bank_ctl__abc_21249_n227_bF_buf1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n422) );
  AND2X2 AND2X2_1070 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n417_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n418), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n419_1) );
  AND2X2 AND2X2_1071 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n421), .B(sdram_resetn_bF_buf0), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n422) );
  AND2X2 AND2X2_1072 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n420_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n422), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_timer0_0__FF_INPUT) );
  AND2X2 AND2X2_1073 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_timer0_1_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_timer0_0_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n426) );
  AND2X2 AND2X2_1074 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n383_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n428_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n429) );
  AND2X2 AND2X2_1075 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n429), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n427_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n430) );
  AND2X2 AND2X2_1076 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n381), .B(\cfg_sdr_trcd_d[1] ), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n431_1) );
  AND2X2 AND2X2_1077 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n434_1), .B(sdram_resetn_bF_buf49), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n435_1) );
  AND2X2 AND2X2_1078 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n433), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n435_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_timer0_1__FF_INPUT) );
  AND2X2 AND2X2_1079 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n424), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_timer0_2_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n439_1) );
  AND2X2 AND2X2_108 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_6_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n424) );
  AND2X2 AND2X2_1080 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n429), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n440_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n441) );
  AND2X2 AND2X2_1081 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n381), .B(\cfg_sdr_trcd_d[2] ), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n442) );
  AND2X2 AND2X2_1082 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n445_1), .B(sdram_resetn_bF_buf48), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n446_1) );
  AND2X2 AND2X2_1083 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n444_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n446_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_timer0_2__FF_INPUT) );
  AND2X2 AND2X2_1084 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n437_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_timer0_3_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n448_1) );
  AND2X2 AND2X2_1085 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n449_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n450), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n451) );
  AND2X2 AND2X2_1086 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n453_1), .B(sdram_resetn_bF_buf47), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n454) );
  AND2X2 AND2X2_1087 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n452), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n454), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_timer0_3__FF_INPUT) );
  AND2X2 AND2X2_1088 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n253_1), .B(u_sdrc_core_r2b_len_0_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n473) );
  AND2X2 AND2X2_1089 ( .A(sdram_resetn_bF_buf46), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_0_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n474) );
  AND2X2 AND2X2_109 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n426), .B(u_sdrc_core_u_bank_ctl__abc_21249_n425), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n427) );
  AND2X2 AND2X2_1090 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf5), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n474), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n475) );
  AND2X2 AND2X2_1091 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n253_1), .B(u_sdrc_core_r2b_len_1_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n477) );
  AND2X2 AND2X2_1092 ( .A(sdram_resetn_bF_buf45), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_1_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n478) );
  AND2X2 AND2X2_1093 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n478), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n479) );
  AND2X2 AND2X2_1094 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n253_1), .B(u_sdrc_core_r2b_len_2_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n481) );
  AND2X2 AND2X2_1095 ( .A(sdram_resetn_bF_buf44), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_2_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n482) );
  AND2X2 AND2X2_1096 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n482), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n483) );
  AND2X2 AND2X2_1097 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n253_1), .B(u_sdrc_core_r2b_len_3_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n485) );
  AND2X2 AND2X2_1098 ( .A(sdram_resetn_bF_buf43), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_3_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n486) );
  AND2X2 AND2X2_1099 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n486), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n487) );
  AND2X2 AND2X2_11 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n224_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n222), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n225_1) );
  AND2X2 AND2X2_110 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n428), .B(u_sdrc_core_u_bank_ctl__abc_21249_n429), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n430) );
  AND2X2 AND2X2_1100 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n253_1), .B(u_sdrc_core_r2b_len_4_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n489) );
  AND2X2 AND2X2_1101 ( .A(sdram_resetn_bF_buf42), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_4_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n490) );
  AND2X2 AND2X2_1102 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n490), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n491) );
  AND2X2 AND2X2_1103 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n253_1), .B(u_sdrc_core_r2b_len_5_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n493) );
  AND2X2 AND2X2_1104 ( .A(sdram_resetn_bF_buf41), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_5_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n494) );
  AND2X2 AND2X2_1105 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n494), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n495) );
  AND2X2 AND2X2_1106 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n253_1), .B(u_sdrc_core_r2b_len_6_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n497) );
  AND2X2 AND2X2_1107 ( .A(sdram_resetn_bF_buf40), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_6_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n498) );
  AND2X2 AND2X2_1108 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf5), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n498), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n499) );
  AND2X2 AND2X2_1109 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_0_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n501) );
  AND2X2 AND2X2_111 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n430), .B(u_sdrc_core_u_bank_ctl__abc_21249_n227_bF_buf0), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n431) );
  AND2X2 AND2X2_1110 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf1), .B(u_sdrc_core_r2b_raddr_0_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n502) );
  AND2X2 AND2X2_1111 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n503), .B(sdram_resetn_bF_buf39), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_0__FF_INPUT) );
  AND2X2 AND2X2_1112 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_1_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n505) );
  AND2X2 AND2X2_1113 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf0), .B(u_sdrc_core_r2b_raddr_1_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n506) );
  AND2X2 AND2X2_1114 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n507), .B(sdram_resetn_bF_buf38), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_1__FF_INPUT) );
  AND2X2 AND2X2_1115 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_2_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n509) );
  AND2X2 AND2X2_1116 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf4), .B(u_sdrc_core_r2b_raddr_2_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n510) );
  AND2X2 AND2X2_1117 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n511), .B(sdram_resetn_bF_buf37), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_2__FF_INPUT) );
  AND2X2 AND2X2_1118 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_3_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n513) );
  AND2X2 AND2X2_1119 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf3), .B(u_sdrc_core_r2b_raddr_3_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n514) );
  AND2X2 AND2X2_112 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_7_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n433) );
  AND2X2 AND2X2_1120 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n515), .B(sdram_resetn_bF_buf36), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_3__FF_INPUT) );
  AND2X2 AND2X2_1121 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_4_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n517) );
  AND2X2 AND2X2_1122 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf2), .B(u_sdrc_core_r2b_raddr_4_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n518) );
  AND2X2 AND2X2_1123 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n519), .B(sdram_resetn_bF_buf35), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_4__FF_INPUT) );
  AND2X2 AND2X2_1124 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf5), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_5_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n521) );
  AND2X2 AND2X2_1125 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf1), .B(u_sdrc_core_r2b_raddr_5_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n522) );
  AND2X2 AND2X2_1126 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n523), .B(sdram_resetn_bF_buf34), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_5__FF_INPUT) );
  AND2X2 AND2X2_1127 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_6_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n525) );
  AND2X2 AND2X2_1128 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf0), .B(u_sdrc_core_r2b_raddr_6_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n526) );
  AND2X2 AND2X2_1129 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n527), .B(sdram_resetn_bF_buf33), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_6__FF_INPUT) );
  AND2X2 AND2X2_113 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n435), .B(u_sdrc_core_u_bank_ctl__abc_21249_n434), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n436) );
  AND2X2 AND2X2_1130 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_7_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n529) );
  AND2X2 AND2X2_1131 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf4), .B(u_sdrc_core_r2b_raddr_7_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n530) );
  AND2X2 AND2X2_1132 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n531), .B(sdram_resetn_bF_buf32), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_7__FF_INPUT) );
  AND2X2 AND2X2_1133 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_8_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n533) );
  AND2X2 AND2X2_1134 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf3), .B(u_sdrc_core_r2b_raddr_8_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n534) );
  AND2X2 AND2X2_1135 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n535), .B(sdram_resetn_bF_buf31), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_8__FF_INPUT) );
  AND2X2 AND2X2_1136 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_9_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n537) );
  AND2X2 AND2X2_1137 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf2), .B(u_sdrc_core_r2b_raddr_9_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n538) );
  AND2X2 AND2X2_1138 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n539), .B(sdram_resetn_bF_buf30), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_9__FF_INPUT) );
  AND2X2 AND2X2_1139 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_10_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n541) );
  AND2X2 AND2X2_114 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n437), .B(u_sdrc_core_u_bank_ctl__abc_21249_n438), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n439) );
  AND2X2 AND2X2_1140 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf1), .B(u_sdrc_core_r2b_raddr_10_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n542) );
  AND2X2 AND2X2_1141 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n543), .B(sdram_resetn_bF_buf29), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_10__FF_INPUT) );
  AND2X2 AND2X2_1142 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf5), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_11_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n545) );
  AND2X2 AND2X2_1143 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf0), .B(u_sdrc_core_r2b_raddr_11_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n546) );
  AND2X2 AND2X2_1144 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n547), .B(sdram_resetn_bF_buf28), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_11__FF_INPUT) );
  AND2X2 AND2X2_1145 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_12_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n549) );
  AND2X2 AND2X2_1146 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf4), .B(u_sdrc_core_r2b_raddr_12_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n550) );
  AND2X2 AND2X2_1147 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n551), .B(sdram_resetn_bF_buf27), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_12__FF_INPUT) );
  AND2X2 AND2X2_1148 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_0_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n553) );
  AND2X2 AND2X2_1149 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf3), .B(u_sdrc_core_r2b_caddr_0_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n554) );
  AND2X2 AND2X2_115 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n439), .B(u_sdrc_core_u_bank_ctl__abc_21249_n227_bF_buf3), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n440) );
  AND2X2 AND2X2_1150 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n555), .B(sdram_resetn_bF_buf26), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_0__FF_INPUT) );
  AND2X2 AND2X2_1151 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_1_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n557) );
  AND2X2 AND2X2_1152 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf2), .B(u_sdrc_core_r2b_caddr_1_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n558) );
  AND2X2 AND2X2_1153 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n559), .B(sdram_resetn_bF_buf25), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_1__FF_INPUT) );
  AND2X2 AND2X2_1154 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_2_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n561) );
  AND2X2 AND2X2_1155 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf1), .B(u_sdrc_core_r2b_caddr_2_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n562) );
  AND2X2 AND2X2_1156 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n563), .B(sdram_resetn_bF_buf24), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_2__FF_INPUT) );
  AND2X2 AND2X2_1157 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_3_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n565) );
  AND2X2 AND2X2_1158 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf0), .B(u_sdrc_core_r2b_caddr_3_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n566) );
  AND2X2 AND2X2_1159 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n567), .B(sdram_resetn_bF_buf23), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_3__FF_INPUT) );
  AND2X2 AND2X2_116 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_8_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n442) );
  AND2X2 AND2X2_1160 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf5), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_4_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n569) );
  AND2X2 AND2X2_1161 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf4), .B(u_sdrc_core_r2b_caddr_4_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n570) );
  AND2X2 AND2X2_1162 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n571), .B(sdram_resetn_bF_buf22), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_4__FF_INPUT) );
  AND2X2 AND2X2_1163 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_5_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n573) );
  AND2X2 AND2X2_1164 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf3), .B(u_sdrc_core_r2b_caddr_5_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n574) );
  AND2X2 AND2X2_1165 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n575), .B(sdram_resetn_bF_buf21), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_5__FF_INPUT) );
  AND2X2 AND2X2_1166 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_6_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n577) );
  AND2X2 AND2X2_1167 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf2), .B(u_sdrc_core_r2b_caddr_6_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n578) );
  AND2X2 AND2X2_1168 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n579), .B(sdram_resetn_bF_buf20), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_6__FF_INPUT) );
  AND2X2 AND2X2_1169 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_7_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n581) );
  AND2X2 AND2X2_117 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n444), .B(u_sdrc_core_u_bank_ctl__abc_21249_n443), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n445) );
  AND2X2 AND2X2_1170 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf1), .B(u_sdrc_core_r2b_caddr_7_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n582) );
  AND2X2 AND2X2_1171 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n583), .B(sdram_resetn_bF_buf19), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_7__FF_INPUT) );
  AND2X2 AND2X2_1172 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_8_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n585) );
  AND2X2 AND2X2_1173 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf0), .B(u_sdrc_core_r2b_caddr_8_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n586) );
  AND2X2 AND2X2_1174 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n587), .B(sdram_resetn_bF_buf18), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_8__FF_INPUT) );
  AND2X2 AND2X2_1175 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_9_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n589) );
  AND2X2 AND2X2_1176 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf4), .B(u_sdrc_core_r2b_caddr_9_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n590) );
  AND2X2 AND2X2_1177 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n591), .B(sdram_resetn_bF_buf17), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_9__FF_INPUT) );
  AND2X2 AND2X2_1178 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf5), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_10_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n593) );
  AND2X2 AND2X2_1179 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf3), .B(u_sdrc_core_r2b_caddr_10_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n594) );
  AND2X2 AND2X2_118 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n446), .B(u_sdrc_core_u_bank_ctl__abc_21249_n447), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n448) );
  AND2X2 AND2X2_1180 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n595), .B(sdram_resetn_bF_buf16), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_10__FF_INPUT) );
  AND2X2 AND2X2_1181 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_11_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n597) );
  AND2X2 AND2X2_1182 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf2), .B(1'b0), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n598) );
  AND2X2 AND2X2_1183 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n599), .B(sdram_resetn_bF_buf15), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_11__FF_INPUT) );
  AND2X2 AND2X2_1184 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_12_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n601) );
  AND2X2 AND2X2_1185 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf1), .B(1'b0), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n602) );
  AND2X2 AND2X2_1186 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n603), .B(sdram_resetn_bF_buf14), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_12__FF_INPUT) );
  AND2X2 AND2X2_1187 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_4_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_0_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n605) );
  AND2X2 AND2X2_1188 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_0_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n607) );
  AND2X2 AND2X2_1189 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n609), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n610), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_0__FF_INPUT) );
  AND2X2 AND2X2_119 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n448), .B(u_sdrc_core_u_bank_ctl__abc_21249_n227_bF_buf2), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n449) );
  AND2X2 AND2X2_1190 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_4_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_1_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n612) );
  AND2X2 AND2X2_1191 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_1_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n613) );
  AND2X2 AND2X2_1192 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n615), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n616), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_1__FF_INPUT) );
  AND2X2 AND2X2_1193 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_4_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_2_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n618) );
  AND2X2 AND2X2_1194 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_2_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n619) );
  AND2X2 AND2X2_1195 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n621), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n622), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_2__FF_INPUT) );
  AND2X2 AND2X2_1196 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_4_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_3_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n624) );
  AND2X2 AND2X2_1197 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_3_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n625) );
  AND2X2 AND2X2_1198 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n627), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n628), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_3__FF_INPUT) );
  AND2X2 AND2X2_1199 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_4_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_4_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n630) );
  AND2X2 AND2X2_12 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n228_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n227_bF_buf3), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n229) );
  AND2X2 AND2X2_120 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_9_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n451) );
  AND2X2 AND2X2_1200 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_4_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n631) );
  AND2X2 AND2X2_1201 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n633), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n634), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_4__FF_INPUT) );
  AND2X2 AND2X2_1202 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_4_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_5_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n636) );
  AND2X2 AND2X2_1203 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_5_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n637) );
  AND2X2 AND2X2_1204 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n639), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n640), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_5__FF_INPUT) );
  AND2X2 AND2X2_1205 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_4_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_6_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n642) );
  AND2X2 AND2X2_1206 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_6_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n643) );
  AND2X2 AND2X2_1207 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n645), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n646), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_6__FF_INPUT) );
  AND2X2 AND2X2_1208 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_4_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_7_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n648) );
  AND2X2 AND2X2_1209 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_7_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n649) );
  AND2X2 AND2X2_121 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n453), .B(u_sdrc_core_u_bank_ctl__abc_21249_n452), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n454) );
  AND2X2 AND2X2_1210 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n651), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n652), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_7__FF_INPUT) );
  AND2X2 AND2X2_1211 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_4_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_8_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n654) );
  AND2X2 AND2X2_1212 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_8_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n655) );
  AND2X2 AND2X2_1213 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n657), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n658), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_8__FF_INPUT) );
  AND2X2 AND2X2_1214 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_4_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_9_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n660) );
  AND2X2 AND2X2_1215 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_9_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n661) );
  AND2X2 AND2X2_1216 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n663), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n664), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_9__FF_INPUT) );
  AND2X2 AND2X2_1217 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_4_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_10_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n666) );
  AND2X2 AND2X2_1218 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n370), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_10_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n667) );
  AND2X2 AND2X2_1219 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n669), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n670), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_10__FF_INPUT) );
  AND2X2 AND2X2_122 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n455), .B(u_sdrc_core_u_bank_ctl__abc_21249_n456), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n457) );
  AND2X2 AND2X2_1220 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_4_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_11_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n672) );
  AND2X2 AND2X2_1221 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_11_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n673) );
  AND2X2 AND2X2_1222 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n675), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n676), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_11__FF_INPUT) );
  AND2X2 AND2X2_1223 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_4_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_12_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n678) );
  AND2X2 AND2X2_1224 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n370), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_12_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n679) );
  AND2X2 AND2X2_1225 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n681), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n682), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_12__FF_INPUT) );
  AND2X2 AND2X2_1226 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n689), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n688), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_last) );
  AND2X2 AND2X2_1227 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n704), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n703), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_len_0_) );
  AND2X2 AND2X2_1228 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n707), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n706), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_len_1_) );
  AND2X2 AND2X2_1229 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n710), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n709), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_len_2_) );
  AND2X2 AND2X2_123 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n457), .B(u_sdrc_core_u_bank_ctl__abc_21249_n227_bF_buf1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n458) );
  AND2X2 AND2X2_1230 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n713), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n712), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_len_3_) );
  AND2X2 AND2X2_1231 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n716), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n715), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_len_4_) );
  AND2X2 AND2X2_1232 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n719), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n718), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_len_5_) );
  AND2X2 AND2X2_1233 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n722), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n721), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_len_6_) );
  AND2X2 AND2X2_1234 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n725), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n724), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_wrap) );
  AND2X2 AND2X2_1235 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_x2b_pre_ok_t), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_tras_ok), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n727) );
  AND2X2 AND2X2_1236 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n368_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n727), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n728) );
  AND2X2 AND2X2_1237 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_2_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_x2b_act_ok_t), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n729) );
  AND2X2 AND2X2_1238 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_4_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_r), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n733) );
  AND2X2 AND2X2_1239 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n732), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n733), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n734) );
  AND2X2 AND2X2_124 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_10_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n460) );
  AND2X2 AND2X2_1240 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n734), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n731), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n735) );
  AND2X2 AND2X2_1241 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n736), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_timer0_tc), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n737) );
  AND2X2 AND2X2_1242 ( .A(sdram_resetn_bF_buf13), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_wrok), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_x2b_wrok_r_FF_INPUT) );
  AND2X2 AND2X2_1243 ( .A(sdram_resetn_bF_buf12), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf2), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_r_FF_INPUT) );
  AND2X2 AND2X2_1244 ( .A(sdram_resetn_bF_buf11), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_rdok), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_x2b_rdok_r_FF_INPUT) );
  AND2X2 AND2X2_1245 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n380), .B(sdram_resetn_bF_buf10), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n743) );
  AND2X2 AND2X2_1246 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n742), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n743), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_timer0_tc_r_FF_INPUT) );
  AND2X2 AND2X2_1247 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n745), .B(sdram_resetn_bF_buf9), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_tras_ok_r_FF_INPUT) );
  AND2X2 AND2X2_1248 ( .A(sdram_resetn_bF_buf8), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_pre_ok), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_x2b_pre_ok_r_FF_INPUT) );
  AND2X2 AND2X2_1249 ( .A(sdram_resetn_bF_buf7), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_act_ok), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_x2b_act_ok_r_FF_INPUT) );
  AND2X2 AND2X2_125 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n462), .B(u_sdrc_core_u_bank_ctl__abc_21249_n461), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n463) );
  AND2X2 AND2X2_1250 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n357), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n336), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n750) );
  AND2X2 AND2X2_1251 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n749), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n750), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_valid_FF_INPUT) );
  AND2X2 AND2X2_1252 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_last), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n756) );
  AND2X2 AND2X2_1253 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf0), .B(u_sdrc_core_r2b_last), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n757) );
  AND2X2 AND2X2_1254 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n758), .B(sdram_resetn_bF_buf6), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_l_last_FF_INPUT) );
  AND2X2 AND2X2_1255 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_wrap), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n760) );
  AND2X2 AND2X2_1256 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf4), .B(u_sdrc_core_r2b_wrap), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n761) );
  AND2X2 AND2X2_1257 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n762), .B(sdram_resetn_bF_buf5), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_l_wrap_FF_INPUT) );
  AND2X2 AND2X2_1258 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_write), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n764) );
  AND2X2 AND2X2_1259 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf3), .B(u_sdrc_core_r2b_write), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n765) );
  AND2X2 AND2X2_126 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n464), .B(u_sdrc_core_u_bank_ctl__abc_21249_n465), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n466) );
  AND2X2 AND2X2_1260 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n766), .B(sdram_resetn_bF_buf4), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_l_write_FF_INPUT) );
  AND2X2 AND2X2_1261 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf5), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_sdr_dma_last), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n768) );
  AND2X2 AND2X2_1262 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf2), .B(1'b0), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n769) );
  AND2X2 AND2X2_1263 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n770), .B(sdram_resetn_bF_buf3), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_l_sdr_dma_last_FF_INPUT) );
  AND2X2 AND2X2_1264 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n168_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n169_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n170_1) );
  AND2X2 AND2X2_1265 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n174_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n176_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n177_1) );
  AND2X2 AND2X2_1266 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n177_1), .B(app_wr_data_0_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n178_1) );
  AND2X2 AND2X2_1267 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf2), .B(app_wr_data_8_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n179_1) );
  AND2X2 AND2X2_1268 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n180_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n181_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n182_1) );
  AND2X2 AND2X2_1269 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n169_1), .B(\cfg_sdr_width[0] ), .Y(u_sdrc_core_u_bs_convert__abc_21684_n184_1) );
  AND2X2 AND2X2_127 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n466), .B(u_sdrc_core_u_bank_ctl__abc_21249_n227_bF_buf0), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n467) );
  AND2X2 AND2X2_1270 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf0), .B(u_sdrc_core_u_bs_convert_wr_xfr_count_1_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n187_1) );
  AND2X2 AND2X2_1271 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n187_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n186_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n188_1) );
  AND2X2 AND2X2_1272 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n189_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n185_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n190_1) );
  AND2X2 AND2X2_1273 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n183_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n190_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n191_1) );
  AND2X2 AND2X2_1274 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf4), .B(u_sdrc_core_u_bs_convert__abc_21684_n193_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n194_1) );
  AND2X2 AND2X2_1275 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n194_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n192_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n195_1) );
  AND2X2 AND2X2_1276 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n197_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n172_1), .Y(u_sdrc_core_a2x_wrdt_0_) );
  AND2X2 AND2X2_1277 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n177_1), .B(app_wr_data_1_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n199) );
  AND2X2 AND2X2_1278 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf3), .B(app_wr_data_9_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n200_1) );
  AND2X2 AND2X2_1279 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n201_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n202), .Y(u_sdrc_core_u_bs_convert__abc_21684_n203_1) );
  AND2X2 AND2X2_128 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_11_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n469) );
  AND2X2 AND2X2_1280 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n187_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n205), .Y(u_sdrc_core_u_bs_convert__abc_21684_n206_1) );
  AND2X2 AND2X2_1281 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n207_1), .B(cfg_sdr_width_1_bF_buf4), .Y(u_sdrc_core_u_bs_convert__abc_21684_n208) );
  AND2X2 AND2X2_1282 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n204_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n208), .Y(u_sdrc_core_u_bs_convert__abc_21684_n209_1) );
  AND2X2 AND2X2_1283 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf3), .B(u_sdrc_core_u_bs_convert__abc_21684_n175_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n210_1) );
  AND2X2 AND2X2_1284 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n211), .B(app_wr_data_1_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n212_1) );
  AND2X2 AND2X2_1285 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf1), .B(app_wr_data_17_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n213_1) );
  AND2X2 AND2X2_1286 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf2), .B(u_sdrc_core_u_bs_convert__abc_21684_n213_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n214) );
  AND2X2 AND2X2_1287 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n177_1), .B(app_wr_data_2_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n217) );
  AND2X2 AND2X2_1288 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n218_1), .B(u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf0), .Y(u_sdrc_core_u_bs_convert__abc_21684_n219) );
  AND2X2 AND2X2_1289 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_1_), .B(app_wr_data_18_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n220_1) );
  AND2X2 AND2X2_129 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n471), .B(u_sdrc_core_u_bank_ctl__abc_21249_n470), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n472) );
  AND2X2 AND2X2_1290 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n187_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n223), .Y(u_sdrc_core_u_bs_convert__abc_21684_n224_1) );
  AND2X2 AND2X2_1291 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n225), .B(cfg_sdr_width_1_bF_buf3), .Y(u_sdrc_core_u_bs_convert__abc_21684_n226_1) );
  AND2X2 AND2X2_1292 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n222_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n226_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n227) );
  AND2X2 AND2X2_1293 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n211), .B(app_wr_data_2_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n228_1) );
  AND2X2 AND2X2_1294 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf4), .B(app_wr_data_18_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n229) );
  AND2X2 AND2X2_1295 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf1), .B(u_sdrc_core_u_bs_convert__abc_21684_n229), .Y(u_sdrc_core_u_bs_convert__abc_21684_n230_1) );
  AND2X2 AND2X2_1296 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n177_1), .B(app_wr_data_3_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n233) );
  AND2X2 AND2X2_1297 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n234_1), .B(u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf3), .Y(u_sdrc_core_u_bs_convert__abc_21684_n235_1) );
  AND2X2 AND2X2_1298 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_1_), .B(app_wr_data_19_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n236_1) );
  AND2X2 AND2X2_1299 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n187_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n239), .Y(u_sdrc_core_u_bs_convert__abc_21684_n240) );
  AND2X2 AND2X2_13 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n226_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n229), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n230_1) );
  AND2X2 AND2X2_130 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n473), .B(u_sdrc_core_u_bank_ctl__abc_21249_n474), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n475) );
  AND2X2 AND2X2_1300 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n241), .B(cfg_sdr_width_1_bF_buf2), .Y(u_sdrc_core_u_bs_convert__abc_21684_n242_1) );
  AND2X2 AND2X2_1301 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n238_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n242_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n243) );
  AND2X2 AND2X2_1302 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n211), .B(app_wr_data_3_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n244_1) );
  AND2X2 AND2X2_1303 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf2), .B(app_wr_data_19_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n245) );
  AND2X2 AND2X2_1304 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf0), .B(u_sdrc_core_u_bs_convert__abc_21684_n245), .Y(u_sdrc_core_u_bs_convert__abc_21684_n246_1) );
  AND2X2 AND2X2_1305 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n177_1), .B(app_wr_data_4_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n249) );
  AND2X2 AND2X2_1306 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n173_1), .B(u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n250) );
  AND2X2 AND2X2_1307 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n250), .B(app_wr_data_12_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n251_1) );
  AND2X2 AND2X2_1308 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_1_), .B(app_wr_data_20_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n252) );
  AND2X2 AND2X2_1309 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n187_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n256), .Y(u_sdrc_core_u_bs_convert__abc_21684_n257) );
  AND2X2 AND2X2_131 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n475), .B(u_sdrc_core_u_bank_ctl__abc_21249_n227_bF_buf3), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n476) );
  AND2X2 AND2X2_1310 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n258_1), .B(cfg_sdr_width_1_bF_buf1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n259) );
  AND2X2 AND2X2_1311 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n255_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n259), .Y(u_sdrc_core_u_bs_convert__abc_21684_n260) );
  AND2X2 AND2X2_1312 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n170_1_bF_buf0), .B(app_wr_data_4_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n261) );
  AND2X2 AND2X2_1313 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf5), .B(u_sdrc_core_u_bs_convert__abc_21684_n263), .Y(u_sdrc_core_u_bs_convert__abc_21684_n264) );
  AND2X2 AND2X2_1314 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n264), .B(u_sdrc_core_u_bs_convert__abc_21684_n262), .Y(u_sdrc_core_u_bs_convert__abc_21684_n265) );
  AND2X2 AND2X2_1315 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n177_1), .B(app_wr_data_5_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n268) );
  AND2X2 AND2X2_1316 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n250), .B(app_wr_data_13_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n269) );
  AND2X2 AND2X2_1317 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_1_), .B(app_wr_data_21_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n270_1) );
  AND2X2 AND2X2_1318 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n187_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n274), .Y(u_sdrc_core_u_bs_convert__abc_21684_n275) );
  AND2X2 AND2X2_1319 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n276), .B(u_sdrc_core_u_bs_convert__abc_21684_n185_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n277) );
  AND2X2 AND2X2_132 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_12_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n478) );
  AND2X2 AND2X2_1320 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n273), .B(u_sdrc_core_u_bs_convert__abc_21684_n277), .Y(u_sdrc_core_u_bs_convert__abc_21684_n278) );
  AND2X2 AND2X2_1321 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf4), .B(u_sdrc_core_u_bs_convert__abc_21684_n280), .Y(u_sdrc_core_u_bs_convert__abc_21684_n281) );
  AND2X2 AND2X2_1322 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n281), .B(u_sdrc_core_u_bs_convert__abc_21684_n279_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n282) );
  AND2X2 AND2X2_1323 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n284), .B(u_sdrc_core_u_bs_convert__abc_21684_n285), .Y(u_sdrc_core_a2x_wrdt_5_) );
  AND2X2 AND2X2_1324 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n177_1), .B(app_wr_data_6_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n287) );
  AND2X2 AND2X2_1325 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n250), .B(app_wr_data_14_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n288_1) );
  AND2X2 AND2X2_1326 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_1_), .B(app_wr_data_22_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n289) );
  AND2X2 AND2X2_1327 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n187_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n293), .Y(u_sdrc_core_u_bs_convert__abc_21684_n294) );
  AND2X2 AND2X2_1328 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n295), .B(cfg_sdr_width_1_bF_buf0), .Y(u_sdrc_core_u_bs_convert__abc_21684_n296) );
  AND2X2 AND2X2_1329 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n292), .B(u_sdrc_core_u_bs_convert__abc_21684_n296), .Y(u_sdrc_core_u_bs_convert__abc_21684_n297_1) );
  AND2X2 AND2X2_133 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n480), .B(u_sdrc_core_u_bank_ctl__abc_21249_n479), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n481) );
  AND2X2 AND2X2_1330 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n211), .B(app_wr_data_6_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n298) );
  AND2X2 AND2X2_1331 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf3), .B(app_wr_data_22_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n299) );
  AND2X2 AND2X2_1332 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf3), .B(u_sdrc_core_u_bs_convert__abc_21684_n299), .Y(u_sdrc_core_u_bs_convert__abc_21684_n300) );
  AND2X2 AND2X2_1333 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n177_1), .B(app_wr_data_7_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n303) );
  AND2X2 AND2X2_1334 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n250), .B(app_wr_data_15_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n304) );
  AND2X2 AND2X2_1335 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_1_), .B(app_wr_data_23_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n305) );
  AND2X2 AND2X2_1336 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n187_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n309), .Y(u_sdrc_core_u_bs_convert__abc_21684_n310) );
  AND2X2 AND2X2_1337 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n311), .B(u_sdrc_core_u_bs_convert__abc_21684_n185_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n312) );
  AND2X2 AND2X2_1338 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n308), .B(u_sdrc_core_u_bs_convert__abc_21684_n312), .Y(u_sdrc_core_u_bs_convert__abc_21684_n313) );
  AND2X2 AND2X2_1339 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf2), .B(u_sdrc_core_u_bs_convert__abc_21684_n315_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n316) );
  AND2X2 AND2X2_134 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n482), .B(u_sdrc_core_u_bank_ctl__abc_21249_n483), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n484) );
  AND2X2 AND2X2_1340 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n316), .B(u_sdrc_core_u_bs_convert__abc_21684_n314), .Y(u_sdrc_core_u_bs_convert__abc_21684_n317) );
  AND2X2 AND2X2_1341 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n319), .B(u_sdrc_core_u_bs_convert__abc_21684_n320), .Y(u_sdrc_core_a2x_wrdt_7_) );
  AND2X2 AND2X2_1342 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n211), .B(app_wr_data_8_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n322) );
  AND2X2 AND2X2_1343 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf1), .B(app_wr_data_24_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n323) );
  AND2X2 AND2X2_1344 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf1), .B(u_sdrc_core_u_bs_convert__abc_21684_n323), .Y(u_sdrc_core_u_bs_convert__abc_21684_n324_1) );
  AND2X2 AND2X2_1345 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n211), .B(app_wr_data_9_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n326) );
  AND2X2 AND2X2_1346 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf0), .B(app_wr_data_25_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n327) );
  AND2X2 AND2X2_1347 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf0), .B(u_sdrc_core_u_bs_convert__abc_21684_n327), .Y(u_sdrc_core_u_bs_convert__abc_21684_n328) );
  AND2X2 AND2X2_1348 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n211), .B(app_wr_data_10_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n330) );
  AND2X2 AND2X2_1349 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf4), .B(app_wr_data_26_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n331) );
  AND2X2 AND2X2_135 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n484), .B(u_sdrc_core_u_bank_ctl__abc_21249_n227_bF_buf2), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n485) );
  AND2X2 AND2X2_1350 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf5), .B(u_sdrc_core_u_bs_convert__abc_21684_n331), .Y(u_sdrc_core_u_bs_convert__abc_21684_n332) );
  AND2X2 AND2X2_1351 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n211), .B(app_wr_data_11_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n334) );
  AND2X2 AND2X2_1352 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf3), .B(app_wr_data_27_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n335) );
  AND2X2 AND2X2_1353 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf4), .B(u_sdrc_core_u_bs_convert__abc_21684_n335), .Y(u_sdrc_core_u_bs_convert__abc_21684_n336) );
  AND2X2 AND2X2_1354 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n211), .B(app_wr_data_12_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n338) );
  AND2X2 AND2X2_1355 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf2), .B(app_wr_data_28_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n339) );
  AND2X2 AND2X2_1356 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf3), .B(u_sdrc_core_u_bs_convert__abc_21684_n339), .Y(u_sdrc_core_u_bs_convert__abc_21684_n340) );
  AND2X2 AND2X2_1357 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n211), .B(app_wr_data_13_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n342) );
  AND2X2 AND2X2_1358 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf1), .B(app_wr_data_29_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n343) );
  AND2X2 AND2X2_1359 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf2), .B(u_sdrc_core_u_bs_convert__abc_21684_n343), .Y(u_sdrc_core_u_bs_convert__abc_21684_n344) );
  AND2X2 AND2X2_136 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_len_0_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n487) );
  AND2X2 AND2X2_1360 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n211), .B(app_wr_data_14_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n346) );
  AND2X2 AND2X2_1361 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf0), .B(app_wr_data_30_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n347) );
  AND2X2 AND2X2_1362 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf1), .B(u_sdrc_core_u_bs_convert__abc_21684_n347), .Y(u_sdrc_core_u_bs_convert__abc_21684_n348) );
  AND2X2 AND2X2_1363 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n211), .B(app_wr_data_15_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n350) );
  AND2X2 AND2X2_1364 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf4), .B(app_wr_data_31_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n351) );
  AND2X2 AND2X2_1365 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf0), .B(u_sdrc_core_u_bs_convert__abc_21684_n351), .Y(u_sdrc_core_u_bs_convert__abc_21684_n352) );
  AND2X2 AND2X2_1366 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n177_1), .B(app_wr_en_n_0_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n354) );
  AND2X2 AND2X2_1367 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n250), .B(app_wr_en_n_1_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n355) );
  AND2X2 AND2X2_1368 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_1_), .B(app_wr_en_n_2_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n356) );
  AND2X2 AND2X2_1369 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n187_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n360), .Y(u_sdrc_core_u_bs_convert__abc_21684_n361_1) );
  AND2X2 AND2X2_137 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n489), .B(u_sdrc_core_u_bank_ctl__abc_21249_n488), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n490) );
  AND2X2 AND2X2_1370 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n362), .B(u_sdrc_core_u_bs_convert__abc_21684_n185_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n363) );
  AND2X2 AND2X2_1371 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n359), .B(u_sdrc_core_u_bs_convert__abc_21684_n363), .Y(u_sdrc_core_u_bs_convert__abc_21684_n364) );
  AND2X2 AND2X2_1372 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf5), .B(u_sdrc_core_u_bs_convert__abc_21684_n366), .Y(u_sdrc_core_u_bs_convert__abc_21684_n367) );
  AND2X2 AND2X2_1373 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n367), .B(u_sdrc_core_u_bs_convert__abc_21684_n365_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n368) );
  AND2X2 AND2X2_1374 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n370), .B(u_sdrc_core_u_bs_convert__abc_21684_n371_1), .Y(u_sdrc_core_a2x_wren_n_0_) );
  AND2X2 AND2X2_1375 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n211), .B(app_wr_en_n_1_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n373) );
  AND2X2 AND2X2_1376 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf2), .B(app_wr_en_n_3_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n374) );
  AND2X2 AND2X2_1377 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf4), .B(u_sdrc_core_u_bs_convert__abc_21684_n374), .Y(u_sdrc_core_u_bs_convert__abc_21684_n375) );
  AND2X2 AND2X2_1378 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n377), .B(u_sdrc_core_u_bs_convert__abc_21684_n169_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n378) );
  AND2X2 AND2X2_1379 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n379), .B(u_sdrc_core_u_bs_convert_x2a_wrnext_bF_buf3), .Y(app_wr_next_req) );
  AND2X2 AND2X2_138 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n491), .B(u_sdrc_core_u_bank_ctl__abc_21249_n492), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n493) );
  AND2X2 AND2X2_1380 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n382), .B(u_sdrc_core_u_bs_convert__abc_21684_n381_1), .Y(app_rd_data_0_) );
  AND2X2 AND2X2_1381 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n385), .B(u_sdrc_core_u_bs_convert__abc_21684_n384), .Y(app_rd_data_1_) );
  AND2X2 AND2X2_1382 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n388), .B(u_sdrc_core_u_bs_convert__abc_21684_n387), .Y(app_rd_data_2_) );
  AND2X2 AND2X2_1383 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n391_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n390), .Y(app_rd_data_3_) );
  AND2X2 AND2X2_1384 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n394), .B(u_sdrc_core_u_bs_convert__abc_21684_n393), .Y(app_rd_data_4_) );
  AND2X2 AND2X2_1385 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n397), .B(u_sdrc_core_u_bs_convert__abc_21684_n396_1), .Y(app_rd_data_5_) );
  AND2X2 AND2X2_1386 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n400), .B(u_sdrc_core_u_bs_convert__abc_21684_n399), .Y(app_rd_data_6_) );
  AND2X2 AND2X2_1387 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n403), .B(u_sdrc_core_u_bs_convert__abc_21684_n402), .Y(app_rd_data_7_) );
  AND2X2 AND2X2_1388 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n406_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n405), .Y(app_rd_data_8_) );
  AND2X2 AND2X2_1389 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n409), .B(u_sdrc_core_u_bs_convert__abc_21684_n408), .Y(app_rd_data_9_) );
  AND2X2 AND2X2_139 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n493), .B(u_sdrc_core_u_bank_ctl__abc_21249_n227_bF_buf1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n494) );
  AND2X2 AND2X2_1390 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n412), .B(u_sdrc_core_u_bs_convert__abc_21684_n411), .Y(app_rd_data_10_) );
  AND2X2 AND2X2_1391 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n415), .B(u_sdrc_core_u_bs_convert__abc_21684_n414), .Y(app_rd_data_11_) );
  AND2X2 AND2X2_1392 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n418), .B(u_sdrc_core_u_bs_convert__abc_21684_n417), .Y(app_rd_data_12_) );
  AND2X2 AND2X2_1393 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n421), .B(u_sdrc_core_u_bs_convert__abc_21684_n420), .Y(app_rd_data_13_) );
  AND2X2 AND2X2_1394 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n424), .B(u_sdrc_core_u_bs_convert__abc_21684_n423), .Y(app_rd_data_14_) );
  AND2X2 AND2X2_1395 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n427), .B(u_sdrc_core_u_bs_convert__abc_21684_n426), .Y(app_rd_data_15_) );
  AND2X2 AND2X2_1396 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf3), .B(u_sdrc_core_pad_sdr_din2_0_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n429) );
  AND2X2 AND2X2_1397 ( .A(cfg_sdr_width_1_bF_buf5), .B(u_sdrc_core_u_bs_convert_saved_rd_data_16_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n430) );
  AND2X2 AND2X2_1398 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf2), .B(u_sdrc_core_pad_sdr_din2_1_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n432) );
  AND2X2 AND2X2_1399 ( .A(cfg_sdr_width_1_bF_buf4), .B(u_sdrc_core_u_bs_convert_saved_rd_data_17_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n433) );
  AND2X2 AND2X2_14 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_xfr_ok), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_req), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n232_1) );
  AND2X2 AND2X2_140 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_len_1_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n496) );
  AND2X2 AND2X2_1400 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf1), .B(u_sdrc_core_pad_sdr_din2_2_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n435) );
  AND2X2 AND2X2_1401 ( .A(cfg_sdr_width_1_bF_buf3), .B(u_sdrc_core_u_bs_convert_saved_rd_data_18_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n436) );
  AND2X2 AND2X2_1402 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf0), .B(u_sdrc_core_pad_sdr_din2_3_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n438) );
  AND2X2 AND2X2_1403 ( .A(cfg_sdr_width_1_bF_buf2), .B(u_sdrc_core_u_bs_convert_saved_rd_data_19_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n439) );
  AND2X2 AND2X2_1404 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf5), .B(u_sdrc_core_pad_sdr_din2_4_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n441) );
  AND2X2 AND2X2_1405 ( .A(cfg_sdr_width_1_bF_buf1), .B(u_sdrc_core_u_bs_convert_saved_rd_data_20_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n442) );
  AND2X2 AND2X2_1406 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf4), .B(u_sdrc_core_pad_sdr_din2_5_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n444) );
  AND2X2 AND2X2_1407 ( .A(cfg_sdr_width_1_bF_buf0), .B(u_sdrc_core_u_bs_convert_saved_rd_data_21_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n445) );
  AND2X2 AND2X2_1408 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf3), .B(u_sdrc_core_pad_sdr_din2_6_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n447) );
  AND2X2 AND2X2_1409 ( .A(cfg_sdr_width_1_bF_buf5), .B(u_sdrc_core_u_bs_convert_saved_rd_data_22_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n448) );
  AND2X2 AND2X2_141 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n498), .B(u_sdrc_core_u_bank_ctl__abc_21249_n497), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n499) );
  AND2X2 AND2X2_1410 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf2), .B(u_sdrc_core_pad_sdr_din2_7_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n450) );
  AND2X2 AND2X2_1411 ( .A(cfg_sdr_width_1_bF_buf4), .B(u_sdrc_core_u_bs_convert_saved_rd_data_23_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n451) );
  AND2X2 AND2X2_1412 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf1), .B(u_sdrc_core_pad_sdr_din2_8_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n453) );
  AND2X2 AND2X2_1413 ( .A(cfg_sdr_width_1_bF_buf3), .B(u_sdrc_core_pad_sdr_din2_0_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n454) );
  AND2X2 AND2X2_1414 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf0), .B(u_sdrc_core_pad_sdr_din2_9_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n456) );
  AND2X2 AND2X2_1415 ( .A(cfg_sdr_width_1_bF_buf2), .B(u_sdrc_core_pad_sdr_din2_1_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n457) );
  AND2X2 AND2X2_1416 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf5), .B(u_sdrc_core_pad_sdr_din2_10_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n459) );
  AND2X2 AND2X2_1417 ( .A(cfg_sdr_width_1_bF_buf1), .B(u_sdrc_core_pad_sdr_din2_2_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n460) );
  AND2X2 AND2X2_1418 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf4), .B(u_sdrc_core_pad_sdr_din2_11_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n462) );
  AND2X2 AND2X2_1419 ( .A(cfg_sdr_width_1_bF_buf0), .B(u_sdrc_core_pad_sdr_din2_3_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n463) );
  AND2X2 AND2X2_142 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n500), .B(u_sdrc_core_u_bank_ctl__abc_21249_n501), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n502) );
  AND2X2 AND2X2_1420 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf3), .B(u_sdrc_core_pad_sdr_din2_12_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n465) );
  AND2X2 AND2X2_1421 ( .A(cfg_sdr_width_1_bF_buf5), .B(u_sdrc_core_pad_sdr_din2_4_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n466) );
  AND2X2 AND2X2_1422 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf2), .B(u_sdrc_core_pad_sdr_din2_13_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n468) );
  AND2X2 AND2X2_1423 ( .A(cfg_sdr_width_1_bF_buf4), .B(u_sdrc_core_pad_sdr_din2_5_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n469) );
  AND2X2 AND2X2_1424 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf1), .B(u_sdrc_core_pad_sdr_din2_14_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n471) );
  AND2X2 AND2X2_1425 ( .A(cfg_sdr_width_1_bF_buf3), .B(u_sdrc_core_pad_sdr_din2_6_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n472) );
  AND2X2 AND2X2_1426 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf0), .B(u_sdrc_core_pad_sdr_din2_15_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n474) );
  AND2X2 AND2X2_1427 ( .A(cfg_sdr_width_1_bF_buf2), .B(u_sdrc_core_pad_sdr_din2_7_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n475) );
  AND2X2 AND2X2_1428 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n478), .B(u_sdrc_core_u_bs_convert_x2a_rdok), .Y(u_sdrc_core_u_bs_convert__abc_21684_n479) );
  AND2X2 AND2X2_1429 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n477), .B(u_sdrc_core_u_bs_convert__abc_21684_n479), .Y(app_rd_valid) );
  AND2X2 AND2X2_143 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n502), .B(u_sdrc_core_u_bank_ctl__abc_21249_n227_bF_buf0), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n503) );
  AND2X2 AND2X2_1430 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n481), .B(sdram_resetn_bF_buf2), .Y(u_sdrc_core_u_bs_convert__abc_21684_n482) );
  AND2X2 AND2X2_1431 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf0), .B(u_sdrc_core_u_bs_convert_x2a_wrnext_bF_buf2), .Y(u_sdrc_core_u_bs_convert__abc_21684_n483) );
  AND2X2 AND2X2_1432 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n484), .B(u_sdrc_core_u_bs_convert__abc_21684_n485), .Y(u_sdrc_core_u_bs_convert__abc_21684_n486) );
  AND2X2 AND2X2_1433 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n486), .B(u_sdrc_core_u_bs_convert__abc_21684_n482), .Y(u_sdrc_core_u_bs_convert_wr_xfr_count_0__FF_INPUT) );
  AND2X2 AND2X2_1434 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n483), .B(u_sdrc_core_u_bs_convert_wr_xfr_count_1_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n488) );
  AND2X2 AND2X2_1435 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n490), .B(u_sdrc_core_u_bs_convert__abc_21684_n482), .Y(u_sdrc_core_u_bs_convert__abc_21684_n491) );
  AND2X2 AND2X2_1436 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n491), .B(u_sdrc_core_u_bs_convert__abc_21684_n489), .Y(u_sdrc_core_u_bs_convert_wr_xfr_count_1__FF_INPUT) );
  AND2X2 AND2X2_1437 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n493), .B(sdram_resetn_bF_buf1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n494) );
  AND2X2 AND2X2_1438 ( .A(u_sdrc_core_u_bs_convert_x2a_rdok), .B(u_sdrc_core_u_bs_convert_rd_xfr_count_0_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n495) );
  AND2X2 AND2X2_1439 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n496), .B(u_sdrc_core_u_bs_convert__abc_21684_n497), .Y(u_sdrc_core_u_bs_convert__abc_21684_n498) );
  AND2X2 AND2X2_144 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_len_2_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n505) );
  AND2X2 AND2X2_1440 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n498), .B(u_sdrc_core_u_bs_convert__abc_21684_n494), .Y(u_sdrc_core_u_bs_convert_rd_xfr_count_0__FF_INPUT) );
  AND2X2 AND2X2_1441 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n495), .B(u_sdrc_core_u_bs_convert_rd_xfr_count_1_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n500) );
  AND2X2 AND2X2_1442 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n502), .B(u_sdrc_core_u_bs_convert__abc_21684_n494), .Y(u_sdrc_core_u_bs_convert__abc_21684_n503) );
  AND2X2 AND2X2_1443 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n503), .B(u_sdrc_core_u_bs_convert__abc_21684_n501), .Y(u_sdrc_core_u_bs_convert_rd_xfr_count_1__FF_INPUT) );
  AND2X2 AND2X2_1444 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n505), .B(u_sdrc_core_u_bs_convert_rd_xfr_count_1_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n506) );
  AND2X2 AND2X2_1445 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n506), .B(u_sdrc_core_u_bs_convert_x2a_rdok), .Y(u_sdrc_core_u_bs_convert__abc_21684_n507) );
  AND2X2 AND2X2_1446 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n507), .B(u_sdrc_core_u_bs_convert__abc_21684_n185_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n508) );
  AND2X2 AND2X2_1447 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n508), .B(u_sdrc_core_pad_sdr_din2_0_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n509) );
  AND2X2 AND2X2_1448 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n510), .B(u_sdrc_core_u_bs_convert_saved_rd_data_16_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n511) );
  AND2X2 AND2X2_1449 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n512), .B(sdram_resetn_bF_buf0), .Y(u_sdrc_core_u_bs_convert_saved_rd_data_16__FF_INPUT) );
  AND2X2 AND2X2_145 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n507), .B(u_sdrc_core_u_bank_ctl__abc_21249_n506), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n508) );
  AND2X2 AND2X2_1450 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n508), .B(u_sdrc_core_pad_sdr_din2_1_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n514) );
  AND2X2 AND2X2_1451 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n510), .B(u_sdrc_core_u_bs_convert_saved_rd_data_17_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n515) );
  AND2X2 AND2X2_1452 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n516), .B(sdram_resetn_bF_buf49), .Y(u_sdrc_core_u_bs_convert_saved_rd_data_17__FF_INPUT) );
  AND2X2 AND2X2_1453 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n508), .B(u_sdrc_core_pad_sdr_din2_2_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n518) );
  AND2X2 AND2X2_1454 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n510), .B(u_sdrc_core_u_bs_convert_saved_rd_data_18_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n519) );
  AND2X2 AND2X2_1455 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n520), .B(sdram_resetn_bF_buf48), .Y(u_sdrc_core_u_bs_convert_saved_rd_data_18__FF_INPUT) );
  AND2X2 AND2X2_1456 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n508), .B(u_sdrc_core_pad_sdr_din2_3_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n522) );
  AND2X2 AND2X2_1457 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n510), .B(u_sdrc_core_u_bs_convert_saved_rd_data_19_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n523) );
  AND2X2 AND2X2_1458 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n524), .B(sdram_resetn_bF_buf47), .Y(u_sdrc_core_u_bs_convert_saved_rd_data_19__FF_INPUT) );
  AND2X2 AND2X2_1459 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n508), .B(u_sdrc_core_pad_sdr_din2_4_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n526) );
  AND2X2 AND2X2_146 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n509), .B(u_sdrc_core_u_bank_ctl__abc_21249_n510), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n511) );
  AND2X2 AND2X2_1460 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n510), .B(u_sdrc_core_u_bs_convert_saved_rd_data_20_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n527) );
  AND2X2 AND2X2_1461 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n528), .B(sdram_resetn_bF_buf46), .Y(u_sdrc_core_u_bs_convert_saved_rd_data_20__FF_INPUT) );
  AND2X2 AND2X2_1462 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n508), .B(u_sdrc_core_pad_sdr_din2_5_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n530) );
  AND2X2 AND2X2_1463 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n510), .B(u_sdrc_core_u_bs_convert_saved_rd_data_21_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n531) );
  AND2X2 AND2X2_1464 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n532), .B(sdram_resetn_bF_buf45), .Y(u_sdrc_core_u_bs_convert_saved_rd_data_21__FF_INPUT) );
  AND2X2 AND2X2_1465 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n508), .B(u_sdrc_core_pad_sdr_din2_6_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n534) );
  AND2X2 AND2X2_1466 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n510), .B(u_sdrc_core_u_bs_convert_saved_rd_data_22_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n535) );
  AND2X2 AND2X2_1467 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n536), .B(sdram_resetn_bF_buf44), .Y(u_sdrc_core_u_bs_convert_saved_rd_data_22__FF_INPUT) );
  AND2X2 AND2X2_1468 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n508), .B(u_sdrc_core_pad_sdr_din2_7_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n538) );
  AND2X2 AND2X2_1469 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n510), .B(u_sdrc_core_u_bs_convert_saved_rd_data_23_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n539) );
  AND2X2 AND2X2_147 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n511), .B(u_sdrc_core_u_bank_ctl__abc_21249_n227_bF_buf3), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n512) );
  AND2X2 AND2X2_1470 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n540), .B(sdram_resetn_bF_buf43), .Y(u_sdrc_core_u_bs_convert_saved_rd_data_23__FF_INPUT) );
  AND2X2 AND2X2_1471 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n185_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n543), .Y(u_sdrc_core_u_bs_convert__abc_21684_n544) );
  AND2X2 AND2X2_1472 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n548), .B(sdram_resetn_bF_buf42), .Y(u_sdrc_core_u_bs_convert__abc_21684_n549) );
  AND2X2 AND2X2_1473 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n549), .B(u_sdrc_core_u_bs_convert__abc_21684_n547), .Y(u_sdrc_core_u_bs_convert_saved_rd_data_0__FF_INPUT) );
  AND2X2 AND2X2_1474 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n552), .B(sdram_resetn_bF_buf41), .Y(u_sdrc_core_u_bs_convert__abc_21684_n553) );
  AND2X2 AND2X2_1475 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n553), .B(u_sdrc_core_u_bs_convert__abc_21684_n551), .Y(u_sdrc_core_u_bs_convert_saved_rd_data_1__FF_INPUT) );
  AND2X2 AND2X2_1476 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n556), .B(sdram_resetn_bF_buf40), .Y(u_sdrc_core_u_bs_convert__abc_21684_n557) );
  AND2X2 AND2X2_1477 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n557), .B(u_sdrc_core_u_bs_convert__abc_21684_n555), .Y(u_sdrc_core_u_bs_convert_saved_rd_data_2__FF_INPUT) );
  AND2X2 AND2X2_1478 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n560), .B(sdram_resetn_bF_buf39), .Y(u_sdrc_core_u_bs_convert__abc_21684_n561) );
  AND2X2 AND2X2_1479 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n561), .B(u_sdrc_core_u_bs_convert__abc_21684_n559), .Y(u_sdrc_core_u_bs_convert_saved_rd_data_3__FF_INPUT) );
  AND2X2 AND2X2_148 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_len_3_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n514) );
  AND2X2 AND2X2_1480 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n564), .B(sdram_resetn_bF_buf38), .Y(u_sdrc_core_u_bs_convert__abc_21684_n565) );
  AND2X2 AND2X2_1481 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n565), .B(u_sdrc_core_u_bs_convert__abc_21684_n563), .Y(u_sdrc_core_u_bs_convert_saved_rd_data_4__FF_INPUT) );
  AND2X2 AND2X2_1482 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n568), .B(sdram_resetn_bF_buf37), .Y(u_sdrc_core_u_bs_convert__abc_21684_n569) );
  AND2X2 AND2X2_1483 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n569), .B(u_sdrc_core_u_bs_convert__abc_21684_n567), .Y(u_sdrc_core_u_bs_convert_saved_rd_data_5__FF_INPUT) );
  AND2X2 AND2X2_1484 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n572), .B(sdram_resetn_bF_buf36), .Y(u_sdrc_core_u_bs_convert__abc_21684_n573) );
  AND2X2 AND2X2_1485 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n573), .B(u_sdrc_core_u_bs_convert__abc_21684_n571), .Y(u_sdrc_core_u_bs_convert_saved_rd_data_6__FF_INPUT) );
  AND2X2 AND2X2_1486 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n576), .B(sdram_resetn_bF_buf35), .Y(u_sdrc_core_u_bs_convert__abc_21684_n577) );
  AND2X2 AND2X2_1487 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n577), .B(u_sdrc_core_u_bs_convert__abc_21684_n575), .Y(u_sdrc_core_u_bs_convert_saved_rd_data_7__FF_INPUT) );
  AND2X2 AND2X2_1488 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n581), .B(u_sdrc_core_u_bs_convert__abc_21684_n582), .Y(u_sdrc_core_u_bs_convert__abc_21684_n583) );
  AND2X2 AND2X2_1489 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n583), .B(u_sdrc_core_u_bs_convert__abc_21684_n185_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n584) );
  AND2X2 AND2X2_149 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n516), .B(u_sdrc_core_u_bank_ctl__abc_21249_n515), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n517) );
  AND2X2 AND2X2_1490 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n587), .B(sdram_resetn_bF_buf34), .Y(u_sdrc_core_u_bs_convert__abc_21684_n588) );
  AND2X2 AND2X2_1491 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n586), .B(u_sdrc_core_u_bs_convert__abc_21684_n588), .Y(u_sdrc_core_u_bs_convert_saved_rd_data_8__FF_INPUT) );
  AND2X2 AND2X2_1492 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n590), .B(u_sdrc_core_u_bs_convert__abc_21684_n591), .Y(u_sdrc_core_u_bs_convert__abc_21684_n592) );
  AND2X2 AND2X2_1493 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n592), .B(u_sdrc_core_u_bs_convert__abc_21684_n185_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n593) );
  AND2X2 AND2X2_1494 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n596), .B(sdram_resetn_bF_buf33), .Y(u_sdrc_core_u_bs_convert__abc_21684_n597) );
  AND2X2 AND2X2_1495 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n595), .B(u_sdrc_core_u_bs_convert__abc_21684_n597), .Y(u_sdrc_core_u_bs_convert_saved_rd_data_9__FF_INPUT) );
  AND2X2 AND2X2_1496 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n599), .B(u_sdrc_core_u_bs_convert__abc_21684_n600), .Y(u_sdrc_core_u_bs_convert__abc_21684_n601) );
  AND2X2 AND2X2_1497 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n601), .B(u_sdrc_core_u_bs_convert__abc_21684_n185_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n602) );
  AND2X2 AND2X2_1498 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n605), .B(sdram_resetn_bF_buf32), .Y(u_sdrc_core_u_bs_convert__abc_21684_n606) );
  AND2X2 AND2X2_1499 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n604), .B(u_sdrc_core_u_bs_convert__abc_21684_n606), .Y(u_sdrc_core_u_bs_convert_saved_rd_data_10__FF_INPUT) );
  AND2X2 AND2X2_15 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_req), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n233_1) );
  AND2X2 AND2X2_150 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n518), .B(u_sdrc_core_u_bank_ctl__abc_21249_n519), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n520) );
  AND2X2 AND2X2_1500 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n608), .B(u_sdrc_core_u_bs_convert__abc_21684_n609), .Y(u_sdrc_core_u_bs_convert__abc_21684_n610) );
  AND2X2 AND2X2_1501 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n610), .B(u_sdrc_core_u_bs_convert__abc_21684_n185_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n611) );
  AND2X2 AND2X2_1502 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n614), .B(sdram_resetn_bF_buf31), .Y(u_sdrc_core_u_bs_convert__abc_21684_n615) );
  AND2X2 AND2X2_1503 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n613), .B(u_sdrc_core_u_bs_convert__abc_21684_n615), .Y(u_sdrc_core_u_bs_convert_saved_rd_data_11__FF_INPUT) );
  AND2X2 AND2X2_1504 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n617), .B(u_sdrc_core_u_bs_convert__abc_21684_n618), .Y(u_sdrc_core_u_bs_convert__abc_21684_n619) );
  AND2X2 AND2X2_1505 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n619), .B(u_sdrc_core_u_bs_convert__abc_21684_n185_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n620) );
  AND2X2 AND2X2_1506 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n623), .B(sdram_resetn_bF_buf30), .Y(u_sdrc_core_u_bs_convert__abc_21684_n624) );
  AND2X2 AND2X2_1507 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n622), .B(u_sdrc_core_u_bs_convert__abc_21684_n624), .Y(u_sdrc_core_u_bs_convert_saved_rd_data_12__FF_INPUT) );
  AND2X2 AND2X2_1508 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n626), .B(u_sdrc_core_u_bs_convert__abc_21684_n627), .Y(u_sdrc_core_u_bs_convert__abc_21684_n628) );
  AND2X2 AND2X2_1509 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n628), .B(u_sdrc_core_u_bs_convert__abc_21684_n185_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n629) );
  AND2X2 AND2X2_151 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n520), .B(u_sdrc_core_u_bank_ctl__abc_21249_n227_bF_buf2), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n521) );
  AND2X2 AND2X2_1510 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n632), .B(sdram_resetn_bF_buf29), .Y(u_sdrc_core_u_bs_convert__abc_21684_n633) );
  AND2X2 AND2X2_1511 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n631), .B(u_sdrc_core_u_bs_convert__abc_21684_n633), .Y(u_sdrc_core_u_bs_convert_saved_rd_data_13__FF_INPUT) );
  AND2X2 AND2X2_1512 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n635), .B(u_sdrc_core_u_bs_convert__abc_21684_n636), .Y(u_sdrc_core_u_bs_convert__abc_21684_n637) );
  AND2X2 AND2X2_1513 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n637), .B(u_sdrc_core_u_bs_convert__abc_21684_n185_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n638) );
  AND2X2 AND2X2_1514 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n641), .B(sdram_resetn_bF_buf28), .Y(u_sdrc_core_u_bs_convert__abc_21684_n642) );
  AND2X2 AND2X2_1515 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n640), .B(u_sdrc_core_u_bs_convert__abc_21684_n642), .Y(u_sdrc_core_u_bs_convert_saved_rd_data_14__FF_INPUT) );
  AND2X2 AND2X2_1516 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n644), .B(u_sdrc_core_u_bs_convert__abc_21684_n645), .Y(u_sdrc_core_u_bs_convert__abc_21684_n646) );
  AND2X2 AND2X2_1517 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n646), .B(u_sdrc_core_u_bs_convert__abc_21684_n185_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n647) );
  AND2X2 AND2X2_1518 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n650), .B(sdram_resetn_bF_buf27), .Y(u_sdrc_core_u_bs_convert__abc_21684_n651) );
  AND2X2 AND2X2_1519 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n649), .B(u_sdrc_core_u_bs_convert__abc_21684_n651), .Y(u_sdrc_core_u_bs_convert_saved_rd_data_15__FF_INPUT) );
  AND2X2 AND2X2_152 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_len_4_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n523) );
  AND2X2 AND2X2_1520 ( .A(u_sdrc_core_u_req_gen__abc_22171_n181), .B(sdram_resetn_bF_buf26), .Y(u_sdrc_core_u_req_gen__abc_22171_n182_1) );
  AND2X2 AND2X2_1521 ( .A(u_sdrc_core_u_req_gen__abc_22171_n182_1), .B(u_sdrc_core_u_req_gen_req_st_1_), .Y(u_sdrc_core_u_req_gen__abc_22171_n183) );
  AND2X2 AND2X2_1522 ( .A(u_sdrc_core_b2r_ack), .B(u_sdrc_core_u_req_gen_req_st_2_), .Y(u_sdrc_core_u_req_gen__abc_22171_n184) );
  AND2X2 AND2X2_1523 ( .A(sdram_resetn_bF_buf25), .B(u_sdrc_core_u_req_gen_page_ovflw_r), .Y(u_sdrc_core_u_req_gen__abc_22171_n185) );
  AND2X2 AND2X2_1524 ( .A(u_sdrc_core_u_req_gen__abc_22171_n184), .B(u_sdrc_core_u_req_gen__abc_22171_n185), .Y(u_sdrc_core_u_req_gen__abc_22171_n186) );
  AND2X2 AND2X2_1525 ( .A(u_sdrc_core_u_req_gen__abc_22171_n182_1), .B(u_sdrc_core_u_req_gen_req_st_2_), .Y(u_sdrc_core_u_req_gen__abc_22171_n188) );
  AND2X2 AND2X2_1526 ( .A(sdram_resetn_bF_buf24), .B(u_sdrc_core_u_req_gen_req_st_0_), .Y(u_sdrc_core_u_req_gen__abc_22171_n189) );
  AND2X2 AND2X2_1527 ( .A(u_sdrc_core_b2r_arb_ok), .B(app_req), .Y(u_sdrc_core_u_req_gen__abc_22171_n190) );
  AND2X2 AND2X2_1528 ( .A(u_sdrc_core_u_req_gen__abc_22171_n189), .B(u_sdrc_core_u_req_gen__abc_22171_n190), .Y(u_sdrc_core_u_req_gen__abc_22171_n191) );
  AND2X2 AND2X2_1529 ( .A(u_sdrc_core_u_req_gen__abc_22171_n193), .B(u_sdrc_core_u_req_gen__abc_22171_n189), .Y(u_sdrc_core_u_req_gen__abc_22171_n194) );
  AND2X2 AND2X2_153 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n525), .B(u_sdrc_core_u_bank_ctl__abc_21249_n524), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n526) );
  AND2X2 AND2X2_1530 ( .A(u_sdrc_core_u_req_gen__abc_22171_n184), .B(u_sdrc_core_u_req_gen__abc_22171_n195_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n196) );
  AND2X2 AND2X2_1531 ( .A(u_sdrc_core_u_req_gen_req_st_1_), .B(u_sdrc_core_b2r_ack), .Y(u_sdrc_core_u_req_gen__abc_22171_n198) );
  AND2X2 AND2X2_1532 ( .A(u_sdrc_core_u_req_gen_page_ovflw_r), .B(u_sdrc_core_r2b_start), .Y(u_sdrc_core_u_req_gen__abc_22171_n202) );
  AND2X2 AND2X2_1533 ( .A(u_sdrc_core_u_req_gen__abc_22171_n202), .B(u_sdrc_core_u_req_gen_max_r2b_len_r_0_), .Y(u_sdrc_core_u_req_gen__abc_22171_n203) );
  AND2X2 AND2X2_1534 ( .A(u_sdrc_core_u_req_gen__abc_22171_n204), .B(u_sdrc_core_u_req_gen_lcl_req_len_0_), .Y(u_sdrc_core_u_req_gen__abc_22171_n205) );
  AND2X2 AND2X2_1535 ( .A(u_sdrc_core_u_req_gen__abc_22171_n202), .B(u_sdrc_core_u_req_gen__abc_22171_n208), .Y(u_sdrc_core_u_req_gen__abc_22171_n209) );
  AND2X2 AND2X2_1536 ( .A(u_sdrc_core_u_req_gen__abc_22171_n210_1), .B(u_sdrc_core_u_req_gen__abc_22171_n207), .Y(u_sdrc_core_r2b_len_1_) );
  AND2X2 AND2X2_1537 ( .A(u_sdrc_core_u_req_gen__abc_22171_n204), .B(u_sdrc_core_u_req_gen__abc_22171_n212), .Y(u_sdrc_core_u_req_gen__abc_22171_n213) );
  AND2X2 AND2X2_1538 ( .A(u_sdrc_core_u_req_gen__abc_22171_n202), .B(u_sdrc_core_u_req_gen__abc_22171_n214), .Y(u_sdrc_core_u_req_gen__abc_22171_n215_1) );
  AND2X2 AND2X2_1539 ( .A(u_sdrc_core_u_req_gen__abc_22171_n204), .B(u_sdrc_core_u_req_gen__abc_22171_n218), .Y(u_sdrc_core_u_req_gen__abc_22171_n219_1) );
  AND2X2 AND2X2_154 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n527), .B(u_sdrc_core_u_bank_ctl__abc_21249_n528), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n529) );
  AND2X2 AND2X2_1540 ( .A(u_sdrc_core_u_req_gen__abc_22171_n202), .B(u_sdrc_core_u_req_gen__abc_22171_n220), .Y(u_sdrc_core_u_req_gen__abc_22171_n221_1) );
  AND2X2 AND2X2_1541 ( .A(u_sdrc_core_u_req_gen__abc_22171_n202), .B(u_sdrc_core_u_req_gen__abc_22171_n225), .Y(u_sdrc_core_u_req_gen__abc_22171_n226_1) );
  AND2X2 AND2X2_1542 ( .A(u_sdrc_core_u_req_gen__abc_22171_n227), .B(u_sdrc_core_u_req_gen__abc_22171_n224), .Y(u_sdrc_core_r2b_len_4_) );
  AND2X2 AND2X2_1543 ( .A(u_sdrc_core_u_req_gen__abc_22171_n202), .B(u_sdrc_core_u_req_gen__abc_22171_n230), .Y(u_sdrc_core_u_req_gen__abc_22171_n231) );
  AND2X2 AND2X2_1544 ( .A(u_sdrc_core_u_req_gen__abc_22171_n232), .B(u_sdrc_core_u_req_gen__abc_22171_n229), .Y(u_sdrc_core_r2b_len_5_) );
  AND2X2 AND2X2_1545 ( .A(u_sdrc_core_u_req_gen__abc_22171_n202), .B(u_sdrc_core_u_req_gen__abc_22171_n235), .Y(u_sdrc_core_u_req_gen__abc_22171_n236_1) );
  AND2X2 AND2X2_1546 ( .A(u_sdrc_core_u_req_gen__abc_22171_n237), .B(u_sdrc_core_u_req_gen__abc_22171_n234_1), .Y(u_sdrc_core_r2b_len_6_) );
  AND2X2 AND2X2_1547 ( .A(u_sdrc_core_u_req_gen__abc_22171_n190), .B(u_sdrc_core_u_req_gen_req_st_0_), .Y(app_req_ack) );
  AND2X2 AND2X2_1548 ( .A(u_sdrc_core_u_req_gen__abc_22171_n240), .B(u_sdrc_core_u_req_gen__abc_22171_n241), .Y(u_sdrc_core_u_req_gen__abc_22171_n242) );
  AND2X2 AND2X2_1549 ( .A(u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf4), .B(app_req_addr_0_), .Y(u_sdrc_core_u_req_gen__abc_22171_n243_1) );
  AND2X2 AND2X2_155 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n529), .B(u_sdrc_core_u_bank_ctl__abc_21249_n227_bF_buf1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n530) );
  AND2X2 AND2X2_1550 ( .A(u_sdrc_core_u_req_gen__abc_22171_n243_1), .B(app_req_ack_bF_buf6), .Y(u_sdrc_core_u_req_gen_max_r2b_len_r_0__FF_INPUT) );
  AND2X2 AND2X2_1551 ( .A(u_sdrc_core_u_req_gen__abc_22171_n241), .B(\cfg_sdr_width[0] ), .Y(u_sdrc_core_u_req_gen__abc_22171_n245_1) );
  AND2X2 AND2X2_1552 ( .A(u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf4), .B(app_req_addr_0_), .Y(u_sdrc_core_u_req_gen__abc_22171_n246) );
  AND2X2 AND2X2_1553 ( .A(u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf3), .B(app_req_addr_1_), .Y(u_sdrc_core_u_req_gen__abc_22171_n247) );
  AND2X2 AND2X2_1554 ( .A(u_sdrc_core_u_req_gen__abc_22171_n243_1), .B(app_req_addr_1_), .Y(u_sdrc_core_u_req_gen__abc_22171_n251) );
  AND2X2 AND2X2_1555 ( .A(u_sdrc_core_u_req_gen__abc_22171_n253), .B(app_req_ack_bF_buf5), .Y(u_sdrc_core_u_req_gen_max_r2b_len_r_1__FF_INPUT) );
  AND2X2 AND2X2_1556 ( .A(u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf2), .B(u_sdrc_core_u_req_gen__abc_22171_n255), .Y(u_sdrc_core_u_req_gen__abc_22171_n256_1) );
  AND2X2 AND2X2_1557 ( .A(u_sdrc_core_u_req_gen__abc_22171_n257), .B(cfg_sdr_width_1_bF_buf0), .Y(u_sdrc_core_u_req_gen__abc_22171_n258) );
  AND2X2 AND2X2_1558 ( .A(u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf3), .B(u_sdrc_core_u_req_gen__abc_22171_n259), .Y(u_sdrc_core_u_req_gen__abc_22171_n260) );
  AND2X2 AND2X2_1559 ( .A(u_sdrc_core_u_req_gen__abc_22171_n250), .B(u_sdrc_core_u_req_gen__abc_22171_n262_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n263_1) );
  AND2X2 AND2X2_156 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_len_5_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n532) );
  AND2X2 AND2X2_1560 ( .A(u_sdrc_core_u_req_gen__abc_22171_n264), .B(u_sdrc_core_u_req_gen__abc_22171_n249), .Y(u_sdrc_core_u_req_gen__abc_22171_n265) );
  AND2X2 AND2X2_1561 ( .A(u_sdrc_core_u_req_gen__abc_22171_n267), .B(app_req_ack_bF_buf4), .Y(u_sdrc_core_u_req_gen_max_r2b_len_r_2__FF_INPUT) );
  AND2X2 AND2X2_1562 ( .A(u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf1), .B(u_sdrc_core_u_req_gen__abc_22171_n269), .Y(u_sdrc_core_u_req_gen__abc_22171_n270) );
  AND2X2 AND2X2_1563 ( .A(u_sdrc_core_u_req_gen__abc_22171_n259), .B(cfg_sdr_width_1_bF_buf5), .Y(u_sdrc_core_u_req_gen__abc_22171_n271) );
  AND2X2 AND2X2_1564 ( .A(u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf2), .B(u_sdrc_core_u_req_gen__abc_22171_n255), .Y(u_sdrc_core_u_req_gen__abc_22171_n272) );
  AND2X2 AND2X2_1565 ( .A(u_sdrc_core_u_req_gen__abc_22171_n263_1), .B(u_sdrc_core_u_req_gen__abc_22171_n274), .Y(u_sdrc_core_u_req_gen__abc_22171_n275) );
  AND2X2 AND2X2_1566 ( .A(u_sdrc_core_u_req_gen__abc_22171_n276), .B(u_sdrc_core_u_req_gen__abc_22171_n277_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n278) );
  AND2X2 AND2X2_1567 ( .A(u_sdrc_core_u_req_gen__abc_22171_n278), .B(app_req_ack_bF_buf3), .Y(u_sdrc_core_u_req_gen_max_r2b_len_r_3__FF_INPUT) );
  AND2X2 AND2X2_1568 ( .A(u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf0), .B(u_sdrc_core_u_req_gen__abc_22171_n280), .Y(u_sdrc_core_u_req_gen__abc_22171_n281_1) );
  AND2X2 AND2X2_1569 ( .A(u_sdrc_core_u_req_gen__abc_22171_n255), .B(cfg_sdr_width_1_bF_buf4), .Y(u_sdrc_core_u_req_gen__abc_22171_n282) );
  AND2X2 AND2X2_157 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n534), .B(u_sdrc_core_u_bank_ctl__abc_21249_n533), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n535) );
  AND2X2 AND2X2_1570 ( .A(u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf1), .B(u_sdrc_core_u_req_gen__abc_22171_n269), .Y(u_sdrc_core_u_req_gen__abc_22171_n283_1) );
  AND2X2 AND2X2_1571 ( .A(u_sdrc_core_u_req_gen__abc_22171_n275), .B(u_sdrc_core_u_req_gen__abc_22171_n285), .Y(u_sdrc_core_u_req_gen__abc_22171_n286) );
  AND2X2 AND2X2_1572 ( .A(u_sdrc_core_u_req_gen__abc_22171_n276), .B(u_sdrc_core_u_req_gen__abc_22171_n287), .Y(u_sdrc_core_u_req_gen__abc_22171_n288) );
  AND2X2 AND2X2_1573 ( .A(u_sdrc_core_u_req_gen__abc_22171_n290_1), .B(app_req_ack_bF_buf2), .Y(u_sdrc_core_u_req_gen_max_r2b_len_r_4__FF_INPUT) );
  AND2X2 AND2X2_1574 ( .A(u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf4), .B(u_sdrc_core_u_req_gen__abc_22171_n292), .Y(u_sdrc_core_u_req_gen__abc_22171_n293) );
  AND2X2 AND2X2_1575 ( .A(u_sdrc_core_u_req_gen__abc_22171_n269), .B(cfg_sdr_width_1_bF_buf3), .Y(u_sdrc_core_u_req_gen__abc_22171_n294_1) );
  AND2X2 AND2X2_1576 ( .A(u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf0), .B(u_sdrc_core_u_req_gen__abc_22171_n280), .Y(u_sdrc_core_u_req_gen__abc_22171_n295) );
  AND2X2 AND2X2_1577 ( .A(u_sdrc_core_u_req_gen__abc_22171_n286), .B(u_sdrc_core_u_req_gen__abc_22171_n297), .Y(u_sdrc_core_u_req_gen__abc_22171_n298_1) );
  AND2X2 AND2X2_1578 ( .A(u_sdrc_core_u_req_gen__abc_22171_n299), .B(u_sdrc_core_u_req_gen__abc_22171_n300), .Y(u_sdrc_core_u_req_gen__abc_22171_n301) );
  AND2X2 AND2X2_1579 ( .A(u_sdrc_core_u_req_gen__abc_22171_n301), .B(app_req_ack_bF_buf1), .Y(u_sdrc_core_u_req_gen_max_r2b_len_r_5__FF_INPUT) );
  AND2X2 AND2X2_158 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n536), .B(u_sdrc_core_u_bank_ctl__abc_21249_n537), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n538) );
  AND2X2 AND2X2_1580 ( .A(u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf3), .B(app_req_addr_6_), .Y(u_sdrc_core_u_req_gen__abc_22171_n303) );
  AND2X2 AND2X2_1581 ( .A(cfg_sdr_width_1_bF_buf2), .B(app_req_addr_4_), .Y(u_sdrc_core_u_req_gen__abc_22171_n304_1) );
  AND2X2 AND2X2_1582 ( .A(u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf4), .B(app_req_addr_5_), .Y(u_sdrc_core_u_req_gen__abc_22171_n305) );
  AND2X2 AND2X2_1583 ( .A(u_sdrc_core_u_req_gen__abc_22171_n298_1), .B(u_sdrc_core_u_req_gen__abc_22171_n308), .Y(u_sdrc_core_u_req_gen__abc_22171_n309) );
  AND2X2 AND2X2_1584 ( .A(u_sdrc_core_u_req_gen__abc_22171_n299), .B(u_sdrc_core_u_req_gen__abc_22171_n307_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n310_1) );
  AND2X2 AND2X2_1585 ( .A(u_sdrc_core_u_req_gen__abc_22171_n312), .B(app_req_ack_bF_buf0), .Y(u_sdrc_core_u_req_gen_max_r2b_len_r_6__FF_INPUT) );
  AND2X2 AND2X2_1586 ( .A(app_req_ack_bF_buf6), .B(app_req_wr_n), .Y(u_sdrc_core_u_req_gen__abc_22171_n314) );
  AND2X2 AND2X2_1587 ( .A(u_sdrc_core_u_req_gen__abc_22171_n315), .B(u_sdrc_core_u_req_gen__abc_22171_n316), .Y(u_sdrc_core_u_req_gen_r2b_write_FF_INPUT) );
  AND2X2 AND2X2_1588 ( .A(u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf4), .B(u_sdrc_core_r2b_wrap), .Y(u_sdrc_core_u_req_gen__abc_22171_n331) );
  AND2X2 AND2X2_1589 ( .A(app_req_ack_bF_buf3), .B(1'b0), .Y(u_sdrc_core_u_req_gen__abc_22171_n332) );
  AND2X2 AND2X2_159 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n538), .B(u_sdrc_core_u_bank_ctl__abc_21249_n227_bF_buf0), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n539) );
  AND2X2 AND2X2_1590 ( .A(u_sdrc_core_r2b_req), .B(u_sdrc_core_b2r_ack), .Y(u_sdrc_core_u_req_gen__abc_22171_n335_1) );
  AND2X2 AND2X2_1591 ( .A(u_sdrc_core_r2b_len_0_), .B(u_sdrc_core_u_req_gen__abc_22171_n335_1_bF_buf3), .Y(u_sdrc_core_u_req_gen__abc_22171_n336) );
  AND2X2 AND2X2_1592 ( .A(u_sdrc_core_u_req_gen__abc_22171_n337_1), .B(u_sdrc_core_u_req_gen_lcl_req_len_0_), .Y(u_sdrc_core_u_req_gen__abc_22171_n338) );
  AND2X2 AND2X2_1593 ( .A(u_sdrc_core_u_req_gen__abc_22171_n336), .B(u_sdrc_core_u_req_gen__abc_22171_n339), .Y(u_sdrc_core_u_req_gen__abc_22171_n340) );
  AND2X2 AND2X2_1594 ( .A(u_sdrc_core_u_req_gen__abc_22171_n341_1), .B(u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf3), .Y(u_sdrc_core_u_req_gen__abc_22171_n342) );
  AND2X2 AND2X2_1595 ( .A(u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf2), .B(app_req_len_0_), .Y(u_sdrc_core_u_req_gen__abc_22171_n343_1) );
  AND2X2 AND2X2_1596 ( .A(u_sdrc_core_u_req_gen__abc_22171_n343_1), .B(app_req_ack_bF_buf2), .Y(u_sdrc_core_u_req_gen__abc_22171_n344) );
  AND2X2 AND2X2_1597 ( .A(u_sdrc_core_u_req_gen__abc_22171_n203), .B(u_sdrc_core_u_req_gen__abc_22171_n339), .Y(u_sdrc_core_u_req_gen__abc_22171_n347) );
  AND2X2 AND2X2_1598 ( .A(u_sdrc_core_u_req_gen__abc_22171_n209), .B(u_sdrc_core_u_req_gen_lcl_req_len_1_), .Y(u_sdrc_core_u_req_gen__abc_22171_n348) );
  AND2X2 AND2X2_1599 ( .A(u_sdrc_core_r2b_len_1_), .B(u_sdrc_core_u_req_gen__abc_22171_n349), .Y(u_sdrc_core_u_req_gen__abc_22171_n350_1) );
  AND2X2 AND2X2_16 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_req), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n235_1) );
  AND2X2 AND2X2_160 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_len_6_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n541) );
  AND2X2 AND2X2_1600 ( .A(u_sdrc_core_u_req_gen__abc_22171_n355), .B(u_sdrc_core_u_req_gen__abc_22171_n352_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n356) );
  AND2X2 AND2X2_1601 ( .A(u_sdrc_core_u_req_gen__abc_22171_n357), .B(u_sdrc_core_u_req_gen__abc_22171_n358_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n359) );
  AND2X2 AND2X2_1602 ( .A(u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf3), .B(app_req_len_0_), .Y(u_sdrc_core_u_req_gen__abc_22171_n361) );
  AND2X2 AND2X2_1603 ( .A(u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf1), .B(app_req_len_1_), .Y(u_sdrc_core_u_req_gen__abc_22171_n362) );
  AND2X2 AND2X2_1604 ( .A(u_sdrc_core_u_req_gen__abc_22171_n360_1), .B(u_sdrc_core_u_req_gen__abc_22171_n364), .Y(u_sdrc_core_u_req_gen_lcl_req_len_1__FF_INPUT) );
  AND2X2 AND2X2_1605 ( .A(u_sdrc_core_u_req_gen__abc_22171_n352_1), .B(u_sdrc_core_u_req_gen__abc_22171_n366), .Y(u_sdrc_core_u_req_gen__abc_22171_n367) );
  AND2X2 AND2X2_1606 ( .A(u_sdrc_core_u_req_gen__abc_22171_n215_1), .B(u_sdrc_core_u_req_gen_lcl_req_len_2_), .Y(u_sdrc_core_u_req_gen__abc_22171_n368) );
  AND2X2 AND2X2_1607 ( .A(u_sdrc_core_r2b_len_2_), .B(u_sdrc_core_u_req_gen__abc_22171_n212), .Y(u_sdrc_core_u_req_gen__abc_22171_n369_1) );
  AND2X2 AND2X2_1608 ( .A(u_sdrc_core_u_req_gen__abc_22171_n374), .B(u_sdrc_core_u_req_gen__abc_22171_n371_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n375) );
  AND2X2 AND2X2_1609 ( .A(u_sdrc_core_u_req_gen__abc_22171_n376), .B(u_sdrc_core_u_req_gen__abc_22171_n377_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n378) );
  AND2X2 AND2X2_161 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n543), .B(u_sdrc_core_u_bank_ctl__abc_21249_n542), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n544) );
  AND2X2 AND2X2_1610 ( .A(u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf0), .B(u_sdrc_core_u_req_gen__abc_22171_n380), .Y(u_sdrc_core_u_req_gen__abc_22171_n381) );
  AND2X2 AND2X2_1611 ( .A(u_sdrc_core_u_req_gen__abc_22171_n382_1), .B(cfg_sdr_width_1_bF_buf1), .Y(u_sdrc_core_u_req_gen__abc_22171_n383) );
  AND2X2 AND2X2_1612 ( .A(u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf2), .B(u_sdrc_core_u_req_gen__abc_22171_n384), .Y(u_sdrc_core_u_req_gen__abc_22171_n385) );
  AND2X2 AND2X2_1613 ( .A(u_sdrc_core_u_req_gen__abc_22171_n379_1), .B(u_sdrc_core_u_req_gen__abc_22171_n389), .Y(u_sdrc_core_u_req_gen_lcl_req_len_2__FF_INPUT) );
  AND2X2 AND2X2_1614 ( .A(u_sdrc_core_u_req_gen__abc_22171_n384), .B(cfg_sdr_width_1_bF_buf0), .Y(u_sdrc_core_u_req_gen__abc_22171_n393) );
  AND2X2 AND2X2_1615 ( .A(u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf1), .B(u_sdrc_core_u_req_gen__abc_22171_n380), .Y(u_sdrc_core_u_req_gen__abc_22171_n394_1) );
  AND2X2 AND2X2_1616 ( .A(u_sdrc_core_u_req_gen__abc_22171_n396_1), .B(u_sdrc_core_u_req_gen__abc_22171_n392), .Y(u_sdrc_core_u_req_gen__abc_22171_n397) );
  AND2X2 AND2X2_1617 ( .A(u_sdrc_core_u_req_gen__abc_22171_n397), .B(app_req_ack_bF_buf6), .Y(u_sdrc_core_u_req_gen__abc_22171_n398) );
  AND2X2 AND2X2_1618 ( .A(u_sdrc_core_u_req_gen__abc_22171_n346_1), .B(u_sdrc_core_u_req_gen_lcl_req_len_3_), .Y(u_sdrc_core_u_req_gen__abc_22171_n399) );
  AND2X2 AND2X2_1619 ( .A(u_sdrc_core_u_req_gen__abc_22171_n371_1), .B(u_sdrc_core_u_req_gen__abc_22171_n400_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n401) );
  AND2X2 AND2X2_162 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n545), .B(u_sdrc_core_u_bank_ctl__abc_21249_n546), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n547) );
  AND2X2 AND2X2_1620 ( .A(u_sdrc_core_u_req_gen__abc_22171_n221_1), .B(u_sdrc_core_u_req_gen_lcl_req_len_3_), .Y(u_sdrc_core_u_req_gen__abc_22171_n403) );
  AND2X2 AND2X2_1621 ( .A(u_sdrc_core_r2b_len_3_), .B(u_sdrc_core_u_req_gen__abc_22171_n218), .Y(u_sdrc_core_u_req_gen__abc_22171_n404_1) );
  AND2X2 AND2X2_1622 ( .A(u_sdrc_core_u_req_gen__abc_22171_n408_1), .B(u_sdrc_core_u_req_gen__abc_22171_n335_1_bF_buf3), .Y(u_sdrc_core_u_req_gen__abc_22171_n409) );
  AND2X2 AND2X2_1623 ( .A(u_sdrc_core_u_req_gen__abc_22171_n409), .B(u_sdrc_core_u_req_gen__abc_22171_n407), .Y(u_sdrc_core_u_req_gen__abc_22171_n410) );
  AND2X2 AND2X2_1624 ( .A(u_sdrc_core_u_req_gen__abc_22171_n411), .B(u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf0), .Y(u_sdrc_core_u_req_gen__abc_22171_n412_1) );
  AND2X2 AND2X2_1625 ( .A(u_sdrc_core_u_req_gen__abc_22171_n417_1), .B(u_sdrc_core_u_req_gen__abc_22171_n415), .Y(u_sdrc_core_u_req_gen__abc_22171_n418) );
  AND2X2 AND2X2_1626 ( .A(u_sdrc_core_u_req_gen__abc_22171_n418), .B(u_sdrc_core_u_req_gen__abc_22171_n414_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n419) );
  AND2X2 AND2X2_1627 ( .A(u_sdrc_core_u_req_gen__abc_22171_n419), .B(app_req_ack_bF_buf5), .Y(u_sdrc_core_u_req_gen__abc_22171_n420) );
  AND2X2 AND2X2_1628 ( .A(u_sdrc_core_u_req_gen__abc_22171_n346_1), .B(u_sdrc_core_u_req_gen_lcl_req_len_4_), .Y(u_sdrc_core_u_req_gen__abc_22171_n421_1) );
  AND2X2 AND2X2_1629 ( .A(u_sdrc_core_u_req_gen__abc_22171_n408_1), .B(u_sdrc_core_u_req_gen__abc_22171_n422), .Y(u_sdrc_core_u_req_gen__abc_22171_n423_1) );
  AND2X2 AND2X2_163 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n547), .B(u_sdrc_core_u_bank_ctl__abc_21249_n227_bF_buf3), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n548) );
  AND2X2 AND2X2_1630 ( .A(u_sdrc_core_u_req_gen__abc_22171_n226_1), .B(u_sdrc_core_u_req_gen_lcl_req_len_4_), .Y(u_sdrc_core_u_req_gen__abc_22171_n425_1) );
  AND2X2 AND2X2_1631 ( .A(u_sdrc_core_u_req_gen__abc_22171_n428), .B(u_sdrc_core_u_req_gen__abc_22171_n426), .Y(u_sdrc_core_u_req_gen__abc_22171_n429_1) );
  AND2X2 AND2X2_1632 ( .A(u_sdrc_core_u_req_gen__abc_22171_n432), .B(u_sdrc_core_u_req_gen__abc_22171_n335_1_bF_buf2), .Y(u_sdrc_core_u_req_gen__abc_22171_n433) );
  AND2X2 AND2X2_1633 ( .A(u_sdrc_core_u_req_gen__abc_22171_n433), .B(u_sdrc_core_u_req_gen__abc_22171_n430), .Y(u_sdrc_core_u_req_gen__abc_22171_n434) );
  AND2X2 AND2X2_1634 ( .A(u_sdrc_core_u_req_gen__abc_22171_n435), .B(u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf4), .Y(u_sdrc_core_u_req_gen__abc_22171_n436_1) );
  AND2X2 AND2X2_1635 ( .A(u_sdrc_core_u_req_gen__abc_22171_n440_1), .B(u_sdrc_core_u_req_gen__abc_22171_n439), .Y(u_sdrc_core_u_req_gen__abc_22171_n441) );
  AND2X2 AND2X2_1636 ( .A(u_sdrc_core_u_req_gen__abc_22171_n441), .B(u_sdrc_core_u_req_gen__abc_22171_n438), .Y(u_sdrc_core_u_req_gen__abc_22171_n442_1) );
  AND2X2 AND2X2_1637 ( .A(u_sdrc_core_u_req_gen__abc_22171_n442_1), .B(app_req_ack_bF_buf4), .Y(u_sdrc_core_u_req_gen__abc_22171_n443) );
  AND2X2 AND2X2_1638 ( .A(u_sdrc_core_u_req_gen__abc_22171_n346_1), .B(u_sdrc_core_u_req_gen_lcl_req_len_5_), .Y(u_sdrc_core_u_req_gen__abc_22171_n444_1) );
  AND2X2 AND2X2_1639 ( .A(u_sdrc_core_u_req_gen__abc_22171_n432), .B(u_sdrc_core_u_req_gen__abc_22171_n426), .Y(u_sdrc_core_u_req_gen__abc_22171_n445) );
  AND2X2 AND2X2_164 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_cmd_0_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n550) );
  AND2X2 AND2X2_1640 ( .A(u_sdrc_core_u_req_gen__abc_22171_n231), .B(u_sdrc_core_u_req_gen_lcl_req_len_5_), .Y(u_sdrc_core_u_req_gen__abc_22171_n447) );
  AND2X2 AND2X2_1641 ( .A(u_sdrc_core_u_req_gen__abc_22171_n450_1), .B(u_sdrc_core_u_req_gen__abc_22171_n448_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n451_1) );
  AND2X2 AND2X2_1642 ( .A(u_sdrc_core_u_req_gen__abc_22171_n454), .B(u_sdrc_core_u_req_gen__abc_22171_n335_1_bF_buf1), .Y(u_sdrc_core_u_req_gen__abc_22171_n455) );
  AND2X2 AND2X2_1643 ( .A(u_sdrc_core_u_req_gen__abc_22171_n455), .B(u_sdrc_core_u_req_gen__abc_22171_n452_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n456) );
  AND2X2 AND2X2_1644 ( .A(u_sdrc_core_u_req_gen__abc_22171_n457), .B(u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf3), .Y(u_sdrc_core_u_req_gen__abc_22171_n458) );
  AND2X2 AND2X2_1645 ( .A(u_sdrc_core_u_req_gen__abc_22171_n462_1), .B(u_sdrc_core_u_req_gen__abc_22171_n461), .Y(u_sdrc_core_u_req_gen__abc_22171_n463) );
  AND2X2 AND2X2_1646 ( .A(u_sdrc_core_u_req_gen__abc_22171_n463), .B(u_sdrc_core_u_req_gen__abc_22171_n460), .Y(u_sdrc_core_u_req_gen__abc_22171_n464_1) );
  AND2X2 AND2X2_1647 ( .A(u_sdrc_core_u_req_gen__abc_22171_n454), .B(u_sdrc_core_u_req_gen__abc_22171_n448_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n467) );
  AND2X2 AND2X2_1648 ( .A(u_sdrc_core_u_req_gen__abc_22171_n467), .B(u_sdrc_core_r2b_len_6_), .Y(u_sdrc_core_u_req_gen__abc_22171_n468_1) );
  AND2X2 AND2X2_1649 ( .A(u_sdrc_core_u_req_gen__abc_22171_n470), .B(u_sdrc_core_u_req_gen__abc_22171_n335_1_bF_buf0), .Y(u_sdrc_core_u_req_gen__abc_22171_n471_1) );
  AND2X2 AND2X2_165 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n552), .B(u_sdrc_core_u_bank_ctl__abc_21249_n551), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n553) );
  AND2X2 AND2X2_1650 ( .A(u_sdrc_core_u_req_gen__abc_22171_n471_1), .B(u_sdrc_core_u_req_gen__abc_22171_n469), .Y(u_sdrc_core_u_req_gen__abc_22171_n472) );
  AND2X2 AND2X2_1651 ( .A(u_sdrc_core_u_req_gen__abc_22171_n474_1), .B(u_sdrc_core_u_req_gen__abc_22171_n475), .Y(u_sdrc_core_u_req_gen__abc_22171_n476) );
  AND2X2 AND2X2_1652 ( .A(u_sdrc_core_u_req_gen__abc_22171_n477_1), .B(u_sdrc_core_u_req_gen__abc_22171_n465), .Y(u_sdrc_core_u_req_gen_lcl_req_len_6__FF_INPUT) );
  AND2X2 AND2X2_1653 ( .A(u_sdrc_core_r2b_len_0_), .B(u_sdrc_core_r2b_caddr_0_), .Y(u_sdrc_core_u_req_gen__abc_22171_n479) );
  AND2X2 AND2X2_1654 ( .A(u_sdrc_core_u_req_gen__abc_22171_n482), .B(u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf1), .Y(u_sdrc_core_u_req_gen__abc_22171_n483_1) );
  AND2X2 AND2X2_1655 ( .A(u_sdrc_core_u_req_gen__abc_22171_n483_1), .B(u_sdrc_core_u_req_gen__abc_22171_n481), .Y(u_sdrc_core_u_req_gen__abc_22171_n484) );
  AND2X2 AND2X2_1656 ( .A(u_sdrc_core_u_req_gen__abc_22171_n204), .B(u_sdrc_core_u_req_gen__abc_22171_n349), .Y(u_sdrc_core_u_req_gen__abc_22171_n487) );
  AND2X2 AND2X2_1657 ( .A(u_sdrc_core_u_req_gen__abc_22171_n489_1), .B(u_sdrc_core_u_req_gen__abc_22171_n490), .Y(u_sdrc_core_u_req_gen__abc_22171_n491) );
  AND2X2 AND2X2_1658 ( .A(u_sdrc_core_u_req_gen__abc_22171_n491), .B(u_sdrc_core_u_req_gen__abc_22171_n479), .Y(u_sdrc_core_u_req_gen__abc_22171_n492_1) );
  AND2X2 AND2X2_1659 ( .A(u_sdrc_core_u_req_gen__abc_22171_n493), .B(u_sdrc_core_u_req_gen__abc_22171_n494), .Y(u_sdrc_core_u_req_gen__abc_22171_n495_1) );
  AND2X2 AND2X2_166 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n554), .B(u_sdrc_core_u_bank_ctl__abc_21249_n555), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n556) );
  AND2X2 AND2X2_1660 ( .A(u_sdrc_core_u_req_gen__abc_22171_n496), .B(u_sdrc_core_u_req_gen__abc_22171_n497), .Y(u_sdrc_core_u_req_gen__abc_22171_n498_1) );
  AND2X2 AND2X2_1661 ( .A(u_sdrc_core_u_req_gen__abc_22171_n499), .B(u_sdrc_core_u_req_gen__abc_22171_n500), .Y(u_sdrc_core_u_req_gen_map_address_1_) );
  AND2X2 AND2X2_1662 ( .A(u_sdrc_core_r2b_len_1_), .B(u_sdrc_core_r2b_caddr_1_), .Y(u_sdrc_core_u_req_gen__abc_22171_n502) );
  AND2X2 AND2X2_1663 ( .A(u_sdrc_core_r2b_len_2_), .B(u_sdrc_core_r2b_caddr_2_), .Y(u_sdrc_core_u_req_gen__abc_22171_n504_1) );
  AND2X2 AND2X2_1664 ( .A(u_sdrc_core_u_req_gen__abc_22171_n505), .B(u_sdrc_core_u_req_gen__abc_22171_n506), .Y(u_sdrc_core_u_req_gen__abc_22171_n507_1) );
  AND2X2 AND2X2_1665 ( .A(u_sdrc_core_u_req_gen__abc_22171_n503), .B(u_sdrc_core_u_req_gen__abc_22171_n507_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n508_1) );
  AND2X2 AND2X2_1666 ( .A(u_sdrc_core_u_req_gen__abc_22171_n509_1), .B(u_sdrc_core_u_req_gen__abc_22171_n510_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n511) );
  AND2X2 AND2X2_1667 ( .A(u_sdrc_core_u_req_gen__abc_22171_n512), .B(u_sdrc_core_u_req_gen__abc_22171_n513), .Y(u_sdrc_core_u_req_gen__abc_22171_n514) );
  AND2X2 AND2X2_1668 ( .A(u_sdrc_core_u_req_gen__abc_22171_n515), .B(u_sdrc_core_u_req_gen__abc_22171_n516), .Y(u_sdrc_core_u_req_gen_map_address_2_) );
  AND2X2 AND2X2_1669 ( .A(u_sdrc_core_u_req_gen__abc_22171_n346_1), .B(u_sdrc_core_r2b_caddr_3_), .Y(u_sdrc_core_u_req_gen__abc_22171_n518) );
  AND2X2 AND2X2_167 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n556), .B(u_sdrc_core_u_bank_ctl__abc_21249_n227_bF_buf2), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n557) );
  AND2X2 AND2X2_1670 ( .A(u_sdrc_core_u_req_gen__abc_22171_n509_1), .B(u_sdrc_core_u_req_gen__abc_22171_n505), .Y(u_sdrc_core_u_req_gen__abc_22171_n519) );
  AND2X2 AND2X2_1671 ( .A(u_sdrc_core_u_req_gen__abc_22171_n222), .B(u_sdrc_core_u_req_gen__abc_22171_n521), .Y(u_sdrc_core_u_req_gen__abc_22171_n523) );
  AND2X2 AND2X2_1672 ( .A(u_sdrc_core_u_req_gen__abc_22171_n524), .B(u_sdrc_core_u_req_gen__abc_22171_n522), .Y(u_sdrc_core_u_req_gen__abc_22171_n525) );
  AND2X2 AND2X2_1673 ( .A(u_sdrc_core_u_req_gen__abc_22171_n526), .B(u_sdrc_core_u_req_gen__abc_22171_n528), .Y(u_sdrc_core_u_req_gen__abc_22171_n529_1) );
  AND2X2 AND2X2_1674 ( .A(u_sdrc_core_u_req_gen__abc_22171_n529_1), .B(u_sdrc_core_u_req_gen__abc_22171_n335_1_bF_buf1), .Y(u_sdrc_core_u_req_gen__abc_22171_n530) );
  AND2X2 AND2X2_1675 ( .A(u_sdrc_core_u_req_gen__abc_22171_n531), .B(u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf3), .Y(u_sdrc_core_u_req_gen__abc_22171_n532) );
  AND2X2 AND2X2_1676 ( .A(u_sdrc_core_u_req_gen__abc_22171_n533), .B(app_req_ack_bF_buf0), .Y(u_sdrc_core_u_req_gen__abc_22171_n534) );
  AND2X2 AND2X2_1677 ( .A(u_sdrc_core_u_req_gen__abc_22171_n287), .B(app_req_ack_bF_buf6), .Y(u_sdrc_core_u_req_gen__abc_22171_n536) );
  AND2X2 AND2X2_1678 ( .A(u_sdrc_core_u_req_gen__abc_22171_n346_1), .B(u_sdrc_core_r2b_caddr_4_), .Y(u_sdrc_core_u_req_gen__abc_22171_n537) );
  AND2X2 AND2X2_1679 ( .A(u_sdrc_core_r2b_len_4_), .B(u_sdrc_core_r2b_caddr_4_), .Y(u_sdrc_core_u_req_gen__abc_22171_n538) );
  AND2X2 AND2X2_168 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_last), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n594) );
  AND2X2 AND2X2_1680 ( .A(u_sdrc_core_u_req_gen__abc_22171_n539), .B(u_sdrc_core_u_req_gen__abc_22171_n540), .Y(u_sdrc_core_u_req_gen__abc_22171_n541) );
  AND2X2 AND2X2_1681 ( .A(u_sdrc_core_u_req_gen__abc_22171_n525), .B(u_sdrc_core_u_req_gen__abc_22171_n504_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n543) );
  AND2X2 AND2X2_1682 ( .A(u_sdrc_core_u_req_gen__abc_22171_n507_1), .B(u_sdrc_core_u_req_gen__abc_22171_n525), .Y(u_sdrc_core_u_req_gen__abc_22171_n545) );
  AND2X2 AND2X2_1683 ( .A(u_sdrc_core_u_req_gen__abc_22171_n503), .B(u_sdrc_core_u_req_gen__abc_22171_n545), .Y(u_sdrc_core_u_req_gen__abc_22171_n546) );
  AND2X2 AND2X2_1684 ( .A(u_sdrc_core_u_req_gen__abc_22171_n547), .B(u_sdrc_core_u_req_gen__abc_22171_n541), .Y(u_sdrc_core_u_req_gen__abc_22171_n549) );
  AND2X2 AND2X2_1685 ( .A(u_sdrc_core_u_req_gen__abc_22171_n550), .B(u_sdrc_core_u_req_gen__abc_22171_n548), .Y(u_sdrc_core_u_req_gen__abc_22171_n551) );
  AND2X2 AND2X2_1686 ( .A(u_sdrc_core_u_req_gen__abc_22171_n551), .B(u_sdrc_core_u_req_gen__abc_22171_n335_1_bF_buf0), .Y(u_sdrc_core_u_req_gen__abc_22171_n552) );
  AND2X2 AND2X2_1687 ( .A(u_sdrc_core_u_req_gen__abc_22171_n553), .B(u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf2), .Y(u_sdrc_core_u_req_gen__abc_22171_n554) );
  AND2X2 AND2X2_1688 ( .A(u_sdrc_core_u_req_gen__abc_22171_n346_1), .B(u_sdrc_core_r2b_caddr_5_), .Y(u_sdrc_core_u_req_gen__abc_22171_n556) );
  AND2X2 AND2X2_1689 ( .A(u_sdrc_core_u_req_gen__abc_22171_n550), .B(u_sdrc_core_u_req_gen__abc_22171_n539), .Y(u_sdrc_core_u_req_gen__abc_22171_n557) );
  AND2X2 AND2X2_169 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_last), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n595) );
  AND2X2 AND2X2_1690 ( .A(u_sdrc_core_r2b_len_5_), .B(u_sdrc_core_r2b_caddr_5_), .Y(u_sdrc_core_u_req_gen__abc_22171_n559) );
  AND2X2 AND2X2_1691 ( .A(u_sdrc_core_u_req_gen__abc_22171_n560), .B(u_sdrc_core_u_req_gen__abc_22171_n561), .Y(u_sdrc_core_u_req_gen__abc_22171_n562) );
  AND2X2 AND2X2_1692 ( .A(u_sdrc_core_u_req_gen__abc_22171_n563), .B(u_sdrc_core_u_req_gen__abc_22171_n565), .Y(u_sdrc_core_u_req_gen__abc_22171_n566) );
  AND2X2 AND2X2_1693 ( .A(u_sdrc_core_u_req_gen__abc_22171_n566), .B(u_sdrc_core_u_req_gen__abc_22171_n335_1_bF_buf3), .Y(u_sdrc_core_u_req_gen__abc_22171_n567) );
  AND2X2 AND2X2_1694 ( .A(u_sdrc_core_u_req_gen__abc_22171_n568), .B(u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf1), .Y(u_sdrc_core_u_req_gen__abc_22171_n569) );
  AND2X2 AND2X2_1695 ( .A(u_sdrc_core_u_req_gen__abc_22171_n570), .B(app_req_ack_bF_buf5), .Y(u_sdrc_core_u_req_gen__abc_22171_n571) );
  AND2X2 AND2X2_1696 ( .A(u_sdrc_core_u_req_gen__abc_22171_n307_1), .B(app_req_ack_bF_buf4), .Y(u_sdrc_core_u_req_gen__abc_22171_n573) );
  AND2X2 AND2X2_1697 ( .A(u_sdrc_core_u_req_gen__abc_22171_n346_1), .B(u_sdrc_core_r2b_caddr_6_), .Y(u_sdrc_core_u_req_gen__abc_22171_n574) );
  AND2X2 AND2X2_1698 ( .A(u_sdrc_core_u_req_gen__abc_22171_n575), .B(u_sdrc_core_u_req_gen__abc_22171_n561), .Y(u_sdrc_core_u_req_gen__abc_22171_n576) );
  AND2X2 AND2X2_1699 ( .A(u_sdrc_core_u_req_gen__abc_22171_n541), .B(u_sdrc_core_u_req_gen__abc_22171_n562), .Y(u_sdrc_core_u_req_gen__abc_22171_n577) );
  AND2X2 AND2X2_17 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_req), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n236) );
  AND2X2 AND2X2_170 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_xfr_ok), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_last), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n597) );
  AND2X2 AND2X2_1700 ( .A(u_sdrc_core_u_req_gen__abc_22171_n547), .B(u_sdrc_core_u_req_gen__abc_22171_n577), .Y(u_sdrc_core_u_req_gen__abc_22171_n578) );
  AND2X2 AND2X2_1701 ( .A(u_sdrc_core_r2b_len_6_), .B(u_sdrc_core_r2b_caddr_6_), .Y(u_sdrc_core_u_req_gen__abc_22171_n580) );
  AND2X2 AND2X2_1702 ( .A(u_sdrc_core_u_req_gen__abc_22171_n581), .B(u_sdrc_core_u_req_gen__abc_22171_n582), .Y(u_sdrc_core_u_req_gen__abc_22171_n583) );
  AND2X2 AND2X2_1703 ( .A(u_sdrc_core_u_req_gen__abc_22171_n579), .B(u_sdrc_core_u_req_gen__abc_22171_n583), .Y(u_sdrc_core_u_req_gen__abc_22171_n585) );
  AND2X2 AND2X2_1704 ( .A(u_sdrc_core_u_req_gen__abc_22171_n586), .B(u_sdrc_core_u_req_gen__abc_22171_n584), .Y(u_sdrc_core_u_req_gen__abc_22171_n587_1) );
  AND2X2 AND2X2_1705 ( .A(u_sdrc_core_u_req_gen__abc_22171_n587_1), .B(u_sdrc_core_u_req_gen__abc_22171_n335_1_bF_buf2), .Y(u_sdrc_core_u_req_gen__abc_22171_n588_1) );
  AND2X2 AND2X2_1706 ( .A(u_sdrc_core_u_req_gen__abc_22171_n589), .B(u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf0), .Y(u_sdrc_core_u_req_gen__abc_22171_n590) );
  AND2X2 AND2X2_1707 ( .A(u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf3), .B(app_req_addr_7_), .Y(u_sdrc_core_u_req_gen__abc_22171_n592) );
  AND2X2 AND2X2_1708 ( .A(cfg_sdr_width_1_bF_buf5), .B(app_req_addr_5_), .Y(u_sdrc_core_u_req_gen__abc_22171_n593) );
  AND2X2 AND2X2_1709 ( .A(u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf4), .B(app_req_addr_6_), .Y(u_sdrc_core_u_req_gen__abc_22171_n594) );
  AND2X2 AND2X2_171 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_last), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n598) );
  AND2X2 AND2X2_1710 ( .A(u_sdrc_core_u_req_gen__abc_22171_n596), .B(app_req_ack_bF_buf3), .Y(u_sdrc_core_u_req_gen__abc_22171_n597) );
  AND2X2 AND2X2_1711 ( .A(u_sdrc_core_u_req_gen__abc_22171_n586), .B(u_sdrc_core_u_req_gen__abc_22171_n581), .Y(u_sdrc_core_u_req_gen__abc_22171_n599) );
  AND2X2 AND2X2_1712 ( .A(u_sdrc_core_u_req_gen__abc_22171_n601), .B(u_sdrc_core_u_req_gen__abc_22171_n598), .Y(u_sdrc_core_u_req_gen__abc_22171_n602) );
  AND2X2 AND2X2_1713 ( .A(u_sdrc_core_u_req_gen__abc_22171_n600), .B(u_sdrc_core_r2b_caddr_7_), .Y(u_sdrc_core_u_req_gen__abc_22171_n603) );
  AND2X2 AND2X2_1714 ( .A(u_sdrc_core_u_req_gen__abc_22171_n604), .B(u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf4), .Y(u_sdrc_core_u_req_gen__abc_22171_n605) );
  AND2X2 AND2X2_1715 ( .A(u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf2), .B(app_req_addr_8_), .Y(u_sdrc_core_u_req_gen__abc_22171_n607) );
  AND2X2 AND2X2_1716 ( .A(cfg_sdr_width_1_bF_buf4), .B(app_req_addr_6_), .Y(u_sdrc_core_u_req_gen__abc_22171_n608) );
  AND2X2 AND2X2_1717 ( .A(u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf3), .B(app_req_addr_7_), .Y(u_sdrc_core_u_req_gen__abc_22171_n609) );
  AND2X2 AND2X2_1718 ( .A(u_sdrc_core_u_req_gen__abc_22171_n611), .B(app_req_ack_bF_buf2), .Y(u_sdrc_core_u_req_gen__abc_22171_n612) );
  AND2X2 AND2X2_1719 ( .A(u_sdrc_core_u_req_gen__abc_22171_n583), .B(u_sdrc_core_r2b_caddr_7_), .Y(u_sdrc_core_u_req_gen__abc_22171_n613) );
  AND2X2 AND2X2_172 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_wrap), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n608) );
  AND2X2 AND2X2_1720 ( .A(u_sdrc_core_u_req_gen__abc_22171_n577), .B(u_sdrc_core_u_req_gen__abc_22171_n613), .Y(u_sdrc_core_u_req_gen__abc_22171_n614) );
  AND2X2 AND2X2_1721 ( .A(u_sdrc_core_u_req_gen__abc_22171_n547), .B(u_sdrc_core_u_req_gen__abc_22171_n614), .Y(u_sdrc_core_u_req_gen__abc_22171_n615) );
  AND2X2 AND2X2_1722 ( .A(u_sdrc_core_u_req_gen__abc_22171_n582), .B(u_sdrc_core_r2b_caddr_7_), .Y(u_sdrc_core_u_req_gen__abc_22171_n617) );
  AND2X2 AND2X2_1723 ( .A(u_sdrc_core_u_req_gen__abc_22171_n616), .B(u_sdrc_core_u_req_gen__abc_22171_n617), .Y(u_sdrc_core_u_req_gen__abc_22171_n618) );
  AND2X2 AND2X2_1724 ( .A(u_sdrc_core_u_req_gen__abc_22171_n619), .B(u_sdrc_core_u_req_gen__abc_22171_n335_1_bF_buf1), .Y(u_sdrc_core_u_req_gen__abc_22171_n620) );
  AND2X2 AND2X2_1725 ( .A(u_sdrc_core_u_req_gen__abc_22171_n620), .B(u_sdrc_core_u_req_gen_curr_sdr_addr_8_), .Y(u_sdrc_core_u_req_gen__abc_22171_n622) );
  AND2X2 AND2X2_1726 ( .A(u_sdrc_core_u_req_gen__abc_22171_n623), .B(u_sdrc_core_u_req_gen__abc_22171_n621), .Y(u_sdrc_core_u_req_gen__abc_22171_n624) );
  AND2X2 AND2X2_1727 ( .A(u_sdrc_core_u_req_gen__abc_22171_n624), .B(u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf3), .Y(u_sdrc_core_u_req_gen__abc_22171_n625) );
  AND2X2 AND2X2_1728 ( .A(u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf1), .B(app_req_addr_9_), .Y(u_sdrc_core_u_req_gen__abc_22171_n627) );
  AND2X2 AND2X2_1729 ( .A(cfg_sdr_width_1_bF_buf3), .B(app_req_addr_7_), .Y(u_sdrc_core_u_req_gen__abc_22171_n628) );
  AND2X2 AND2X2_173 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_wrap), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n609) );
  AND2X2 AND2X2_1730 ( .A(u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf2), .B(app_req_addr_8_), .Y(u_sdrc_core_u_req_gen__abc_22171_n629) );
  AND2X2 AND2X2_1731 ( .A(u_sdrc_core_u_req_gen__abc_22171_n631), .B(app_req_ack_bF_buf1), .Y(u_sdrc_core_u_req_gen__abc_22171_n632) );
  AND2X2 AND2X2_1732 ( .A(u_sdrc_core_u_req_gen_curr_sdr_addr_8_), .B(u_sdrc_core_u_req_gen_curr_sdr_addr_9_), .Y(u_sdrc_core_u_req_gen__abc_22171_n634) );
  AND2X2 AND2X2_1733 ( .A(u_sdrc_core_u_req_gen__abc_22171_n620), .B(u_sdrc_core_u_req_gen__abc_22171_n634), .Y(u_sdrc_core_u_req_gen__abc_22171_n635) );
  AND2X2 AND2X2_1734 ( .A(u_sdrc_core_u_req_gen__abc_22171_n636), .B(u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf2), .Y(u_sdrc_core_u_req_gen__abc_22171_n637) );
  AND2X2 AND2X2_1735 ( .A(u_sdrc_core_u_req_gen__abc_22171_n637), .B(u_sdrc_core_u_req_gen__abc_22171_n633), .Y(u_sdrc_core_u_req_gen__abc_22171_n638) );
  AND2X2 AND2X2_1736 ( .A(u_sdrc_core_u_req_gen__abc_22171_n642), .B(u_sdrc_core_u_req_gen__abc_22171_n641), .Y(u_sdrc_core_u_req_gen__abc_22171_n643) );
  AND2X2 AND2X2_1737 ( .A(u_sdrc_core_u_req_gen__abc_22171_n643), .B(u_sdrc_core_u_req_gen__abc_22171_n640), .Y(u_sdrc_core_u_req_gen__abc_22171_n644) );
  AND2X2 AND2X2_1738 ( .A(u_sdrc_core_u_req_gen__abc_22171_n644), .B(app_req_ack_bF_buf0), .Y(u_sdrc_core_u_req_gen__abc_22171_n645) );
  AND2X2 AND2X2_1739 ( .A(u_sdrc_core_u_req_gen__abc_22171_n635), .B(u_sdrc_core_u_req_gen_curr_sdr_addr_10_), .Y(u_sdrc_core_u_req_gen__abc_22171_n646) );
  AND2X2 AND2X2_174 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_xfr_ok), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_wrap), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n611) );
  AND2X2 AND2X2_1740 ( .A(u_sdrc_core_u_req_gen__abc_22171_n648), .B(u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf1), .Y(u_sdrc_core_u_req_gen__abc_22171_n649) );
  AND2X2 AND2X2_1741 ( .A(u_sdrc_core_u_req_gen__abc_22171_n649), .B(u_sdrc_core_u_req_gen__abc_22171_n647), .Y(u_sdrc_core_u_req_gen__abc_22171_n650) );
  AND2X2 AND2X2_1742 ( .A(u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf0), .B(app_req_addr_11_), .Y(u_sdrc_core_u_req_gen__abc_22171_n652) );
  AND2X2 AND2X2_1743 ( .A(u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf1), .B(app_req_addr_10_), .Y(u_sdrc_core_u_req_gen__abc_22171_n653) );
  AND2X2 AND2X2_1744 ( .A(cfg_sdr_width_1_bF_buf2), .B(app_req_addr_9_), .Y(u_sdrc_core_u_req_gen__abc_22171_n654) );
  AND2X2 AND2X2_1745 ( .A(u_sdrc_core_u_req_gen__abc_22171_n656), .B(app_req_ack_bF_buf6), .Y(u_sdrc_core_u_req_gen__abc_22171_n657) );
  AND2X2 AND2X2_1746 ( .A(u_sdrc_core_u_req_gen_curr_sdr_addr_10_), .B(u_sdrc_core_u_req_gen_curr_sdr_addr_11_), .Y(u_sdrc_core_u_req_gen__abc_22171_n658) );
  AND2X2 AND2X2_1747 ( .A(u_sdrc_core_u_req_gen__abc_22171_n634), .B(u_sdrc_core_u_req_gen__abc_22171_n658), .Y(u_sdrc_core_u_req_gen__abc_22171_n659) );
  AND2X2 AND2X2_1748 ( .A(u_sdrc_core_u_req_gen__abc_22171_n620), .B(u_sdrc_core_u_req_gen__abc_22171_n659), .Y(u_sdrc_core_u_req_gen__abc_22171_n660) );
  AND2X2 AND2X2_1749 ( .A(u_sdrc_core_u_req_gen__abc_22171_n662), .B(u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf0), .Y(u_sdrc_core_u_req_gen__abc_22171_n663) );
  AND2X2 AND2X2_175 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_wrap), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n612) );
  AND2X2 AND2X2_1750 ( .A(u_sdrc_core_u_req_gen__abc_22171_n663), .B(u_sdrc_core_u_req_gen__abc_22171_n661), .Y(u_sdrc_core_u_req_gen__abc_22171_n664) );
  AND2X2 AND2X2_1751 ( .A(u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf4), .B(app_req_addr_12_), .Y(u_sdrc_core_u_req_gen__abc_22171_n666) );
  AND2X2 AND2X2_1752 ( .A(cfg_sdr_width_1_bF_buf1), .B(app_req_addr_10_), .Y(u_sdrc_core_u_req_gen__abc_22171_n667) );
  AND2X2 AND2X2_1753 ( .A(u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf0), .B(app_req_addr_11_), .Y(u_sdrc_core_u_req_gen__abc_22171_n668) );
  AND2X2 AND2X2_1754 ( .A(u_sdrc_core_u_req_gen__abc_22171_n670), .B(app_req_ack_bF_buf5), .Y(u_sdrc_core_u_req_gen__abc_22171_n671) );
  AND2X2 AND2X2_1755 ( .A(u_sdrc_core_u_req_gen__abc_22171_n660), .B(u_sdrc_core_u_req_gen_curr_sdr_addr_12_), .Y(u_sdrc_core_u_req_gen__abc_22171_n672) );
  AND2X2 AND2X2_1756 ( .A(u_sdrc_core_u_req_gen__abc_22171_n673), .B(u_sdrc_core_u_req_gen__abc_22171_n674), .Y(u_sdrc_core_u_req_gen__abc_22171_n675) );
  AND2X2 AND2X2_1757 ( .A(u_sdrc_core_u_req_gen__abc_22171_n675), .B(u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf4), .Y(u_sdrc_core_u_req_gen__abc_22171_n676) );
  AND2X2 AND2X2_1758 ( .A(u_sdrc_core_u_req_gen_curr_sdr_addr_12_), .B(u_sdrc_core_u_req_gen_curr_sdr_addr_13_), .Y(u_sdrc_core_u_req_gen__abc_22171_n679) );
  AND2X2 AND2X2_1759 ( .A(u_sdrc_core_u_req_gen__abc_22171_n659), .B(u_sdrc_core_u_req_gen__abc_22171_n679), .Y(u_sdrc_core_u_req_gen__abc_22171_n680) );
  AND2X2 AND2X2_176 ( .A(u_sdrc_core_u_bank_ctl_rank_cnt_1_), .B(\cfg_req_depth[1] ), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n615) );
  AND2X2 AND2X2_1760 ( .A(u_sdrc_core_u_req_gen__abc_22171_n620), .B(u_sdrc_core_u_req_gen__abc_22171_n680), .Y(u_sdrc_core_u_req_gen__abc_22171_n681) );
  AND2X2 AND2X2_1761 ( .A(u_sdrc_core_u_req_gen__abc_22171_n678), .B(u_sdrc_core_u_req_gen__abc_22171_n682), .Y(u_sdrc_core_u_req_gen__abc_22171_n683) );
  AND2X2 AND2X2_1762 ( .A(u_sdrc_core_u_req_gen__abc_22171_n683), .B(u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf3), .Y(u_sdrc_core_u_req_gen__abc_22171_n684) );
  AND2X2 AND2X2_1763 ( .A(u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf3), .B(app_req_addr_13_), .Y(u_sdrc_core_u_req_gen__abc_22171_n685) );
  AND2X2 AND2X2_1764 ( .A(cfg_sdr_width_1_bF_buf0), .B(app_req_addr_11_), .Y(u_sdrc_core_u_req_gen__abc_22171_n686) );
  AND2X2 AND2X2_1765 ( .A(u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf4), .B(app_req_addr_12_), .Y(u_sdrc_core_u_req_gen__abc_22171_n687) );
  AND2X2 AND2X2_1766 ( .A(u_sdrc_core_u_req_gen__abc_22171_n689), .B(app_req_ack_bF_buf4), .Y(u_sdrc_core_u_req_gen__abc_22171_n690) );
  AND2X2 AND2X2_1767 ( .A(u_sdrc_core_u_req_gen__abc_22171_n681), .B(u_sdrc_core_u_req_gen_curr_sdr_addr_14_), .Y(u_sdrc_core_u_req_gen__abc_22171_n693) );
  AND2X2 AND2X2_1768 ( .A(u_sdrc_core_u_req_gen__abc_22171_n694), .B(u_sdrc_core_u_req_gen__abc_22171_n692), .Y(u_sdrc_core_u_req_gen__abc_22171_n695) );
  AND2X2 AND2X2_1769 ( .A(u_sdrc_core_u_req_gen__abc_22171_n695), .B(u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf2), .Y(u_sdrc_core_u_req_gen__abc_22171_n696) );
  AND2X2 AND2X2_177 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n616), .B(u_sdrc_core_u_bank_ctl__abc_21249_n617), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n618) );
  AND2X2 AND2X2_1770 ( .A(u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf2), .B(app_req_addr_14_), .Y(u_sdrc_core_u_req_gen__abc_22171_n697) );
  AND2X2 AND2X2_1771 ( .A(cfg_sdr_width_1_bF_buf5), .B(app_req_addr_12_), .Y(u_sdrc_core_u_req_gen__abc_22171_n698) );
  AND2X2 AND2X2_1772 ( .A(u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf3), .B(app_req_addr_13_), .Y(u_sdrc_core_u_req_gen__abc_22171_n699) );
  AND2X2 AND2X2_1773 ( .A(u_sdrc_core_u_req_gen__abc_22171_n701), .B(app_req_ack_bF_buf3), .Y(u_sdrc_core_u_req_gen__abc_22171_n702) );
  AND2X2 AND2X2_1774 ( .A(u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf1), .B(app_req_addr_15_), .Y(u_sdrc_core_u_req_gen__abc_22171_n704) );
  AND2X2 AND2X2_1775 ( .A(u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf2), .B(app_req_addr_14_), .Y(u_sdrc_core_u_req_gen__abc_22171_n705) );
  AND2X2 AND2X2_1776 ( .A(cfg_sdr_width_1_bF_buf4), .B(app_req_addr_13_), .Y(u_sdrc_core_u_req_gen__abc_22171_n706) );
  AND2X2 AND2X2_1777 ( .A(u_sdrc_core_u_req_gen__abc_22171_n708), .B(app_req_ack_bF_buf2), .Y(u_sdrc_core_u_req_gen__abc_22171_n709) );
  AND2X2 AND2X2_1778 ( .A(u_sdrc_core_u_req_gen_curr_sdr_addr_14_), .B(u_sdrc_core_u_req_gen_curr_sdr_addr_15_), .Y(u_sdrc_core_u_req_gen__abc_22171_n711) );
  AND2X2 AND2X2_1779 ( .A(u_sdrc_core_u_req_gen__abc_22171_n680), .B(u_sdrc_core_u_req_gen__abc_22171_n711), .Y(u_sdrc_core_u_req_gen__abc_22171_n712) );
  AND2X2 AND2X2_178 ( .A(u_sdrc_core_u_bank_ctl_rank_cnt_0_), .B(\cfg_req_depth[0] ), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n619) );
  AND2X2 AND2X2_1780 ( .A(u_sdrc_core_u_req_gen__abc_22171_n619), .B(u_sdrc_core_u_req_gen__abc_22171_n712), .Y(u_sdrc_core_u_req_gen__abc_22171_n713) );
  AND2X2 AND2X2_1781 ( .A(u_sdrc_core_u_req_gen__abc_22171_n713), .B(u_sdrc_core_u_req_gen__abc_22171_n335_1_bF_buf0), .Y(u_sdrc_core_u_req_gen__abc_22171_n714) );
  AND2X2 AND2X2_1782 ( .A(u_sdrc_core_u_req_gen__abc_22171_n715), .B(u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf1), .Y(u_sdrc_core_u_req_gen__abc_22171_n716) );
  AND2X2 AND2X2_1783 ( .A(u_sdrc_core_u_req_gen__abc_22171_n710), .B(u_sdrc_core_u_req_gen__abc_22171_n716), .Y(u_sdrc_core_u_req_gen__abc_22171_n717) );
  AND2X2 AND2X2_1784 ( .A(u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf0), .B(app_req_addr_16_), .Y(u_sdrc_core_u_req_gen__abc_22171_n719) );
  AND2X2 AND2X2_1785 ( .A(cfg_sdr_width_1_bF_buf3), .B(app_req_addr_14_), .Y(u_sdrc_core_u_req_gen__abc_22171_n720) );
  AND2X2 AND2X2_1786 ( .A(u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf1), .B(app_req_addr_15_), .Y(u_sdrc_core_u_req_gen__abc_22171_n721) );
  AND2X2 AND2X2_1787 ( .A(u_sdrc_core_u_req_gen__abc_22171_n723), .B(app_req_ack_bF_buf1), .Y(u_sdrc_core_u_req_gen__abc_22171_n724) );
  AND2X2 AND2X2_1788 ( .A(u_sdrc_core_u_req_gen__abc_22171_n714), .B(u_sdrc_core_u_req_gen_curr_sdr_addr_16_), .Y(u_sdrc_core_u_req_gen__abc_22171_n725) );
  AND2X2 AND2X2_1789 ( .A(u_sdrc_core_u_req_gen__abc_22171_n726), .B(u_sdrc_core_u_req_gen__abc_22171_n727), .Y(u_sdrc_core_u_req_gen__abc_22171_n728) );
  AND2X2 AND2X2_179 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n620), .B(u_sdrc_core_u_bank_ctl__abc_21249_n621), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n622) );
  AND2X2 AND2X2_1790 ( .A(u_sdrc_core_u_req_gen__abc_22171_n728), .B(u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf0), .Y(u_sdrc_core_u_req_gen__abc_22171_n729) );
  AND2X2 AND2X2_1791 ( .A(u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf4), .B(app_req_addr_17_), .Y(u_sdrc_core_u_req_gen__abc_22171_n731) );
  AND2X2 AND2X2_1792 ( .A(u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf0), .B(app_req_addr_16_), .Y(u_sdrc_core_u_req_gen__abc_22171_n732) );
  AND2X2 AND2X2_1793 ( .A(cfg_sdr_width_1_bF_buf2), .B(app_req_addr_15_), .Y(u_sdrc_core_u_req_gen__abc_22171_n733) );
  AND2X2 AND2X2_1794 ( .A(u_sdrc_core_u_req_gen__abc_22171_n735), .B(app_req_ack_bF_buf0), .Y(u_sdrc_core_u_req_gen__abc_22171_n736) );
  AND2X2 AND2X2_1795 ( .A(u_sdrc_core_u_req_gen_curr_sdr_addr_16_), .B(u_sdrc_core_u_req_gen_curr_sdr_addr_17_), .Y(u_sdrc_core_u_req_gen__abc_22171_n737) );
  AND2X2 AND2X2_1796 ( .A(u_sdrc_core_u_req_gen__abc_22171_n714), .B(u_sdrc_core_u_req_gen__abc_22171_n737), .Y(u_sdrc_core_u_req_gen__abc_22171_n738) );
  AND2X2 AND2X2_1797 ( .A(u_sdrc_core_u_req_gen__abc_22171_n740), .B(u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf4), .Y(u_sdrc_core_u_req_gen__abc_22171_n741) );
  AND2X2 AND2X2_1798 ( .A(u_sdrc_core_u_req_gen__abc_22171_n741), .B(u_sdrc_core_u_req_gen__abc_22171_n739), .Y(u_sdrc_core_u_req_gen__abc_22171_n742) );
  AND2X2 AND2X2_1799 ( .A(u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf3), .B(app_req_addr_18_), .Y(u_sdrc_core_u_req_gen__abc_22171_n744) );
  AND2X2 AND2X2_18 ( .A(u_sdrc_core_b2x_req), .B(u_sdrc_core_u_bank_ctl_x2b_ack_bF_buf3), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n240_1) );
  AND2X2 AND2X2_180 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n623), .B(u_sdrc_core_u_bank_ctl__abc_21249_n216_1), .Y(u_sdrc_core_b2r_arb_ok) );
  AND2X2 AND2X2_1800 ( .A(u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf4), .B(app_req_addr_17_), .Y(u_sdrc_core_u_req_gen__abc_22171_n745) );
  AND2X2 AND2X2_1801 ( .A(cfg_sdr_width_1_bF_buf1), .B(app_req_addr_16_), .Y(u_sdrc_core_u_req_gen__abc_22171_n746) );
  AND2X2 AND2X2_1802 ( .A(u_sdrc_core_u_req_gen__abc_22171_n748), .B(app_req_ack_bF_buf6), .Y(u_sdrc_core_u_req_gen__abc_22171_n749) );
  AND2X2 AND2X2_1803 ( .A(u_sdrc_core_u_req_gen__abc_22171_n739), .B(u_sdrc_core_u_req_gen_curr_sdr_addr_18_), .Y(u_sdrc_core_u_req_gen__abc_22171_n750) );
  AND2X2 AND2X2_1804 ( .A(u_sdrc_core_u_req_gen__abc_22171_n738), .B(u_sdrc_core_u_req_gen__abc_22171_n751), .Y(u_sdrc_core_u_req_gen__abc_22171_n752) );
  AND2X2 AND2X2_1805 ( .A(u_sdrc_core_u_req_gen__abc_22171_n753), .B(u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf3), .Y(u_sdrc_core_u_req_gen__abc_22171_n754) );
  AND2X2 AND2X2_1806 ( .A(u_sdrc_core_u_req_gen__abc_22171_n737), .B(u_sdrc_core_u_req_gen_curr_sdr_addr_18_), .Y(u_sdrc_core_u_req_gen__abc_22171_n756) );
  AND2X2 AND2X2_1807 ( .A(u_sdrc_core_u_req_gen__abc_22171_n714), .B(u_sdrc_core_u_req_gen__abc_22171_n756), .Y(u_sdrc_core_u_req_gen__abc_22171_n757) );
  AND2X2 AND2X2_1808 ( .A(u_sdrc_core_u_req_gen__abc_22171_n756), .B(u_sdrc_core_u_req_gen_curr_sdr_addr_19_), .Y(u_sdrc_core_u_req_gen__abc_22171_n759) );
  AND2X2 AND2X2_1809 ( .A(u_sdrc_core_u_req_gen__abc_22171_n713), .B(u_sdrc_core_u_req_gen__abc_22171_n759), .Y(u_sdrc_core_u_req_gen__abc_22171_n760) );
  AND2X2 AND2X2_181 ( .A(u_sdrc_core_b2r_arb_ok), .B(u_sdrc_core_r2b_req), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n627) );
  AND2X2 AND2X2_1810 ( .A(u_sdrc_core_u_req_gen__abc_22171_n760), .B(u_sdrc_core_u_req_gen__abc_22171_n335_1_bF_buf3), .Y(u_sdrc_core_u_req_gen__abc_22171_n761) );
  AND2X2 AND2X2_1811 ( .A(u_sdrc_core_u_req_gen__abc_22171_n758), .B(u_sdrc_core_u_req_gen__abc_22171_n762), .Y(u_sdrc_core_u_req_gen__abc_22171_n763) );
  AND2X2 AND2X2_1812 ( .A(u_sdrc_core_u_req_gen__abc_22171_n763), .B(u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf2), .Y(u_sdrc_core_u_req_gen__abc_22171_n764) );
  AND2X2 AND2X2_1813 ( .A(u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf2), .B(app_req_addr_19_), .Y(u_sdrc_core_u_req_gen__abc_22171_n765) );
  AND2X2 AND2X2_1814 ( .A(cfg_sdr_width_1_bF_buf0), .B(app_req_addr_17_), .Y(u_sdrc_core_u_req_gen__abc_22171_n766) );
  AND2X2 AND2X2_1815 ( .A(u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf3), .B(app_req_addr_18_), .Y(u_sdrc_core_u_req_gen__abc_22171_n767) );
  AND2X2 AND2X2_1816 ( .A(u_sdrc_core_u_req_gen__abc_22171_n769), .B(app_req_ack_bF_buf5), .Y(u_sdrc_core_u_req_gen__abc_22171_n770) );
  AND2X2 AND2X2_1817 ( .A(u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf1), .B(app_req_addr_20_), .Y(u_sdrc_core_u_req_gen__abc_22171_n772) );
  AND2X2 AND2X2_1818 ( .A(u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf2), .B(app_req_addr_19_), .Y(u_sdrc_core_u_req_gen__abc_22171_n773) );
  AND2X2 AND2X2_1819 ( .A(cfg_sdr_width_1_bF_buf5), .B(app_req_addr_18_), .Y(u_sdrc_core_u_req_gen__abc_22171_n774) );
  AND2X2 AND2X2_182 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n627), .B(u_sdrc_core_u_bank_ctl__abc_21249_n626), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n628) );
  AND2X2 AND2X2_1820 ( .A(u_sdrc_core_u_req_gen__abc_22171_n776), .B(app_req_ack_bF_buf4), .Y(u_sdrc_core_u_req_gen__abc_22171_n777) );
  AND2X2 AND2X2_1821 ( .A(u_sdrc_core_u_req_gen__abc_22171_n759), .B(u_sdrc_core_u_req_gen_curr_sdr_addr_20_), .Y(u_sdrc_core_u_req_gen__abc_22171_n779) );
  AND2X2 AND2X2_1822 ( .A(u_sdrc_core_u_req_gen__abc_22171_n714), .B(u_sdrc_core_u_req_gen__abc_22171_n779), .Y(u_sdrc_core_u_req_gen__abc_22171_n780) );
  AND2X2 AND2X2_1823 ( .A(u_sdrc_core_u_req_gen__abc_22171_n781), .B(u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf1), .Y(u_sdrc_core_u_req_gen__abc_22171_n782) );
  AND2X2 AND2X2_1824 ( .A(u_sdrc_core_u_req_gen__abc_22171_n782), .B(u_sdrc_core_u_req_gen__abc_22171_n778), .Y(u_sdrc_core_u_req_gen__abc_22171_n783) );
  AND2X2 AND2X2_1825 ( .A(cfg_sdr_width_1_bF_buf4), .B(app_req_addr_19_), .Y(u_sdrc_core_u_req_gen__abc_22171_n785) );
  AND2X2 AND2X2_1826 ( .A(app_req_ack_bF_buf3), .B(u_sdrc_core_u_req_gen__abc_22171_n786), .Y(u_sdrc_core_u_req_gen__abc_22171_n787) );
  AND2X2 AND2X2_1827 ( .A(u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf0), .B(app_req_addr_21_), .Y(u_sdrc_core_u_req_gen__abc_22171_n788) );
  AND2X2 AND2X2_1828 ( .A(u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf1), .B(app_req_addr_20_), .Y(u_sdrc_core_u_req_gen__abc_22171_n789) );
  AND2X2 AND2X2_1829 ( .A(u_sdrc_core_u_req_gen__abc_22171_n791), .B(u_sdrc_core_u_req_gen__abc_22171_n787), .Y(u_sdrc_core_u_req_gen__abc_22171_n792) );
  AND2X2 AND2X2_183 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n628), .B(u_sdrc_core_u_bank_ctl__abc_21249_n625), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_r2b_req) );
  AND2X2 AND2X2_1830 ( .A(u_sdrc_core_u_req_gen__abc_22171_n780), .B(u_sdrc_core_u_req_gen_curr_sdr_addr_21_), .Y(u_sdrc_core_u_req_gen__abc_22171_n795) );
  AND2X2 AND2X2_1831 ( .A(u_sdrc_core_u_req_gen__abc_22171_n796), .B(u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf0), .Y(u_sdrc_core_u_req_gen__abc_22171_n797) );
  AND2X2 AND2X2_1832 ( .A(u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf4), .B(app_req_addr_22_), .Y(u_sdrc_core_u_req_gen__abc_22171_n800) );
  AND2X2 AND2X2_1833 ( .A(cfg_sdr_width_1_bF_buf3), .B(app_req_addr_20_), .Y(u_sdrc_core_u_req_gen__abc_22171_n801) );
  AND2X2 AND2X2_1834 ( .A(u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf0), .B(app_req_addr_21_), .Y(u_sdrc_core_u_req_gen__abc_22171_n802) );
  AND2X2 AND2X2_1835 ( .A(u_sdrc_core_u_req_gen__abc_22171_n805), .B(app_req_ack_bF_buf2), .Y(u_sdrc_core_u_req_gen__abc_22171_n806) );
  AND2X2 AND2X2_1836 ( .A(u_sdrc_core_u_req_gen__abc_22171_n795), .B(u_sdrc_core_u_req_gen__abc_22171_n807), .Y(u_sdrc_core_u_req_gen__abc_22171_n808) );
  AND2X2 AND2X2_1837 ( .A(u_sdrc_core_u_req_gen__abc_22171_n810), .B(u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf4), .Y(u_sdrc_core_u_req_gen__abc_22171_n811) );
  AND2X2 AND2X2_1838 ( .A(u_sdrc_core_u_req_gen__abc_22171_n811), .B(u_sdrc_core_u_req_gen__abc_22171_n809), .Y(u_sdrc_core_u_req_gen__abc_22171_n812) );
  AND2X2 AND2X2_1839 ( .A(u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf3), .B(app_req_addr_23_), .Y(u_sdrc_core_u_req_gen__abc_22171_n815) );
  AND2X2 AND2X2_184 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n628), .B(u_sdrc_core_r2b_ba_0_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_r2b_req) );
  AND2X2 AND2X2_1840 ( .A(u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf4), .B(app_req_addr_22_), .Y(u_sdrc_core_u_req_gen__abc_22171_n816) );
  AND2X2 AND2X2_1841 ( .A(cfg_sdr_width_1_bF_buf2), .B(app_req_addr_21_), .Y(u_sdrc_core_u_req_gen__abc_22171_n817) );
  AND2X2 AND2X2_1842 ( .A(u_sdrc_core_u_req_gen__abc_22171_n819), .B(app_req_ack_bF_buf1), .Y(u_sdrc_core_u_req_gen__abc_22171_n820) );
  AND2X2 AND2X2_1843 ( .A(u_sdrc_core_u_req_gen_curr_sdr_addr_20_), .B(u_sdrc_core_u_req_gen_curr_sdr_addr_21_), .Y(u_sdrc_core_u_req_gen__abc_22171_n823) );
  AND2X2 AND2X2_1844 ( .A(u_sdrc_core_u_req_gen__abc_22171_n823), .B(u_sdrc_core_u_req_gen_curr_sdr_addr_22_), .Y(u_sdrc_core_u_req_gen__abc_22171_n824) );
  AND2X2 AND2X2_1845 ( .A(u_sdrc_core_u_req_gen__abc_22171_n761), .B(u_sdrc_core_u_req_gen__abc_22171_n824), .Y(u_sdrc_core_u_req_gen__abc_22171_n825) );
  AND2X2 AND2X2_1846 ( .A(u_sdrc_core_u_req_gen__abc_22171_n826), .B(u_sdrc_core_u_req_gen__abc_22171_n822), .Y(u_sdrc_core_u_req_gen__abc_22171_n827) );
  AND2X2 AND2X2_1847 ( .A(u_sdrc_core_u_req_gen__abc_22171_n825), .B(u_sdrc_core_u_req_gen_curr_sdr_addr_23_), .Y(u_sdrc_core_u_req_gen__abc_22171_n828) );
  AND2X2 AND2X2_1848 ( .A(u_sdrc_core_u_req_gen__abc_22171_n830), .B(u_sdrc_core_u_req_gen__abc_22171_n821), .Y(u_sdrc_core_u_req_gen__abc_22171_n831) );
  AND2X2 AND2X2_1849 ( .A(u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf2), .B(app_req_addr_24_), .Y(u_sdrc_core_u_req_gen__abc_22171_n833) );
  AND2X2 AND2X2_185 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n627), .B(u_sdrc_core_r2b_ba_1_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n631) );
  AND2X2 AND2X2_1850 ( .A(u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf3), .B(app_req_addr_23_), .Y(u_sdrc_core_u_req_gen__abc_22171_n834) );
  AND2X2 AND2X2_1851 ( .A(cfg_sdr_width_1_bF_buf1), .B(app_req_addr_22_), .Y(u_sdrc_core_u_req_gen__abc_22171_n835) );
  AND2X2 AND2X2_1852 ( .A(u_sdrc_core_u_req_gen__abc_22171_n837), .B(app_req_ack_bF_buf6), .Y(u_sdrc_core_u_req_gen__abc_22171_n838) );
  AND2X2 AND2X2_1853 ( .A(u_sdrc_core_u_req_gen_curr_sdr_addr_22_), .B(u_sdrc_core_u_req_gen_curr_sdr_addr_23_), .Y(u_sdrc_core_u_req_gen__abc_22171_n841) );
  AND2X2 AND2X2_1854 ( .A(u_sdrc_core_u_req_gen__abc_22171_n823), .B(u_sdrc_core_u_req_gen__abc_22171_n841), .Y(u_sdrc_core_u_req_gen__abc_22171_n842) );
  AND2X2 AND2X2_1855 ( .A(u_sdrc_core_u_req_gen__abc_22171_n760), .B(u_sdrc_core_u_req_gen__abc_22171_n842), .Y(u_sdrc_core_u_req_gen__abc_22171_n843) );
  AND2X2 AND2X2_1856 ( .A(u_sdrc_core_u_req_gen__abc_22171_n843), .B(u_sdrc_core_u_req_gen__abc_22171_n335_1_bF_buf2), .Y(u_sdrc_core_u_req_gen__abc_22171_n844) );
  AND2X2 AND2X2_1857 ( .A(u_sdrc_core_u_req_gen__abc_22171_n845), .B(u_sdrc_core_u_req_gen__abc_22171_n840), .Y(u_sdrc_core_u_req_gen__abc_22171_n846) );
  AND2X2 AND2X2_1858 ( .A(u_sdrc_core_u_req_gen__abc_22171_n844), .B(u_sdrc_core_u_req_gen_curr_sdr_addr_24_), .Y(u_sdrc_core_u_req_gen__abc_22171_n847) );
  AND2X2 AND2X2_1859 ( .A(u_sdrc_core_u_req_gen__abc_22171_n849), .B(u_sdrc_core_u_req_gen__abc_22171_n839), .Y(u_sdrc_core_u_req_gen__abc_22171_n850) );
  AND2X2 AND2X2_186 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n631), .B(u_sdrc_core_u_bank_ctl__abc_21249_n625), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_r2b_req) );
  AND2X2 AND2X2_1860 ( .A(u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf1), .B(app_req_addr_25_), .Y(u_sdrc_core_u_req_gen__abc_22171_n852) );
  AND2X2 AND2X2_1861 ( .A(u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf2), .B(app_req_addr_24_), .Y(u_sdrc_core_u_req_gen__abc_22171_n853) );
  AND2X2 AND2X2_1862 ( .A(cfg_sdr_width_1_bF_buf0), .B(app_req_addr_23_), .Y(u_sdrc_core_u_req_gen__abc_22171_n854) );
  AND2X2 AND2X2_1863 ( .A(u_sdrc_core_u_req_gen__abc_22171_n856), .B(app_req_ack_bF_buf4), .Y(u_sdrc_core_u_req_gen__abc_22171_n857) );
  AND2X2 AND2X2_1864 ( .A(u_sdrc_core_u_req_gen_curr_sdr_addr_23_), .B(u_sdrc_core_u_req_gen_curr_sdr_addr_24_), .Y(u_sdrc_core_u_req_gen__abc_22171_n860) );
  AND2X2 AND2X2_1865 ( .A(u_sdrc_core_u_req_gen__abc_22171_n335_1_bF_buf1), .B(u_sdrc_core_u_req_gen__abc_22171_n860), .Y(u_sdrc_core_u_req_gen__abc_22171_n861) );
  AND2X2 AND2X2_1866 ( .A(u_sdrc_core_u_req_gen__abc_22171_n861), .B(u_sdrc_core_u_req_gen__abc_22171_n824), .Y(u_sdrc_core_u_req_gen__abc_22171_n862) );
  AND2X2 AND2X2_1867 ( .A(u_sdrc_core_u_req_gen__abc_22171_n760), .B(u_sdrc_core_u_req_gen__abc_22171_n862), .Y(u_sdrc_core_u_req_gen__abc_22171_n863) );
  AND2X2 AND2X2_1868 ( .A(u_sdrc_core_u_req_gen__abc_22171_n866), .B(u_sdrc_core_u_req_gen__abc_22171_n864), .Y(u_sdrc_core_u_req_gen__abc_22171_n867) );
  AND2X2 AND2X2_1869 ( .A(u_sdrc_core_u_req_gen__abc_22171_n868), .B(u_sdrc_core_u_req_gen__abc_22171_n858), .Y(u_sdrc_core_u_req_gen__abc_22171_n869) );
  AND2X2 AND2X2_187 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n631), .B(u_sdrc_core_r2b_ba_0_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_r2b_req) );
  AND2X2 AND2X2_1870 ( .A(\cfg_colbits[0] ), .B(\cfg_colbits[1] ), .Y(u_sdrc_core_u_req_gen__abc_22171_n871) );
  AND2X2 AND2X2_1871 ( .A(u_sdrc_core_u_req_gen_map_address_11_), .B(u_sdrc_core_u_req_gen__abc_22171_n871), .Y(u_sdrc_core_u_req_gen__abc_22171_n872) );
  AND2X2 AND2X2_1872 ( .A(u_sdrc_core_u_req_gen__abc_22171_n873), .B(\cfg_colbits[1] ), .Y(u_sdrc_core_u_req_gen__abc_22171_n874) );
  AND2X2 AND2X2_1873 ( .A(u_sdrc_core_u_req_gen_map_address_10_), .B(u_sdrc_core_u_req_gen__abc_22171_n874), .Y(u_sdrc_core_u_req_gen__abc_22171_n875) );
  AND2X2 AND2X2_1874 ( .A(u_sdrc_core_u_req_gen__abc_22171_n873), .B(u_sdrc_core_u_req_gen__abc_22171_n876), .Y(u_sdrc_core_u_req_gen__abc_22171_n877) );
  AND2X2 AND2X2_1875 ( .A(u_sdrc_core_u_req_gen_map_address_8_), .B(u_sdrc_core_u_req_gen__abc_22171_n877), .Y(u_sdrc_core_u_req_gen__abc_22171_n878) );
  AND2X2 AND2X2_1876 ( .A(u_sdrc_core_u_req_gen__abc_22171_n876), .B(\cfg_colbits[0] ), .Y(u_sdrc_core_u_req_gen__abc_22171_n879) );
  AND2X2 AND2X2_1877 ( .A(u_sdrc_core_u_req_gen_map_address_9_), .B(u_sdrc_core_u_req_gen__abc_22171_n879), .Y(u_sdrc_core_u_req_gen__abc_22171_n880) );
  AND2X2 AND2X2_1878 ( .A(u_sdrc_core_u_req_gen_map_address_11_), .B(u_sdrc_core_u_req_gen__abc_22171_n874), .Y(u_sdrc_core_u_req_gen__abc_22171_n884) );
  AND2X2 AND2X2_1879 ( .A(u_sdrc_core_u_req_gen_map_address_10_), .B(u_sdrc_core_u_req_gen__abc_22171_n876), .Y(u_sdrc_core_u_req_gen__abc_22171_n885) );
  AND2X2 AND2X2_188 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_xfr_ok), .B(u_sdrc_core_u_bank_ctl_x2b_ack_bF_buf2), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_ack) );
  AND2X2 AND2X2_1880 ( .A(u_sdrc_core_u_req_gen__abc_22171_n886), .B(u_sdrc_core_u_req_gen__abc_22171_n887), .Y(u_sdrc_core_u_req_gen__abc_22171_n888) );
  AND2X2 AND2X2_1881 ( .A(u_sdrc_core_u_req_gen_map_address_12_), .B(u_sdrc_core_u_req_gen__abc_22171_n888), .Y(u_sdrc_core_u_req_gen__abc_22171_n889) );
  AND2X2 AND2X2_1882 ( .A(u_sdrc_core_u_req_gen__abc_22171_n892), .B(u_sdrc_core_u_req_gen__abc_22171_n894), .Y(u_sdrc_core_u_req_gen_r2b_ba_1__FF_INPUT) );
  AND2X2 AND2X2_1883 ( .A(u_sdrc_core_u_req_gen_map_address_8_), .B(u_sdrc_core_u_req_gen__abc_22171_n893_bF_buf2), .Y(u_sdrc_core_u_req_gen_r2b_caddr_8__FF_INPUT) );
  AND2X2 AND2X2_1884 ( .A(u_sdrc_core_u_req_gen_map_address_9_), .B(\cfg_colbits[1] ), .Y(u_sdrc_core_u_req_gen_r2b_caddr_9__FF_INPUT) );
  AND2X2 AND2X2_1885 ( .A(u_sdrc_core_u_req_gen_map_address_10_), .B(u_sdrc_core_u_req_gen__abc_22171_n871), .Y(u_sdrc_core_u_req_gen_r2b_caddr_10__FF_INPUT) );
  AND2X2 AND2X2_1886 ( .A(u_sdrc_core_u_req_gen_map_address_11_), .B(u_sdrc_core_u_req_gen__abc_22171_n876), .Y(u_sdrc_core_u_req_gen__abc_22171_n899) );
  AND2X2 AND2X2_1887 ( .A(u_sdrc_core_u_req_gen_map_address_13_), .B(u_sdrc_core_u_req_gen__abc_22171_n888), .Y(u_sdrc_core_u_req_gen__abc_22171_n900) );
  AND2X2 AND2X2_1888 ( .A(u_sdrc_core_u_req_gen_map_address_12_), .B(u_sdrc_core_u_req_gen__abc_22171_n874), .Y(u_sdrc_core_u_req_gen__abc_22171_n901) );
  AND2X2 AND2X2_1889 ( .A(u_sdrc_core_u_req_gen__abc_22171_n904), .B(u_sdrc_core_u_req_gen__abc_22171_n905), .Y(u_sdrc_core_u_req_gen_r2b_raddr_0__FF_INPUT) );
  AND2X2 AND2X2_189 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf3), .B(u_sdrc_core_u_bank_ctl_x2b_ack_bF_buf1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_x2b_ack) );
  AND2X2 AND2X2_1890 ( .A(u_sdrc_core_u_req_gen_map_address_13_), .B(u_sdrc_core_u_req_gen__abc_22171_n873), .Y(u_sdrc_core_u_req_gen__abc_22171_n907) );
  AND2X2 AND2X2_1891 ( .A(u_sdrc_core_u_req_gen_map_address_14_), .B(u_sdrc_core_u_req_gen__abc_22171_n888), .Y(u_sdrc_core_u_req_gen__abc_22171_n908) );
  AND2X2 AND2X2_1892 ( .A(u_sdrc_core_u_req_gen_map_address_12_), .B(u_sdrc_core_u_req_gen__abc_22171_n876), .Y(u_sdrc_core_u_req_gen__abc_22171_n909) );
  AND2X2 AND2X2_1893 ( .A(u_sdrc_core_u_req_gen__abc_22171_n912), .B(u_sdrc_core_u_req_gen__abc_22171_n913), .Y(u_sdrc_core_u_req_gen_r2b_raddr_1__FF_INPUT) );
  AND2X2 AND2X2_1894 ( .A(u_sdrc_core_u_req_gen_map_address_13_), .B(u_sdrc_core_u_req_gen__abc_22171_n876), .Y(u_sdrc_core_u_req_gen__abc_22171_n915) );
  AND2X2 AND2X2_1895 ( .A(u_sdrc_core_u_req_gen_map_address_15_), .B(u_sdrc_core_u_req_gen__abc_22171_n888), .Y(u_sdrc_core_u_req_gen__abc_22171_n916) );
  AND2X2 AND2X2_1896 ( .A(u_sdrc_core_u_req_gen_map_address_14_), .B(u_sdrc_core_u_req_gen__abc_22171_n874), .Y(u_sdrc_core_u_req_gen__abc_22171_n917) );
  AND2X2 AND2X2_1897 ( .A(u_sdrc_core_u_req_gen__abc_22171_n920), .B(u_sdrc_core_u_req_gen__abc_22171_n921), .Y(u_sdrc_core_u_req_gen_r2b_raddr_2__FF_INPUT) );
  AND2X2 AND2X2_1898 ( .A(u_sdrc_core_u_req_gen_map_address_13_), .B(u_sdrc_core_u_req_gen__abc_22171_n877), .Y(u_sdrc_core_u_req_gen__abc_22171_n923) );
  AND2X2 AND2X2_1899 ( .A(u_sdrc_core_u_req_gen_map_address_16_), .B(u_sdrc_core_u_req_gen__abc_22171_n871), .Y(u_sdrc_core_u_req_gen__abc_22171_n924) );
  AND2X2 AND2X2_19 ( .A(u_sdrc_core_b2x_cmd_1_), .B(u_sdrc_core_u_bank_ctl__abc_21249_n240_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n241) );
  AND2X2 AND2X2_190 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf3), .B(u_sdrc_core_u_bank_ctl_x2b_ack_bF_buf0), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_x2b_ack) );
  AND2X2 AND2X2_1900 ( .A(u_sdrc_core_u_req_gen_map_address_15_), .B(u_sdrc_core_u_req_gen__abc_22171_n874), .Y(u_sdrc_core_u_req_gen__abc_22171_n925) );
  AND2X2 AND2X2_1901 ( .A(u_sdrc_core_u_req_gen_map_address_14_), .B(u_sdrc_core_u_req_gen__abc_22171_n879), .Y(u_sdrc_core_u_req_gen__abc_22171_n926) );
  AND2X2 AND2X2_1902 ( .A(u_sdrc_core_u_req_gen_map_address_17_), .B(u_sdrc_core_u_req_gen__abc_22171_n888), .Y(u_sdrc_core_u_req_gen__abc_22171_n930) );
  AND2X2 AND2X2_1903 ( .A(u_sdrc_core_u_req_gen_map_address_15_), .B(u_sdrc_core_u_req_gen__abc_22171_n876), .Y(u_sdrc_core_u_req_gen__abc_22171_n931) );
  AND2X2 AND2X2_1904 ( .A(u_sdrc_core_u_req_gen_map_address_16_), .B(u_sdrc_core_u_req_gen__abc_22171_n874), .Y(u_sdrc_core_u_req_gen__abc_22171_n932) );
  AND2X2 AND2X2_1905 ( .A(u_sdrc_core_u_req_gen__abc_22171_n935), .B(u_sdrc_core_u_req_gen__abc_22171_n936), .Y(u_sdrc_core_u_req_gen_r2b_raddr_4__FF_INPUT) );
  AND2X2 AND2X2_1906 ( .A(u_sdrc_core_u_req_gen_map_address_18_), .B(u_sdrc_core_u_req_gen__abc_22171_n888), .Y(u_sdrc_core_u_req_gen__abc_22171_n938) );
  AND2X2 AND2X2_1907 ( .A(u_sdrc_core_u_req_gen_map_address_17_), .B(u_sdrc_core_u_req_gen__abc_22171_n874), .Y(u_sdrc_core_u_req_gen__abc_22171_n939) );
  AND2X2 AND2X2_1908 ( .A(u_sdrc_core_u_req_gen_map_address_16_), .B(u_sdrc_core_u_req_gen__abc_22171_n876), .Y(u_sdrc_core_u_req_gen__abc_22171_n940) );
  AND2X2 AND2X2_1909 ( .A(u_sdrc_core_u_req_gen__abc_22171_n943), .B(u_sdrc_core_u_req_gen__abc_22171_n944), .Y(u_sdrc_core_u_req_gen_r2b_raddr_5__FF_INPUT) );
  AND2X2 AND2X2_191 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf3), .B(u_sdrc_core_u_bank_ctl_x2b_ack_bF_buf3), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_x2b_ack) );
  AND2X2 AND2X2_1910 ( .A(u_sdrc_core_u_req_gen_map_address_18_), .B(u_sdrc_core_u_req_gen__abc_22171_n874), .Y(u_sdrc_core_u_req_gen__abc_22171_n946) );
  AND2X2 AND2X2_1911 ( .A(u_sdrc_core_u_req_gen_map_address_17_), .B(u_sdrc_core_u_req_gen__abc_22171_n876), .Y(u_sdrc_core_u_req_gen__abc_22171_n948) );
  AND2X2 AND2X2_1912 ( .A(u_sdrc_core_u_req_gen_map_address_19_), .B(u_sdrc_core_u_req_gen__abc_22171_n888), .Y(u_sdrc_core_u_req_gen__abc_22171_n949) );
  AND2X2 AND2X2_1913 ( .A(u_sdrc_core_u_req_gen__abc_22171_n951), .B(u_sdrc_core_u_req_gen__abc_22171_n952), .Y(u_sdrc_core_u_req_gen_r2b_raddr_6__FF_INPUT) );
  AND2X2 AND2X2_1914 ( .A(u_sdrc_core_u_req_gen_map_address_18_), .B(u_sdrc_core_u_req_gen__abc_22171_n876), .Y(u_sdrc_core_u_req_gen__abc_22171_n954) );
  AND2X2 AND2X2_1915 ( .A(u_sdrc_core_u_req_gen_map_address_19_), .B(u_sdrc_core_u_req_gen__abc_22171_n874), .Y(u_sdrc_core_u_req_gen__abc_22171_n955) );
  AND2X2 AND2X2_1916 ( .A(u_sdrc_core_u_req_gen_map_address_20_), .B(u_sdrc_core_u_req_gen__abc_22171_n888), .Y(u_sdrc_core_u_req_gen__abc_22171_n956) );
  AND2X2 AND2X2_1917 ( .A(u_sdrc_core_u_req_gen__abc_22171_n959), .B(u_sdrc_core_u_req_gen__abc_22171_n960), .Y(u_sdrc_core_u_req_gen_r2b_raddr_7__FF_INPUT) );
  AND2X2 AND2X2_1918 ( .A(u_sdrc_core_u_req_gen_map_address_21_), .B(u_sdrc_core_u_req_gen__abc_22171_n888), .Y(u_sdrc_core_u_req_gen__abc_22171_n962) );
  AND2X2 AND2X2_1919 ( .A(u_sdrc_core_u_req_gen_map_address_19_), .B(u_sdrc_core_u_req_gen__abc_22171_n876), .Y(u_sdrc_core_u_req_gen__abc_22171_n963) );
  AND2X2 AND2X2_192 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n249_1), .B(sdram_resetn_bF_buf38), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n250_1) );
  AND2X2 AND2X2_1920 ( .A(u_sdrc_core_u_req_gen_map_address_20_), .B(u_sdrc_core_u_req_gen__abc_22171_n874), .Y(u_sdrc_core_u_req_gen__abc_22171_n964) );
  AND2X2 AND2X2_1921 ( .A(u_sdrc_core_u_req_gen__abc_22171_n967), .B(u_sdrc_core_u_req_gen__abc_22171_n968), .Y(u_sdrc_core_u_req_gen_r2b_raddr_8__FF_INPUT) );
  AND2X2 AND2X2_1922 ( .A(u_sdrc_core_u_req_gen_map_address_20_), .B(u_sdrc_core_u_req_gen__abc_22171_n879), .Y(u_sdrc_core_u_req_gen__abc_22171_n970) );
  AND2X2 AND2X2_1923 ( .A(u_sdrc_core_u_req_gen_map_address_21_), .B(u_sdrc_core_u_req_gen__abc_22171_n874), .Y(u_sdrc_core_u_req_gen__abc_22171_n971) );
  AND2X2 AND2X2_1924 ( .A(u_sdrc_core_u_req_gen_map_address_22_), .B(u_sdrc_core_u_req_gen__abc_22171_n871), .Y(u_sdrc_core_u_req_gen__abc_22171_n973) );
  AND2X2 AND2X2_1925 ( .A(u_sdrc_core_u_req_gen_map_address_19_), .B(u_sdrc_core_u_req_gen__abc_22171_n877), .Y(u_sdrc_core_u_req_gen__abc_22171_n974) );
  AND2X2 AND2X2_1926 ( .A(u_sdrc_core_u_req_gen__abc_22171_n977), .B(u_sdrc_core_u_req_gen__abc_22171_n893_bF_buf1), .Y(u_sdrc_core_u_req_gen__abc_22171_n978) );
  AND2X2 AND2X2_1927 ( .A(u_sdrc_core_u_req_gen__abc_22171_n979), .B(u_sdrc_core_u_req_gen__abc_22171_n981), .Y(u_sdrc_core_u_req_gen__abc_22171_n982) );
  AND2X2 AND2X2_1928 ( .A(u_sdrc_core_u_req_gen__abc_22171_n982), .B(u_sdrc_core_u_req_gen__abc_22171_n978), .Y(u_sdrc_core_u_req_gen__abc_22171_n983) );
  AND2X2 AND2X2_1929 ( .A(u_sdrc_core_u_req_gen__abc_22171_n984), .B(u_sdrc_core_u_req_gen__abc_22171_n985), .Y(u_sdrc_core_u_req_gen_r2b_raddr_10__FF_INPUT) );
  AND2X2 AND2X2_193 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n250_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_3_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n251) );
  AND2X2 AND2X2_1930 ( .A(u_sdrc_core_u_req_gen__abc_22171_n988), .B(u_sdrc_core_u_req_gen__abc_22171_n989), .Y(u_sdrc_core_u_req_gen__abc_22171_n990) );
  AND2X2 AND2X2_1931 ( .A(u_sdrc_core_u_req_gen__abc_22171_n991), .B(u_sdrc_core_u_req_gen__abc_22171_n893_bF_buf2), .Y(u_sdrc_core_u_req_gen__abc_22171_n992) );
  AND2X2 AND2X2_1932 ( .A(u_sdrc_core_u_req_gen__abc_22171_n990), .B(u_sdrc_core_u_req_gen__abc_22171_n992), .Y(u_sdrc_core_u_req_gen__abc_22171_n993) );
  AND2X2 AND2X2_1933 ( .A(u_sdrc_core_u_req_gen__abc_22171_n994), .B(u_sdrc_core_u_req_gen__abc_22171_n987), .Y(u_sdrc_core_u_req_gen_r2b_raddr_11__FF_INPUT) );
  AND2X2 AND2X2_1934 ( .A(u_sdrc_core_u_req_gen__abc_22171_n996), .B(u_sdrc_core_u_req_gen__abc_22171_n893_bF_buf1), .Y(u_sdrc_core_u_req_gen__abc_22171_n997) );
  AND2X2 AND2X2_1935 ( .A(u_sdrc_core_u_req_gen__abc_22171_n998), .B(u_sdrc_core_u_req_gen__abc_22171_n999), .Y(u_sdrc_core_u_req_gen__abc_22171_n1000) );
  AND2X2 AND2X2_1936 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1000), .B(u_sdrc_core_u_req_gen__abc_22171_n997), .Y(u_sdrc_core_u_req_gen__abc_22171_n1001) );
  AND2X2 AND2X2_1937 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1002), .B(u_sdrc_core_u_req_gen__abc_22171_n1003), .Y(u_sdrc_core_u_req_gen_r2b_raddr_12__FF_INPUT) );
  AND2X2 AND2X2_1938 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1005), .B(u_sdrc_core_u_req_gen_req_st_0_), .Y(u_sdrc_core_r2x_idle) );
  AND2X2 AND2X2_1939 ( .A(u_sdrc_core_u_req_gen__abc_22171_n195_1), .B(u_sdrc_core_r2b_start), .Y(u_sdrc_core_u_req_gen__abc_22171_n1007) );
  AND2X2 AND2X2_194 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_r2b_req), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_0_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack) );
  AND2X2 AND2X2_1940 ( .A(u_sdrc_core_u_req_gen__abc_22171_n309), .B(u_sdrc_core_u_req_gen__abc_22171_n1009), .Y(u_sdrc_core_u_req_gen__abc_22171_n1010) );
  AND2X2 AND2X2_1941 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1011), .B(u_sdrc_core_u_req_gen__abc_22171_n1012), .Y(u_sdrc_core_u_req_gen__abc_22171_n1013) );
  AND2X2 AND2X2_1942 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1016), .B(u_sdrc_core_u_req_gen__abc_22171_n1015), .Y(u_sdrc_core_u_req_gen__abc_22171_n1017) );
  AND2X2 AND2X2_1943 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1017), .B(u_sdrc_core_u_req_gen__abc_22171_n1014), .Y(u_sdrc_core_u_req_gen__abc_22171_n1018) );
  AND2X2 AND2X2_1944 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1013), .B(u_sdrc_core_u_req_gen__abc_22171_n1019), .Y(u_sdrc_core_u_req_gen__abc_22171_n1020) );
  AND2X2 AND2X2_1945 ( .A(u_sdrc_core_u_req_gen__abc_22171_n311), .B(u_sdrc_core_u_req_gen__abc_22171_n464_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n1022) );
  AND2X2 AND2X2_1946 ( .A(u_sdrc_core_u_req_gen__abc_22171_n278), .B(u_sdrc_core_u_req_gen__abc_22171_n1023), .Y(u_sdrc_core_u_req_gen__abc_22171_n1024) );
  AND2X2 AND2X2_1947 ( .A(u_sdrc_core_u_req_gen__abc_22171_n267), .B(u_sdrc_core_u_req_gen__abc_22171_n387), .Y(u_sdrc_core_u_req_gen__abc_22171_n1025) );
  AND2X2 AND2X2_1948 ( .A(u_sdrc_core_u_req_gen__abc_22171_n343_1), .B(u_sdrc_core_u_req_gen__abc_22171_n257), .Y(u_sdrc_core_u_req_gen__abc_22171_n1027) );
  AND2X2 AND2X2_1949 ( .A(u_sdrc_core_u_req_gen__abc_22171_n243_1), .B(u_sdrc_core_u_req_gen__abc_22171_n382_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n1028) );
  AND2X2 AND2X2_195 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf3), .B(sdram_resetn_bF_buf37), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n253_1) );
  AND2X2 AND2X2_1950 ( .A(u_sdrc_core_u_req_gen__abc_22171_n253), .B(u_sdrc_core_u_req_gen__abc_22171_n1029), .Y(u_sdrc_core_u_req_gen__abc_22171_n1030) );
  AND2X2 AND2X2_1951 ( .A(u_sdrc_core_u_req_gen__abc_22171_n252), .B(u_sdrc_core_u_req_gen__abc_22171_n363), .Y(u_sdrc_core_u_req_gen__abc_22171_n1031) );
  AND2X2 AND2X2_1952 ( .A(u_sdrc_core_u_req_gen__abc_22171_n266), .B(u_sdrc_core_u_req_gen__abc_22171_n388_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n1037) );
  AND2X2 AND2X2_1953 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1038), .B(u_sdrc_core_u_req_gen__abc_22171_n1042), .Y(u_sdrc_core_u_req_gen__abc_22171_n1043) );
  AND2X2 AND2X2_1954 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1046), .B(u_sdrc_core_u_req_gen__abc_22171_n1044), .Y(u_sdrc_core_u_req_gen__abc_22171_n1047) );
  AND2X2 AND2X2_1955 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1048), .B(u_sdrc_core_u_req_gen__abc_22171_n1041), .Y(u_sdrc_core_u_req_gen__abc_22171_n1049) );
  AND2X2 AND2X2_1956 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1049), .B(u_sdrc_core_u_req_gen__abc_22171_n1040), .Y(u_sdrc_core_u_req_gen__abc_22171_n1050) );
  AND2X2 AND2X2_1957 ( .A(u_sdrc_core_u_req_gen__abc_22171_n289), .B(u_sdrc_core_u_req_gen__abc_22171_n419), .Y(u_sdrc_core_u_req_gen__abc_22171_n1051) );
  AND2X2 AND2X2_1958 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1052), .B(u_sdrc_core_u_req_gen__abc_22171_n442_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n1053) );
  AND2X2 AND2X2_1959 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1056), .B(u_sdrc_core_u_req_gen__abc_22171_n1057), .Y(u_sdrc_core_u_req_gen__abc_22171_n1058) );
  AND2X2 AND2X2_196 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n257), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n259_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n260) );
  AND2X2 AND2X2_1960 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1055), .B(u_sdrc_core_u_req_gen__abc_22171_n1058), .Y(u_sdrc_core_u_req_gen__abc_22171_n1059) );
  AND2X2 AND2X2_1961 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1060), .B(u_sdrc_core_u_req_gen__abc_22171_n1021), .Y(u_sdrc_core_u_req_gen__abc_22171_n1061) );
  AND2X2 AND2X2_1962 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1062), .B(u_sdrc_core_u_req_gen__abc_22171_n1018), .Y(u_sdrc_core_u_req_gen__abc_22171_n1063) );
  AND2X2 AND2X2_1963 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1064), .B(u_sdrc_core_u_req_gen__abc_22171_n893_bF_buf3), .Y(u_sdrc_core_u_req_gen__abc_22171_n1065) );
  AND2X2 AND2X2_1964 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1010), .B(u_sdrc_core_u_req_gen__abc_22171_n1065), .Y(u_sdrc_core_u_req_gen__abc_22171_n1066) );
  AND2X2 AND2X2_1965 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1011), .B(u_sdrc_core_u_req_gen__abc_22171_n1067), .Y(u_sdrc_core_u_req_gen__abc_22171_n1068) );
  AND2X2 AND2X2_1966 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1072), .B(u_sdrc_core_u_req_gen__abc_22171_n1071), .Y(u_sdrc_core_u_req_gen__abc_22171_n1073) );
  AND2X2 AND2X2_1967 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1073), .B(u_sdrc_core_u_req_gen__abc_22171_n1070), .Y(u_sdrc_core_u_req_gen__abc_22171_n1074) );
  AND2X2 AND2X2_1968 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1069), .B(u_sdrc_core_u_req_gen__abc_22171_n1074), .Y(u_sdrc_core_u_req_gen__abc_22171_n1075) );
  AND2X2 AND2X2_1969 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1010), .B(u_sdrc_core_u_req_gen__abc_22171_n1064), .Y(u_sdrc_core_u_req_gen__abc_22171_n1079) );
  AND2X2 AND2X2_197 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n260), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n255_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n261_1) );
  AND2X2 AND2X2_1970 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1079), .B(u_sdrc_core_u_req_gen__abc_22171_n1078), .Y(u_sdrc_core_u_req_gen__abc_22171_n1080) );
  AND2X2 AND2X2_1971 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1080), .B(u_sdrc_core_u_req_gen__abc_22171_n1081), .Y(u_sdrc_core_u_req_gen__abc_22171_n1082) );
  AND2X2 AND2X2_1972 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1083), .B(u_sdrc_core_u_req_gen__abc_22171_n1084), .Y(u_sdrc_core_u_req_gen__abc_22171_n1085) );
  AND2X2 AND2X2_1973 ( .A(app_req_ack_bF_buf2), .B(u_sdrc_core_u_req_gen__abc_22171_n1087), .Y(u_sdrc_core_u_req_gen__abc_22171_n1088) );
  AND2X2 AND2X2_1974 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1089), .B(u_sdrc_core_u_req_gen__abc_22171_n871), .Y(u_sdrc_core_u_req_gen__abc_22171_n1090) );
  AND2X2 AND2X2_1975 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1080), .B(u_sdrc_core_u_req_gen__abc_22171_n1090), .Y(u_sdrc_core_u_req_gen__abc_22171_n1091) );
  AND2X2 AND2X2_1976 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1092), .B(u_sdrc_core_u_req_gen__abc_22171_n1088), .Y(u_sdrc_core_u_req_gen__abc_22171_n1093) );
  AND2X2 AND2X2_1977 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1078), .B(\cfg_colbits[1] ), .Y(u_sdrc_core_u_req_gen__abc_22171_n1095) );
  AND2X2 AND2X2_1978 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1094), .B(u_sdrc_core_u_req_gen__abc_22171_n1096), .Y(u_sdrc_core_u_req_gen__abc_22171_n1097) );
  AND2X2 AND2X2_1979 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1079), .B(u_sdrc_core_u_req_gen__abc_22171_n1095), .Y(u_sdrc_core_u_req_gen__abc_22171_n1098) );
  AND2X2 AND2X2_198 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n263), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n265_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n266) );
  AND2X2 AND2X2_1980 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1100), .B(u_sdrc_core_u_req_gen__abc_22171_n1099), .Y(u_sdrc_core_u_req_gen__abc_22171_n1101) );
  AND2X2 AND2X2_1981 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1101), .B(u_sdrc_core_u_req_gen__abc_22171_n1093), .Y(u_sdrc_core_u_req_gen__abc_22171_n1102) );
  AND2X2 AND2X2_1982 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1102), .B(u_sdrc_core_u_req_gen__abc_22171_n1086), .Y(u_sdrc_core_u_req_gen__abc_22171_n1103) );
  AND2X2 AND2X2_1983 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1077), .B(u_sdrc_core_u_req_gen__abc_22171_n1103), .Y(u_sdrc_core_u_req_gen_page_ovflw_r_FF_INPUT) );
  AND2X2 AND2X2_1984 ( .A(u_sdrc_core_u_req_gen__abc_22171_n181), .B(u_sdrc_core_r2b_start), .Y(u_sdrc_core_u_req_gen__abc_22171_n1105) );
  AND2X2 AND2X2_1985 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n357), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n358_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n359) );
  AND2X2 AND2X2_1986 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n359), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n356_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n360) );
  AND2X2 AND2X2_1987 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n360), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n355), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n361) );
  AND2X2 AND2X2_1988 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n354), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n361), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n362_1) );
  AND2X2 AND2X2_1989 ( .A(sdram_resetn_bF_buf22), .B(u_sdrc_core_u_xfr_ctl_mgmt_st_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n363) );
  AND2X2 AND2X2_199 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n268_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n270_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n271_1) );
  AND2X2 AND2X2_1990 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n363), .B(_auto_iopadmap_cc_313_execute_24701), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n364) );
  AND2X2 AND2X2_1991 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n362_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n364), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n365_1) );
  AND2X2 AND2X2_1992 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n366), .B(\cfg_sdr_rfmax[2] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n367_1) );
  AND2X2 AND2X2_1993 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n368), .B(\cfg_sdr_rfmax[1] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n369_1) );
  AND2X2 AND2X2_1994 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n370), .B(\cfg_sdr_rfmax[0] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n371) );
  AND2X2 AND2X2_1995 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n373), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n374_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n375) );
  AND2X2 AND2X2_1996 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n372_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n375), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n376) );
  AND2X2 AND2X2_1997 ( .A(sdram_resetn_bF_buf21), .B(cfg_sdr_en), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n378) );
  AND2X2 AND2X2_1998 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n378), .B(u_sdrc_core_u_xfr_ctl_mgmt_st_7_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n379) );
  AND2X2 AND2X2_1999 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n377_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n379), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n380_1) );
  AND2X2 AND2X2_2 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_tras_ok), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_tras_ok), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n205_1) );
  AND2X2 AND2X2_20 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n241), .B(u_sdrc_core_u_bank_ctl__abc_21249_n239_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n243) );
  AND2X2 AND2X2_200 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n266), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n271_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n272) );
  AND2X2 AND2X2_2000 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n354), .B(sdram_resetn_bF_buf20), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n381) );
  AND2X2 AND2X2_2001 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n381), .B(u_sdrc_core_u_xfr_ctl_mgmt_st_3_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n382_1) );
  AND2X2 AND2X2_2002 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n385), .B(u_sdrc_core_u_xfr_ctl_xfr_st_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n386) );
  AND2X2 AND2X2_2003 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n388), .B(u_sdrc_core_u_xfr_ctl_xfr_st_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n389_1) );
  AND2X2 AND2X2_2004 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n387_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n390), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_pre_ok) );
  AND2X2 AND2X2_2005 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n392), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n393_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n394) );
  AND2X2 AND2X2_2006 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n397), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n398_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n399_1) );
  AND2X2 AND2X2_2007 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n399_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n396_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n400_1) );
  AND2X2 AND2X2_2008 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n403_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_pre_ok), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n404_1) );
  AND2X2 AND2X2_2009 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n405_1_bF_buf3), .B(sdram_resetn_bF_buf19), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n406_1) );
  AND2X2 AND2X2_201 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n272), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n261_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n273_1) );
  AND2X2 AND2X2_2010 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n406_1), .B(u_sdrc_core_u_xfr_ctl_mgmt_st_6_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n407_1) );
  AND2X2 AND2X2_2011 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n381), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n395), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n410_1) );
  AND2X2 AND2X2_2012 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n410_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n409_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n411_1) );
  AND2X2 AND2X2_2013 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n415), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n414_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n416_1) );
  AND2X2 AND2X2_2014 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n353_1), .B(sdram_resetn_bF_buf17), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n418_1) );
  AND2X2 AND2X2_2015 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n418_1), .B(u_sdrc_core_u_xfr_ctl_mgmt_st_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n419) );
  AND2X2 AND2X2_2016 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n404_1), .B(sdram_resetn_bF_buf16), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n420_1) );
  AND2X2 AND2X2_2017 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n420_1), .B(u_sdrc_core_u_xfr_ctl_mgmt_st_6_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n421) );
  AND2X2 AND2X2_2018 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n406_1), .B(u_sdrc_core_u_xfr_ctl_mgmt_st_5_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n423) );
  AND2X2 AND2X2_2019 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n363), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n424), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n425_1) );
  AND2X2 AND2X2_202 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n275), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n277_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n278) );
  AND2X2 AND2X2_2020 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n362_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n425_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n426) );
  AND2X2 AND2X2_2021 ( .A(sdram_resetn_bF_buf15), .B(u_sdrc_core_u_xfr_ctl_mgmt_st_4_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n428_1) );
  AND2X2 AND2X2_2022 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_pre_ok), .B(u_sdrc_core_b2x_tras_ok), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n429) );
  AND2X2 AND2X2_2023 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n403_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n429), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n430) );
  AND2X2 AND2X2_2024 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n431), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n428_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n432_1) );
  AND2X2 AND2X2_2025 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n433), .B(u_sdrc_core_u_xfr_ctl_mgmt_st_7_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n434_1) );
  AND2X2 AND2X2_2026 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n435), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n378), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n436_1) );
  AND2X2 AND2X2_2027 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n418_1), .B(u_sdrc_core_u_xfr_ctl_mgmt_st_3_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n438_1) );
  AND2X2 AND2X2_2028 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n420_1), .B(u_sdrc_core_u_xfr_ctl_mgmt_st_5_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n439) );
  AND2X2 AND2X2_2029 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n430), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n428_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n441) );
  AND2X2 AND2X2_203 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n280_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n282_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n283_1) );
  AND2X2 AND2X2_2030 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n418_1), .B(u_sdrc_core_u_xfr_ctl_mgmt_st_2_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n442_1) );
  AND2X2 AND2X2_2031 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n444_1), .B(u_sdrc_core_b2x_req), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n445) );
  AND2X2 AND2X2_2032 ( .A(u_sdrc_core_u_xfr_ctl_xfr_st_1_), .B(u_sdrc_core_u_xfr_ctl_xfr_st_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n446_1) );
  AND2X2 AND2X2_2033 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n447), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n448_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n449_1) );
  AND2X2 AND2X2_2034 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n450_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n451_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n452_1) );
  AND2X2 AND2X2_2035 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n449_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n452_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n453_1) );
  AND2X2 AND2X2_2036 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n454_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n455_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n456_1) );
  AND2X2 AND2X2_2037 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n453_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n456_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n457) );
  AND2X2 AND2X2_2038 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n457), .B(u_sdrc_core_u_xfr_ctl_l_len_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n458) );
  AND2X2 AND2X2_2039 ( .A(u_sdrc_core_b2x_cmd_0_), .B(u_sdrc_core_b2x_cmd_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n459_1) );
  AND2X2 AND2X2_204 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n278), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n283_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n284_1) );
  AND2X2 AND2X2_2040 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n461_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n462_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n463_1) );
  AND2X2 AND2X2_2041 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n464_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n460_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n465_1) );
  AND2X2 AND2X2_2042 ( .A(u_sdrc_core_b2x_ba_1_), .B(u_sdrc_core_u_bank_ctl_xfr_bank_sel_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n467_1) );
  AND2X2 AND2X2_2043 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n468_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n466_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n469_1) );
  AND2X2 AND2X2_2044 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n471_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n461_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n472) );
  AND2X2 AND2X2_2045 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n473), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n474), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n475) );
  AND2X2 AND2X2_2046 ( .A(u_sdrc_core_u_bank_ctl_xfr_bank_sel_0_), .B(u_sdrc_core_b2x_ba_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n476) );
  AND2X2 AND2X2_2047 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n477), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n472), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n478) );
  AND2X2 AND2X2_2048 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n478), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n470_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n479) );
  AND2X2 AND2X2_2049 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n479), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n462_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n480) );
  AND2X2 AND2X2_205 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n286_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n288_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n289) );
  AND2X2 AND2X2_2050 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n481), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n386), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n482) );
  AND2X2 AND2X2_2051 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n479), .B(u_sdrc_core_u_xfr_ctl_l_wrap), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n483) );
  AND2X2 AND2X2_2052 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n464_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n389_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n485_1) );
  AND2X2 AND2X2_2053 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n484_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n485_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n486) );
  AND2X2 AND2X2_2054 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n487), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n458), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n488_1) );
  AND2X2 AND2X2_2055 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n489_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n445), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n490_1) );
  AND2X2 AND2X2_2056 ( .A(u_sdrc_core_u_xfr_ctl_xfr_caddr_1_), .B(u_sdrc_core_u_xfr_ctl_xfr_caddr_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n492_1) );
  AND2X2 AND2X2_2057 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n492_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n462_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n493_1) );
  AND2X2 AND2X2_2058 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n494_1), .B(u_sdrc_core_b2x_req), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n495_1) );
  AND2X2 AND2X2_2059 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n444_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n389_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n496_1) );
  AND2X2 AND2X2_206 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n291_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n293), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n294_1) );
  AND2X2 AND2X2_2060 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n497_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n495_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n498_1) );
  AND2X2 AND2X2_2061 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n498_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n491_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n499_1) );
  AND2X2 AND2X2_2062 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n388), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n385), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n500_1) );
  AND2X2 AND2X2_2063 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n500_1), .B(_auto_iopadmap_cc_313_execute_24701), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n501_1) );
  AND2X2 AND2X2_2064 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n445), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n501_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n502) );
  AND2X2 AND2X2_2065 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n510), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n509), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n511_1) );
  AND2X2 AND2X2_2066 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n514), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n507), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n515) );
  AND2X2 AND2X2_2067 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n516_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n517_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n518_1) );
  AND2X2 AND2X2_2068 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n519), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n506_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n520_1) );
  AND2X2 AND2X2_2069 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n521_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n522), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n523_1) );
  AND2X2 AND2X2_207 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n289), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n294_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n295_1) );
  AND2X2 AND2X2_2070 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n458), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n462_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n524_1) );
  AND2X2 AND2X2_2071 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n525), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n494_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n526_1) );
  AND2X2 AND2X2_2072 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n525), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n390), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n528) );
  AND2X2 AND2X2_2073 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n523_1_bF_buf3), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n529_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n530_1) );
  AND2X2 AND2X2_2074 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n508), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n460_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n531) );
  AND2X2 AND2X2_2075 ( .A(u_sdrc_core_u_bank_ctl_x2b_ack_bF_buf2), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n531), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n532) );
  AND2X2 AND2X2_2076 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n533_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n405_1_bF_buf2), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n534_1) );
  AND2X2 AND2X2_2077 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n535), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n401_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n536_1) );
  AND2X2 AND2X2_2078 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n404_1), .B(u_sdrc_core_u_xfr_ctl_mgmt_st_6_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n539_1) );
  AND2X2 AND2X2_2079 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n541), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n544), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_refresh) );
  AND2X2 AND2X2_208 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n284_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n295_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n296_1) );
  AND2X2 AND2X2_2080 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n491_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n389_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n546_1) );
  AND2X2 AND2X2_2081 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n547), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n390), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n548_1) );
  AND2X2 AND2X2_2082 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n445), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n459_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n550) );
  AND2X2 AND2X2_2083 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n550), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n549), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n551_1) );
  AND2X2 AND2X2_2084 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n471_1), .B(u_sdrc_core_b2x_cmd_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n553) );
  AND2X2 AND2X2_2085 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n445), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n553), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n554_1) );
  AND2X2 AND2X2_2086 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n558_1), .B(\cfg_sdr_cas[0] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n559) );
  AND2X2 AND2X2_2087 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n559), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n557_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n560_1) );
  AND2X2 AND2X2_2088 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n557_1), .B(\cfg_sdr_cas[1] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n562) );
  AND2X2 AND2X2_2089 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n558_1), .B(\cfg_sdr_cas[2] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n565) );
  AND2X2 AND2X2_209 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n296_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n273_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n297) );
  AND2X2 AND2X2_2090 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n565), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n564_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n566_1) );
  AND2X2 AND2X2_2091 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n567), .B(u_sdrc_core_u_xfr_ctl_l_rd_next_5_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n568) );
  AND2X2 AND2X2_2092 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n569_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n563_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n570_1) );
  AND2X2 AND2X2_2093 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n562), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n564_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n571) );
  AND2X2 AND2X2_2094 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n572_1), .B(u_sdrc_core_u_xfr_ctl_l_rd_next_3_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n573) );
  AND2X2 AND2X2_2095 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n575_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n561), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n576_1) );
  AND2X2 AND2X2_2096 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n577), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n446_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n578_1) );
  AND2X2 AND2X2_2097 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n386), .B(_auto_iopadmap_cc_313_execute_24701), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n579) );
  AND2X2 AND2X2_2098 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n458), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n579), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n580) );
  AND2X2 AND2X2_2099 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n550), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n446_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n581_1) );
  AND2X2 AND2X2_21 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n244_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n242_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n245_1) );
  AND2X2 AND2X2_210 ( .A(u_sdrc_core_r2b_raddr_10_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_10_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n298_1) );
  AND2X2 AND2X2_2100 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n583), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n555), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n584_1) );
  AND2X2 AND2X2_2101 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n585), .B(sdram_resetn_bF_buf14), .Y(u_sdrc_core_u_xfr_ctl_xfr_st_0__FF_INPUT) );
  AND2X2 AND2X2_2102 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n587_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n386), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n588_1) );
  AND2X2 AND2X2_2103 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n458), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n389_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n589) );
  AND2X2 AND2X2_2104 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n554_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n590_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n591) );
  AND2X2 AND2X2_2105 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n502), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n553), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n592) );
  AND2X2 AND2X2_2106 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n595), .B(sdram_resetn_bF_buf13), .Y(u_sdrc_core_u_xfr_ctl_xfr_st_1__FF_INPUT) );
  AND2X2 AND2X2_2107 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n601), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n598), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n602) );
  AND2X2 AND2X2_2108 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n555), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n458), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n604_1) );
  AND2X2 AND2X2_2109 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n603_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n605), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n606_1) );
  AND2X2 AND2X2_211 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n299_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n300_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n301) );
  AND2X2 AND2X2_2110 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n602_bF_buf3), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n606_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n607) );
  AND2X2 AND2X2_2111 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n611), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf4), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n612) );
  AND2X2 AND2X2_2112 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n612), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n608), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n613) );
  AND2X2 AND2X2_2113 ( .A(u_sdrc_core_u_bank_ctl_x2b_ack_bF_buf1), .B(u_sdrc_core_b2x_cmd_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n614) );
  AND2X2 AND2X2_2114 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n614_bF_buf3), .B(u_sdrc_core_b2x_addr_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n615) );
  AND2X2 AND2X2_2115 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n616), .B(sdram_resetn_bF_buf12), .Y(u_sdrc_core_u_xfr_ctl_xfr_caddr_0__FF_INPUT) );
  AND2X2 AND2X2_2116 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n619), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n620_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n621) );
  AND2X2 AND2X2_2117 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n622), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf3), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n623) );
  AND2X2 AND2X2_2118 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n623), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n618_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n624) );
  AND2X2 AND2X2_2119 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n614_bF_buf2), .B(u_sdrc_core_b2x_addr_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n625_1) );
  AND2X2 AND2X2_212 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_8_), .B(u_sdrc_core_r2b_raddr_8_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n303_1) );
  AND2X2 AND2X2_2120 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n626), .B(sdram_resetn_bF_buf11), .Y(u_sdrc_core_u_xfr_ctl_xfr_caddr_1__FF_INPUT) );
  AND2X2 AND2X2_2121 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n492_1), .B(u_sdrc_core_u_xfr_ctl_xfr_caddr_2_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n629) );
  AND2X2 AND2X2_2122 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n630_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n631), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n632) );
  AND2X2 AND2X2_2123 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n633), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf2), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n634) );
  AND2X2 AND2X2_2124 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n634), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n628_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n635_1) );
  AND2X2 AND2X2_2125 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n614_bF_buf1), .B(u_sdrc_core_b2x_addr_2_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n636) );
  AND2X2 AND2X2_2126 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n637), .B(sdram_resetn_bF_buf10), .Y(u_sdrc_core_u_xfr_ctl_xfr_caddr_2__FF_INPUT) );
  AND2X2 AND2X2_2127 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n629), .B(u_sdrc_core_u_xfr_ctl_xfr_caddr_3_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n640) );
  AND2X2 AND2X2_2128 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n641_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n642), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n643) );
  AND2X2 AND2X2_2129 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n644), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n645) );
  AND2X2 AND2X2_213 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n304_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n305), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n306_1) );
  AND2X2 AND2X2_2130 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n645), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n639_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n646_1) );
  AND2X2 AND2X2_2131 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n614_bF_buf0), .B(u_sdrc_core_b2x_addr_3_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n647) );
  AND2X2 AND2X2_2132 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n648), .B(sdram_resetn_bF_buf9), .Y(u_sdrc_core_u_xfr_ctl_xfr_caddr_3__FF_INPUT) );
  AND2X2 AND2X2_2133 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n640), .B(u_sdrc_core_u_xfr_ctl_xfr_caddr_4_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n651) );
  AND2X2 AND2X2_2134 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n652_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n653_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n654) );
  AND2X2 AND2X2_2135 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n655), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf0), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n656) );
  AND2X2 AND2X2_2136 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n656), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n650), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n657_1) );
  AND2X2 AND2X2_2137 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n614_bF_buf3), .B(u_sdrc_core_b2x_addr_4_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n658) );
  AND2X2 AND2X2_2138 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n659), .B(sdram_resetn_bF_buf8), .Y(u_sdrc_core_u_xfr_ctl_xfr_caddr_4__FF_INPUT) );
  AND2X2 AND2X2_2139 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n651), .B(u_sdrc_core_u_xfr_ctl_xfr_caddr_5_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n662) );
  AND2X2 AND2X2_214 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n302_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n307_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n308_1) );
  AND2X2 AND2X2_2140 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n663), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n664), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n665) );
  AND2X2 AND2X2_2141 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n666), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf4), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n667_1) );
  AND2X2 AND2X2_2142 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n667_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n661), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n668) );
  AND2X2 AND2X2_2143 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n614_bF_buf2), .B(u_sdrc_core_b2x_addr_5_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n669) );
  AND2X2 AND2X2_2144 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n670), .B(sdram_resetn_bF_buf7), .Y(u_sdrc_core_u_xfr_ctl_xfr_caddr_5__FF_INPUT) );
  AND2X2 AND2X2_2145 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n662), .B(u_sdrc_core_u_xfr_ctl_xfr_caddr_6_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n673) );
  AND2X2 AND2X2_2146 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n674), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n675), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n676) );
  AND2X2 AND2X2_2147 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n677_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf3), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n678) );
  AND2X2 AND2X2_2148 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n678), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n672_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n679) );
  AND2X2 AND2X2_2149 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n614_bF_buf1), .B(u_sdrc_core_b2x_addr_6_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n680) );
  AND2X2 AND2X2_215 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n310_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n312_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n313) );
  AND2X2 AND2X2_2150 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n681), .B(sdram_resetn_bF_buf6), .Y(u_sdrc_core_u_xfr_ctl_xfr_caddr_6__FF_INPUT) );
  AND2X2 AND2X2_2151 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n673), .B(u_sdrc_core_u_xfr_ctl_xfr_caddr_7_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n684_1) );
  AND2X2 AND2X2_2152 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n685_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n686_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n687) );
  AND2X2 AND2X2_2153 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n688_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf2), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n689_1) );
  AND2X2 AND2X2_2154 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n689_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n683), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n690) );
  AND2X2 AND2X2_2155 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n614_bF_buf0), .B(u_sdrc_core_b2x_addr_7_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n691) );
  AND2X2 AND2X2_2156 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n692_1), .B(sdram_resetn_bF_buf5), .Y(u_sdrc_core_u_xfr_ctl_xfr_caddr_7__FF_INPUT) );
  AND2X2 AND2X2_2157 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n684_1), .B(u_sdrc_core_u_xfr_ctl_xfr_caddr_8_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n695_1) );
  AND2X2 AND2X2_2158 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n696_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n697), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n698) );
  AND2X2 AND2X2_2159 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n699), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n700_1) );
  AND2X2 AND2X2_216 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n315_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n317), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n318_1) );
  AND2X2 AND2X2_2160 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n700_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n694), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n701_1) );
  AND2X2 AND2X2_2161 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n614_bF_buf3), .B(u_sdrc_core_b2x_addr_8_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n702) );
  AND2X2 AND2X2_2162 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n703_1), .B(sdram_resetn_bF_buf4), .Y(u_sdrc_core_u_xfr_ctl_xfr_caddr_8__FF_INPUT) );
  AND2X2 AND2X2_2163 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n695_1), .B(u_sdrc_core_u_xfr_ctl_xfr_caddr_9_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n706) );
  AND2X2 AND2X2_2164 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n707_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n708_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n709) );
  AND2X2 AND2X2_2165 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n710_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf0), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n711_1) );
  AND2X2 AND2X2_2166 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n711_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n705), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n712) );
  AND2X2 AND2X2_2167 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n614_bF_buf2), .B(u_sdrc_core_b2x_addr_9_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n713) );
  AND2X2 AND2X2_2168 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n714), .B(sdram_resetn_bF_buf3), .Y(u_sdrc_core_u_xfr_ctl_xfr_caddr_9__FF_INPUT) );
  AND2X2 AND2X2_2169 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n706), .B(u_sdrc_core_u_xfr_ctl_xfr_caddr_10_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n717) );
  AND2X2 AND2X2_217 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n313), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n318_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n319_1) );
  AND2X2 AND2X2_2170 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n718_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n719_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n720) );
  AND2X2 AND2X2_2171 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n721), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf4), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n722_1) );
  AND2X2 AND2X2_2172 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n722_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n716_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n723_1) );
  AND2X2 AND2X2_2173 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n614_bF_buf1), .B(u_sdrc_core_b2x_addr_10_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n724) );
  AND2X2 AND2X2_2174 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n725_1), .B(sdram_resetn_bF_buf2), .Y(u_sdrc_core_u_xfr_ctl_xfr_caddr_10__FF_INPUT) );
  AND2X2 AND2X2_2175 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n717), .B(u_sdrc_core_u_xfr_ctl_xfr_caddr_11_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n728) );
  AND2X2 AND2X2_2176 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n729), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n730), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n731) );
  AND2X2 AND2X2_2177 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n732), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf3), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n733_1) );
  AND2X2 AND2X2_2178 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n733_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n727), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n734) );
  AND2X2 AND2X2_2179 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n614_bF_buf0), .B(u_sdrc_core_b2x_addr_11_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n735) );
  AND2X2 AND2X2_218 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n321), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n323_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n324_1) );
  AND2X2 AND2X2_2180 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n736_1), .B(sdram_resetn_bF_buf1), .Y(u_sdrc_core_u_xfr_ctl_xfr_caddr_11__FF_INPUT) );
  AND2X2 AND2X2_2181 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n728), .B(u_sdrc_core_u_xfr_ctl_xfr_caddr_12_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n740_1) );
  AND2X2 AND2X2_2182 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n741), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n739), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n742) );
  AND2X2 AND2X2_2183 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n743), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf2), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n744_1) );
  AND2X2 AND2X2_2184 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n744_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n738), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n745) );
  AND2X2 AND2X2_2185 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n614_bF_buf3), .B(u_sdrc_core_b2x_addr_12_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n746) );
  AND2X2 AND2X2_2186 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n747), .B(sdram_resetn_bF_buf0), .Y(u_sdrc_core_u_xfr_ctl_xfr_caddr_12__FF_INPUT) );
  AND2X2 AND2X2_2187 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf1), .B(u_sdrc_core_u_bank_ctl_xfr_bank_sel_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n765) );
  AND2X2 AND2X2_2188 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n614_bF_buf2), .B(u_sdrc_core_b2x_ba_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n766) );
  AND2X2 AND2X2_2189 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n767), .B(sdram_resetn_bF_buf49), .Y(u_sdrc_core_u_xfr_ctl_l_ba_0__FF_INPUT) );
  AND2X2 AND2X2_219 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n326_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_valid), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n327_1) );
  AND2X2 AND2X2_2190 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf0), .B(u_sdrc_core_u_bank_ctl_xfr_bank_sel_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n769) );
  AND2X2 AND2X2_2191 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n614_bF_buf1), .B(u_sdrc_core_b2x_ba_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n770) );
  AND2X2 AND2X2_2192 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n771_1), .B(sdram_resetn_bF_buf48), .Y(u_sdrc_core_u_xfr_ctl_l_ba_1__FF_INPUT) );
  AND2X2 AND2X2_2193 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n776), .B(sdram_resetn_bF_buf47), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n777) );
  AND2X2 AND2X2_2194 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n777), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n775_1), .Y(u_sdrc_core_u_xfr_ctl_l_len_0__FF_INPUT) );
  AND2X2 AND2X2_2195 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n773), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n448_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n780) );
  AND2X2 AND2X2_2196 ( .A(u_sdrc_core_u_xfr_ctl_l_len_0_), .B(u_sdrc_core_u_xfr_ctl_l_len_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n781_1) );
  AND2X2 AND2X2_2197 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n783), .B(sdram_resetn_bF_buf46), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n784_1) );
  AND2X2 AND2X2_2198 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n784_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n779), .Y(u_sdrc_core_u_xfr_ctl_l_len_1__FF_INPUT) );
  AND2X2 AND2X2_2199 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n780), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n451_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n786) );
  AND2X2 AND2X2_22 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n247_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n248), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n249_1) );
  AND2X2 AND2X2_220 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n324_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n327_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n328_1) );
  AND2X2 AND2X2_2200 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n787), .B(u_sdrc_core_u_xfr_ctl_l_len_2_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n788_1) );
  AND2X2 AND2X2_2201 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n791), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n790), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n792) );
  AND2X2 AND2X2_2202 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n792), .B(sdram_resetn_bF_buf45), .Y(u_sdrc_core_u_xfr_ctl_l_len_2__FF_INPUT) );
  AND2X2 AND2X2_2203 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n452_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n780), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n794_1) );
  AND2X2 AND2X2_2204 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n795), .B(u_sdrc_core_u_xfr_ctl_l_len_3_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n796) );
  AND2X2 AND2X2_2205 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n797), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n798_1) );
  AND2X2 AND2X2_2206 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n614_bF_buf1), .B(u_sdrc_core_b2x_len_3_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n799_1) );
  AND2X2 AND2X2_2207 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n800), .B(sdram_resetn_bF_buf44), .Y(u_sdrc_core_u_xfr_ctl_l_len_3__FF_INPUT) );
  AND2X2 AND2X2_2208 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n794_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n447), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n802) );
  AND2X2 AND2X2_2209 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n803_1), .B(u_sdrc_core_u_xfr_ctl_l_len_4_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n804_1) );
  AND2X2 AND2X2_221 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n319_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n328_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n329) );
  AND2X2 AND2X2_2210 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf0), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n805_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n806_1) );
  AND2X2 AND2X2_2211 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n614_bF_buf0), .B(u_sdrc_core_b2x_len_4_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n807_1) );
  AND2X2 AND2X2_2212 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n808_1), .B(sdram_resetn_bF_buf43), .Y(u_sdrc_core_u_xfr_ctl_l_len_4__FF_INPUT) );
  AND2X2 AND2X2_2213 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n802), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n455_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n810_1) );
  AND2X2 AND2X2_2214 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n811_1), .B(u_sdrc_core_u_xfr_ctl_l_len_5_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n812_1) );
  AND2X2 AND2X2_2215 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf4), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n813_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n814_1) );
  AND2X2 AND2X2_2216 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n614_bF_buf3), .B(u_sdrc_core_b2x_len_5_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n815_1) );
  AND2X2 AND2X2_2217 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n816_1), .B(sdram_resetn_bF_buf42), .Y(u_sdrc_core_u_xfr_ctl_l_len_5__FF_INPUT) );
  AND2X2 AND2X2_2218 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n614_bF_buf2), .B(u_sdrc_core_b2x_len_6_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n818_1) );
  AND2X2 AND2X2_2219 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n819_1), .B(u_sdrc_core_u_xfr_ctl_l_len_6_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n820_1) );
  AND2X2 AND2X2_222 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n329), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n308_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n330_1) );
  AND2X2 AND2X2_2220 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n802), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n456_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n821_1) );
  AND2X2 AND2X2_2221 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf3), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n822_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n823_1) );
  AND2X2 AND2X2_2222 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n824_1), .B(sdram_resetn_bF_buf41), .Y(u_sdrc_core_u_xfr_ctl_l_len_6__FF_INPUT) );
  AND2X2 AND2X2_2223 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n826_1), .B(sdram_resetn_bF_buf40), .Y(u_sdrc_core_u_xfr_ctl_l_rd_next_0__FF_INPUT) );
  AND2X2 AND2X2_2224 ( .A(sdram_resetn_bF_buf39), .B(u_sdrc_core_u_xfr_ctl_l_rd_next_0_), .Y(u_sdrc_core_u_xfr_ctl_l_rd_next_1__FF_INPUT) );
  AND2X2 AND2X2_2225 ( .A(sdram_resetn_bF_buf38), .B(u_sdrc_core_u_xfr_ctl_l_rd_next_1_), .Y(u_sdrc_core_u_xfr_ctl_l_rd_next_2__FF_INPUT) );
  AND2X2 AND2X2_2226 ( .A(sdram_resetn_bF_buf37), .B(u_sdrc_core_u_xfr_ctl_l_rd_next_2_), .Y(u_sdrc_core_u_xfr_ctl_l_rd_next_3__FF_INPUT) );
  AND2X2 AND2X2_2227 ( .A(sdram_resetn_bF_buf36), .B(u_sdrc_core_u_xfr_ctl_l_rd_next_3_), .Y(u_sdrc_core_u_xfr_ctl_l_rd_next_4__FF_INPUT) );
  AND2X2 AND2X2_2228 ( .A(sdram_resetn_bF_buf35), .B(u_sdrc_core_u_xfr_ctl_l_rd_next_4_), .Y(u_sdrc_core_u_xfr_ctl_l_rd_next_5__FF_INPUT) );
  AND2X2 AND2X2_2229 ( .A(sdram_resetn_bF_buf34), .B(u_sdrc_core_u_xfr_ctl_l_rd_next_5_), .Y(u_sdrc_core_u_xfr_ctl_l_rd_next_6__FF_INPUT) );
  AND2X2 AND2X2_223 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n297), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n330_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n331_1) );
  AND2X2 AND2X2_2230 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n844_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n843_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n845_1) );
  AND2X2 AND2X2_2231 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n846_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n847_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n848_1) );
  AND2X2 AND2X2_2232 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n849_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n774), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n850_1) );
  AND2X2 AND2X2_2233 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n845_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n850_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n851_1) );
  AND2X2 AND2X2_2234 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n852_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n853), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n854) );
  AND2X2 AND2X2_2235 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n856_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n857_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n858) );
  AND2X2 AND2X2_2236 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n855_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n859_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n860) );
  AND2X2 AND2X2_2237 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n851_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n860), .Y(app_last_wr) );
  AND2X2 AND2X2_2238 ( .A(app_last_wr), .B(u_sdrc_core_u_xfr_ctl_l_rd_next_0__FF_INPUT), .Y(u_sdrc_core_u_xfr_ctl_l_rd_last_0__FF_INPUT) );
  AND2X2 AND2X2_2239 ( .A(sdram_resetn_bF_buf33), .B(u_sdrc_core_u_xfr_ctl_l_rd_last_0_), .Y(u_sdrc_core_u_xfr_ctl_l_rd_last_1__FF_INPUT) );
  AND2X2 AND2X2_224 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n332_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n253_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n333) );
  AND2X2 AND2X2_2240 ( .A(sdram_resetn_bF_buf32), .B(u_sdrc_core_u_xfr_ctl_l_rd_last_1_), .Y(u_sdrc_core_u_xfr_ctl_l_rd_last_2__FF_INPUT) );
  AND2X2 AND2X2_2241 ( .A(sdram_resetn_bF_buf31), .B(u_sdrc_core_u_xfr_ctl_l_rd_last_2_), .Y(u_sdrc_core_u_xfr_ctl_l_rd_last_3__FF_INPUT) );
  AND2X2 AND2X2_2242 ( .A(sdram_resetn_bF_buf30), .B(u_sdrc_core_u_xfr_ctl_l_rd_last_3_), .Y(u_sdrc_core_u_xfr_ctl_l_rd_last_4__FF_INPUT) );
  AND2X2 AND2X2_2243 ( .A(sdram_resetn_bF_buf29), .B(u_sdrc_core_u_xfr_ctl_l_rd_last_4_), .Y(u_sdrc_core_u_xfr_ctl_l_rd_last_5__FF_INPUT) );
  AND2X2 AND2X2_2244 ( .A(sdram_resetn_bF_buf28), .B(u_sdrc_core_u_xfr_ctl_l_rd_last_5_), .Y(u_sdrc_core_u_xfr_ctl_l_rd_last_6__FF_INPUT) );
  AND2X2 AND2X2_2245 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n444_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n869_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_rdok) );
  AND2X2 AND2X2_2246 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n444_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n871_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n872) );
  AND2X2 AND2X2_2247 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n872), .B(sdram_resetn_bF_buf27), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n873) );
  AND2X2 AND2X2_2248 ( .A(u_sdrc_core_r2x_idle), .B(u_sdrc_core_b2x_idle), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n876) );
  AND2X2 AND2X2_2249 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n527), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n405_1_bF_buf3), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n881) );
  AND2X2 AND2X2_225 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n250_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_prech_page_closed), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n335) );
  AND2X2 AND2X2_2250 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n523_1_bF_buf1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n881), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n882) );
  AND2X2 AND2X2_2251 ( .A(u_sdrc_core_u_bank_ctl_x2b_ack_bF_buf0), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n461_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n885) );
  AND2X2 AND2X2_2252 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n886), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n537), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n887) );
  AND2X2 AND2X2_2253 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n887), .B(sdram_resetn_bF_buf26), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n888) );
  AND2X2 AND2X2_2254 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n543), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n890), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n891) );
  AND2X2 AND2X2_2255 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf3), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n891), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n892) );
  AND2X2 AND2X2_2256 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n895), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n446_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n896) );
  AND2X2 AND2X2_2257 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n896), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n550), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n897) );
  AND2X2 AND2X2_2258 ( .A(u_sdrc_core_u_bs_convert_x2a_wrnext_bF_buf0), .B(u_sdrc_core_a2x_wren_n_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n899) );
  AND2X2 AND2X2_2259 ( .A(u_sdrc_core_u_bs_convert_x2a_wrnext_bF_buf3), .B(u_sdrc_core_a2x_wren_n_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n901) );
  AND2X2 AND2X2_226 ( .A(sdram_resetn_bF_buf36), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_4_bF_buf3), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n337) );
  AND2X2 AND2X2_2260 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n883_bF_buf2), .B(_auto_iopadmap_cc_313_execute_24689_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n904) );
  AND2X2 AND2X2_2261 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n908), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n907), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n909) );
  AND2X2 AND2X2_2262 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n909), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n906), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n910) );
  AND2X2 AND2X2_2263 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n404_1), .B(u_sdrc_core_u_xfr_ctl_mgmt_st_5_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n912) );
  AND2X2 AND2X2_2264 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n912), .B(\cfg_sdr_mode_reg[11] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n913) );
  AND2X2 AND2X2_2265 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n911), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n913), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n914) );
  AND2X2 AND2X2_2266 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n883_bF_buf0), .B(_auto_iopadmap_cc_313_execute_24689_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n917) );
  AND2X2 AND2X2_2267 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n919), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n918), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n920) );
  AND2X2 AND2X2_2268 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n920), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n906), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n921) );
  AND2X2 AND2X2_2269 ( .A(u_sdrc_core_u_bank_ctl_x2b_ack_bF_buf0), .B(u_sdrc_core_b2x_addr_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n923) );
  AND2X2 AND2X2_227 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n337), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n336), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n338_1) );
  AND2X2 AND2X2_2270 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n523_1_bF_buf2), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n597), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n924) );
  AND2X2 AND2X2_2271 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n925), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n405_1_bF_buf2), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n926) );
  AND2X2 AND2X2_2272 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n912), .B(\cfg_sdr_mode_reg[0] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n927) );
  AND2X2 AND2X2_2273 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n929), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n930), .Y(u_sdrc_core_u_xfr_ctl_sdr_addr_0__FF_INPUT) );
  AND2X2 AND2X2_2274 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n523_1_bF_buf1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n621), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n932) );
  AND2X2 AND2X2_2275 ( .A(u_sdrc_core_u_bank_ctl_x2b_ack_bF_buf3), .B(u_sdrc_core_b2x_addr_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n933) );
  AND2X2 AND2X2_2276 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n934), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n405_1_bF_buf1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n935) );
  AND2X2 AND2X2_2277 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n912), .B(\cfg_sdr_mode_reg[1] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n936) );
  AND2X2 AND2X2_2278 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n938), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n939), .Y(u_sdrc_core_u_xfr_ctl_sdr_addr_1__FF_INPUT) );
  AND2X2 AND2X2_2279 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n523_1_bF_buf0), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n632), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n941) );
  AND2X2 AND2X2_228 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n338_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_ack), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n339_1) );
  AND2X2 AND2X2_2280 ( .A(u_sdrc_core_u_bank_ctl_x2b_ack_bF_buf2), .B(u_sdrc_core_b2x_addr_2_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n942) );
  AND2X2 AND2X2_2281 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n943), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n405_1_bF_buf0), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n944) );
  AND2X2 AND2X2_2282 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n912), .B(\cfg_sdr_mode_reg[2] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n945) );
  AND2X2 AND2X2_2283 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n947), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n948), .Y(u_sdrc_core_u_xfr_ctl_sdr_addr_2__FF_INPUT) );
  AND2X2 AND2X2_2284 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n523_1_bF_buf3), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n643), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n950) );
  AND2X2 AND2X2_2285 ( .A(u_sdrc_core_u_bank_ctl_x2b_ack_bF_buf1), .B(u_sdrc_core_b2x_addr_3_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n951) );
  AND2X2 AND2X2_2286 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n952), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n405_1_bF_buf3), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n953) );
  AND2X2 AND2X2_2287 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n912), .B(\cfg_sdr_mode_reg[3] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n954) );
  AND2X2 AND2X2_2288 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n956), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n957), .Y(u_sdrc_core_u_xfr_ctl_sdr_addr_3__FF_INPUT) );
  AND2X2 AND2X2_2289 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n523_1_bF_buf2), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n654), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n959) );
  AND2X2 AND2X2_229 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n339_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_sdr_dma_last), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n340) );
  AND2X2 AND2X2_2290 ( .A(u_sdrc_core_u_bank_ctl_x2b_ack_bF_buf0), .B(u_sdrc_core_b2x_addr_4_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n960) );
  AND2X2 AND2X2_2291 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n961), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n405_1_bF_buf2), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n962) );
  AND2X2 AND2X2_2292 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n912), .B(\cfg_sdr_mode_reg[4] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n963) );
  AND2X2 AND2X2_2293 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n965), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n966), .Y(u_sdrc_core_u_xfr_ctl_sdr_addr_4__FF_INPUT) );
  AND2X2 AND2X2_2294 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n523_1_bF_buf1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n665), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n968) );
  AND2X2 AND2X2_2295 ( .A(u_sdrc_core_u_bank_ctl_x2b_ack_bF_buf3), .B(u_sdrc_core_b2x_addr_5_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n969) );
  AND2X2 AND2X2_2296 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n970), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n405_1_bF_buf1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n971) );
  AND2X2 AND2X2_2297 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n912), .B(\cfg_sdr_mode_reg[5] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n972) );
  AND2X2 AND2X2_2298 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n974), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n975), .Y(u_sdrc_core_u_xfr_ctl_sdr_addr_5__FF_INPUT) );
  AND2X2 AND2X2_2299 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n523_1_bF_buf0), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n676), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n977) );
  AND2X2 AND2X2_23 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n249_1), .B(sdram_resetn_bF_buf49), .Y(u_sdrc_core_u_bank_ctl_rank_cnt_0__FF_INPUT) );
  AND2X2 AND2X2_230 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n250_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_2_bF_buf3), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n342) );
  AND2X2 AND2X2_2300 ( .A(u_sdrc_core_u_bank_ctl_x2b_ack_bF_buf2), .B(u_sdrc_core_b2x_addr_6_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n978) );
  AND2X2 AND2X2_2301 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n979), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n405_1_bF_buf0), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n980) );
  AND2X2 AND2X2_2302 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n912), .B(\cfg_sdr_mode_reg[6] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n981) );
  AND2X2 AND2X2_2303 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n983), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n984), .Y(u_sdrc_core_u_xfr_ctl_sdr_addr_6__FF_INPUT) );
  AND2X2 AND2X2_2304 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n523_1_bF_buf3), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n687), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n986) );
  AND2X2 AND2X2_2305 ( .A(u_sdrc_core_u_bank_ctl_x2b_ack_bF_buf1), .B(u_sdrc_core_b2x_addr_7_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n987) );
  AND2X2 AND2X2_2306 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n988), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n405_1_bF_buf3), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n989) );
  AND2X2 AND2X2_2307 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n912), .B(\cfg_sdr_mode_reg[7] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n990) );
  AND2X2 AND2X2_2308 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n992), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n993), .Y(u_sdrc_core_u_xfr_ctl_sdr_addr_7__FF_INPUT) );
  AND2X2 AND2X2_2309 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n523_1_bF_buf2), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n698), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n995) );
  AND2X2 AND2X2_231 ( .A(sdram_resetn_bF_buf35), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_ack), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n343_1) );
  AND2X2 AND2X2_2310 ( .A(u_sdrc_core_u_bank_ctl_x2b_ack_bF_buf0), .B(u_sdrc_core_b2x_addr_8_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n996) );
  AND2X2 AND2X2_2311 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n997), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n405_1_bF_buf2), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n998) );
  AND2X2 AND2X2_2312 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n912), .B(\cfg_sdr_mode_reg[8] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n999) );
  AND2X2 AND2X2_2313 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1001), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1002), .Y(u_sdrc_core_u_xfr_ctl_sdr_addr_8__FF_INPUT) );
  AND2X2 AND2X2_2314 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n523_1_bF_buf1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n709), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1004) );
  AND2X2 AND2X2_2315 ( .A(u_sdrc_core_u_bank_ctl_x2b_ack_bF_buf3), .B(u_sdrc_core_b2x_addr_9_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1005) );
  AND2X2 AND2X2_2316 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1006), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n405_1_bF_buf1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1007) );
  AND2X2 AND2X2_2317 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n912), .B(\cfg_sdr_mode_reg[9] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1008) );
  AND2X2 AND2X2_2318 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1010), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1011), .Y(u_sdrc_core_u_xfr_ctl_sdr_addr_9__FF_INPUT) );
  AND2X2 AND2X2_2319 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1016), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1015), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1017) );
  AND2X2 AND2X2_232 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n343_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_3_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n344_1) );
  AND2X2 AND2X2_2320 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1018), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1014), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1019) );
  AND2X2 AND2X2_2321 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1020), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1021), .Y(u_sdrc_core_u_xfr_ctl_sdr_addr_10__FF_INPUT) );
  AND2X2 AND2X2_2322 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1024), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n405_1_bF_buf0), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1025) );
  AND2X2 AND2X2_2323 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1025), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1023), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1026) );
  AND2X2 AND2X2_2324 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1026), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n911), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1027) );
  AND2X2 AND2X2_2325 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n883_bF_buf0), .B(_auto_iopadmap_cc_313_execute_24675_11_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1028) );
  AND2X2 AND2X2_2326 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1032), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n405_1_bF_buf3), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1033) );
  AND2X2 AND2X2_2327 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1033), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1031), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1034) );
  AND2X2 AND2X2_2328 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n912), .B(\cfg_sdr_mode_reg[12] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1035) );
  AND2X2 AND2X2_2329 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1037), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1038), .Y(u_sdrc_core_u_xfr_ctl_sdr_addr_12__FF_INPUT) );
  AND2X2 AND2X2_233 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n337), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_refresh), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n345) );
  AND2X2 AND2X2_2330 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n404_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n401_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1040) );
  AND2X2 AND2X2_2331 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n392), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n397), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1041) );
  AND2X2 AND2X2_2332 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n396_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n393_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1042) );
  AND2X2 AND2X2_2333 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1042), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n871_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1043) );
  AND2X2 AND2X2_2334 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1043), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1041), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1044) );
  AND2X2 AND2X2_2335 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1045), .B(\cfg_sdr_trcar_d[0] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1046) );
  AND2X2 AND2X2_2336 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1047), .B(\cfg_sdr_trp_d[0] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1048) );
  AND2X2 AND2X2_2337 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1040), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1050), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1051) );
  AND2X2 AND2X2_2338 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n353_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1053), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1054) );
  AND2X2 AND2X2_2339 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1052), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1054), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1055) );
  AND2X2 AND2X2_234 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n343_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_2_bF_buf2), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n348_1) );
  AND2X2 AND2X2_2340 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1056), .B(sdram_resetn_bF_buf25), .Y(u_sdrc_core_u_xfr_ctl_tmr0_0__FF_INPUT) );
  AND2X2 AND2X2_2341 ( .A(u_sdrc_core_u_xfr_ctl_tmr0_0_), .B(u_sdrc_core_u_xfr_ctl_tmr0_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1059) );
  AND2X2 AND2X2_2342 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n353_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1060), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1061) );
  AND2X2 AND2X2_2343 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1052), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1061), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1062) );
  AND2X2 AND2X2_2344 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1045), .B(\cfg_sdr_trcar_d[1] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1063) );
  AND2X2 AND2X2_2345 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1047), .B(\cfg_sdr_trp_d[1] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1064) );
  AND2X2 AND2X2_2346 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1040), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1066), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1067) );
  AND2X2 AND2X2_2347 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1068), .B(sdram_resetn_bF_buf24), .Y(u_sdrc_core_u_xfr_ctl_tmr0_1__FF_INPUT) );
  AND2X2 AND2X2_2348 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n351_1), .B(u_sdrc_core_u_xfr_ctl_tmr0_2_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1070) );
  AND2X2 AND2X2_2349 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1071), .B(u_sdrc_core_u_xfr_ctl_tmr0_3_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1072) );
  AND2X2 AND2X2_235 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n338_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n249_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n349_1) );
  AND2X2 AND2X2_2350 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1052), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1073), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1074) );
  AND2X2 AND2X2_2351 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1047), .B(\cfg_sdr_trp_d[2] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1075) );
  AND2X2 AND2X2_2352 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1045), .B(\cfg_sdr_trcar_d[2] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1076) );
  AND2X2 AND2X2_2353 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1040), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1078), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1079) );
  AND2X2 AND2X2_2354 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1080), .B(sdram_resetn_bF_buf23), .Y(u_sdrc_core_u_xfr_ctl_tmr0_2__FF_INPUT) );
  AND2X2 AND2X2_2355 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1045), .B(\cfg_sdr_trcar_d[3] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1082) );
  AND2X2 AND2X2_2356 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1047), .B(\cfg_sdr_trp_d[3] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1083) );
  AND2X2 AND2X2_2357 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1040), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1084), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1085) );
  AND2X2 AND2X2_2358 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n352), .B(u_sdrc_core_u_xfr_ctl_tmr0_3_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1086) );
  AND2X2 AND2X2_2359 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1052), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1086), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1087) );
  AND2X2 AND2X2_236 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n331_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n253_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n351) );
  AND2X2 AND2X2_2360 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1088), .B(sdram_resetn_bF_buf22), .Y(u_sdrc_core_u_xfr_ctl_tmr0_3__FF_INPUT) );
  AND2X2 AND2X2_2361 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n444_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n433), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1090) );
  AND2X2 AND2X2_2362 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1093), .B(u_sdrc_core_u_xfr_ctl_cntr1_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1094) );
  AND2X2 AND2X2_2363 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n539_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n357), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1095) );
  AND2X2 AND2X2_2364 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1096), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1092), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1097) );
  AND2X2 AND2X2_2365 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n393_1), .B(u_sdrc_core_u_xfr_ctl_rfsh_row_cnt_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1100) );
  AND2X2 AND2X2_2366 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1091), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1101), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1102) );
  AND2X2 AND2X2_2367 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1105), .B(u_sdrc_core_u_xfr_ctl_cntr1_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1106) );
  AND2X2 AND2X2_2368 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1095), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n358_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1107) );
  AND2X2 AND2X2_2369 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1108), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1092), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1109) );
  AND2X2 AND2X2_237 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n339_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n353_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n354_1) );
  AND2X2 AND2X2_2370 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n393_1), .B(u_sdrc_core_u_xfr_ctl_rfsh_row_cnt_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1110) );
  AND2X2 AND2X2_2371 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1091), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1111), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1112) );
  AND2X2 AND2X2_2372 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1115), .B(u_sdrc_core_u_xfr_ctl_cntr1_2_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1116) );
  AND2X2 AND2X2_2373 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1107), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n356_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1117) );
  AND2X2 AND2X2_2374 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1118), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1092), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1119) );
  AND2X2 AND2X2_2375 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n393_1), .B(u_sdrc_core_u_xfr_ctl_rfsh_row_cnt_2_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1120) );
  AND2X2 AND2X2_2376 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1091), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1121), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1122) );
  AND2X2 AND2X2_2377 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1125), .B(u_sdrc_core_u_xfr_ctl_cntr1_3_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1126) );
  AND2X2 AND2X2_2378 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n539_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n361), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1127) );
  AND2X2 AND2X2_2379 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1128), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1092), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1129) );
  AND2X2 AND2X2_238 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n356), .B(sdram_resetn_bF_buf34), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n357) );
  AND2X2 AND2X2_2380 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1130), .B(sdram_resetn_bF_buf21), .Y(u_sdrc_core_u_xfr_ctl_cntr1_3__FF_INPUT) );
  AND2X2 AND2X2_2381 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1134), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1136), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1137) );
  AND2X2 AND2X2_2382 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1139), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1141), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1142) );
  AND2X2 AND2X2_2383 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1137), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1142), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1143) );
  AND2X2 AND2X2_2384 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1145), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1147), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1148) );
  AND2X2 AND2X2_2385 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1143), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1148), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1149) );
  AND2X2 AND2X2_2386 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1151), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1153), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1154) );
  AND2X2 AND2X2_2387 ( .A(\cfg_sdr_rfsh[9] ), .B(u_sdrc_core_u_xfr_ctl_rfsh_timer_9_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1156) );
  AND2X2 AND2X2_2388 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1157), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1155), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1158) );
  AND2X2 AND2X2_2389 ( .A(\cfg_sdr_rfsh[8] ), .B(u_sdrc_core_u_xfr_ctl_rfsh_timer_8_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1160) );
  AND2X2 AND2X2_239 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n355), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n358_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n359_1) );
  AND2X2 AND2X2_2390 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1161), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1162), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1163) );
  AND2X2 AND2X2_2391 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1159), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1164), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1165) );
  AND2X2 AND2X2_2392 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1165), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1154), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1166) );
  AND2X2 AND2X2_2393 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1166), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1149), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1167) );
  AND2X2 AND2X2_2394 ( .A(\cfg_sdr_rfsh[3] ), .B(u_sdrc_core_u_xfr_ctl_rfsh_timer_3_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1169) );
  AND2X2 AND2X2_2395 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1170), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1168), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1171) );
  AND2X2 AND2X2_2396 ( .A(\cfg_sdr_rfsh[1] ), .B(u_sdrc_core_u_xfr_ctl_rfsh_timer_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1174) );
  AND2X2 AND2X2_2397 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1175), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1173), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1176) );
  AND2X2 AND2X2_2398 ( .A(\cfg_sdr_rfsh[0] ), .B(u_sdrc_core_u_xfr_ctl_rfsh_timer_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1178) );
  AND2X2 AND2X2_2399 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1179), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1132), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1180) );
  AND2X2 AND2X2_24 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n245_1), .B(u_sdrc_core_u_bank_ctl_rank_cnt_1_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n251_1) );
  AND2X2 AND2X2_240 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n360), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_0_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n361) );
  AND2X2 AND2X2_2400 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1177), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1181), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1182) );
  AND2X2 AND2X2_2401 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1182), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1172), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1183) );
  AND2X2 AND2X2_2402 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1185), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1187), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1188) );
  AND2X2 AND2X2_2403 ( .A(\cfg_sdr_rfsh[10] ), .B(u_sdrc_core_u_xfr_ctl_rfsh_timer_10_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1189) );
  AND2X2 AND2X2_2404 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1190), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1191), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1192) );
  AND2X2 AND2X2_2405 ( .A(\cfg_sdr_rfsh[6] ), .B(u_sdrc_core_u_xfr_ctl_rfsh_timer_6_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1194) );
  AND2X2 AND2X2_2406 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1195), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1196), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1197) );
  AND2X2 AND2X2_2407 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1193), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1198), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1199) );
  AND2X2 AND2X2_2408 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1199), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1188), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1200) );
  AND2X2 AND2X2_2409 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1183), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1200), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1201) );
  AND2X2 AND2X2_241 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_4_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_write), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n364_1) );
  AND2X2 AND2X2_2410 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1201), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1167), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1202) );
  AND2X2 AND2X2_2411 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1203), .B(sdram_resetn_bF_buf20), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1204) );
  AND2X2 AND2X2_2412 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1204), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1132), .Y(u_sdrc_core_u_xfr_ctl_rfsh_timer_0__FF_INPUT) );
  AND2X2 AND2X2_2413 ( .A(u_sdrc_core_u_xfr_ctl_rfsh_timer_0_), .B(u_sdrc_core_u_xfr_ctl_rfsh_timer_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1207) );
  AND2X2 AND2X2_2414 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1208), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1206), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1209) );
  AND2X2 AND2X2_2415 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1204), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1209), .Y(u_sdrc_core_u_xfr_ctl_rfsh_timer_1__FF_INPUT) );
  AND2X2 AND2X2_2416 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1207), .B(u_sdrc_core_u_xfr_ctl_rfsh_timer_2_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1212) );
  AND2X2 AND2X2_2417 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1213), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1211), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1214) );
  AND2X2 AND2X2_2418 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1204), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1214), .Y(u_sdrc_core_u_xfr_ctl_rfsh_timer_2__FF_INPUT) );
  AND2X2 AND2X2_2419 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1212), .B(u_sdrc_core_u_xfr_ctl_rfsh_timer_3_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1217) );
  AND2X2 AND2X2_242 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n369_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n367), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n370) );
  AND2X2 AND2X2_2420 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1218), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1216), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1219) );
  AND2X2 AND2X2_2421 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1204), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1219), .Y(u_sdrc_core_u_xfr_ctl_rfsh_timer_3__FF_INPUT) );
  AND2X2 AND2X2_2422 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1217), .B(u_sdrc_core_u_xfr_ctl_rfsh_timer_4_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1222) );
  AND2X2 AND2X2_2423 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1223), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1221), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1224) );
  AND2X2 AND2X2_2424 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1204), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1224), .Y(u_sdrc_core_u_xfr_ctl_rfsh_timer_4__FF_INPUT) );
  AND2X2 AND2X2_2425 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1222), .B(u_sdrc_core_u_xfr_ctl_rfsh_timer_5_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1227) );
  AND2X2 AND2X2_2426 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1228), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1226), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1229) );
  AND2X2 AND2X2_2427 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1204), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1229), .Y(u_sdrc_core_u_xfr_ctl_rfsh_timer_5__FF_INPUT) );
  AND2X2 AND2X2_2428 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1227), .B(u_sdrc_core_u_xfr_ctl_rfsh_timer_6_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1232) );
  AND2X2 AND2X2_2429 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1233), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1231), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1234) );
  AND2X2 AND2X2_243 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n370), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n371) );
  AND2X2 AND2X2_2430 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1204), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1234), .Y(u_sdrc_core_u_xfr_ctl_rfsh_timer_6__FF_INPUT) );
  AND2X2 AND2X2_2431 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1232), .B(u_sdrc_core_u_xfr_ctl_rfsh_timer_7_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1236) );
  AND2X2 AND2X2_2432 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1204), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1238), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1239) );
  AND2X2 AND2X2_2433 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1239), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1237), .Y(u_sdrc_core_u_xfr_ctl_rfsh_timer_7__FF_INPUT) );
  AND2X2 AND2X2_2434 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1236), .B(u_sdrc_core_u_xfr_ctl_rfsh_timer_8_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1241) );
  AND2X2 AND2X2_2435 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1204), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1243), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1244) );
  AND2X2 AND2X2_2436 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1244), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1242), .Y(u_sdrc_core_u_xfr_ctl_rfsh_timer_8__FF_INPUT) );
  AND2X2 AND2X2_2437 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1241), .B(u_sdrc_core_u_xfr_ctl_rfsh_timer_9_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1246) );
  AND2X2 AND2X2_2438 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1248), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1204), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1249) );
  AND2X2 AND2X2_2439 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1249), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1247), .Y(u_sdrc_core_u_xfr_ctl_rfsh_timer_9__FF_INPUT) );
  AND2X2 AND2X2_244 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n371), .B(u_sdrc_core_r2b_write), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n372) );
  AND2X2 AND2X2_2440 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1246), .B(u_sdrc_core_u_xfr_ctl_rfsh_timer_10_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1251) );
  AND2X2 AND2X2_2441 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1253), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1204), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1254) );
  AND2X2 AND2X2_2442 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1254), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1252), .Y(u_sdrc_core_u_xfr_ctl_rfsh_timer_10__FF_INPUT) );
  AND2X2 AND2X2_2443 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1252), .B(u_sdrc_core_u_xfr_ctl_rfsh_timer_11_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1256) );
  AND2X2 AND2X2_2444 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1251), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1152), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1257) );
  AND2X2 AND2X2_2445 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1258), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1204), .Y(u_sdrc_core_u_xfr_ctl_rfsh_timer_11__FF_INPUT) );
  AND2X2 AND2X2_2446 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1202), .B(u_sdrc_core_u_xfr_ctl_rfsh_row_cnt_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1260) );
  AND2X2 AND2X2_2447 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1262), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n873), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1263) );
  AND2X2 AND2X2_2448 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1263), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1261), .Y(u_sdrc_core_u_xfr_ctl_rfsh_row_cnt_0__FF_INPUT) );
  AND2X2 AND2X2_2449 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1260), .B(u_sdrc_core_u_xfr_ctl_rfsh_row_cnt_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1265) );
  AND2X2 AND2X2_245 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n331_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n372), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n373_1) );
  AND2X2 AND2X2_2450 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1267), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n873), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1268) );
  AND2X2 AND2X2_2451 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1268), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1266), .Y(u_sdrc_core_u_xfr_ctl_rfsh_row_cnt_1__FF_INPUT) );
  AND2X2 AND2X2_2452 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1265), .B(u_sdrc_core_u_xfr_ctl_rfsh_row_cnt_2_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1270) );
  AND2X2 AND2X2_2453 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1272), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n873), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1273) );
  AND2X2 AND2X2_2454 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1273), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1271), .Y(u_sdrc_core_u_xfr_ctl_rfsh_row_cnt_2__FF_INPUT) );
  AND2X2 AND2X2_2455 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1275), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1276), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1277) );
  AND2X2 AND2X2_2456 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1281), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1279), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1282) );
  AND2X2 AND2X2_2457 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1278), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1282), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1283) );
  AND2X2 AND2X2_2458 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1284), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1285), .Y(u_sdrc_core_u_bs_convert_x2a_rdok) );
  AND2X2 AND2X2_2459 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1288), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1280), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1289) );
  AND2X2 AND2X2_246 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n374_1), .B(sdram_resetn_bF_buf33), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_cmd_r_0__FF_INPUT) );
  AND2X2 AND2X2_2460 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1289), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1287), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1290) );
  AND2X2 AND2X2_2461 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n562), .B(u_sdrc_core_u_xfr_ctl_l_rd_last_4_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1291) );
  AND2X2 AND2X2_2462 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1294), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n561), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1295) );
  AND2X2 AND2X2_2463 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1293), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1295), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1296) );
  AND2X2 AND2X2_2464 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n560_1), .B(u_sdrc_core_u_xfr_ctl_l_rd_last_2_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1297) );
  AND2X2 AND2X2_2465 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1312), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1311), .Y(u_sdrc_core_u_xfr_ctl_sdr_dout_0__FF_INPUT) );
  AND2X2 AND2X2_2466 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1315), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1314), .Y(u_sdrc_core_u_xfr_ctl_sdr_dout_1__FF_INPUT) );
  AND2X2 AND2X2_2467 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1318), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1317), .Y(u_sdrc_core_u_xfr_ctl_sdr_dout_2__FF_INPUT) );
  AND2X2 AND2X2_2468 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1321), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1320), .Y(u_sdrc_core_u_xfr_ctl_sdr_dout_3__FF_INPUT) );
  AND2X2 AND2X2_2469 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1324), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1323), .Y(u_sdrc_core_u_xfr_ctl_sdr_dout_4__FF_INPUT) );
  AND2X2 AND2X2_247 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n371), .B(sdram_resetn_bF_buf32), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n376) );
  AND2X2 AND2X2_2470 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1327), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1326), .Y(u_sdrc_core_u_xfr_ctl_sdr_dout_5__FF_INPUT) );
  AND2X2 AND2X2_2471 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1330), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1329), .Y(u_sdrc_core_u_xfr_ctl_sdr_dout_6__FF_INPUT) );
  AND2X2 AND2X2_2472 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1333), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1332), .Y(u_sdrc_core_u_xfr_ctl_sdr_dout_7__FF_INPUT) );
  AND2X2 AND2X2_2473 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1336), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1335), .Y(u_sdrc_core_u_xfr_ctl_sdr_dout_8__FF_INPUT) );
  AND2X2 AND2X2_2474 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1339), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1338), .Y(u_sdrc_core_u_xfr_ctl_sdr_dout_9__FF_INPUT) );
  AND2X2 AND2X2_2475 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1342), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1341), .Y(u_sdrc_core_u_xfr_ctl_sdr_dout_10__FF_INPUT) );
  AND2X2 AND2X2_2476 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1345), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1344), .Y(u_sdrc_core_u_xfr_ctl_sdr_dout_11__FF_INPUT) );
  AND2X2 AND2X2_2477 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1348), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1347), .Y(u_sdrc_core_u_xfr_ctl_sdr_dout_12__FF_INPUT) );
  AND2X2 AND2X2_2478 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1351), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1350), .Y(u_sdrc_core_u_xfr_ctl_sdr_dout_13__FF_INPUT) );
  AND2X2 AND2X2_2479 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1354), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1353), .Y(u_sdrc_core_u_xfr_ctl_sdr_dout_14__FF_INPUT) );
  AND2X2 AND2X2_248 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n331_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n376), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n377) );
  AND2X2 AND2X2_2480 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1357), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1356), .Y(u_sdrc_core_u_xfr_ctl_sdr_dout_15__FF_INPUT) );
  AND2X2 AND2X2_2481 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1360), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n444_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_wrok) );
  AND2X2 AND2X2_2482 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n845_1), .B(sdram_resetn_bF_buf19), .Y(u_sdrc_core_u_xfr_ctl_l_last_FF_INPUT) );
  AND2X2 AND2X2_2483 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n614_bF_buf0), .B(u_sdrc_core_b2x_wrap), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1363) );
  AND2X2 AND2X2_2484 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf2), .B(u_sdrc_core_u_xfr_ctl_l_wrap), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1364) );
  AND2X2 AND2X2_2485 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1365), .B(sdram_resetn_bF_buf18), .Y(u_sdrc_core_u_xfr_ctl_l_wrap_FF_INPUT) );
  AND2X2 AND2X2_2486 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n888), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n892), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1367) );
  AND2X2 AND2X2_2487 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1367), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n541), .Y(u_sdrc_core_u_xfr_ctl_act_cmd_FF_INPUT) );
  AND2X2 AND2X2_2488 ( .A(sdram_resetn_bF_buf17), .B(u_sdrc_core_u_xfr_ctl_act_cmd), .Y(u_sdrc_core_u_xfr_ctl_d_act_cmd_FF_INPUT) );
  AND2X2 AND2X2_2489 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1370), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n378), .Y(u_sdrc_core_u_xfr_ctl_sdr_init_done_FF_INPUT) );
  AND2X2 AND2X2_249 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n381), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_cmd_0_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n382) );
  AND2X2 AND2X2_2490 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1374), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1375), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_act_ok) );
  AND2X2 AND2X2_2491 ( .A(wb_cyc_i), .B(wb_stb_i), .Y(u_wb2sdrc__abc_24125_n29_1) );
  AND2X2 AND2X2_2492 ( .A(u_wb2sdrc__abc_24125_n29_1), .B(u_wb2sdrc__abc_24125_n28_1), .Y(u_wb2sdrc__abc_24125_n30) );
  AND2X2 AND2X2_2493 ( .A(u_wb2sdrc__abc_24125_n31), .B(wb_we_i), .Y(u_wb2sdrc__abc_24125_n32) );
  AND2X2 AND2X2_2494 ( .A(u_wb2sdrc__abc_24125_n30), .B(u_wb2sdrc__abc_24125_n32), .Y(u_wb2sdrc_u_wrdatafifo_wr_en) );
  AND2X2 AND2X2_2495 ( .A(u_wb2sdrc_u_cmdfifo_wr_data_26_), .B(u_wb2sdrc__abc_24125_n39_1), .Y(u_wb2sdrc__abc_24125_n40) );
  AND2X2 AND2X2_2496 ( .A(u_wb2sdrc__abc_24125_n30), .B(u_wb2sdrc__abc_24125_n40), .Y(u_wb2sdrc__abc_24125_n41) );
  AND2X2 AND2X2_2497 ( .A(u_wb2sdrc__abc_24125_n36_1), .B(u_wb2sdrc_pending_read), .Y(u_wb2sdrc__abc_24125_n47) );
  AND2X2 AND2X2_2498 ( .A(u_wb2sdrc_u_cmdfifo_sync_rd_ptr_1_1_), .B(u_wb2sdrc_u_cmdfifo_sync_rd_ptr_2_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n400_1) );
  AND2X2 AND2X2_2499 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n401_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n399), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n402) );
  AND2X2 AND2X2_25 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n217_1), .B(u_sdrc_core_u_bank_ctl_rank_cnt_1_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n253_1) );
  AND2X2 AND2X2_250 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n383_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n386_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n387_1) );
  AND2X2 AND2X2_2500 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n403_1), .B(u_wb2sdrc_u_cmdfifo_wr_ptr_1_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n404_1) );
  AND2X2 AND2X2_2501 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n403_1), .B(u_wb2sdrc_u_cmdfifo_sync_rd_ptr_1_0_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n407_1) );
  AND2X2 AND2X2_2502 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n402), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n408), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n409_1) );
  AND2X2 AND2X2_2503 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n410_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n406_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n411) );
  AND2X2 AND2X2_2504 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n402), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n412_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n413_1) );
  AND2X2 AND2X2_2505 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n415_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n405), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n416_1) );
  AND2X2 AND2X2_2506 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n417), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n418_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n419_1) );
  AND2X2 AND2X2_2507 ( .A(u_wb2sdrc_u_cmdfifo_sync_rd_ptr_2_), .B(u_wb2sdrc_u_cmdfifo_wr_ptr_2_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n420) );
  AND2X2 AND2X2_2508 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n416_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n422_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n423) );
  AND2X2 AND2X2_2509 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n424_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n421_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n425_1) );
  AND2X2 AND2X2_251 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n387_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n379_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n388) );
  AND2X2 AND2X2_2510 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n427_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n428_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n429) );
  AND2X2 AND2X2_2511 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n414), .B(u_wb2sdrc_u_cmdfifo_wr_ptr_0_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n432) );
  AND2X2 AND2X2_2512 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n433_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n431_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n434_1) );
  AND2X2 AND2X2_2513 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n426), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n434_1), .Y(u_wb2sdrc_u_cmdfifo_afull) );
  AND2X2 AND2X2_2514 ( .A(u_wb2sdrc_u_cmdfifo_sync_wr_ptr_1_1_), .B(u_wb2sdrc_u_cmdfifo_sync_wr_ptr_2_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n438) );
  AND2X2 AND2X2_2515 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n439_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n437_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n440_1) );
  AND2X2 AND2X2_2516 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n440_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf5), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n441) );
  AND2X2 AND2X2_2517 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n443_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n444), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n445_1) );
  AND2X2 AND2X2_2518 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n446_1), .B(u_wb2sdrc_u_cmdfifo_sync_wr_ptr_1_0_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n447) );
  AND2X2 AND2X2_2519 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n440_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n448_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n449_1) );
  AND2X2 AND2X2_252 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n382), .B(\cfg_sdr_tras_d[0] ), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n389) );
  AND2X2 AND2X2_2520 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n446_1), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf4), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n452_1) );
  AND2X2 AND2X2_2521 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n451_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n454_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n455) );
  AND2X2 AND2X2_2522 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n457_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n459_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n460_1) );
  AND2X2 AND2X2_2523 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n456_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n460_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n461_1) );
  AND2X2 AND2X2_2524 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n464_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n463_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n465_1) );
  AND2X2 AND2X2_2525 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n465_1), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf6), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n466_1) );
  AND2X2 AND2X2_2526 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n467_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n462_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n468_1) );
  AND2X2 AND2X2_2527 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n468_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n469_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n470_1) );
  AND2X2 AND2X2_2528 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n466_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n453), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n472_1) );
  AND2X2 AND2X2_2529 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n450), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf6), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n474_1) );
  AND2X2 AND2X2_253 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n390), .B(sdram_resetn_bF_buf31), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_tras_cntr_0__FF_INPUT) );
  AND2X2 AND2X2_2530 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n473_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n475_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n476_1) );
  AND2X2 AND2X2_2531 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n471_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n476_1), .Y(u_wb2sdrc_u_cmdfifo_aempty) );
  AND2X2 AND2X2_2532 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n406_1), .B(u_wb2sdrc_cmdfifo_wr), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n478_1) );
  AND2X2 AND2X2_2533 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n478_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n412_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1) );
  AND2X2 AND2X2_2534 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n482_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n480_1), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n99) );
  AND2X2 AND2X2_2535 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n485_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n484_1), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n102) );
  AND2X2 AND2X2_2536 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n488_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n487_1), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n105) );
  AND2X2 AND2X2_2537 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n491_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n490_1), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n108) );
  AND2X2 AND2X2_2538 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n494_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n493_1), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n111) );
  AND2X2 AND2X2_2539 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n497_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n496_1), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n114) );
  AND2X2 AND2X2_254 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n382), .B(\cfg_sdr_tras_d[1] ), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n392_1) );
  AND2X2 AND2X2_2540 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n500_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n499_1), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n117) );
  AND2X2 AND2X2_2541 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n503_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n502_1), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n120) );
  AND2X2 AND2X2_2542 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n506_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n505_1), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n123) );
  AND2X2 AND2X2_2543 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n509_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n508_1), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n126) );
  AND2X2 AND2X2_2544 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n512_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n511_1), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n129) );
  AND2X2 AND2X2_2545 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n515_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n514_1), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n132) );
  AND2X2 AND2X2_2546 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n518_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n517_1), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n135) );
  AND2X2 AND2X2_2547 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n521_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n520_1), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n138) );
  AND2X2 AND2X2_2548 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n524_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n523_1), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n141) );
  AND2X2 AND2X2_2549 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n527_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n526_1), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n144) );
  AND2X2 AND2X2_255 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_tras_cntr_0_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_tras_cntr_1_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n394_1) );
  AND2X2 AND2X2_2550 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n530_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n529), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n147) );
  AND2X2 AND2X2_2551 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n533_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n532_1), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n150) );
  AND2X2 AND2X2_2552 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n536_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n535_1), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n153) );
  AND2X2 AND2X2_2553 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n539_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n538_1), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n156) );
  AND2X2 AND2X2_2554 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n542_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n541_1), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n159) );
  AND2X2 AND2X2_2555 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n545_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n544_1), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n162) );
  AND2X2 AND2X2_2556 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n548_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n547_1), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n165) );
  AND2X2 AND2X2_2557 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n551_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n550_1), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n168) );
  AND2X2 AND2X2_2558 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n554_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n553_1), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n171) );
  AND2X2 AND2X2_2559 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n557_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n556_1), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n174) );
  AND2X2 AND2X2_256 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n387_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n395_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n396_1) );
  AND2X2 AND2X2_2560 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n560_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n559_1), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n177) );
  AND2X2 AND2X2_2561 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n563_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n562_1), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n180) );
  AND2X2 AND2X2_2562 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n566), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n565_1), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n183) );
  AND2X2 AND2X2_2563 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n569), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n568), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n186) );
  AND2X2 AND2X2_2564 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n572), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n571), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n189) );
  AND2X2 AND2X2_2565 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n575), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n574), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n192) );
  AND2X2 AND2X2_2566 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n578), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n577), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n195) );
  AND2X2 AND2X2_2567 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n581), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n580), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n198) );
  AND2X2 AND2X2_2568 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n584), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n583), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n201) );
  AND2X2 AND2X2_2569 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n587), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n586), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n204) );
  AND2X2 AND2X2_257 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n397_1), .B(sdram_resetn_bF_buf30), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_tras_cntr_1__FF_INPUT) );
  AND2X2 AND2X2_2570 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf4), .B(app_req_ack_bF_buf0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n589) );
  AND2X2 AND2X2_2571 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n590), .B(u_wb2sdrc_u_cmdfifo_grey_rd_ptr_0_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n591) );
  AND2X2 AND2X2_2572 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf5), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n593) );
  AND2X2 AND2X2_2573 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf3), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf5), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n594) );
  AND2X2 AND2X2_2574 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n593), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_2_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n596) );
  AND2X2 AND2X2_2575 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n597), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n598), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n599) );
  AND2X2 AND2X2_2576 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n599), .B(app_req_ack_bF_buf5), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n600) );
  AND2X2 AND2X2_2577 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n600), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n595), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n601) );
  AND2X2 AND2X2_2578 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n590), .B(u_wb2sdrc_u_cmdfifo_grey_rd_ptr_1_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n602) );
  AND2X2 AND2X2_2579 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n603), .B(app_req_ack_bF_buf4), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n604) );
  AND2X2 AND2X2_258 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n382), .B(\cfg_sdr_tras_d[2] ), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n399_1) );
  AND2X2 AND2X2_2580 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n604), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n458_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n605) );
  AND2X2 AND2X2_2581 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n590), .B(u_wb2sdrc_u_cmdfifo_grey_rd_ptr_2_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n608) );
  AND2X2 AND2X2_2582 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf4), .B(app_req_ack_bF_buf3), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n610) );
  AND2X2 AND2X2_2583 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n590), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf4), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n611) );
  AND2X2 AND2X2_2584 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n590), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf2), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n613) );
  AND2X2 AND2X2_2585 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n590), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_2_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n615) );
  AND2X2 AND2X2_2586 ( .A(u_wb2sdrc_u_cmdfifo_aempty), .B(app_req_ack_bF_buf2), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n617) );
  AND2X2 AND2X2_2587 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n473_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n619), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n620) );
  AND2X2 AND2X2_2588 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n471_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n620), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n621) );
  AND2X2 AND2X2_2589 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n618), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n622), .Y(u_wb2sdrc_u_cmdfifo_empty_q_FF_INPUT) );
  AND2X2 AND2X2_259 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n384_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_tras_cntr_2_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n401_1) );
  AND2X2 AND2X2_2590 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n624), .B(u_wb2sdrc_u_cmdfifo_wr_ptr_0_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n625) );
  AND2X2 AND2X2_2591 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n478_1), .B(u_wb2sdrc_u_cmdfifo_wr_ptr_1_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n627) );
  AND2X2 AND2X2_2592 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n624), .B(u_wb2sdrc_u_cmdfifo_wr_ptr_1_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n628) );
  AND2X2 AND2X2_2593 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n412_1), .B(u_wb2sdrc_cmdfifo_wr), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n629) );
  AND2X2 AND2X2_2594 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n629), .B(u_wb2sdrc_u_cmdfifo_wr_ptr_0_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n630) );
  AND2X2 AND2X2_2595 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n624), .B(u_wb2sdrc_u_cmdfifo_wr_ptr_2_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n633) );
  AND2X2 AND2X2_2596 ( .A(u_wb2sdrc_u_cmdfifo_wr_ptr_1_), .B(u_wb2sdrc_u_cmdfifo_wr_ptr_0_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n634) );
  AND2X2 AND2X2_2597 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n634), .B(u_wb2sdrc_u_cmdfifo_wr_ptr_2_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n635) );
  AND2X2 AND2X2_2598 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n637), .B(u_wb2sdrc_cmdfifo_wr), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n638) );
  AND2X2 AND2X2_2599 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n638), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n636), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n639) );
  AND2X2 AND2X2_26 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n218_1), .B(u_sdrc_core_u_bank_ctl_rank_cnt_0_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n255) );
  AND2X2 AND2X2_260 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n387_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n402_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n403_1) );
  AND2X2 AND2X2_2600 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n624), .B(u_wb2sdrc_u_cmdfifo_grey_wr_ptr_0_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n641) );
  AND2X2 AND2X2_2601 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n412_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n406_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n644) );
  AND2X2 AND2X2_2602 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n646), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n647), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n648) );
  AND2X2 AND2X2_2603 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n649), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n643), .Y(u_wb2sdrc_u_cmdfifo_grey_wr_ptr_1__FF_INPUT) );
  AND2X2 AND2X2_2604 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n624), .B(u_wb2sdrc_u_cmdfifo_grey_wr_ptr_2_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n651) );
  AND2X2 AND2X2_2605 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n653), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n655), .Y(u_wb2sdrc_u_cmdfifo_full_q_FF_INPUT) );
  AND2X2 AND2X2_2606 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n658), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n657), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n659) );
  AND2X2 AND2X2_2607 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n659), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf2), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n660) );
  AND2X2 AND2X2_2608 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n662), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n663) );
  AND2X2 AND2X2_2609 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n663), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n661), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n664) );
  AND2X2 AND2X2_261 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n404_1), .B(sdram_resetn_bF_buf29), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_tras_cntr_2__FF_INPUT) );
  AND2X2 AND2X2_2610 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n667), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n666), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n668) );
  AND2X2 AND2X2_2611 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n668), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n669) );
  AND2X2 AND2X2_2612 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n671), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n672) );
  AND2X2 AND2X2_2613 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n672), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n670), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n673) );
  AND2X2 AND2X2_2614 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n676), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n675), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n677) );
  AND2X2 AND2X2_2615 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n677), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n678) );
  AND2X2 AND2X2_2616 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n680), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf5), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n681) );
  AND2X2 AND2X2_2617 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n681), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n679), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n682) );
  AND2X2 AND2X2_2618 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n685), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n684), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n686) );
  AND2X2 AND2X2_2619 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n686), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf5), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n687) );
  AND2X2 AND2X2_262 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n385), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_tras_cntr_3_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n406_1) );
  AND2X2 AND2X2_2620 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n689), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf4), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n690) );
  AND2X2 AND2X2_2621 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n690), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n688), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n691) );
  AND2X2 AND2X2_2622 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n694), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n693), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n695) );
  AND2X2 AND2X2_2623 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n695), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf4), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n696) );
  AND2X2 AND2X2_2624 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n698), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf3), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n699) );
  AND2X2 AND2X2_2625 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n699), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n697), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n700) );
  AND2X2 AND2X2_2626 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n703), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n702), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n704) );
  AND2X2 AND2X2_2627 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n704), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf3), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n705) );
  AND2X2 AND2X2_2628 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n707), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf2), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n708) );
  AND2X2 AND2X2_2629 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n708), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n706), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n709) );
  AND2X2 AND2X2_263 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n408_1), .B(sdram_resetn_bF_buf28), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n409_1) );
  AND2X2 AND2X2_2630 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n712), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n711), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n713) );
  AND2X2 AND2X2_2631 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n713), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf2), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n714) );
  AND2X2 AND2X2_2632 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n716), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n717) );
  AND2X2 AND2X2_2633 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n717), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n715), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n718) );
  AND2X2 AND2X2_2634 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n721), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n720), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n722) );
  AND2X2 AND2X2_2635 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n722), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n723) );
  AND2X2 AND2X2_2636 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n725), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n726) );
  AND2X2 AND2X2_2637 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n726), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n724), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n727) );
  AND2X2 AND2X2_2638 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n730), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n729), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n731) );
  AND2X2 AND2X2_2639 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n731), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n732) );
  AND2X2 AND2X2_264 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n409_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n407_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_tras_cntr_3__FF_INPUT) );
  AND2X2 AND2X2_2640 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n734), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf5), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n735) );
  AND2X2 AND2X2_2641 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n735), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n733), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n736) );
  AND2X2 AND2X2_2642 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n739), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n738), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n740) );
  AND2X2 AND2X2_2643 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n740), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf5), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n741) );
  AND2X2 AND2X2_2644 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n743), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf4), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n744) );
  AND2X2 AND2X2_2645 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n744), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n742), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n745) );
  AND2X2 AND2X2_2646 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n748), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n747), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n749) );
  AND2X2 AND2X2_2647 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n749), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf4), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n750) );
  AND2X2 AND2X2_2648 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n752), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf3), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n753) );
  AND2X2 AND2X2_2649 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n753), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n751), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n754) );
  AND2X2 AND2X2_265 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n415_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n413_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n416) );
  AND2X2 AND2X2_2650 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n757), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n756), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n758) );
  AND2X2 AND2X2_2651 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n758), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf3), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n759) );
  AND2X2 AND2X2_2652 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n761), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf2), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n762) );
  AND2X2 AND2X2_2653 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n762), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n760), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n763) );
  AND2X2 AND2X2_2654 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n766), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n765), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n767) );
  AND2X2 AND2X2_2655 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n767), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf2), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n768) );
  AND2X2 AND2X2_2656 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n770), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n771) );
  AND2X2 AND2X2_2657 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n771), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n769), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n772) );
  AND2X2 AND2X2_2658 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n775), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n774), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n776) );
  AND2X2 AND2X2_2659 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n776), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n777) );
  AND2X2 AND2X2_266 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n417_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n418), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n419_1) );
  AND2X2 AND2X2_2660 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n779), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n780) );
  AND2X2 AND2X2_2661 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n780), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n778), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n781) );
  AND2X2 AND2X2_2662 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n784), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n783), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n785) );
  AND2X2 AND2X2_2663 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n785), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n786) );
  AND2X2 AND2X2_2664 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n788), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf5), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n789) );
  AND2X2 AND2X2_2665 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n789), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n787), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n790) );
  AND2X2 AND2X2_2666 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n793), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n792), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n794) );
  AND2X2 AND2X2_2667 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n794), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf5), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n795) );
  AND2X2 AND2X2_2668 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n797), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf4), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n798) );
  AND2X2 AND2X2_2669 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n798), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n796), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n799) );
  AND2X2 AND2X2_267 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n421), .B(sdram_resetn_bF_buf27), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n422) );
  AND2X2 AND2X2_2670 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n802), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n801), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n803) );
  AND2X2 AND2X2_2671 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n803), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf4), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n804) );
  AND2X2 AND2X2_2672 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n806), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf3), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n807) );
  AND2X2 AND2X2_2673 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n807), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n805), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n808) );
  AND2X2 AND2X2_2674 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n811), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n810), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n812) );
  AND2X2 AND2X2_2675 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n812), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf3), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n813) );
  AND2X2 AND2X2_2676 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n815), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf2), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n816) );
  AND2X2 AND2X2_2677 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n816), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n814), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n817) );
  AND2X2 AND2X2_2678 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n820), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n819), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n821) );
  AND2X2 AND2X2_2679 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n821), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf2), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n822) );
  AND2X2 AND2X2_268 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n420_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n422), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_timer0_0__FF_INPUT) );
  AND2X2 AND2X2_2680 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n824), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n825) );
  AND2X2 AND2X2_2681 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n825), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n823), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n826) );
  AND2X2 AND2X2_2682 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n829), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n828), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n830) );
  AND2X2 AND2X2_2683 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n830), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n831) );
  AND2X2 AND2X2_2684 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n833), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n834) );
  AND2X2 AND2X2_2685 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n834), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n832), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n835) );
  AND2X2 AND2X2_2686 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n838), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n837), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n839) );
  AND2X2 AND2X2_2687 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n839), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n840) );
  AND2X2 AND2X2_2688 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n842), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf5), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n843) );
  AND2X2 AND2X2_2689 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n843), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n841), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n844) );
  AND2X2 AND2X2_269 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_timer0_1_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_timer0_0_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n426) );
  AND2X2 AND2X2_2690 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n847), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n846), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n848) );
  AND2X2 AND2X2_2691 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n848), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf5), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n849) );
  AND2X2 AND2X2_2692 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n851), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf4), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n852) );
  AND2X2 AND2X2_2693 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n852), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n850), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n853) );
  AND2X2 AND2X2_2694 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n856), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n855), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n857) );
  AND2X2 AND2X2_2695 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n857), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf4), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n858) );
  AND2X2 AND2X2_2696 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n860), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf3), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n861) );
  AND2X2 AND2X2_2697 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n861), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n859), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n862) );
  AND2X2 AND2X2_2698 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n865), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n864), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n866) );
  AND2X2 AND2X2_2699 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n866), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf3), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n867) );
  AND2X2 AND2X2_27 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n254_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n256_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n257) );
  AND2X2 AND2X2_270 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n383_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n428_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n429) );
  AND2X2 AND2X2_2700 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n869), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf2), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n870) );
  AND2X2 AND2X2_2701 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n870), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n868), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n871) );
  AND2X2 AND2X2_2702 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n874), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n873), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n875) );
  AND2X2 AND2X2_2703 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n875), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf2), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n876) );
  AND2X2 AND2X2_2704 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n878), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n879) );
  AND2X2 AND2X2_2705 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n879), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n877), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n880) );
  AND2X2 AND2X2_2706 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n883), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n882), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n884) );
  AND2X2 AND2X2_2707 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n884), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n885) );
  AND2X2 AND2X2_2708 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n887), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n888) );
  AND2X2 AND2X2_2709 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n888), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n886), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n889) );
  AND2X2 AND2X2_271 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n429), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n427_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n430) );
  AND2X2 AND2X2_2710 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n892), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n891), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n893) );
  AND2X2 AND2X2_2711 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n893), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n894) );
  AND2X2 AND2X2_2712 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n896), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf5), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n897) );
  AND2X2 AND2X2_2713 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n897), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n895), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n898) );
  AND2X2 AND2X2_2714 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n901), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n900), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n902) );
  AND2X2 AND2X2_2715 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n902), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf5), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n903) );
  AND2X2 AND2X2_2716 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n905), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf4), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n906) );
  AND2X2 AND2X2_2717 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n906), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n904), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n907) );
  AND2X2 AND2X2_2718 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n910), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n909), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n911) );
  AND2X2 AND2X2_2719 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n911), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf4), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n912) );
  AND2X2 AND2X2_272 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n381), .B(\cfg_sdr_trcd_d[1] ), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n431_1) );
  AND2X2 AND2X2_2720 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n914), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf3), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n915) );
  AND2X2 AND2X2_2721 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n915), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n913), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n916) );
  AND2X2 AND2X2_2722 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n919), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n918), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n920) );
  AND2X2 AND2X2_2723 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n920), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf3), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n921) );
  AND2X2 AND2X2_2724 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n923), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf2), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n924) );
  AND2X2 AND2X2_2725 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n924), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n922), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n925) );
  AND2X2 AND2X2_2726 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n928), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n927), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n929) );
  AND2X2 AND2X2_2727 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n929), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf2), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n930) );
  AND2X2 AND2X2_2728 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n932), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n933) );
  AND2X2 AND2X2_2729 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n933), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n931), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n934) );
  AND2X2 AND2X2_273 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n434_1), .B(sdram_resetn_bF_buf26), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n435_1) );
  AND2X2 AND2X2_2730 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n937), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n936), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n938) );
  AND2X2 AND2X2_2731 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n938), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n939) );
  AND2X2 AND2X2_2732 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n941), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n942) );
  AND2X2 AND2X2_2733 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n942), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n940), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n943) );
  AND2X2 AND2X2_2734 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n946), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n945), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n947) );
  AND2X2 AND2X2_2735 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n947), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n948) );
  AND2X2 AND2X2_2736 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n950), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf5), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n951) );
  AND2X2 AND2X2_2737 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n951), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n949), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n952) );
  AND2X2 AND2X2_2738 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n955), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n954), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n956) );
  AND2X2 AND2X2_2739 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n956), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf5), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n957) );
  AND2X2 AND2X2_274 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n433), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n435_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_timer0_1__FF_INPUT) );
  AND2X2 AND2X2_2740 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n959), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf4), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n960) );
  AND2X2 AND2X2_2741 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n960), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n958), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n961) );
  AND2X2 AND2X2_2742 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n964), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n963), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n965) );
  AND2X2 AND2X2_2743 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n965), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf4), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n966) );
  AND2X2 AND2X2_2744 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n968), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf3), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n969) );
  AND2X2 AND2X2_2745 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n969), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n967), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n970) );
  AND2X2 AND2X2_2746 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n973), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n972), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n974) );
  AND2X2 AND2X2_2747 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n974), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf3), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n975) );
  AND2X2 AND2X2_2748 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n977), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf2), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n978) );
  AND2X2 AND2X2_2749 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n978), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n976), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n979) );
  AND2X2 AND2X2_275 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n424), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_timer0_2_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n439_1) );
  AND2X2 AND2X2_2750 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n634), .B(u_wb2sdrc_cmdfifo_wr), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n981) );
  AND2X2 AND2X2_2751 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_3__0_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n983) );
  AND2X2 AND2X2_2752 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf4), .B(\wb_addr_i[0] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n984) );
  AND2X2 AND2X2_2753 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_3__1_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n986) );
  AND2X2 AND2X2_2754 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf3), .B(\wb_addr_i[1] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n987) );
  AND2X2 AND2X2_2755 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_3__2_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n989) );
  AND2X2 AND2X2_2756 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf2), .B(\wb_addr_i[2] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n990) );
  AND2X2 AND2X2_2757 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_3__3_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n992) );
  AND2X2 AND2X2_2758 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf1), .B(\wb_addr_i[3] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n993) );
  AND2X2 AND2X2_2759 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_3__4_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n995) );
  AND2X2 AND2X2_276 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n429), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n440_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n441) );
  AND2X2 AND2X2_2760 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf0), .B(\wb_addr_i[4] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n996) );
  AND2X2 AND2X2_2761 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_3__5_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n998) );
  AND2X2 AND2X2_2762 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf5), .B(\wb_addr_i[5] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n999) );
  AND2X2 AND2X2_2763 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_3__6_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1001) );
  AND2X2 AND2X2_2764 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf4), .B(\wb_addr_i[6] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1002) );
  AND2X2 AND2X2_2765 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_3__7_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1004) );
  AND2X2 AND2X2_2766 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf3), .B(\wb_addr_i[7] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1005) );
  AND2X2 AND2X2_2767 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_3__8_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1007) );
  AND2X2 AND2X2_2768 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf2), .B(\wb_addr_i[8] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1008) );
  AND2X2 AND2X2_2769 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_3__9_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1010) );
  AND2X2 AND2X2_277 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n381), .B(\cfg_sdr_trcd_d[2] ), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n442) );
  AND2X2 AND2X2_2770 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf1), .B(\wb_addr_i[9] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1011) );
  AND2X2 AND2X2_2771 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_3__10_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1013) );
  AND2X2 AND2X2_2772 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf0), .B(\wb_addr_i[10] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1014) );
  AND2X2 AND2X2_2773 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_3__11_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1016) );
  AND2X2 AND2X2_2774 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf5), .B(\wb_addr_i[11] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1017) );
  AND2X2 AND2X2_2775 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_3__12_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1019) );
  AND2X2 AND2X2_2776 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf4), .B(\wb_addr_i[12] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1020) );
  AND2X2 AND2X2_2777 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_3__13_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1022) );
  AND2X2 AND2X2_2778 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf3), .B(\wb_addr_i[13] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1023) );
  AND2X2 AND2X2_2779 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_3__14_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1025) );
  AND2X2 AND2X2_278 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n445_1), .B(sdram_resetn_bF_buf25), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n446_1) );
  AND2X2 AND2X2_2780 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf2), .B(\wb_addr_i[14] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1026) );
  AND2X2 AND2X2_2781 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_3__15_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1028) );
  AND2X2 AND2X2_2782 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf1), .B(\wb_addr_i[15] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1029) );
  AND2X2 AND2X2_2783 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_3__16_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1031) );
  AND2X2 AND2X2_2784 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf0), .B(\wb_addr_i[16] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1032) );
  AND2X2 AND2X2_2785 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_3__17_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1034) );
  AND2X2 AND2X2_2786 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf5), .B(\wb_addr_i[17] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1035) );
  AND2X2 AND2X2_2787 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_3__18_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1037) );
  AND2X2 AND2X2_2788 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf4), .B(\wb_addr_i[18] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1038) );
  AND2X2 AND2X2_2789 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_3__19_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1040) );
  AND2X2 AND2X2_279 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n444_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n446_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_timer0_2__FF_INPUT) );
  AND2X2 AND2X2_2790 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf3), .B(\wb_addr_i[19] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1041) );
  AND2X2 AND2X2_2791 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_3__20_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1043) );
  AND2X2 AND2X2_2792 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf2), .B(\wb_addr_i[20] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1044) );
  AND2X2 AND2X2_2793 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_3__21_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1046) );
  AND2X2 AND2X2_2794 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf1), .B(\wb_addr_i[21] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1047) );
  AND2X2 AND2X2_2795 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_3__22_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1049) );
  AND2X2 AND2X2_2796 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf0), .B(\wb_addr_i[22] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1050) );
  AND2X2 AND2X2_2797 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_3__23_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1052) );
  AND2X2 AND2X2_2798 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf5), .B(\wb_addr_i[23] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1053) );
  AND2X2 AND2X2_2799 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_3__24_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1055) );
  AND2X2 AND2X2_28 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n258_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n260_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n261_1) );
  AND2X2 AND2X2_280 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n437_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_timer0_3_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n448_1) );
  AND2X2 AND2X2_2800 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf4), .B(\wb_addr_i[24] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1056) );
  AND2X2 AND2X2_2801 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_3__25_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1058) );
  AND2X2 AND2X2_2802 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf3), .B(\wb_addr_i[25] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1059) );
  AND2X2 AND2X2_2803 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_3__26_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1061) );
  AND2X2 AND2X2_2804 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_wr_data_26_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1062) );
  AND2X2 AND2X2_2805 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_3__27_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1064) );
  AND2X2 AND2X2_2806 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf1), .B(1'b1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1065) );
  AND2X2 AND2X2_2807 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_3__28_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1067) );
  AND2X2 AND2X2_2808 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf0), .B(1'b0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1068) );
  AND2X2 AND2X2_2809 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_3__29_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1070) );
  AND2X2 AND2X2_281 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n449_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n450), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n451) );
  AND2X2 AND2X2_2810 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf5), .B(1'b0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1071) );
  AND2X2 AND2X2_2811 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_3__30_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1073) );
  AND2X2 AND2X2_2812 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf4), .B(1'b0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1074) );
  AND2X2 AND2X2_2813 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_3__31_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1076) );
  AND2X2 AND2X2_2814 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf3), .B(1'b0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1077) );
  AND2X2 AND2X2_2815 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_3__32_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1079) );
  AND2X2 AND2X2_2816 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf2), .B(1'b0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1080) );
  AND2X2 AND2X2_2817 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_3__33_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1082) );
  AND2X2 AND2X2_2818 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf1), .B(1'b0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1083) );
  AND2X2 AND2X2_2819 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_3__34_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1085) );
  AND2X2 AND2X2_282 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n453_1), .B(sdram_resetn_bF_buf24), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n454) );
  AND2X2 AND2X2_2820 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf0), .B(1'b0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1086) );
  AND2X2 AND2X2_2821 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_3__35_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1088) );
  AND2X2 AND2X2_2822 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf5), .B(1'b0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1089) );
  AND2X2 AND2X2_2823 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1093), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1091), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n494) );
  AND2X2 AND2X2_2824 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1096), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1095), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n495) );
  AND2X2 AND2X2_2825 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1099), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1098), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n496) );
  AND2X2 AND2X2_2826 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1102), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1101), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n497) );
  AND2X2 AND2X2_2827 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1105), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1104), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n498) );
  AND2X2 AND2X2_2828 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1108), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1107), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n499) );
  AND2X2 AND2X2_2829 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1111), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1110), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n500) );
  AND2X2 AND2X2_283 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n452), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n454), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_timer0_3__FF_INPUT) );
  AND2X2 AND2X2_2830 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1114), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1113), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n501) );
  AND2X2 AND2X2_2831 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1117), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1116), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n502) );
  AND2X2 AND2X2_2832 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1120), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1119), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n503) );
  AND2X2 AND2X2_2833 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1123), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1122), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n504) );
  AND2X2 AND2X2_2834 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1126), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1125), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n505) );
  AND2X2 AND2X2_2835 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1129), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1128), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n506) );
  AND2X2 AND2X2_2836 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1132), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1131), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n507) );
  AND2X2 AND2X2_2837 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1135), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1134), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n508) );
  AND2X2 AND2X2_2838 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1138), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1137), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n509) );
  AND2X2 AND2X2_2839 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1141), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1140), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n510) );
  AND2X2 AND2X2_284 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n253_1), .B(u_sdrc_core_r2b_len_0_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n473) );
  AND2X2 AND2X2_2840 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1144), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1143), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n511) );
  AND2X2 AND2X2_2841 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1147), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1146), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n512) );
  AND2X2 AND2X2_2842 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1150), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1149), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n513) );
  AND2X2 AND2X2_2843 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1153), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1152), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n514) );
  AND2X2 AND2X2_2844 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1156), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1155), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n515) );
  AND2X2 AND2X2_2845 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1159), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1158), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n516) );
  AND2X2 AND2X2_2846 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1162), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1161), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n517) );
  AND2X2 AND2X2_2847 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1165), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1164), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n518) );
  AND2X2 AND2X2_2848 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1168), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1167), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n519) );
  AND2X2 AND2X2_2849 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1171), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1170), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n520) );
  AND2X2 AND2X2_285 ( .A(sdram_resetn_bF_buf23), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_0_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n474) );
  AND2X2 AND2X2_2850 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1174), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1173), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n521) );
  AND2X2 AND2X2_2851 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1177), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1176), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n522) );
  AND2X2 AND2X2_2852 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1180), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1179), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n523) );
  AND2X2 AND2X2_2853 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1183), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1182), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n524) );
  AND2X2 AND2X2_2854 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1186), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1185), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n525) );
  AND2X2 AND2X2_2855 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1189), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1188), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n526) );
  AND2X2 AND2X2_2856 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1192), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1191), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n527) );
  AND2X2 AND2X2_2857 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1195), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1194), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n528) );
  AND2X2 AND2X2_2858 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1198), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1197), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n529) );
  AND2X2 AND2X2_2859 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1202), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1200), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n532) );
  AND2X2 AND2X2_286 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf5), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n474), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n475) );
  AND2X2 AND2X2_2860 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1205), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1204), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n534) );
  AND2X2 AND2X2_2861 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1208), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1207), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n536) );
  AND2X2 AND2X2_2862 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1211), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1210), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n538) );
  AND2X2 AND2X2_2863 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1214), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1213), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n540) );
  AND2X2 AND2X2_2864 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1217), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1216), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n542) );
  AND2X2 AND2X2_2865 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1220), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1219), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n544) );
  AND2X2 AND2X2_2866 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1223), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1222), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n546) );
  AND2X2 AND2X2_2867 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1226), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1225), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n548) );
  AND2X2 AND2X2_2868 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1229), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1228), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n550) );
  AND2X2 AND2X2_2869 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1232), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1231), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n552) );
  AND2X2 AND2X2_287 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n253_1), .B(u_sdrc_core_r2b_len_1_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n477) );
  AND2X2 AND2X2_2870 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1235), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1234), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n554) );
  AND2X2 AND2X2_2871 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1238), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1237), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n556) );
  AND2X2 AND2X2_2872 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1241), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1240), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n558) );
  AND2X2 AND2X2_2873 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1244), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1243), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n560) );
  AND2X2 AND2X2_2874 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1247), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1246), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n562) );
  AND2X2 AND2X2_2875 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1250), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1249), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n564) );
  AND2X2 AND2X2_2876 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1253), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1252), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n566) );
  AND2X2 AND2X2_2877 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1256), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1255), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n568) );
  AND2X2 AND2X2_2878 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1259), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1258), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n570) );
  AND2X2 AND2X2_2879 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1262), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1261), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n572) );
  AND2X2 AND2X2_288 ( .A(sdram_resetn_bF_buf22), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_1_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n478) );
  AND2X2 AND2X2_2880 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1265), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1264), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n574) );
  AND2X2 AND2X2_2881 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1268), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1267), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n576) );
  AND2X2 AND2X2_2882 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1271), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1270), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n578) );
  AND2X2 AND2X2_2883 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1274), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1273), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n580) );
  AND2X2 AND2X2_2884 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1277), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1276), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n582) );
  AND2X2 AND2X2_2885 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1280), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1279), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n584) );
  AND2X2 AND2X2_2886 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1283), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1282), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n586) );
  AND2X2 AND2X2_2887 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1286), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1285), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n588) );
  AND2X2 AND2X2_2888 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1289), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1288), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n590) );
  AND2X2 AND2X2_2889 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1292), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1291), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n592) );
  AND2X2 AND2X2_289 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n478), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n479) );
  AND2X2 AND2X2_2890 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1295), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1294), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n594) );
  AND2X2 AND2X2_2891 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1298), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1297), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n596) );
  AND2X2 AND2X2_2892 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1301), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1300), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n598) );
  AND2X2 AND2X2_2893 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1304), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1303), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n600) );
  AND2X2 AND2X2_2894 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1307), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1306), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n602) );
  AND2X2 AND2X2_2895 ( .A(u_wb2sdrc_u_rddatafifo_sync_wr_ptr_1_1_), .B(u_wb2sdrc_u_rddatafifo_sync_wr_ptr_2_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n411_1) );
  AND2X2 AND2X2_2896 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n412_1), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n410), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n413) );
  AND2X2 AND2X2_2897 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n413), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf4), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n414) );
  AND2X2 AND2X2_2898 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n415_1), .B(u_wb2sdrc_u_rddatafifo_rd_ptr_1_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n416_1) );
  AND2X2 AND2X2_2899 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n415_1), .B(u_wb2sdrc_u_rddatafifo_sync_wr_ptr_1_0_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n420_1) );
  AND2X2 AND2X2_29 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n262), .B(sdram_resetn_bF_buf48), .Y(u_sdrc_core_u_bank_ctl_rank_cnt_1__FF_INPUT) );
  AND2X2 AND2X2_290 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n253_1), .B(u_sdrc_core_r2b_len_2_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n481) );
  AND2X2 AND2X2_2900 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n413), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n421), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n422) );
  AND2X2 AND2X2_2901 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n424_1), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n418), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n425) );
  AND2X2 AND2X2_2902 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n427_1), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n429), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n430) );
  AND2X2 AND2X2_2903 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n423_1), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf4), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n431_1) );
  AND2X2 AND2X2_2904 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n432_1), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n430), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n433) );
  AND2X2 AND2X2_2905 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n433), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n425), .Y(u_wb2sdrc_rddatafifo_empty) );
  AND2X2 AND2X2_2906 ( .A(u_wb2sdrc_u_rddatafifo_wr_ptr_1_), .B(u_wb2sdrc_u_rddatafifo_wr_ptr_0_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n446) );
  AND2X2 AND2X2_2907 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n446), .B(app_rd_valid), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1) );
  AND2X2 AND2X2_2908 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf4), .B(app_rd_data_0_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n448) );
  AND2X2 AND2X2_2909 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_3__0_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n450_1) );
  AND2X2 AND2X2_291 ( .A(sdram_resetn_bF_buf21), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_2_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n482) );
  AND2X2 AND2X2_2910 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf2), .B(app_rd_data_1_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n452_1) );
  AND2X2 AND2X2_2911 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_3__1_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n453_1) );
  AND2X2 AND2X2_2912 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf1), .B(app_rd_data_2_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n455_1) );
  AND2X2 AND2X2_2913 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_3__2_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n456_1) );
  AND2X2 AND2X2_2914 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf0), .B(app_rd_data_3_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n458_1) );
  AND2X2 AND2X2_2915 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_3__3_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n459_1) );
  AND2X2 AND2X2_2916 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf4), .B(app_rd_data_4_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n461_1) );
  AND2X2 AND2X2_2917 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_3__4_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n462_1) );
  AND2X2 AND2X2_2918 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf3), .B(app_rd_data_5_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n464_1) );
  AND2X2 AND2X2_2919 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_3__5_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n465_1) );
  AND2X2 AND2X2_292 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n482), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n483) );
  AND2X2 AND2X2_2920 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf2), .B(app_rd_data_6_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n467_1) );
  AND2X2 AND2X2_2921 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_3__6_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n468_1) );
  AND2X2 AND2X2_2922 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf1), .B(app_rd_data_7_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n470_1) );
  AND2X2 AND2X2_2923 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_3__7_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n471_1) );
  AND2X2 AND2X2_2924 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf0), .B(app_rd_data_8_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n473_1) );
  AND2X2 AND2X2_2925 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_3__8_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n474_1) );
  AND2X2 AND2X2_2926 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf4), .B(app_rd_data_9_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n476_1) );
  AND2X2 AND2X2_2927 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_3__9_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n477_1) );
  AND2X2 AND2X2_2928 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf3), .B(app_rd_data_10_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n479_1) );
  AND2X2 AND2X2_2929 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_3__10_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n480_1) );
  AND2X2 AND2X2_293 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n253_1), .B(u_sdrc_core_r2b_len_3_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n485) );
  AND2X2 AND2X2_2930 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf2), .B(app_rd_data_11_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n482_1) );
  AND2X2 AND2X2_2931 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_3__11_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n483_1) );
  AND2X2 AND2X2_2932 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf1), .B(app_rd_data_12_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n485) );
  AND2X2 AND2X2_2933 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_3__12_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n486_1) );
  AND2X2 AND2X2_2934 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf0), .B(app_rd_data_13_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n488) );
  AND2X2 AND2X2_2935 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_3__13_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n489_1) );
  AND2X2 AND2X2_2936 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf4), .B(app_rd_data_14_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n491) );
  AND2X2 AND2X2_2937 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_3__14_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n492) );
  AND2X2 AND2X2_2938 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf3), .B(app_rd_data_15_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n494) );
  AND2X2 AND2X2_2939 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_3__15_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n495_1) );
  AND2X2 AND2X2_294 ( .A(sdram_resetn_bF_buf20), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_3_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n486) );
  AND2X2 AND2X2_2940 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf2), .B(app_rd_data_16_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n497) );
  AND2X2 AND2X2_2941 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_3__16_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n498) );
  AND2X2 AND2X2_2942 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf1), .B(app_rd_data_17_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n500_1) );
  AND2X2 AND2X2_2943 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_3__17_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n501_1) );
  AND2X2 AND2X2_2944 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf0), .B(app_rd_data_18_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n503_1) );
  AND2X2 AND2X2_2945 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_3__18_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n504) );
  AND2X2 AND2X2_2946 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf4), .B(app_rd_data_19_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n506) );
  AND2X2 AND2X2_2947 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_3__19_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n507) );
  AND2X2 AND2X2_2948 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf3), .B(app_rd_data_20_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n509_1) );
  AND2X2 AND2X2_2949 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_3__20_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n510_1) );
  AND2X2 AND2X2_295 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n486), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n487) );
  AND2X2 AND2X2_2950 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf2), .B(app_rd_data_21_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n512) );
  AND2X2 AND2X2_2951 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_3__21_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n513) );
  AND2X2 AND2X2_2952 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf1), .B(app_rd_data_22_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n515) );
  AND2X2 AND2X2_2953 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_3__22_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n516) );
  AND2X2 AND2X2_2954 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf0), .B(app_rd_data_23_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n518) );
  AND2X2 AND2X2_2955 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_3__23_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n519) );
  AND2X2 AND2X2_2956 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf4), .B(app_rd_data_24_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n521_1) );
  AND2X2 AND2X2_2957 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_3__24_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n522_1) );
  AND2X2 AND2X2_2958 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf3), .B(app_rd_data_25_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n524_1) );
  AND2X2 AND2X2_2959 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_3__25_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n525) );
  AND2X2 AND2X2_296 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n253_1), .B(u_sdrc_core_r2b_len_4_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n489) );
  AND2X2 AND2X2_2960 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf2), .B(app_rd_data_26_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n527_1) );
  AND2X2 AND2X2_2961 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_3__26_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n528) );
  AND2X2 AND2X2_2962 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf1), .B(app_rd_data_27_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n530) );
  AND2X2 AND2X2_2963 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_3__27_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n531) );
  AND2X2 AND2X2_2964 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf0), .B(app_rd_data_28_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n533) );
  AND2X2 AND2X2_2965 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_3__28_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n534) );
  AND2X2 AND2X2_2966 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf4), .B(app_rd_data_29_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n536) );
  AND2X2 AND2X2_2967 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_3__29_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n537) );
  AND2X2 AND2X2_2968 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf3), .B(app_rd_data_30_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n539) );
  AND2X2 AND2X2_2969 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_3__30_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n540) );
  AND2X2 AND2X2_297 ( .A(sdram_resetn_bF_buf19), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_4_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n490) );
  AND2X2 AND2X2_2970 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf2), .B(app_rd_data_31_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n542) );
  AND2X2 AND2X2_2971 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_3__31_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n543) );
  AND2X2 AND2X2_2972 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n375_1), .B(app_rd_valid), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n548) );
  AND2X2 AND2X2_2973 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n548), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n384_1), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n549) );
  AND2X2 AND2X2_2974 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n552), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n550), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n197) );
  AND2X2 AND2X2_2975 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n555), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n554), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n199) );
  AND2X2 AND2X2_2976 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n558), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n557), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n201) );
  AND2X2 AND2X2_2977 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n561), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n560), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n203) );
  AND2X2 AND2X2_2978 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n564), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n563), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n205) );
  AND2X2 AND2X2_2979 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n567), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n566), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n207) );
  AND2X2 AND2X2_298 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n490), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n491) );
  AND2X2 AND2X2_2980 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n570), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n569), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n209) );
  AND2X2 AND2X2_2981 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n573), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n572), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n211) );
  AND2X2 AND2X2_2982 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n576), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n575), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n213) );
  AND2X2 AND2X2_2983 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n579), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n578), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n215) );
  AND2X2 AND2X2_2984 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n582), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n581), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n217) );
  AND2X2 AND2X2_2985 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n585), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n584), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n219) );
  AND2X2 AND2X2_2986 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n588), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n587), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n221) );
  AND2X2 AND2X2_2987 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n591), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n590), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n223) );
  AND2X2 AND2X2_2988 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n594), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n593), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n225) );
  AND2X2 AND2X2_2989 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n597), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n596), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n227) );
  AND2X2 AND2X2_299 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n253_1), .B(u_sdrc_core_r2b_len_5_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n493) );
  AND2X2 AND2X2_2990 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n600), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n599), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n229) );
  AND2X2 AND2X2_2991 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n603), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n602), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n231) );
  AND2X2 AND2X2_2992 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n606), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n605), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n233) );
  AND2X2 AND2X2_2993 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n609), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n608), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n235) );
  AND2X2 AND2X2_2994 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n612), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n611), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n237) );
  AND2X2 AND2X2_2995 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n615), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n614), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n239) );
  AND2X2 AND2X2_2996 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n618), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n617), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n241) );
  AND2X2 AND2X2_2997 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n621), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n620), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n243) );
  AND2X2 AND2X2_2998 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n624), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n623), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n245) );
  AND2X2 AND2X2_2999 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n627), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n626), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n247) );
  AND2X2 AND2X2_3 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n204_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n205_1), .Y(u_sdrc_core_b2x_tras_ok) );
  AND2X2 AND2X2_30 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n242_1), .B(u_sdrc_core_u_bank_ctl_rank_cnt_2_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n266_1) );
  AND2X2 AND2X2_300 ( .A(sdram_resetn_bF_buf18), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_5_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n494) );
  AND2X2 AND2X2_3000 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n630), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n629), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n249) );
  AND2X2 AND2X2_3001 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n633), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n632), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n251) );
  AND2X2 AND2X2_3002 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n636), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n635), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n253) );
  AND2X2 AND2X2_3003 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n639), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n638), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n255) );
  AND2X2 AND2X2_3004 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n642), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n641), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n257) );
  AND2X2 AND2X2_3005 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n645), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n644), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n259) );
  AND2X2 AND2X2_3006 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n548), .B(u_wb2sdrc_u_rddatafifo_wr_ptr_1_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n650) );
  AND2X2 AND2X2_3007 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n653), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n651), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n264) );
  AND2X2 AND2X2_3008 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n656), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n655), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n266) );
  AND2X2 AND2X2_3009 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n659), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n658), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n268) );
  AND2X2 AND2X2_301 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n494), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n495) );
  AND2X2 AND2X2_3010 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n662), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n661), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n270) );
  AND2X2 AND2X2_3011 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n665), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n664), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n272) );
  AND2X2 AND2X2_3012 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n668), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n667), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n274) );
  AND2X2 AND2X2_3013 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n671), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n670), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n276) );
  AND2X2 AND2X2_3014 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n674), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n673), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n278) );
  AND2X2 AND2X2_3015 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n677), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n676), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n280) );
  AND2X2 AND2X2_3016 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n680), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n679), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n282) );
  AND2X2 AND2X2_3017 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n683), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n682), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n284) );
  AND2X2 AND2X2_3018 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n686), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n685), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n286) );
  AND2X2 AND2X2_3019 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n689), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n688), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n288) );
  AND2X2 AND2X2_302 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n253_1), .B(u_sdrc_core_r2b_len_6_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n497) );
  AND2X2 AND2X2_3020 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n692), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n691), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n290) );
  AND2X2 AND2X2_3021 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n695), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n694), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n292) );
  AND2X2 AND2X2_3022 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n698), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n697), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n294) );
  AND2X2 AND2X2_3023 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n701), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n700), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n296) );
  AND2X2 AND2X2_3024 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n704), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n703), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n298) );
  AND2X2 AND2X2_3025 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n707), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n706), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n300) );
  AND2X2 AND2X2_3026 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n710), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n709), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n302) );
  AND2X2 AND2X2_3027 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n713), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n712), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n304) );
  AND2X2 AND2X2_3028 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n716), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n715), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n306) );
  AND2X2 AND2X2_3029 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n719), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n718), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n308) );
  AND2X2 AND2X2_303 ( .A(sdram_resetn_bF_buf17), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_6_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n498) );
  AND2X2 AND2X2_3030 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n722), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n721), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n310) );
  AND2X2 AND2X2_3031 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n725), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n724), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n312) );
  AND2X2 AND2X2_3032 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n728), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n727), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n314) );
  AND2X2 AND2X2_3033 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n731), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n730), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n316) );
  AND2X2 AND2X2_3034 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n734), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n733), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n318) );
  AND2X2 AND2X2_3035 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n737), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n736), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n320) );
  AND2X2 AND2X2_3036 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n740), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n739), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n322) );
  AND2X2 AND2X2_3037 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n743), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n742), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n324) );
  AND2X2 AND2X2_3038 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n746), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n745), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n326) );
  AND2X2 AND2X2_3039 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_0__0_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n751) );
  AND2X2 AND2X2_304 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf5), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n498), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n499) );
  AND2X2 AND2X2_3040 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_1__0_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n752) );
  AND2X2 AND2X2_3041 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n753), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf3), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n754) );
  AND2X2 AND2X2_3042 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_1_), .B(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf3), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n755) );
  AND2X2 AND2X2_3043 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_3__0_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n756) );
  AND2X2 AND2X2_3044 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_rd_ptr_1_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n757) );
  AND2X2 AND2X2_3045 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_2__0_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n758) );
  AND2X2 AND2X2_3046 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_0__1_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n761) );
  AND2X2 AND2X2_3047 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_1__1_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n762) );
  AND2X2 AND2X2_3048 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n763), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf2), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n764) );
  AND2X2 AND2X2_3049 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_3__1_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n765) );
  AND2X2 AND2X2_305 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_0_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n501) );
  AND2X2 AND2X2_3050 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_2__1_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n766) );
  AND2X2 AND2X2_3051 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_0__2_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n769) );
  AND2X2 AND2X2_3052 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_1__2_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n770) );
  AND2X2 AND2X2_3053 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n771), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf1), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n772) );
  AND2X2 AND2X2_3054 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_3__2_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n773) );
  AND2X2 AND2X2_3055 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_2__2_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n774) );
  AND2X2 AND2X2_3056 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf5), .B(u_wb2sdrc_u_rddatafifo_mem_0__3_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n777) );
  AND2X2 AND2X2_3057 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_1__3_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n778) );
  AND2X2 AND2X2_3058 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n779), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf0), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n780) );
  AND2X2 AND2X2_3059 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_3__3_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n781) );
  AND2X2 AND2X2_306 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf1), .B(u_sdrc_core_r2b_raddr_0_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n502) );
  AND2X2 AND2X2_3060 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_2__3_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n782) );
  AND2X2 AND2X2_3061 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_0__4_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n785) );
  AND2X2 AND2X2_3062 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf5), .B(u_wb2sdrc_u_rddatafifo_mem_1__4_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n786) );
  AND2X2 AND2X2_3063 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n787), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf4), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n788) );
  AND2X2 AND2X2_3064 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_3__4_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n789) );
  AND2X2 AND2X2_3065 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_2__4_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n790) );
  AND2X2 AND2X2_3066 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_0__5_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n793) );
  AND2X2 AND2X2_3067 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_1__5_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n794) );
  AND2X2 AND2X2_3068 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n795), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf3), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n796) );
  AND2X2 AND2X2_3069 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_3__5_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n797) );
  AND2X2 AND2X2_307 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n503), .B(sdram_resetn_bF_buf16), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_0__FF_INPUT) );
  AND2X2 AND2X2_3070 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_2__5_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n798) );
  AND2X2 AND2X2_3071 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_0__6_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n801) );
  AND2X2 AND2X2_3072 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_1__6_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n802) );
  AND2X2 AND2X2_3073 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n803), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf2), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n804) );
  AND2X2 AND2X2_3074 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_3__6_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n805) );
  AND2X2 AND2X2_3075 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_2__6_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n806) );
  AND2X2 AND2X2_3076 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_0__7_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n809) );
  AND2X2 AND2X2_3077 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_1__7_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n810) );
  AND2X2 AND2X2_3078 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n811), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf1), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n812) );
  AND2X2 AND2X2_3079 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_3__7_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n813) );
  AND2X2 AND2X2_308 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_1_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n505) );
  AND2X2 AND2X2_3080 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_2__7_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n814) );
  AND2X2 AND2X2_3081 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_0__8_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n817) );
  AND2X2 AND2X2_3082 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_1__8_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n818) );
  AND2X2 AND2X2_3083 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n819), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf0), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n820) );
  AND2X2 AND2X2_3084 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_3__8_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n821) );
  AND2X2 AND2X2_3085 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_2__8_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n822) );
  AND2X2 AND2X2_3086 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf5), .B(u_wb2sdrc_u_rddatafifo_mem_0__9_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n825) );
  AND2X2 AND2X2_3087 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_1__9_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n826) );
  AND2X2 AND2X2_3088 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n827), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf4), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n828) );
  AND2X2 AND2X2_3089 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_3__9_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n829) );
  AND2X2 AND2X2_309 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf0), .B(u_sdrc_core_r2b_raddr_1_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n506) );
  AND2X2 AND2X2_3090 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_2__9_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n830) );
  AND2X2 AND2X2_3091 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_0__10_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n833) );
  AND2X2 AND2X2_3092 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf5), .B(u_wb2sdrc_u_rddatafifo_mem_1__10_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n834) );
  AND2X2 AND2X2_3093 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n835), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf3), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n836) );
  AND2X2 AND2X2_3094 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_3__10_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n837) );
  AND2X2 AND2X2_3095 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_2__10_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n838) );
  AND2X2 AND2X2_3096 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_0__11_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n841) );
  AND2X2 AND2X2_3097 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_1__11_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n842) );
  AND2X2 AND2X2_3098 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n843), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf2), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n844) );
  AND2X2 AND2X2_3099 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_3__11_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n845) );
  AND2X2 AND2X2_31 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n265_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n266_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n267_1) );
  AND2X2 AND2X2_310 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n507), .B(sdram_resetn_bF_buf15), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_1__FF_INPUT) );
  AND2X2 AND2X2_3100 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_2__11_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n846) );
  AND2X2 AND2X2_3101 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_0__12_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n849) );
  AND2X2 AND2X2_3102 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_1__12_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n850) );
  AND2X2 AND2X2_3103 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n851), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf1), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n852) );
  AND2X2 AND2X2_3104 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_3__12_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n853) );
  AND2X2 AND2X2_3105 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_2__12_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n854) );
  AND2X2 AND2X2_3106 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_0__13_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n857) );
  AND2X2 AND2X2_3107 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_1__13_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n858) );
  AND2X2 AND2X2_3108 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n859), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf0), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n860) );
  AND2X2 AND2X2_3109 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_3__13_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n861) );
  AND2X2 AND2X2_311 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_2_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n509) );
  AND2X2 AND2X2_3110 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_2__13_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n862) );
  AND2X2 AND2X2_3111 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_0__14_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n865) );
  AND2X2 AND2X2_3112 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_1__14_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n866) );
  AND2X2 AND2X2_3113 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n867), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf4), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n868) );
  AND2X2 AND2X2_3114 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_3__14_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n869) );
  AND2X2 AND2X2_3115 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_2__14_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n870) );
  AND2X2 AND2X2_3116 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf5), .B(u_wb2sdrc_u_rddatafifo_mem_0__15_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n873) );
  AND2X2 AND2X2_3117 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_1__15_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n874) );
  AND2X2 AND2X2_3118 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n875), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf3), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n876) );
  AND2X2 AND2X2_3119 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_3__15_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n877) );
  AND2X2 AND2X2_312 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf4), .B(u_sdrc_core_r2b_raddr_2_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n510) );
  AND2X2 AND2X2_3120 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_2__15_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n878) );
  AND2X2 AND2X2_3121 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_0__16_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n881) );
  AND2X2 AND2X2_3122 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf5), .B(u_wb2sdrc_u_rddatafifo_mem_1__16_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n882) );
  AND2X2 AND2X2_3123 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n883), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf2), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n884) );
  AND2X2 AND2X2_3124 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_3__16_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n885) );
  AND2X2 AND2X2_3125 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_2__16_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n886) );
  AND2X2 AND2X2_3126 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_0__17_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n889) );
  AND2X2 AND2X2_3127 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_1__17_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n890) );
  AND2X2 AND2X2_3128 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n891), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf1), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n892) );
  AND2X2 AND2X2_3129 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_3__17_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n893) );
  AND2X2 AND2X2_313 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n511), .B(sdram_resetn_bF_buf14), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_2__FF_INPUT) );
  AND2X2 AND2X2_3130 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_2__17_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n894) );
  AND2X2 AND2X2_3131 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_0__18_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n897) );
  AND2X2 AND2X2_3132 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_1__18_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n898) );
  AND2X2 AND2X2_3133 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n899), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf0), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n900) );
  AND2X2 AND2X2_3134 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_3__18_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n901) );
  AND2X2 AND2X2_3135 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_2__18_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n902) );
  AND2X2 AND2X2_3136 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_0__19_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n905) );
  AND2X2 AND2X2_3137 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_1__19_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n906) );
  AND2X2 AND2X2_3138 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n907), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf4), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n908) );
  AND2X2 AND2X2_3139 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_3__19_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n909) );
  AND2X2 AND2X2_314 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_3_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n513) );
  AND2X2 AND2X2_3140 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_2__19_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n910) );
  AND2X2 AND2X2_3141 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_0__20_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n913) );
  AND2X2 AND2X2_3142 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_1__20_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n914) );
  AND2X2 AND2X2_3143 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n915), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf3), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n916) );
  AND2X2 AND2X2_3144 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_3__20_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n917) );
  AND2X2 AND2X2_3145 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_2__20_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n918) );
  AND2X2 AND2X2_3146 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf5), .B(u_wb2sdrc_u_rddatafifo_mem_0__21_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n921) );
  AND2X2 AND2X2_3147 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_1__21_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n922) );
  AND2X2 AND2X2_3148 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n923), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf2), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n924) );
  AND2X2 AND2X2_3149 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_3__21_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n925) );
  AND2X2 AND2X2_315 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf3), .B(u_sdrc_core_r2b_raddr_3_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n514) );
  AND2X2 AND2X2_3150 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_2__21_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n926) );
  AND2X2 AND2X2_3151 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_0__22_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n929) );
  AND2X2 AND2X2_3152 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf5), .B(u_wb2sdrc_u_rddatafifo_mem_1__22_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n930) );
  AND2X2 AND2X2_3153 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n931), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf1), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n932) );
  AND2X2 AND2X2_3154 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_3__22_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n933) );
  AND2X2 AND2X2_3155 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_2__22_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n934) );
  AND2X2 AND2X2_3156 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_0__23_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n937) );
  AND2X2 AND2X2_3157 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_1__23_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n938) );
  AND2X2 AND2X2_3158 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n939), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf0), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n940) );
  AND2X2 AND2X2_3159 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_3__23_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n941) );
  AND2X2 AND2X2_316 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n515), .B(sdram_resetn_bF_buf13), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_3__FF_INPUT) );
  AND2X2 AND2X2_3160 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_2__23_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n942) );
  AND2X2 AND2X2_3161 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_0__24_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n945) );
  AND2X2 AND2X2_3162 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_1__24_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n946) );
  AND2X2 AND2X2_3163 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n947), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf4), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n948) );
  AND2X2 AND2X2_3164 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_3__24_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n949) );
  AND2X2 AND2X2_3165 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_2__24_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n950) );
  AND2X2 AND2X2_3166 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_0__25_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n953) );
  AND2X2 AND2X2_3167 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_1__25_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n954) );
  AND2X2 AND2X2_3168 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n955), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf3), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n956) );
  AND2X2 AND2X2_3169 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_3__25_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n957) );
  AND2X2 AND2X2_317 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_4_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n517) );
  AND2X2 AND2X2_3170 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_2__25_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n958) );
  AND2X2 AND2X2_3171 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_0__26_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n961) );
  AND2X2 AND2X2_3172 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_1__26_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n962) );
  AND2X2 AND2X2_3173 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n963), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf2), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n964) );
  AND2X2 AND2X2_3174 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_3__26_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n965) );
  AND2X2 AND2X2_3175 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_2__26_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n966) );
  AND2X2 AND2X2_3176 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf5), .B(u_wb2sdrc_u_rddatafifo_mem_0__27_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n969) );
  AND2X2 AND2X2_3177 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_1__27_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n970) );
  AND2X2 AND2X2_3178 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n971), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf1), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n972) );
  AND2X2 AND2X2_3179 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_3__27_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n973) );
  AND2X2 AND2X2_318 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf2), .B(u_sdrc_core_r2b_raddr_4_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n518) );
  AND2X2 AND2X2_3180 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_2__27_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n974) );
  AND2X2 AND2X2_3181 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_0__28_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n977) );
  AND2X2 AND2X2_3182 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf5), .B(u_wb2sdrc_u_rddatafifo_mem_1__28_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n978) );
  AND2X2 AND2X2_3183 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n979), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf0), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n980) );
  AND2X2 AND2X2_3184 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_3__28_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n981) );
  AND2X2 AND2X2_3185 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_2__28_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n982) );
  AND2X2 AND2X2_3186 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_0__29_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n985) );
  AND2X2 AND2X2_3187 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_1__29_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n986) );
  AND2X2 AND2X2_3188 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n987), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf4), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n988) );
  AND2X2 AND2X2_3189 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_3__29_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n989) );
  AND2X2 AND2X2_319 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n519), .B(sdram_resetn_bF_buf12), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_4__FF_INPUT) );
  AND2X2 AND2X2_3190 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_2__29_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n990) );
  AND2X2 AND2X2_3191 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_0__30_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n993) );
  AND2X2 AND2X2_3192 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_1__30_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n994) );
  AND2X2 AND2X2_3193 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n995), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf3), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n996) );
  AND2X2 AND2X2_3194 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_3__30_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n997) );
  AND2X2 AND2X2_3195 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_2__30_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n998) );
  AND2X2 AND2X2_3196 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_0__31_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1001) );
  AND2X2 AND2X2_3197 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_1__31_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1002) );
  AND2X2 AND2X2_3198 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1003), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf2), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1004) );
  AND2X2 AND2X2_3199 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_3__31_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1005) );
  AND2X2 AND2X2_32 ( .A(u_sdrc_core_u_bank_ctl_rank_cnt_0_), .B(u_sdrc_core_u_bank_ctl_rank_cnt_1_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n268_1) );
  AND2X2 AND2X2_320 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf5), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_5_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n521) );
  AND2X2 AND2X2_3200 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_2__31_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1006) );
  AND2X2 AND2X2_3201 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n384_1), .B(app_rd_valid), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1017) );
  AND2X2 AND2X2_3202 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1017), .B(u_wb2sdrc_u_rddatafifo_wr_ptr_0_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1018) );
  AND2X2 AND2X2_3203 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1021), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1019), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n464) );
  AND2X2 AND2X2_3204 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1024), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1023), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n465) );
  AND2X2 AND2X2_3205 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1027), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1026), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n466) );
  AND2X2 AND2X2_3206 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1030), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1029), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n467) );
  AND2X2 AND2X2_3207 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1033), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1032), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n468) );
  AND2X2 AND2X2_3208 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1036), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1035), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n469) );
  AND2X2 AND2X2_3209 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1039), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1038), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n470) );
  AND2X2 AND2X2_321 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf1), .B(u_sdrc_core_r2b_raddr_5_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n522) );
  AND2X2 AND2X2_3210 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1042), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1041), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n471) );
  AND2X2 AND2X2_3211 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1045), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1044), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n472) );
  AND2X2 AND2X2_3212 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1048), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1047), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n473) );
  AND2X2 AND2X2_3213 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1051), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1050), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n474) );
  AND2X2 AND2X2_3214 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1054), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1053), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n475) );
  AND2X2 AND2X2_3215 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1057), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1056), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n476) );
  AND2X2 AND2X2_3216 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1060), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1059), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n477) );
  AND2X2 AND2X2_3217 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1063), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1062), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n478) );
  AND2X2 AND2X2_3218 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1066), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1065), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n479) );
  AND2X2 AND2X2_3219 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1069), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1068), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n480) );
  AND2X2 AND2X2_322 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n523), .B(sdram_resetn_bF_buf11), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_5__FF_INPUT) );
  AND2X2 AND2X2_3220 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1072), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1071), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n481) );
  AND2X2 AND2X2_3221 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1075), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1074), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n482) );
  AND2X2 AND2X2_3222 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1078), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1077), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n483) );
  AND2X2 AND2X2_3223 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1081), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1080), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n484) );
  AND2X2 AND2X2_3224 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1084), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1083), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n485) );
  AND2X2 AND2X2_3225 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1087), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1086), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n486) );
  AND2X2 AND2X2_3226 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1090), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1089), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n487) );
  AND2X2 AND2X2_3227 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1093), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1092), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n488) );
  AND2X2 AND2X2_3228 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1096), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1095), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n489) );
  AND2X2 AND2X2_3229 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1099), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1098), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n490) );
  AND2X2 AND2X2_323 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_6_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n525) );
  AND2X2 AND2X2_3230 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1102), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1101), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n491) );
  AND2X2 AND2X2_3231 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1105), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1104), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n492) );
  AND2X2 AND2X2_3232 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1108), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1107), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n493) );
  AND2X2 AND2X2_3233 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1111), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1110), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n494) );
  AND2X2 AND2X2_3234 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1114), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1113), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n495) );
  AND2X2 AND2X2_3235 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1119), .B(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf1), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1120) );
  AND2X2 AND2X2_3236 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf0), .B(u_wb2sdrc_rddatafifo_rd), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1121) );
  AND2X2 AND2X2_3237 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1119), .B(u_wb2sdrc_u_rddatafifo_rd_ptr_1_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1123) );
  AND2X2 AND2X2_3238 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf0), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1124) );
  AND2X2 AND2X2_3239 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1125), .B(u_wb2sdrc_rddatafifo_rd), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1126) );
  AND2X2 AND2X2_324 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf0), .B(u_sdrc_core_r2b_raddr_6_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n526) );
  AND2X2 AND2X2_3240 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1119), .B(u_wb2sdrc_u_rddatafifo_rd_ptr_2_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1128) );
  AND2X2 AND2X2_3241 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_rd_ptr_2_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1130) );
  AND2X2 AND2X2_3242 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1131), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1129), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1132) );
  AND2X2 AND2X2_3243 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1132), .B(u_wb2sdrc_rddatafifo_rd), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1133) );
  AND2X2 AND2X2_3244 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1151), .B(u_wb2sdrc_u_rddatafifo_grey_wr_ptr_0_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1152) );
  AND2X2 AND2X2_3245 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n384_1), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n375_1), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1154) );
  AND2X2 AND2X2_3246 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n446), .B(u_wb2sdrc_u_rddatafifo_wr_ptr_2_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1156) );
  AND2X2 AND2X2_3247 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1157), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1158), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1159) );
  AND2X2 AND2X2_3248 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1159), .B(app_rd_valid), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1160) );
  AND2X2 AND2X2_3249 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1160), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1155), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1161) );
  AND2X2 AND2X2_325 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n527), .B(sdram_resetn_bF_buf10), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_6__FF_INPUT) );
  AND2X2 AND2X2_3250 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1151), .B(u_wb2sdrc_u_rddatafifo_grey_wr_ptr_1_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1162) );
  AND2X2 AND2X2_3251 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1163), .B(app_rd_valid), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1164) );
  AND2X2 AND2X2_3252 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1164), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n389), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1165) );
  AND2X2 AND2X2_3253 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1151), .B(u_wb2sdrc_u_rddatafifo_grey_wr_ptr_2_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1168) );
  AND2X2 AND2X2_3254 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1151), .B(u_wb2sdrc_u_rddatafifo_wr_ptr_0_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1170) );
  AND2X2 AND2X2_3255 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1151), .B(u_wb2sdrc_u_rddatafifo_wr_ptr_1_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1172) );
  AND2X2 AND2X2_3256 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1151), .B(u_wb2sdrc_u_rddatafifo_wr_ptr_2_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1174) );
  AND2X2 AND2X2_3257 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n696_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n697_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n698) );
  AND2X2 AND2X2_3258 ( .A(u_wb2sdrc_u_wrdatafifo_sync_rd_ptr_1_2_), .B(u_wb2sdrc_u_wrdatafifo_sync_rd_ptr_1_3_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n699_1) );
  AND2X2 AND2X2_3259 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n700), .B(u_wb2sdrc_u_wrdatafifo_wr_ptr_2_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n701) );
  AND2X2 AND2X2_326 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_7_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n529) );
  AND2X2 AND2X2_3260 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n704_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n703), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n705_1) );
  AND2X2 AND2X2_3261 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n707), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n706), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n708_1) );
  AND2X2 AND2X2_3262 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n708_1), .B(u_wb2sdrc_u_wrdatafifo_wr_ptr_1_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n709_1) );
  AND2X2 AND2X2_3263 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n710), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n702_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n711_1) );
  AND2X2 AND2X2_3264 ( .A(u_wb2sdrc_u_wrdatafifo_sync_rd_ptr_1_0_), .B(u_wb2sdrc_u_wrdatafifo_sync_rd_ptr_1_1_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n712) );
  AND2X2 AND2X2_3265 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n716_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n715), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n717_1) );
  AND2X2 AND2X2_3266 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n714_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n718), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n719) );
  AND2X2 AND2X2_3267 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n720_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n721_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n722) );
  AND2X2 AND2X2_3268 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n705_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n724), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n725) );
  AND2X2 AND2X2_3269 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n723_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n727), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n728_1) );
  AND2X2 AND2X2_327 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf4), .B(u_sdrc_core_r2b_raddr_7_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n530) );
  AND2X2 AND2X2_3270 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n730), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n732_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n733_1) );
  AND2X2 AND2X2_3271 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n700), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n717_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n739) );
  AND2X2 AND2X2_3272 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n713), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n705_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n740_1) );
  AND2X2 AND2X2_3273 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n741_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n738_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n742) );
  AND2X2 AND2X2_3274 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n700), .B(u_wb2sdrc_u_wrdatafifo_sync_rd_ptr_1_1_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n744_1) );
  AND2X2 AND2X2_3275 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n705_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n702_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n745_1) );
  AND2X2 AND2X2_3276 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n746), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n743), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n747_1) );
  AND2X2 AND2X2_3277 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n748), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n737), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n749) );
  AND2X2 AND2X2_3278 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n750_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n736), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n751) );
  AND2X2 AND2X2_3279 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n735_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n752_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n753_1) );
  AND2X2 AND2X2_328 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n531), .B(sdram_resetn_bF_buf9), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_7__FF_INPUT) );
  AND2X2 AND2X2_3280 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n737), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n721_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n754) );
  AND2X2 AND2X2_3281 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n750_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n755), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n756_1) );
  AND2X2 AND2X2_3282 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n757_1), .B(u_wb2sdrc_u_wrdatafifo_wr_ptr_0_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n758) );
  AND2X2 AND2X2_3283 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n759_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n760), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n761) );
  AND2X2 AND2X2_3284 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n761), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n756_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n762_1) );
  AND2X2 AND2X2_3285 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n753_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n762_1), .Y(u_wb2sdrc_u_wrdatafifo_afull) );
  AND2X2 AND2X2_3286 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n738_1), .B(u_wb2sdrc_u_wrdatafifo_wr_en), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n817_1) );
  AND2X2 AND2X2_3287 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n743), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n724), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n818_1) );
  AND2X2 AND2X2_3288 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n818_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n817_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1) );
  AND2X2 AND2X2_3289 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n822_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n820_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n154) );
  AND2X2 AND2X2_329 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_8_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n533) );
  AND2X2 AND2X2_3290 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n825_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n824_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n157) );
  AND2X2 AND2X2_3291 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n828_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n827_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n160) );
  AND2X2 AND2X2_3292 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n831_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n830_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n163) );
  AND2X2 AND2X2_3293 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n834_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n833_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n166) );
  AND2X2 AND2X2_3294 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n837_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n836_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n169) );
  AND2X2 AND2X2_3295 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n840_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n839_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n172) );
  AND2X2 AND2X2_3296 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n843), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n842_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n175) );
  AND2X2 AND2X2_3297 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n846_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n845_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n178) );
  AND2X2 AND2X2_3298 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n849_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n848_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n181) );
  AND2X2 AND2X2_3299 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n852_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n851_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n184) );
  AND2X2 AND2X2_33 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n268_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n216_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n269) );
  AND2X2 AND2X2_330 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf3), .B(u_sdrc_core_r2b_raddr_8_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n534) );
  AND2X2 AND2X2_3300 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n855_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n854_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n187) );
  AND2X2 AND2X2_3301 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n858_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n857_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n190) );
  AND2X2 AND2X2_3302 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n861_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n860_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n193) );
  AND2X2 AND2X2_3303 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n864_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n863_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n196) );
  AND2X2 AND2X2_3304 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n867_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n866_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n199) );
  AND2X2 AND2X2_3305 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n870_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n869_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n202) );
  AND2X2 AND2X2_3306 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n873_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n872_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n205) );
  AND2X2 AND2X2_3307 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n876_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n875_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n208) );
  AND2X2 AND2X2_3308 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n879_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n878_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n211) );
  AND2X2 AND2X2_3309 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n882_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n881_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n214) );
  AND2X2 AND2X2_331 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n535), .B(sdram_resetn_bF_buf8), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_8__FF_INPUT) );
  AND2X2 AND2X2_3310 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n885_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n884_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n217) );
  AND2X2 AND2X2_3311 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n888_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n887_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n220) );
  AND2X2 AND2X2_3312 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n891_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n890_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n223) );
  AND2X2 AND2X2_3313 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n894_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n893_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n226) );
  AND2X2 AND2X2_3314 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n897_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n896_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n229) );
  AND2X2 AND2X2_3315 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n900_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n899_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n232) );
  AND2X2 AND2X2_3316 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n903_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n902_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n235) );
  AND2X2 AND2X2_3317 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n906_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n905_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n238) );
  AND2X2 AND2X2_3318 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n909_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n908_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n241) );
  AND2X2 AND2X2_3319 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n912_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n911_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n244) );
  AND2X2 AND2X2_332 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_9_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n537) );
  AND2X2 AND2X2_3320 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n915_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n914_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n247) );
  AND2X2 AND2X2_3321 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n918_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n917), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n250) );
  AND2X2 AND2X2_3322 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n921_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n920_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n253) );
  AND2X2 AND2X2_3323 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n924_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n923_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n256) );
  AND2X2 AND2X2_3324 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n927_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n926_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n259) );
  AND2X2 AND2X2_3325 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n743), .B(u_wb2sdrc_u_wrdatafifo_wr_ptr_2_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n929_1) );
  AND2X2 AND2X2_3326 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n817_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n929_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1) );
  AND2X2 AND2X2_3327 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n933_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n931_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n513) );
  AND2X2 AND2X2_3328 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n936_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n935_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n515) );
  AND2X2 AND2X2_3329 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n939_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n938_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n517) );
  AND2X2 AND2X2_333 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf2), .B(u_sdrc_core_r2b_raddr_9_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n538) );
  AND2X2 AND2X2_3330 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n942_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n941_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n519) );
  AND2X2 AND2X2_3331 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n945_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n944_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n521) );
  AND2X2 AND2X2_3332 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n948_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n947_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n523) );
  AND2X2 AND2X2_3333 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n951_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n950_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n525) );
  AND2X2 AND2X2_3334 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n954_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n953_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n527) );
  AND2X2 AND2X2_3335 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n957_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n956), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n529) );
  AND2X2 AND2X2_3336 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n960), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n959), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n531) );
  AND2X2 AND2X2_3337 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n963), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n962), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n533) );
  AND2X2 AND2X2_3338 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n966_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n965_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n535) );
  AND2X2 AND2X2_3339 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n969), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n968), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n537) );
  AND2X2 AND2X2_334 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n539), .B(sdram_resetn_bF_buf7), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_9__FF_INPUT) );
  AND2X2 AND2X2_3340 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n972), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n971_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n539) );
  AND2X2 AND2X2_3341 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n975), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n974), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n541) );
  AND2X2 AND2X2_3342 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n978_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n977_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n543) );
  AND2X2 AND2X2_3343 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n981), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n980), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n545) );
  AND2X2 AND2X2_3344 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n984_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n983), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n547) );
  AND2X2 AND2X2_3345 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n987), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n986), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n549) );
  AND2X2 AND2X2_3346 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n990), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n989_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n551) );
  AND2X2 AND2X2_3347 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n993_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n992), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n553) );
  AND2X2 AND2X2_3348 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n996), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n995), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n555) );
  AND2X2 AND2X2_3349 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n999_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n998_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n557) );
  AND2X2 AND2X2_335 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_10_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n541) );
  AND2X2 AND2X2_3350 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1002), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1001), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n559) );
  AND2X2 AND2X2_3351 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1005_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1004), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n561) );
  AND2X2 AND2X2_3352 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1008), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1007), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n563) );
  AND2X2 AND2X2_3353 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1011_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1010), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n565) );
  AND2X2 AND2X2_3354 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1014), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1013_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n567) );
  AND2X2 AND2X2_3355 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1017), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1016), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n569) );
  AND2X2 AND2X2_3356 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1020), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1019), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n571) );
  AND2X2 AND2X2_3357 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1023_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1022_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n573) );
  AND2X2 AND2X2_3358 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1026), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1025), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n575) );
  AND2X2 AND2X2_3359 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1029), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1028_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n577) );
  AND2X2 AND2X2_336 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf1), .B(u_sdrc_core_r2b_raddr_10_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n542) );
  AND2X2 AND2X2_3360 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1032), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1031_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n579) );
  AND2X2 AND2X2_3361 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1035_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1034), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n581) );
  AND2X2 AND2X2_3362 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1038_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1037_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n583) );
  AND2X2 AND2X2_3363 ( .A(u_wb2sdrc_u_wrdatafifo_wr_ptr_0_), .B(u_wb2sdrc_u_wrdatafifo_wr_en), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1040_1) );
  AND2X2 AND2X2_3364 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n724), .B(u_wb2sdrc_u_wrdatafifo_wr_ptr_1_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1041_1) );
  AND2X2 AND2X2_3365 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1041_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1040_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1) );
  AND2X2 AND2X2_3366 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1045_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1043_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n586) );
  AND2X2 AND2X2_3367 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1048_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1047_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n588) );
  AND2X2 AND2X2_3368 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1051_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1050_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n590) );
  AND2X2 AND2X2_3369 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1054_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1053_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n592) );
  AND2X2 AND2X2_337 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n543), .B(sdram_resetn_bF_buf6), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_10__FF_INPUT) );
  AND2X2 AND2X2_3370 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1057_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1056_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n594) );
  AND2X2 AND2X2_3371 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1060_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1059_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n596) );
  AND2X2 AND2X2_3372 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1063_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1062_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n598) );
  AND2X2 AND2X2_3373 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1066_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1065_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n600) );
  AND2X2 AND2X2_3374 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1069_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1068_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n602) );
  AND2X2 AND2X2_3375 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1072), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1071), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n604) );
  AND2X2 AND2X2_3376 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1075), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1074), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n606) );
  AND2X2 AND2X2_3377 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1078), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1077), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n608) );
  AND2X2 AND2X2_3378 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1081), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1080), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n610) );
  AND2X2 AND2X2_3379 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1084), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1083), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n612) );
  AND2X2 AND2X2_338 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf5), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_11_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n545) );
  AND2X2 AND2X2_3380 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1087), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1086), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n614) );
  AND2X2 AND2X2_3381 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1090), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1089), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n616) );
  AND2X2 AND2X2_3382 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1093), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1092), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n618) );
  AND2X2 AND2X2_3383 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1096), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1095), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n620) );
  AND2X2 AND2X2_3384 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1099), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1098), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n622) );
  AND2X2 AND2X2_3385 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1102), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1101), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n624) );
  AND2X2 AND2X2_3386 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1105), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1104), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n626) );
  AND2X2 AND2X2_3387 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1108), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1107), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n628) );
  AND2X2 AND2X2_3388 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1111), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1110), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n630) );
  AND2X2 AND2X2_3389 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1114), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1113), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n632) );
  AND2X2 AND2X2_339 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf0), .B(u_sdrc_core_r2b_raddr_11_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n546) );
  AND2X2 AND2X2_3390 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1117), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1116), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n634) );
  AND2X2 AND2X2_3391 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1120), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1119), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n636) );
  AND2X2 AND2X2_3392 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1123), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1122), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n638) );
  AND2X2 AND2X2_3393 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1126), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1125), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n640) );
  AND2X2 AND2X2_3394 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1129), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1128), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n642) );
  AND2X2 AND2X2_3395 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1132), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1131), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n644) );
  AND2X2 AND2X2_3396 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1135), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1134), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n646) );
  AND2X2 AND2X2_3397 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1138), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1137), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n648) );
  AND2X2 AND2X2_3398 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1141), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1140), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n650) );
  AND2X2 AND2X2_3399 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1144), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1143), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n652) );
  AND2X2 AND2X2_34 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n270_1), .B(u_sdrc_core_u_bank_ctl_rank_cnt_2_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n271) );
  AND2X2 AND2X2_340 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n547), .B(sdram_resetn_bF_buf5), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_11__FF_INPUT) );
  AND2X2 AND2X2_3400 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1147), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1146), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n654) );
  AND2X2 AND2X2_3401 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1150), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1149), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n656) );
  AND2X2 AND2X2_3402 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_mem_1__0_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1152) );
  AND2X2 AND2X2_3403 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo_mem_0__0_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1153) );
  AND2X2 AND2X2_3404 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1154), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf7), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1155) );
  AND2X2 AND2X2_3405 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_1_), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf5), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156) );
  AND2X2 AND2X2_3406 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo_mem_3__0_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1157) );
  AND2X2 AND2X2_3407 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_1_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158) );
  AND2X2 AND2X2_3408 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo_mem_2__0_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1159) );
  AND2X2 AND2X2_3409 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_5__0_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1163) );
  AND2X2 AND2X2_341 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_12_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n549) );
  AND2X2 AND2X2_3410 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_4__0_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1164) );
  AND2X2 AND2X2_3411 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1165), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf6), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1166) );
  AND2X2 AND2X2_3412 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_mem_7__0_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1167) );
  AND2X2 AND2X2_3413 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_mem_6__0_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1168) );
  AND2X2 AND2X2_3414 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1162), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1171), .Y(app_wr_data_0_) );
  AND2X2 AND2X2_3415 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_5__1_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1173) );
  AND2X2 AND2X2_3416 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_4__1_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1174) );
  AND2X2 AND2X2_3417 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1175), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf5), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1176) );
  AND2X2 AND2X2_3418 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_6__1_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1177) );
  AND2X2 AND2X2_3419 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_7__1_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1178) );
  AND2X2 AND2X2_342 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf4), .B(u_sdrc_core_r2b_raddr_12_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n550) );
  AND2X2 AND2X2_3420 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_1__1_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1182) );
  AND2X2 AND2X2_3421 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_0__1_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1183) );
  AND2X2 AND2X2_3422 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1184), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf4), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1185) );
  AND2X2 AND2X2_3423 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_2__1_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1186) );
  AND2X2 AND2X2_3424 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_3__1_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1187) );
  AND2X2 AND2X2_3425 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1181), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1190), .Y(app_wr_data_1_) );
  AND2X2 AND2X2_3426 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_1__2_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1192) );
  AND2X2 AND2X2_3427 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_0__2_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1193) );
  AND2X2 AND2X2_3428 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1194), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf3), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1195) );
  AND2X2 AND2X2_3429 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_2__2_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1196) );
  AND2X2 AND2X2_343 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n551), .B(sdram_resetn_bF_buf4), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_12__FF_INPUT) );
  AND2X2 AND2X2_3430 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_3__2_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1197) );
  AND2X2 AND2X2_3431 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_5__2_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1201) );
  AND2X2 AND2X2_3432 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_4__2_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1202) );
  AND2X2 AND2X2_3433 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1203), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf2), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1204) );
  AND2X2 AND2X2_3434 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_7__2_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1205) );
  AND2X2 AND2X2_3435 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_6__2_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1206) );
  AND2X2 AND2X2_3436 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1209), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1200), .Y(app_wr_data_2_) );
  AND2X2 AND2X2_3437 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo_mem_5__3_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1211) );
  AND2X2 AND2X2_3438 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_4__3_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1212) );
  AND2X2 AND2X2_3439 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1213), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1214) );
  AND2X2 AND2X2_344 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_0_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n553) );
  AND2X2 AND2X2_3440 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_6__3_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1215) );
  AND2X2 AND2X2_3441 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_7__3_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1216) );
  AND2X2 AND2X2_3442 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_mem_1__3_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1220) );
  AND2X2 AND2X2_3443 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo_mem_0__3_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1221) );
  AND2X2 AND2X2_3444 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1222), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf0), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1223) );
  AND2X2 AND2X2_3445 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_2__3_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1224) );
  AND2X2 AND2X2_3446 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_3__3_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1225) );
  AND2X2 AND2X2_3447 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1219), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1228), .Y(app_wr_data_3_) );
  AND2X2 AND2X2_3448 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_5__4_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1230) );
  AND2X2 AND2X2_3449 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_mem_4__4_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1231) );
  AND2X2 AND2X2_345 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf3), .B(u_sdrc_core_r2b_caddr_0_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n554) );
  AND2X2 AND2X2_3450 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1232), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf7), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1233) );
  AND2X2 AND2X2_3451 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo_mem_6__4_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1234) );
  AND2X2 AND2X2_3452 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo_mem_7__4_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1235) );
  AND2X2 AND2X2_3453 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_1__4_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1239) );
  AND2X2 AND2X2_3454 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_0__4_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1240) );
  AND2X2 AND2X2_3455 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1241), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf6), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1242) );
  AND2X2 AND2X2_3456 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_mem_3__4_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1243) );
  AND2X2 AND2X2_3457 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_mem_2__4_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1244) );
  AND2X2 AND2X2_3458 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1247), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1238), .Y(app_wr_data_4_) );
  AND2X2 AND2X2_3459 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_5__5_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1249) );
  AND2X2 AND2X2_346 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n555), .B(sdram_resetn_bF_buf3), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_0__FF_INPUT) );
  AND2X2 AND2X2_3460 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_4__5_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1250) );
  AND2X2 AND2X2_3461 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1251), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf5), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1252) );
  AND2X2 AND2X2_3462 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_6__5_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1253) );
  AND2X2 AND2X2_3463 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_7__5_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1254) );
  AND2X2 AND2X2_3464 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_1__5_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1258) );
  AND2X2 AND2X2_3465 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_0__5_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1259) );
  AND2X2 AND2X2_3466 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1260), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf4), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1261) );
  AND2X2 AND2X2_3467 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_3__5_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1262) );
  AND2X2 AND2X2_3468 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_2__5_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1263) );
  AND2X2 AND2X2_3469 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1266), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1257), .Y(app_wr_data_5_) );
  AND2X2 AND2X2_347 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_1_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n557) );
  AND2X2 AND2X2_3470 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_5__6_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1268) );
  AND2X2 AND2X2_3471 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_4__6_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1269) );
  AND2X2 AND2X2_3472 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1270), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf3), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1271) );
  AND2X2 AND2X2_3473 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_6__6_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1272) );
  AND2X2 AND2X2_3474 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_7__6_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1273) );
  AND2X2 AND2X2_3475 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_1__6_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1277) );
  AND2X2 AND2X2_3476 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_0__6_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1278) );
  AND2X2 AND2X2_3477 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1279), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf2), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1280) );
  AND2X2 AND2X2_3478 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_2__6_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1281) );
  AND2X2 AND2X2_3479 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_3__6_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1282) );
  AND2X2 AND2X2_348 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf2), .B(u_sdrc_core_r2b_caddr_1_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n558) );
  AND2X2 AND2X2_3480 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1276), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1285), .Y(app_wr_data_6_) );
  AND2X2 AND2X2_3481 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo_mem_5__7_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1287) );
  AND2X2 AND2X2_3482 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_4__7_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1288) );
  AND2X2 AND2X2_3483 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1289), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1290) );
  AND2X2 AND2X2_3484 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_6__7_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1291) );
  AND2X2 AND2X2_3485 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_7__7_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1292) );
  AND2X2 AND2X2_3486 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_mem_1__7_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1296) );
  AND2X2 AND2X2_3487 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo_mem_0__7_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1297) );
  AND2X2 AND2X2_3488 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1298), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf0), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1299) );
  AND2X2 AND2X2_3489 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_2__7_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1300) );
  AND2X2 AND2X2_349 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n559), .B(sdram_resetn_bF_buf2), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_1__FF_INPUT) );
  AND2X2 AND2X2_3490 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_3__7_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1301) );
  AND2X2 AND2X2_3491 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1295), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1304), .Y(app_wr_data_7_) );
  AND2X2 AND2X2_3492 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_1__8_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1306) );
  AND2X2 AND2X2_3493 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_mem_0__8_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1307) );
  AND2X2 AND2X2_3494 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1308), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf7), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1309) );
  AND2X2 AND2X2_3495 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo_mem_3__8_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1310) );
  AND2X2 AND2X2_3496 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo_mem_2__8_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1311) );
  AND2X2 AND2X2_3497 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_5__8_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1315) );
  AND2X2 AND2X2_3498 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_4__8_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1316) );
  AND2X2 AND2X2_3499 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1317), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf6), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1318) );
  AND2X2 AND2X2_35 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n252_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n272_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n273_1) );
  AND2X2 AND2X2_350 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_2_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n561) );
  AND2X2 AND2X2_3500 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_mem_7__8_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1319) );
  AND2X2 AND2X2_3501 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_mem_6__8_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1320) );
  AND2X2 AND2X2_3502 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1314), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1323), .Y(app_wr_data_8_) );
  AND2X2 AND2X2_3503 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_1__9_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1325) );
  AND2X2 AND2X2_3504 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_0__9_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1326) );
  AND2X2 AND2X2_3505 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1327), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf5), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1328) );
  AND2X2 AND2X2_3506 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_2__9_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1329) );
  AND2X2 AND2X2_3507 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_3__9_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1330) );
  AND2X2 AND2X2_3508 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_5__9_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1334) );
  AND2X2 AND2X2_3509 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_4__9_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1335) );
  AND2X2 AND2X2_351 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf1), .B(u_sdrc_core_r2b_caddr_2_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n562) );
  AND2X2 AND2X2_3510 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1336), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf4), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1337) );
  AND2X2 AND2X2_3511 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_7__9_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1338) );
  AND2X2 AND2X2_3512 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_6__9_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1339) );
  AND2X2 AND2X2_3513 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1342), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1333), .Y(app_wr_data_9_) );
  AND2X2 AND2X2_3514 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_5__10_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1344) );
  AND2X2 AND2X2_3515 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_4__10_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1345) );
  AND2X2 AND2X2_3516 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1346), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf3), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1347) );
  AND2X2 AND2X2_3517 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_6__10_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1348) );
  AND2X2 AND2X2_3518 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_7__10_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1349) );
  AND2X2 AND2X2_3519 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_1__10_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1353) );
  AND2X2 AND2X2_352 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n563), .B(sdram_resetn_bF_buf1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_2__FF_INPUT) );
  AND2X2 AND2X2_3520 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_0__10_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1354) );
  AND2X2 AND2X2_3521 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1355), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf2), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1356) );
  AND2X2 AND2X2_3522 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_2__10_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1357) );
  AND2X2 AND2X2_3523 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_3__10_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1358) );
  AND2X2 AND2X2_3524 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1352), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1361), .Y(app_wr_data_10_) );
  AND2X2 AND2X2_3525 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo_mem_5__11_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1363) );
  AND2X2 AND2X2_3526 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_4__11_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1364) );
  AND2X2 AND2X2_3527 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1365), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1366) );
  AND2X2 AND2X2_3528 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_6__11_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1367) );
  AND2X2 AND2X2_3529 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_7__11_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1369) );
  AND2X2 AND2X2_353 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_3_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n565) );
  AND2X2 AND2X2_3530 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_mem_1__11_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1372) );
  AND2X2 AND2X2_3531 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo_mem_0__11_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1373) );
  AND2X2 AND2X2_3532 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1374), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf0), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1375) );
  AND2X2 AND2X2_3533 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_3__11_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1376) );
  AND2X2 AND2X2_3534 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_2__11_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1377) );
  AND2X2 AND2X2_3535 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1380), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1371), .Y(app_wr_data_11_) );
  AND2X2 AND2X2_3536 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_1__12_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1382) );
  AND2X2 AND2X2_3537 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_mem_0__12_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1383) );
  AND2X2 AND2X2_3538 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1384), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf7), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1385) );
  AND2X2 AND2X2_3539 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo_mem_2__12_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1386) );
  AND2X2 AND2X2_354 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf0), .B(u_sdrc_core_r2b_caddr_3_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n566) );
  AND2X2 AND2X2_3540 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo_mem_3__12_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1387) );
  AND2X2 AND2X2_3541 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_5__12_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1391) );
  AND2X2 AND2X2_3542 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_4__12_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1392) );
  AND2X2 AND2X2_3543 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1393), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf6), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1394) );
  AND2X2 AND2X2_3544 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_mem_7__12_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1395) );
  AND2X2 AND2X2_3545 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_mem_6__12_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1396) );
  AND2X2 AND2X2_3546 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1399), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1390), .Y(app_wr_data_12_) );
  AND2X2 AND2X2_3547 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_5__13_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1401) );
  AND2X2 AND2X2_3548 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_4__13_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1402) );
  AND2X2 AND2X2_3549 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1403), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf5), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1404) );
  AND2X2 AND2X2_355 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n567), .B(sdram_resetn_bF_buf0), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_3__FF_INPUT) );
  AND2X2 AND2X2_3550 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_6__13_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1405) );
  AND2X2 AND2X2_3551 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_7__13_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1406) );
  AND2X2 AND2X2_3552 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_1__13_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1410) );
  AND2X2 AND2X2_3553 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_0__13_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1411) );
  AND2X2 AND2X2_3554 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1412), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf4), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1413) );
  AND2X2 AND2X2_3555 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_3__13_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1414) );
  AND2X2 AND2X2_3556 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_2__13_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1415) );
  AND2X2 AND2X2_3557 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1418), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1409), .Y(app_wr_data_13_) );
  AND2X2 AND2X2_3558 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_5__14_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1420) );
  AND2X2 AND2X2_3559 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_4__14_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1421) );
  AND2X2 AND2X2_356 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf5), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_4_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n569) );
  AND2X2 AND2X2_3560 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1422), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf3), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1423) );
  AND2X2 AND2X2_3561 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_6__14_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1424) );
  AND2X2 AND2X2_3562 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_7__14_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1425) );
  AND2X2 AND2X2_3563 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_1__14_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1429) );
  AND2X2 AND2X2_3564 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_0__14_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1430) );
  AND2X2 AND2X2_3565 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1431), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf2), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1432) );
  AND2X2 AND2X2_3566 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_2__14_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1433) );
  AND2X2 AND2X2_3567 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_3__14_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1434) );
  AND2X2 AND2X2_3568 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1428), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1437), .Y(app_wr_data_14_) );
  AND2X2 AND2X2_3569 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo_mem_1__15_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1439) );
  AND2X2 AND2X2_357 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf4), .B(u_sdrc_core_r2b_caddr_4_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n570) );
  AND2X2 AND2X2_3570 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_0__15_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1440) );
  AND2X2 AND2X2_3571 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1441), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1442) );
  AND2X2 AND2X2_3572 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_3__15_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1443) );
  AND2X2 AND2X2_3573 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_2__15_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1444) );
  AND2X2 AND2X2_3574 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_mem_5__15_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1448) );
  AND2X2 AND2X2_3575 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo_mem_4__15_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1449) );
  AND2X2 AND2X2_3576 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1450), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf0), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1451) );
  AND2X2 AND2X2_3577 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_6__15_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1452) );
  AND2X2 AND2X2_3578 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_7__15_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1453) );
  AND2X2 AND2X2_3579 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1447), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1456), .Y(app_wr_data_15_) );
  AND2X2 AND2X2_358 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n571), .B(sdram_resetn_bF_buf49), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_4__FF_INPUT) );
  AND2X2 AND2X2_3580 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_1__16_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1458) );
  AND2X2 AND2X2_3581 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_mem_0__16_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1459) );
  AND2X2 AND2X2_3582 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1460), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf7), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1461) );
  AND2X2 AND2X2_3583 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo_mem_3__16_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1462) );
  AND2X2 AND2X2_3584 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo_mem_2__16_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1463) );
  AND2X2 AND2X2_3585 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_5__16_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1467) );
  AND2X2 AND2X2_3586 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_4__16_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1468) );
  AND2X2 AND2X2_3587 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1469), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf6), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1470) );
  AND2X2 AND2X2_3588 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_mem_7__16_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1471) );
  AND2X2 AND2X2_3589 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_mem_6__16_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1472) );
  AND2X2 AND2X2_359 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_5_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n573) );
  AND2X2 AND2X2_3590 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1466), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1475), .Y(app_wr_data_16_) );
  AND2X2 AND2X2_3591 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_5__17_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1477) );
  AND2X2 AND2X2_3592 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_4__17_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1478) );
  AND2X2 AND2X2_3593 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1479), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf5), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1480) );
  AND2X2 AND2X2_3594 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_6__17_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1481) );
  AND2X2 AND2X2_3595 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_7__17_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1482) );
  AND2X2 AND2X2_3596 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_1__17_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1486) );
  AND2X2 AND2X2_3597 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_0__17_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1487) );
  AND2X2 AND2X2_3598 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1488), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf4), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1489) );
  AND2X2 AND2X2_3599 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_2__17_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1490) );
  AND2X2 AND2X2_36 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n243), .B(u_sdrc_core_b2x_idle), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n274_1) );
  AND2X2 AND2X2_360 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf3), .B(u_sdrc_core_r2b_caddr_5_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n574) );
  AND2X2 AND2X2_3600 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_3__17_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1491) );
  AND2X2 AND2X2_3601 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1485), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1494), .Y(app_wr_data_17_) );
  AND2X2 AND2X2_3602 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_1__18_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1496) );
  AND2X2 AND2X2_3603 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_0__18_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1497) );
  AND2X2 AND2X2_3604 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1498), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf3), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1499) );
  AND2X2 AND2X2_3605 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_2__18_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1500) );
  AND2X2 AND2X2_3606 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_3__18_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1501) );
  AND2X2 AND2X2_3607 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_5__18_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1505) );
  AND2X2 AND2X2_3608 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_4__18_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1506) );
  AND2X2 AND2X2_3609 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1507), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf2), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1508) );
  AND2X2 AND2X2_361 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n575), .B(sdram_resetn_bF_buf48), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_5__FF_INPUT) );
  AND2X2 AND2X2_3610 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_7__18_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1509) );
  AND2X2 AND2X2_3611 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_6__18_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1510) );
  AND2X2 AND2X2_3612 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1513), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1504), .Y(app_wr_data_18_) );
  AND2X2 AND2X2_3613 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo_mem_1__19_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1515) );
  AND2X2 AND2X2_3614 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_0__19_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1516) );
  AND2X2 AND2X2_3615 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1517), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1518) );
  AND2X2 AND2X2_3616 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_3__19_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1519) );
  AND2X2 AND2X2_3617 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_2__19_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1520) );
  AND2X2 AND2X2_3618 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_mem_5__19_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1524) );
  AND2X2 AND2X2_3619 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo_mem_4__19_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1525) );
  AND2X2 AND2X2_362 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_6_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n577) );
  AND2X2 AND2X2_3620 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1526), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf0), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1527) );
  AND2X2 AND2X2_3621 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_7__19_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1528) );
  AND2X2 AND2X2_3622 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_6__19_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1529) );
  AND2X2 AND2X2_3623 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1523), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1532), .Y(app_wr_data_19_) );
  AND2X2 AND2X2_3624 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_5__20_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1534) );
  AND2X2 AND2X2_3625 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_mem_4__20_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1535) );
  AND2X2 AND2X2_3626 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1536), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf7), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1537) );
  AND2X2 AND2X2_3627 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo_mem_6__20_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1538) );
  AND2X2 AND2X2_3628 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo_mem_7__20_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1539) );
  AND2X2 AND2X2_3629 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_1__20_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1543) );
  AND2X2 AND2X2_363 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf2), .B(u_sdrc_core_r2b_caddr_6_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n578) );
  AND2X2 AND2X2_3630 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_0__20_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1544) );
  AND2X2 AND2X2_3631 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1545), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf6), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1546) );
  AND2X2 AND2X2_3632 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_mem_2__20_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1547) );
  AND2X2 AND2X2_3633 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_mem_3__20_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1548) );
  AND2X2 AND2X2_3634 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1542), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1551), .Y(app_wr_data_20_) );
  AND2X2 AND2X2_3635 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_1__21_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1553) );
  AND2X2 AND2X2_3636 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_0__21_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1554) );
  AND2X2 AND2X2_3637 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1555), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf5), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1556) );
  AND2X2 AND2X2_3638 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_3__21_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1557) );
  AND2X2 AND2X2_3639 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_2__21_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1558) );
  AND2X2 AND2X2_364 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n579), .B(sdram_resetn_bF_buf47), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_6__FF_INPUT) );
  AND2X2 AND2X2_3640 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_5__21_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1562) );
  AND2X2 AND2X2_3641 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_4__21_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1563) );
  AND2X2 AND2X2_3642 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1564), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf4), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1565) );
  AND2X2 AND2X2_3643 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_7__21_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1566) );
  AND2X2 AND2X2_3644 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_6__21_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1567) );
  AND2X2 AND2X2_3645 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1561), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1570), .Y(app_wr_data_21_) );
  AND2X2 AND2X2_3646 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_1__22_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1572) );
  AND2X2 AND2X2_3647 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_0__22_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1573) );
  AND2X2 AND2X2_3648 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1574), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf3), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1575) );
  AND2X2 AND2X2_3649 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_2__22_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1576) );
  AND2X2 AND2X2_365 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_7_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n581) );
  AND2X2 AND2X2_3650 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_3__22_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1578) );
  AND2X2 AND2X2_3651 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_5__22_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1581) );
  AND2X2 AND2X2_3652 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_4__22_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1582) );
  AND2X2 AND2X2_3653 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1583), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf2), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1584) );
  AND2X2 AND2X2_3654 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_7__22_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1585) );
  AND2X2 AND2X2_3655 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_6__22_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1586) );
  AND2X2 AND2X2_3656 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1589), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1580), .Y(app_wr_data_22_) );
  AND2X2 AND2X2_3657 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo_mem_5__23_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1591) );
  AND2X2 AND2X2_3658 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_4__23_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1592) );
  AND2X2 AND2X2_3659 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1593), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1594) );
  AND2X2 AND2X2_366 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf1), .B(u_sdrc_core_r2b_caddr_7_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n582) );
  AND2X2 AND2X2_3660 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_6__23_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1595) );
  AND2X2 AND2X2_3661 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_7__23_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1596) );
  AND2X2 AND2X2_3662 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_mem_1__23_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1600) );
  AND2X2 AND2X2_3663 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo_mem_0__23_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1601) );
  AND2X2 AND2X2_3664 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1602), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf0), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1603) );
  AND2X2 AND2X2_3665 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_2__23_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1604) );
  AND2X2 AND2X2_3666 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_3__23_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1605) );
  AND2X2 AND2X2_3667 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1599), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1608), .Y(app_wr_data_23_) );
  AND2X2 AND2X2_3668 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_1__24_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1610) );
  AND2X2 AND2X2_3669 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_mem_0__24_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1611) );
  AND2X2 AND2X2_367 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n583), .B(sdram_resetn_bF_buf46), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_7__FF_INPUT) );
  AND2X2 AND2X2_3670 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1612), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf7), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1613) );
  AND2X2 AND2X2_3671 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo_mem_3__24_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1614) );
  AND2X2 AND2X2_3672 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo_mem_2__24_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1615) );
  AND2X2 AND2X2_3673 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_5__24_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1619) );
  AND2X2 AND2X2_3674 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_4__24_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1620) );
  AND2X2 AND2X2_3675 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1621), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf6), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1622) );
  AND2X2 AND2X2_3676 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_mem_7__24_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1623) );
  AND2X2 AND2X2_3677 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_mem_6__24_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1624) );
  AND2X2 AND2X2_3678 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1618), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1627), .Y(app_wr_data_24_) );
  AND2X2 AND2X2_3679 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_5__25_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1629) );
  AND2X2 AND2X2_368 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_8_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n585) );
  AND2X2 AND2X2_3680 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_4__25_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1630) );
  AND2X2 AND2X2_3681 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1631), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf5), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1632) );
  AND2X2 AND2X2_3682 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_6__25_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1633) );
  AND2X2 AND2X2_3683 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_7__25_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1634) );
  AND2X2 AND2X2_3684 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_1__25_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1638) );
  AND2X2 AND2X2_3685 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_0__25_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1639) );
  AND2X2 AND2X2_3686 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1640), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf4), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1641) );
  AND2X2 AND2X2_3687 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_2__25_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1642) );
  AND2X2 AND2X2_3688 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_3__25_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1643) );
  AND2X2 AND2X2_3689 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1637), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1646), .Y(app_wr_data_25_) );
  AND2X2 AND2X2_369 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf0), .B(u_sdrc_core_r2b_caddr_8_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n586) );
  AND2X2 AND2X2_3690 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_5__26_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1648) );
  AND2X2 AND2X2_3691 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_4__26_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1649) );
  AND2X2 AND2X2_3692 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1650), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf3), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1651) );
  AND2X2 AND2X2_3693 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_6__26_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1652) );
  AND2X2 AND2X2_3694 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_7__26_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1653) );
  AND2X2 AND2X2_3695 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_1__26_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1657) );
  AND2X2 AND2X2_3696 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_0__26_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1658) );
  AND2X2 AND2X2_3697 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1659), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf2), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1660) );
  AND2X2 AND2X2_3698 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_2__26_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1661) );
  AND2X2 AND2X2_3699 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_3__26_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1662) );
  AND2X2 AND2X2_37 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n276), .B(sdram_resetn_bF_buf47), .Y(u_sdrc_core_u_bank_ctl_rank_cnt_2__FF_INPUT) );
  AND2X2 AND2X2_370 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n587), .B(sdram_resetn_bF_buf45), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_8__FF_INPUT) );
  AND2X2 AND2X2_3700 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1656), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1665), .Y(app_wr_data_26_) );
  AND2X2 AND2X2_3701 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo_mem_1__27_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1667) );
  AND2X2 AND2X2_3702 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_0__27_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1668) );
  AND2X2 AND2X2_3703 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1669), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1670) );
  AND2X2 AND2X2_3704 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_3__27_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1671) );
  AND2X2 AND2X2_3705 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_2__27_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1672) );
  AND2X2 AND2X2_3706 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_mem_5__27_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1676) );
  AND2X2 AND2X2_3707 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo_mem_4__27_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1677) );
  AND2X2 AND2X2_3708 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1678), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf0), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1679) );
  AND2X2 AND2X2_3709 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_6__27_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1680) );
  AND2X2 AND2X2_371 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_9_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n589) );
  AND2X2 AND2X2_3710 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_7__27_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1681) );
  AND2X2 AND2X2_3711 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1675), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1684), .Y(app_wr_data_27_) );
  AND2X2 AND2X2_3712 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_1__28_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1686) );
  AND2X2 AND2X2_3713 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_mem_0__28_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1687) );
  AND2X2 AND2X2_3714 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1688), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf7), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1689) );
  AND2X2 AND2X2_3715 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo_mem_2__28_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1690) );
  AND2X2 AND2X2_3716 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo_mem_3__28_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1692) );
  AND2X2 AND2X2_3717 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_5__28_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1695) );
  AND2X2 AND2X2_3718 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_4__28_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1696) );
  AND2X2 AND2X2_3719 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1697), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf6), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1698) );
  AND2X2 AND2X2_372 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf4), .B(u_sdrc_core_r2b_caddr_9_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n590) );
  AND2X2 AND2X2_3720 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_mem_7__28_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1699) );
  AND2X2 AND2X2_3721 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_mem_6__28_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1700) );
  AND2X2 AND2X2_3722 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1703), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1694), .Y(app_wr_data_28_) );
  AND2X2 AND2X2_3723 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_5__29_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1705) );
  AND2X2 AND2X2_3724 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_4__29_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1706) );
  AND2X2 AND2X2_3725 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1707), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf5), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1708) );
  AND2X2 AND2X2_3726 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_6__29_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1709) );
  AND2X2 AND2X2_3727 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_7__29_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1711) );
  AND2X2 AND2X2_3728 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_1__29_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1714) );
  AND2X2 AND2X2_3729 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_0__29_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1715) );
  AND2X2 AND2X2_373 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n591), .B(sdram_resetn_bF_buf44), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_9__FF_INPUT) );
  AND2X2 AND2X2_3730 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1716), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf4), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1717) );
  AND2X2 AND2X2_3731 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_3__29_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1718) );
  AND2X2 AND2X2_3732 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_2__29_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1719) );
  AND2X2 AND2X2_3733 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1722), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1713), .Y(app_wr_data_29_) );
  AND2X2 AND2X2_3734 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_5__30_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1724) );
  AND2X2 AND2X2_3735 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_4__30_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1725) );
  AND2X2 AND2X2_3736 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1726), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf3), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1727) );
  AND2X2 AND2X2_3737 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_6__30_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1728) );
  AND2X2 AND2X2_3738 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_7__30_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1729) );
  AND2X2 AND2X2_3739 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_1__30_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1733) );
  AND2X2 AND2X2_374 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf5), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_10_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n593) );
  AND2X2 AND2X2_3740 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_0__30_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1734) );
  AND2X2 AND2X2_3741 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1735), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf2), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1736) );
  AND2X2 AND2X2_3742 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_2__30_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1737) );
  AND2X2 AND2X2_3743 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_3__30_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1738) );
  AND2X2 AND2X2_3744 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1732), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1741), .Y(app_wr_data_30_) );
  AND2X2 AND2X2_3745 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo_mem_1__31_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1743) );
  AND2X2 AND2X2_3746 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_0__31_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1744) );
  AND2X2 AND2X2_3747 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1745), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1746) );
  AND2X2 AND2X2_3748 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_2__31_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1747) );
  AND2X2 AND2X2_3749 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_3__31_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1748) );
  AND2X2 AND2X2_375 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf3), .B(u_sdrc_core_r2b_caddr_10_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n594) );
  AND2X2 AND2X2_3750 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_mem_5__31_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1752) );
  AND2X2 AND2X2_3751 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo_mem_4__31_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1753) );
  AND2X2 AND2X2_3752 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1754), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf0), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1755) );
  AND2X2 AND2X2_3753 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_6__31_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1756) );
  AND2X2 AND2X2_3754 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_7__31_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1757) );
  AND2X2 AND2X2_3755 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1751), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1760), .Y(app_wr_data_31_) );
  AND2X2 AND2X2_3756 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_5__32_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1762) );
  AND2X2 AND2X2_3757 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_mem_4__32_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1763) );
  AND2X2 AND2X2_3758 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1764), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf7), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1765) );
  AND2X2 AND2X2_3759 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo_mem_6__32_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1766) );
  AND2X2 AND2X2_376 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n595), .B(sdram_resetn_bF_buf43), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_10__FF_INPUT) );
  AND2X2 AND2X2_3760 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo_mem_7__32_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1767) );
  AND2X2 AND2X2_3761 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_1__32_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1771) );
  AND2X2 AND2X2_3762 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_0__32_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1772) );
  AND2X2 AND2X2_3763 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1773), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf6), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1774) );
  AND2X2 AND2X2_3764 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_mem_3__32_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1775) );
  AND2X2 AND2X2_3765 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_mem_2__32_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1776) );
  AND2X2 AND2X2_3766 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1779), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1770), .Y(app_wr_en_n_0_) );
  AND2X2 AND2X2_3767 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_5__33_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1781) );
  AND2X2 AND2X2_3768 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_4__33_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1782) );
  AND2X2 AND2X2_3769 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1783), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf5), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1784) );
  AND2X2 AND2X2_377 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_11_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n597) );
  AND2X2 AND2X2_3770 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_6__33_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1785) );
  AND2X2 AND2X2_3771 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_7__33_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1786) );
  AND2X2 AND2X2_3772 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_1__33_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1790) );
  AND2X2 AND2X2_3773 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_0__33_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1791) );
  AND2X2 AND2X2_3774 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1792), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf4), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1793) );
  AND2X2 AND2X2_3775 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_2__33_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1794) );
  AND2X2 AND2X2_3776 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_3__33_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1795) );
  AND2X2 AND2X2_3777 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1789), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1798), .Y(app_wr_en_n_1_) );
  AND2X2 AND2X2_3778 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_1__34_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1800) );
  AND2X2 AND2X2_3779 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_0__34_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1801) );
  AND2X2 AND2X2_378 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf2), .B(1'b0), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n598) );
  AND2X2 AND2X2_3780 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1802), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf3), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1803) );
  AND2X2 AND2X2_3781 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_3__34_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1804) );
  AND2X2 AND2X2_3782 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_2__34_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1805) );
  AND2X2 AND2X2_3783 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_5__34_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1809) );
  AND2X2 AND2X2_3784 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_4__34_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1810) );
  AND2X2 AND2X2_3785 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1811), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf2), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1812) );
  AND2X2 AND2X2_3786 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_7__34_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1813) );
  AND2X2 AND2X2_3787 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_6__34_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1814) );
  AND2X2 AND2X2_3788 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1808), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1817), .Y(app_wr_en_n_2_) );
  AND2X2 AND2X2_3789 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo_mem_1__35_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1819) );
  AND2X2 AND2X2_379 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n599), .B(sdram_resetn_bF_buf42), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_11__FF_INPUT) );
  AND2X2 AND2X2_3790 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_0__35_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1820) );
  AND2X2 AND2X2_3791 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1821), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1822) );
  AND2X2 AND2X2_3792 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_2__35_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1823) );
  AND2X2 AND2X2_3793 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_3__35_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1824) );
  AND2X2 AND2X2_3794 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_mem_5__35_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1828) );
  AND2X2 AND2X2_3795 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo_mem_4__35_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1829) );
  AND2X2 AND2X2_3796 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1830), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf0), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1831) );
  AND2X2 AND2X2_3797 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_6__35_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1832) );
  AND2X2 AND2X2_3798 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_7__35_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1834) );
  AND2X2 AND2X2_3799 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1836), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1827), .Y(app_wr_en_n_3_) );
  AND2X2 AND2X2_38 ( .A(u_sdrc_core_b2x_idle), .B(u_sdrc_core_b2r_ack), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n278) );
  AND2X2 AND2X2_380 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_12_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n601) );
  AND2X2 AND2X2_3800 ( .A(u_wb2sdrc_u_wrdatafifo_wr_ptr_1_), .B(u_wb2sdrc_u_wrdatafifo_wr_ptr_2_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1838) );
  AND2X2 AND2X2_3801 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n817_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1838), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839) );
  AND2X2 AND2X2_3802 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1842), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1840), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n767) );
  AND2X2 AND2X2_3803 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1845), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1844), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n768) );
  AND2X2 AND2X2_3804 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1848), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1847), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n769) );
  AND2X2 AND2X2_3805 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1851), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1850), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n770) );
  AND2X2 AND2X2_3806 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1854), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1853), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n771) );
  AND2X2 AND2X2_3807 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1857), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1856), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n772) );
  AND2X2 AND2X2_3808 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1860), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1859), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n773) );
  AND2X2 AND2X2_3809 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1863), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1862), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n774) );
  AND2X2 AND2X2_381 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf1), .B(1'b0), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n602) );
  AND2X2 AND2X2_3810 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1866), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1865), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n775) );
  AND2X2 AND2X2_3811 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1869), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1868), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n776) );
  AND2X2 AND2X2_3812 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1872), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1871), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n777) );
  AND2X2 AND2X2_3813 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1875), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1874), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n778) );
  AND2X2 AND2X2_3814 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1878), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1877), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n779) );
  AND2X2 AND2X2_3815 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1881), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1880), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n780) );
  AND2X2 AND2X2_3816 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1884), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1883), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n781) );
  AND2X2 AND2X2_3817 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1887), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1886), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n782) );
  AND2X2 AND2X2_3818 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1890), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1889), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n783) );
  AND2X2 AND2X2_3819 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1893), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1892), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n784) );
  AND2X2 AND2X2_382 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n603), .B(sdram_resetn_bF_buf41), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_12__FF_INPUT) );
  AND2X2 AND2X2_3820 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1896), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1895), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n785) );
  AND2X2 AND2X2_3821 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1899), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1898), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n786) );
  AND2X2 AND2X2_3822 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1902), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1901), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n787) );
  AND2X2 AND2X2_3823 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1905), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1904), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n788) );
  AND2X2 AND2X2_3824 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1908), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1907), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n789) );
  AND2X2 AND2X2_3825 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1911), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1910), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n790) );
  AND2X2 AND2X2_3826 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1914), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1913), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n791) );
  AND2X2 AND2X2_3827 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1917), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1916), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n792) );
  AND2X2 AND2X2_3828 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1920), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1919), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n793) );
  AND2X2 AND2X2_3829 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1923), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1922), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n794) );
  AND2X2 AND2X2_383 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_4_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_0_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n605) );
  AND2X2 AND2X2_3830 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1926), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1925), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n795) );
  AND2X2 AND2X2_3831 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1929), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1928), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n796) );
  AND2X2 AND2X2_3832 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1932), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1931), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n797) );
  AND2X2 AND2X2_3833 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1935), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1934), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n798) );
  AND2X2 AND2X2_3834 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1938), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1937), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n799) );
  AND2X2 AND2X2_3835 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1941), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1940), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n800) );
  AND2X2 AND2X2_3836 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1944), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1943), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n801) );
  AND2X2 AND2X2_3837 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1947), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1946), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n802) );
  AND2X2 AND2X2_3838 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n818_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1040_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949) );
  AND2X2 AND2X2_3839 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1952), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1950), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n876) );
  AND2X2 AND2X2_384 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_0_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n607) );
  AND2X2 AND2X2_3840 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1955), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1954), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n877) );
  AND2X2 AND2X2_3841 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1958), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1957), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n878) );
  AND2X2 AND2X2_3842 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1961), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1960), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n879) );
  AND2X2 AND2X2_3843 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1964), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1963), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n880) );
  AND2X2 AND2X2_3844 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1967), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1966), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n881) );
  AND2X2 AND2X2_3845 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1970), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1969), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n882) );
  AND2X2 AND2X2_3846 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1973), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1972), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n883) );
  AND2X2 AND2X2_3847 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1976), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1975), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n884) );
  AND2X2 AND2X2_3848 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1979), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1978), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n885) );
  AND2X2 AND2X2_3849 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1982), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1981), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n886) );
  AND2X2 AND2X2_385 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n609), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n610), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_0__FF_INPUT) );
  AND2X2 AND2X2_3850 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1985), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1984), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n887) );
  AND2X2 AND2X2_3851 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1988), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1987), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n888) );
  AND2X2 AND2X2_3852 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1991), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1990), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n889) );
  AND2X2 AND2X2_3853 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1994), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1993), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n890) );
  AND2X2 AND2X2_3854 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1997), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1996), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n891) );
  AND2X2 AND2X2_3855 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2000), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1999), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n892) );
  AND2X2 AND2X2_3856 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2003), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2002), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n893) );
  AND2X2 AND2X2_3857 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2006), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2005), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n894) );
  AND2X2 AND2X2_3858 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2009), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2008), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n895) );
  AND2X2 AND2X2_3859 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2012), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2011), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n896) );
  AND2X2 AND2X2_386 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_4_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_1_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n612) );
  AND2X2 AND2X2_3860 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2015), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2014), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n897) );
  AND2X2 AND2X2_3861 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2018), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2017), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n898) );
  AND2X2 AND2X2_3862 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2021), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2020), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n899) );
  AND2X2 AND2X2_3863 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2024), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2023), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n900) );
  AND2X2 AND2X2_3864 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2027), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2026), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n901) );
  AND2X2 AND2X2_3865 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2030), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2029), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n902) );
  AND2X2 AND2X2_3866 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2033), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2032), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n903) );
  AND2X2 AND2X2_3867 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2036), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2035), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n904) );
  AND2X2 AND2X2_3868 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2039), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2038), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n905) );
  AND2X2 AND2X2_3869 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2042), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2041), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n906) );
  AND2X2 AND2X2_387 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_1_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n613) );
  AND2X2 AND2X2_3870 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2045), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2044), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n907) );
  AND2X2 AND2X2_3871 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2048), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2047), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n908) );
  AND2X2 AND2X2_3872 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2051), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2050), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n909) );
  AND2X2 AND2X2_3873 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2054), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2053), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n910) );
  AND2X2 AND2X2_3874 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2057), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2056), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n911) );
  AND2X2 AND2X2_3875 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n817_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1041_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059) );
  AND2X2 AND2X2_3876 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2062), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2060), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n914) );
  AND2X2 AND2X2_3877 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2065), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2064), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n916) );
  AND2X2 AND2X2_3878 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2068), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2067), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n918) );
  AND2X2 AND2X2_3879 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2071), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2070), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n920) );
  AND2X2 AND2X2_388 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n615), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n616), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_1__FF_INPUT) );
  AND2X2 AND2X2_3880 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2074), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2073), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n922) );
  AND2X2 AND2X2_3881 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2077), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2076), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n924) );
  AND2X2 AND2X2_3882 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2080), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2079), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n926) );
  AND2X2 AND2X2_3883 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2083), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2082), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n928) );
  AND2X2 AND2X2_3884 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2086), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2085), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n930) );
  AND2X2 AND2X2_3885 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2089), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2088), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n932) );
  AND2X2 AND2X2_3886 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2092), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2091), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n934) );
  AND2X2 AND2X2_3887 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2095), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2094), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n936) );
  AND2X2 AND2X2_3888 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2098), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2097), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n938) );
  AND2X2 AND2X2_3889 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2101), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2100), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n940) );
  AND2X2 AND2X2_389 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_4_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_2_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n618) );
  AND2X2 AND2X2_3890 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2104), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2103), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n942) );
  AND2X2 AND2X2_3891 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2107), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2106), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n944) );
  AND2X2 AND2X2_3892 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2110), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2109), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n946) );
  AND2X2 AND2X2_3893 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2113), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2112), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n948) );
  AND2X2 AND2X2_3894 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2116), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2115), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n950) );
  AND2X2 AND2X2_3895 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2119), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2118), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n952) );
  AND2X2 AND2X2_3896 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2122), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2121), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n954) );
  AND2X2 AND2X2_3897 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2125), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2124), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n956) );
  AND2X2 AND2X2_3898 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2128), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2127), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n958) );
  AND2X2 AND2X2_3899 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2131), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2130), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n960) );
  AND2X2 AND2X2_39 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n255), .B(u_sdrc_core_u_bank_ctl__abc_21249_n216_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n280_1) );
  AND2X2 AND2X2_390 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_2_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n619) );
  AND2X2 AND2X2_3900 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2134), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2133), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n962) );
  AND2X2 AND2X2_3901 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2137), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2136), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n964) );
  AND2X2 AND2X2_3902 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2140), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2139), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n966) );
  AND2X2 AND2X2_3903 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2143), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2142), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n968) );
  AND2X2 AND2X2_3904 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2146), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2145), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n970) );
  AND2X2 AND2X2_3905 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2149), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2148), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n972) );
  AND2X2 AND2X2_3906 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2152), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2151), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n974) );
  AND2X2 AND2X2_3907 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2155), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2154), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n976) );
  AND2X2 AND2X2_3908 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2158), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2157), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n978) );
  AND2X2 AND2X2_3909 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2161), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2160), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n980) );
  AND2X2 AND2X2_391 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n621), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n622), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_2__FF_INPUT) );
  AND2X2 AND2X2_3910 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2164), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2163), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n982) );
  AND2X2 AND2X2_3911 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2167), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2166), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n984) );
  AND2X2 AND2X2_3912 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n929_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1040_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169) );
  AND2X2 AND2X2_3913 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2172), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2170), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n986) );
  AND2X2 AND2X2_3914 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2175), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2174), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n987) );
  AND2X2 AND2X2_3915 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2178), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2177), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n988) );
  AND2X2 AND2X2_3916 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2181), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2180), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n989) );
  AND2X2 AND2X2_3917 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2184), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2183), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n990) );
  AND2X2 AND2X2_3918 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2187), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2186), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n991) );
  AND2X2 AND2X2_3919 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2190), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2189), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n992) );
  AND2X2 AND2X2_392 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_4_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_3_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n624) );
  AND2X2 AND2X2_3920 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2193), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2192), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n993) );
  AND2X2 AND2X2_3921 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2196), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2195), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n994) );
  AND2X2 AND2X2_3922 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2199), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2198), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n995) );
  AND2X2 AND2X2_3923 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2202), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2201), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n996) );
  AND2X2 AND2X2_3924 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2205), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2204), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n997) );
  AND2X2 AND2X2_3925 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2208), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2207), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n998) );
  AND2X2 AND2X2_3926 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2211), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2210), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n999) );
  AND2X2 AND2X2_3927 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2214), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2213), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1000) );
  AND2X2 AND2X2_3928 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2217), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2216), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1001) );
  AND2X2 AND2X2_3929 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2220), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2219), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1002) );
  AND2X2 AND2X2_393 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_3_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n625) );
  AND2X2 AND2X2_3930 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2223), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2222), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1003) );
  AND2X2 AND2X2_3931 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2226), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2225), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1004) );
  AND2X2 AND2X2_3932 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2229), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2228), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1005) );
  AND2X2 AND2X2_3933 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2232), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2231), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1006) );
  AND2X2 AND2X2_3934 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2235), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2234), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1007) );
  AND2X2 AND2X2_3935 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2238), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2237), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1008) );
  AND2X2 AND2X2_3936 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2241), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2240), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1009) );
  AND2X2 AND2X2_3937 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2244), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2243), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1010) );
  AND2X2 AND2X2_3938 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2247), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2246), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1011) );
  AND2X2 AND2X2_3939 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2250), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2249), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1012) );
  AND2X2 AND2X2_394 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n627), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n628), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_3__FF_INPUT) );
  AND2X2 AND2X2_3940 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2253), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2252), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1013) );
  AND2X2 AND2X2_3941 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2256), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2255), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1014) );
  AND2X2 AND2X2_3942 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2259), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2258), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1015) );
  AND2X2 AND2X2_3943 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2262), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2261), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1016) );
  AND2X2 AND2X2_3944 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2265), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2264), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1017) );
  AND2X2 AND2X2_3945 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2268), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2267), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1018) );
  AND2X2 AND2X2_3946 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2271), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2270), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1019) );
  AND2X2 AND2X2_3947 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2274), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2273), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1020) );
  AND2X2 AND2X2_3948 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2277), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2276), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1021) );
  AND2X2 AND2X2_3949 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2279), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf5), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2280) );
  AND2X2 AND2X2_395 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_4_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_4_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n630) );
  AND2X2 AND2X2_3950 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf6), .B(app_wr_next_req), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2281) );
  AND2X2 AND2X2_3951 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2279), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_1_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2283) );
  AND2X2 AND2X2_3952 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf7), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf5), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2284) );
  AND2X2 AND2X2_3953 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2279), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf4), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2289) );
  AND2X2 AND2X2_3954 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf6), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf3), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2290) );
  AND2X2 AND2X2_3955 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2291), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2292), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2293) );
  AND2X2 AND2X2_3956 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2293), .B(app_wr_next_req), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2294) );
  AND2X2 AND2X2_3957 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2279), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_3_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2296) );
  AND2X2 AND2X2_3958 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2291), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_3_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2297) );
  AND2X2 AND2X2_3959 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2290), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n792_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2298) );
  AND2X2 AND2X2_396 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_4_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n631) );
  AND2X2 AND2X2_3960 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2299), .B(app_wr_next_req), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2300) );
  AND2X2 AND2X2_3961 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf6), .B(app_wr_next_req), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2302) );
  AND2X2 AND2X2_3962 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2279), .B(u_wb2sdrc_u_wrdatafifo_grey_rd_ptr_0_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2303) );
  AND2X2 AND2X2_3963 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2294), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2286), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2305) );
  AND2X2 AND2X2_3964 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2279), .B(u_wb2sdrc_u_wrdatafifo_grey_rd_ptr_1_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2306) );
  AND2X2 AND2X2_3965 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2287), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf5), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2307) );
  AND2X2 AND2X2_3966 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2300), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2310), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2311) );
  AND2X2 AND2X2_3967 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2279), .B(u_wb2sdrc_u_wrdatafifo_grey_rd_ptr_2_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2312) );
  AND2X2 AND2X2_3968 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2294), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n792_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2313) );
  AND2X2 AND2X2_3969 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2279), .B(u_wb2sdrc_u_wrdatafifo_grey_rd_ptr_3_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2316) );
  AND2X2 AND2X2_397 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n633), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n634), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_4__FF_INPUT) );
  AND2X2 AND2X2_3970 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2318), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2320), .Y(u_wb2sdrc_u_wrdatafifo_full_q_FF_INPUT) );
  AND2X2 AND2X2_3971 ( .A(u_wb2sdrc_u_wrdatafifo_wr_ptr_0_), .B(u_wb2sdrc_u_wrdatafifo_wr_ptr_1_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2326) );
  AND2X2 AND2X2_3972 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2326), .B(u_wb2sdrc_u_wrdatafifo_wr_ptr_2_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2328) );
  AND2X2 AND2X2_3973 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2329), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2327), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2330) );
  AND2X2 AND2X2_3974 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2330), .B(u_wb2sdrc_u_wrdatafifo_wr_en), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2331) );
  AND2X2 AND2X2_3975 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n738_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n743), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2332) );
  AND2X2 AND2X2_3976 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2328), .B(u_wb2sdrc_u_wrdatafifo_wr_ptr_3_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2342) );
  AND2X2 AND2X2_3977 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2344), .B(u_wb2sdrc_u_wrdatafifo_wr_en), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2345) );
  AND2X2 AND2X2_3978 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2345), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2343), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2346) );
  AND2X2 AND2X2_3979 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2323), .B(u_wb2sdrc_u_wrdatafifo_wr_ptr_0_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2354) );
  AND2X2 AND2X2_398 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_4_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_5_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n636) );
  AND2X2 AND2X2_3980 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2323), .B(u_wb2sdrc_u_wrdatafifo_wr_ptr_1_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2356) );
  AND2X2 AND2X2_3981 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2323), .B(u_wb2sdrc_u_wrdatafifo_wr_ptr_2_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2358) );
  AND2X2 AND2X2_3982 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2323), .B(u_wb2sdrc_u_wrdatafifo_wr_ptr_3_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2360) );
  AND2X2 AND2X2_3983 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1040_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1838), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362) );
  AND2X2 AND2X2_3984 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_7__0_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2364) );
  AND2X2 AND2X2_3985 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf4), .B(\wb_dat_i[0] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2365) );
  AND2X2 AND2X2_3986 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_7__1_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2367) );
  AND2X2 AND2X2_3987 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf3), .B(\wb_dat_i[1] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2368) );
  AND2X2 AND2X2_3988 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_7__2_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2370) );
  AND2X2 AND2X2_3989 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf2), .B(\wb_dat_i[2] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2371) );
  AND2X2 AND2X2_399 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_5_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n637) );
  AND2X2 AND2X2_3990 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_7__3_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2373) );
  AND2X2 AND2X2_3991 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf1), .B(\wb_dat_i[3] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2374) );
  AND2X2 AND2X2_3992 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_7__4_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2376) );
  AND2X2 AND2X2_3993 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf0), .B(\wb_dat_i[4] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2377) );
  AND2X2 AND2X2_3994 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_7__5_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2379) );
  AND2X2 AND2X2_3995 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf5), .B(\wb_dat_i[5] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2380) );
  AND2X2 AND2X2_3996 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_7__6_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2382) );
  AND2X2 AND2X2_3997 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf4), .B(\wb_dat_i[6] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2383) );
  AND2X2 AND2X2_3998 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_7__7_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2385) );
  AND2X2 AND2X2_3999 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf3), .B(\wb_dat_i[7] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2386) );
  AND2X2 AND2X2_4 ( .A(u_sdrc_core_b2x_ba_1_), .B(u_sdrc_core_b2x_ba_0_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok) );
  AND2X2 AND2X2_40 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n223_1_bF_buf2), .B(u_sdrc_core_u_bank_ctl__abc_21249_n284_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n285) );
  AND2X2 AND2X2_400 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n639), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n640), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_5__FF_INPUT) );
  AND2X2 AND2X2_4000 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_7__8_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2388) );
  AND2X2 AND2X2_4001 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf2), .B(\wb_dat_i[8] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2389) );
  AND2X2 AND2X2_4002 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_7__9_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2391) );
  AND2X2 AND2X2_4003 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf1), .B(\wb_dat_i[9] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2392) );
  AND2X2 AND2X2_4004 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_7__10_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2394) );
  AND2X2 AND2X2_4005 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf0), .B(\wb_dat_i[10] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2395) );
  AND2X2 AND2X2_4006 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_7__11_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2397) );
  AND2X2 AND2X2_4007 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf5), .B(\wb_dat_i[11] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2398) );
  AND2X2 AND2X2_4008 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_7__12_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2400) );
  AND2X2 AND2X2_4009 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf4), .B(\wb_dat_i[12] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2401) );
  AND2X2 AND2X2_401 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_4_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_6_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n642) );
  AND2X2 AND2X2_4010 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_7__13_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2403) );
  AND2X2 AND2X2_4011 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf3), .B(\wb_dat_i[13] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2404) );
  AND2X2 AND2X2_4012 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_7__14_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2406) );
  AND2X2 AND2X2_4013 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf2), .B(\wb_dat_i[14] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2407) );
  AND2X2 AND2X2_4014 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_7__15_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2409) );
  AND2X2 AND2X2_4015 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf1), .B(\wb_dat_i[15] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2410) );
  AND2X2 AND2X2_4016 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_7__16_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2412) );
  AND2X2 AND2X2_4017 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf0), .B(\wb_dat_i[16] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2413) );
  AND2X2 AND2X2_4018 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_7__17_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2415) );
  AND2X2 AND2X2_4019 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf5), .B(\wb_dat_i[17] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2416) );
  AND2X2 AND2X2_402 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_6_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n643) );
  AND2X2 AND2X2_4020 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_7__18_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2418) );
  AND2X2 AND2X2_4021 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf4), .B(\wb_dat_i[18] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2419) );
  AND2X2 AND2X2_4022 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_7__19_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2421) );
  AND2X2 AND2X2_4023 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf3), .B(\wb_dat_i[19] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2422) );
  AND2X2 AND2X2_4024 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_7__20_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2424) );
  AND2X2 AND2X2_4025 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf2), .B(\wb_dat_i[20] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2425) );
  AND2X2 AND2X2_4026 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_7__21_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2427) );
  AND2X2 AND2X2_4027 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf1), .B(\wb_dat_i[21] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2428) );
  AND2X2 AND2X2_4028 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_7__22_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2430) );
  AND2X2 AND2X2_4029 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf0), .B(\wb_dat_i[22] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2431) );
  AND2X2 AND2X2_403 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n645), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n646), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_6__FF_INPUT) );
  AND2X2 AND2X2_4030 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_7__23_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2433) );
  AND2X2 AND2X2_4031 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf5), .B(\wb_dat_i[23] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2434) );
  AND2X2 AND2X2_4032 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_7__24_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2436) );
  AND2X2 AND2X2_4033 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf4), .B(\wb_dat_i[24] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2437) );
  AND2X2 AND2X2_4034 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_7__25_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2439) );
  AND2X2 AND2X2_4035 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf3), .B(\wb_dat_i[25] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2440) );
  AND2X2 AND2X2_4036 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_7__26_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2442) );
  AND2X2 AND2X2_4037 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf2), .B(\wb_dat_i[26] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2443) );
  AND2X2 AND2X2_4038 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_7__27_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2445) );
  AND2X2 AND2X2_4039 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf1), .B(\wb_dat_i[27] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2446) );
  AND2X2 AND2X2_404 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_4_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_7_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n648) );
  AND2X2 AND2X2_4040 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_7__28_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2448) );
  AND2X2 AND2X2_4041 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf0), .B(\wb_dat_i[28] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2449) );
  AND2X2 AND2X2_4042 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_7__29_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2451) );
  AND2X2 AND2X2_4043 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf5), .B(\wb_dat_i[29] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2452) );
  AND2X2 AND2X2_4044 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_7__30_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2454) );
  AND2X2 AND2X2_4045 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf4), .B(\wb_dat_i[30] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2455) );
  AND2X2 AND2X2_4046 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_7__31_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2457) );
  AND2X2 AND2X2_4047 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf3), .B(\wb_dat_i[31] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2458) );
  AND2X2 AND2X2_4048 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_7__32_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2460) );
  AND2X2 AND2X2_4049 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_wr_data_32_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2461) );
  AND2X2 AND2X2_405 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_7_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n649) );
  AND2X2 AND2X2_4050 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_7__33_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2463) );
  AND2X2 AND2X2_4051 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_wr_data_33_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2464) );
  AND2X2 AND2X2_4052 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_7__34_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2466) );
  AND2X2 AND2X2_4053 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_wr_data_34_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2467) );
  AND2X2 AND2X2_4054 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_7__35_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2469) );
  AND2X2 AND2X2_4055 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_wr_data_35_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2470) );
  AND2X2 AND2X2_406 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n651), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n652), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_7__FF_INPUT) );
  AND2X2 AND2X2_407 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_4_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_8_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n654) );
  AND2X2 AND2X2_408 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_8_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n655) );
  AND2X2 AND2X2_409 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n657), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n658), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_8__FF_INPUT) );
  AND2X2 AND2X2_41 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf2), .B(u_sdrc_core_u_bank_ctl__abc_21249_n286_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n287_1) );
  AND2X2 AND2X2_410 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_4_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_9_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n660) );
  AND2X2 AND2X2_411 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_9_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n661) );
  AND2X2 AND2X2_412 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n663), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n664), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_9__FF_INPUT) );
  AND2X2 AND2X2_413 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_4_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_10_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n666) );
  AND2X2 AND2X2_414 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n370), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_10_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n667) );
  AND2X2 AND2X2_415 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n669), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n670), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_10__FF_INPUT) );
  AND2X2 AND2X2_416 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_4_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_11_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n672) );
  AND2X2 AND2X2_417 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_11_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n673) );
  AND2X2 AND2X2_418 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n675), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n676), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_11__FF_INPUT) );
  AND2X2 AND2X2_419 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_4_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_12_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n678) );
  AND2X2 AND2X2_42 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n288_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n283_bF_buf3), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n289_1) );
  AND2X2 AND2X2_420 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n370), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_12_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n679) );
  AND2X2 AND2X2_421 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n681), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n682), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_12__FF_INPUT) );
  AND2X2 AND2X2_422 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n689), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n688), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_last) );
  AND2X2 AND2X2_423 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n704), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n703), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_len_0_) );
  AND2X2 AND2X2_424 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n707), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n706), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_len_1_) );
  AND2X2 AND2X2_425 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n710), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n709), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_len_2_) );
  AND2X2 AND2X2_426 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n713), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n712), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_len_3_) );
  AND2X2 AND2X2_427 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n716), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n715), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_len_4_) );
  AND2X2 AND2X2_428 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n719), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n718), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_len_5_) );
  AND2X2 AND2X2_429 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n722), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n721), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_len_6_) );
  AND2X2 AND2X2_43 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n291_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n282_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n292_1) );
  AND2X2 AND2X2_430 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n725), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n724), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_wrap) );
  AND2X2 AND2X2_431 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_pre_ok_t), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_tras_ok), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n727) );
  AND2X2 AND2X2_432 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n368_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n727), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n728) );
  AND2X2 AND2X2_433 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_2_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_act_ok_t), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n729) );
  AND2X2 AND2X2_434 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_4_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_xfr_ok_r), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n733) );
  AND2X2 AND2X2_435 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n732), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n733), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n734) );
  AND2X2 AND2X2_436 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n734), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n731), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n735) );
  AND2X2 AND2X2_437 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n736), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_timer0_tc), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n737) );
  AND2X2 AND2X2_438 ( .A(sdram_resetn_bF_buf40), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_wrok), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_wrok_r_FF_INPUT) );
  AND2X2 AND2X2_439 ( .A(sdram_resetn_bF_buf39), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_xfr_ok), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_xfr_ok_r_FF_INPUT) );
  AND2X2 AND2X2_44 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n296_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n279_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n297) );
  AND2X2 AND2X2_440 ( .A(sdram_resetn_bF_buf38), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_rdok), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_rdok_r_FF_INPUT) );
  AND2X2 AND2X2_441 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n380), .B(sdram_resetn_bF_buf37), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n743) );
  AND2X2 AND2X2_442 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n742), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n743), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_timer0_tc_r_FF_INPUT) );
  AND2X2 AND2X2_443 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n745), .B(sdram_resetn_bF_buf36), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_tras_ok_r_FF_INPUT) );
  AND2X2 AND2X2_444 ( .A(sdram_resetn_bF_buf35), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_pre_ok), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_pre_ok_r_FF_INPUT) );
  AND2X2 AND2X2_445 ( .A(sdram_resetn_bF_buf34), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_act_ok), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_act_ok_r_FF_INPUT) );
  AND2X2 AND2X2_446 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n357), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n336), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n750) );
  AND2X2 AND2X2_447 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n749), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n750), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_valid_FF_INPUT) );
  AND2X2 AND2X2_448 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_last), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n756) );
  AND2X2 AND2X2_449 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf0), .B(u_sdrc_core_r2b_last), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n757) );
  AND2X2 AND2X2_45 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n241), .B(u_sdrc_core_u_bank_ctl_rank_ba_2_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n298_1) );
  AND2X2 AND2X2_450 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n758), .B(sdram_resetn_bF_buf33), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_l_last_FF_INPUT) );
  AND2X2 AND2X2_451 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_wrap), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n760) );
  AND2X2 AND2X2_452 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf4), .B(u_sdrc_core_r2b_wrap), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n761) );
  AND2X2 AND2X2_453 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n762), .B(sdram_resetn_bF_buf32), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_l_wrap_FF_INPUT) );
  AND2X2 AND2X2_454 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_write), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n764) );
  AND2X2 AND2X2_455 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf3), .B(u_sdrc_core_r2b_write), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n765) );
  AND2X2 AND2X2_456 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n766), .B(sdram_resetn_bF_buf31), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_l_write_FF_INPUT) );
  AND2X2 AND2X2_457 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf5), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_sdr_dma_last), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n768) );
  AND2X2 AND2X2_458 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf2), .B(1'b0), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n769) );
  AND2X2 AND2X2_459 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n770), .B(sdram_resetn_bF_buf30), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_l_sdr_dma_last_FF_INPUT) );
  AND2X2 AND2X2_46 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n294_1), .B(u_sdrc_core_b2x_ba_0_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n299_1) );
  AND2X2 AND2X2_460 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n249_1), .B(sdram_resetn_bF_buf29), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n250_1) );
  AND2X2 AND2X2_461 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n250_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_3_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n251) );
  AND2X2 AND2X2_462 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_r2b_req), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_0_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack) );
  AND2X2 AND2X2_463 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf3), .B(sdram_resetn_bF_buf28), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n253_1) );
  AND2X2 AND2X2_464 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n257), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n259_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n260) );
  AND2X2 AND2X2_465 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n260), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n255_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n261_1) );
  AND2X2 AND2X2_466 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n263), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n265_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n266) );
  AND2X2 AND2X2_467 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n268_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n270_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n271_1) );
  AND2X2 AND2X2_468 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n266), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n271_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n272) );
  AND2X2 AND2X2_469 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n272), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n261_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n273_1) );
  AND2X2 AND2X2_47 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n297), .B(u_sdrc_core_u_bank_ctl__abc_21249_n300), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n301_1) );
  AND2X2 AND2X2_470 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n275), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n277_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n278) );
  AND2X2 AND2X2_471 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n280_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n282_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n283_1) );
  AND2X2 AND2X2_472 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n278), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n283_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n284_1) );
  AND2X2 AND2X2_473 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n286_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n288_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n289) );
  AND2X2 AND2X2_474 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n291_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n293), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n294_1) );
  AND2X2 AND2X2_475 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n289), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n294_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n295_1) );
  AND2X2 AND2X2_476 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n284_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n295_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n296_1) );
  AND2X2 AND2X2_477 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n296_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n273_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n297) );
  AND2X2 AND2X2_478 ( .A(u_sdrc_core_r2b_raddr_10_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_10_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n298_1) );
  AND2X2 AND2X2_479 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n299_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n300_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n301) );
  AND2X2 AND2X2_48 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n241), .B(u_sdrc_core_b2r_ack), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n302_1) );
  AND2X2 AND2X2_480 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_8_), .B(u_sdrc_core_r2b_raddr_8_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n303_1) );
  AND2X2 AND2X2_481 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n304_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n305), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n306_1) );
  AND2X2 AND2X2_482 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n302_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n307_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n308_1) );
  AND2X2 AND2X2_483 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n310_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n312_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n313) );
  AND2X2 AND2X2_484 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n315_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n317), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n318_1) );
  AND2X2 AND2X2_485 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n313), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n318_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n319_1) );
  AND2X2 AND2X2_486 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n321), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n323_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n324_1) );
  AND2X2 AND2X2_487 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n326_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_valid), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n327_1) );
  AND2X2 AND2X2_488 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n324_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n327_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n328_1) );
  AND2X2 AND2X2_489 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n319_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n328_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n329) );
  AND2X2 AND2X2_49 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n302_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n280_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n303_1) );
  AND2X2 AND2X2_490 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n329), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n308_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n330_1) );
  AND2X2 AND2X2_491 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n297), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n330_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n331_1) );
  AND2X2 AND2X2_492 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n332_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n253_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n333) );
  AND2X2 AND2X2_493 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n250_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_prech_page_closed), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n335) );
  AND2X2 AND2X2_494 ( .A(sdram_resetn_bF_buf27), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_4_bF_buf3), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n337) );
  AND2X2 AND2X2_495 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n337), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n336), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n338_1) );
  AND2X2 AND2X2_496 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n338_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_x2b_ack), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n339_1) );
  AND2X2 AND2X2_497 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n339_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_sdr_dma_last), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n340) );
  AND2X2 AND2X2_498 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n250_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_2_bF_buf3), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n342) );
  AND2X2 AND2X2_499 ( .A(sdram_resetn_bF_buf26), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_x2b_ack), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n343_1) );
  AND2X2 AND2X2_5 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n211_1), .B(u_sdrc_core_b2x_ba_1_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok) );
  AND2X2 AND2X2_50 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n304), .B(u_sdrc_core_r2b_ba_0_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n305_1) );
  AND2X2 AND2X2_500 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n343_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_3_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n344_1) );
  AND2X2 AND2X2_501 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n337), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_refresh), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n345) );
  AND2X2 AND2X2_502 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n343_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_2_bF_buf2), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n348_1) );
  AND2X2 AND2X2_503 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n338_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n249_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n349_1) );
  AND2X2 AND2X2_504 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n331_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n253_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n351) );
  AND2X2 AND2X2_505 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n339_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n353_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n354_1) );
  AND2X2 AND2X2_506 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n356), .B(sdram_resetn_bF_buf25), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n357) );
  AND2X2 AND2X2_507 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n355), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n358_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n359_1) );
  AND2X2 AND2X2_508 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n360), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_0_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n361) );
  AND2X2 AND2X2_509 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_4_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_write), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n364_1) );
  AND2X2 AND2X2_51 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n306_1), .B(sdram_resetn_bF_buf46), .Y(u_sdrc_core_u_bank_ctl_rank_ba_0__FF_INPUT) );
  AND2X2 AND2X2_510 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n369_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n367), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n370) );
  AND2X2 AND2X2_511 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n370), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n371) );
  AND2X2 AND2X2_512 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n371), .B(u_sdrc_core_r2b_write), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n372) );
  AND2X2 AND2X2_513 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n331_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n372), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n373_1) );
  AND2X2 AND2X2_514 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n374_1), .B(sdram_resetn_bF_buf24), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_cmd_r_0__FF_INPUT) );
  AND2X2 AND2X2_515 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n371), .B(sdram_resetn_bF_buf23), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n376) );
  AND2X2 AND2X2_516 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n331_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n376), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n377) );
  AND2X2 AND2X2_517 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n381), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_cmd_0_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n382) );
  AND2X2 AND2X2_518 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n383_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n386_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n387_1) );
  AND2X2 AND2X2_519 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n387_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n379_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n388) );
  AND2X2 AND2X2_52 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n241), .B(u_sdrc_core_u_bank_ctl_rank_ba_3_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n308_1) );
  AND2X2 AND2X2_520 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n382), .B(\cfg_sdr_tras_d[0] ), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n389) );
  AND2X2 AND2X2_521 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n390), .B(sdram_resetn_bF_buf22), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_tras_cntr_0__FF_INPUT) );
  AND2X2 AND2X2_522 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n382), .B(\cfg_sdr_tras_d[1] ), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n392_1) );
  AND2X2 AND2X2_523 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_tras_cntr_0_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_tras_cntr_1_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n394_1) );
  AND2X2 AND2X2_524 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n387_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n395_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n396_1) );
  AND2X2 AND2X2_525 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n397_1), .B(sdram_resetn_bF_buf21), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_tras_cntr_1__FF_INPUT) );
  AND2X2 AND2X2_526 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n382), .B(\cfg_sdr_tras_d[2] ), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n399_1) );
  AND2X2 AND2X2_527 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n384_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_tras_cntr_2_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n401_1) );
  AND2X2 AND2X2_528 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n387_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n402_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n403_1) );
  AND2X2 AND2X2_529 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n404_1), .B(sdram_resetn_bF_buf20), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_tras_cntr_2__FF_INPUT) );
  AND2X2 AND2X2_53 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n294_1), .B(u_sdrc_core_b2x_ba_1_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n309_1) );
  AND2X2 AND2X2_530 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n385), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_tras_cntr_3_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n406_1) );
  AND2X2 AND2X2_531 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n408_1), .B(sdram_resetn_bF_buf19), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n409_1) );
  AND2X2 AND2X2_532 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n409_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n407_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_tras_cntr_3__FF_INPUT) );
  AND2X2 AND2X2_533 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n415_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n413_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n416) );
  AND2X2 AND2X2_534 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n417_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n418), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n419_1) );
  AND2X2 AND2X2_535 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n421), .B(sdram_resetn_bF_buf18), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n422) );
  AND2X2 AND2X2_536 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n420_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n422), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_timer0_0__FF_INPUT) );
  AND2X2 AND2X2_537 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_timer0_1_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_timer0_0_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n426) );
  AND2X2 AND2X2_538 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n383_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n428_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n429) );
  AND2X2 AND2X2_539 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n429), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n427_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n430) );
  AND2X2 AND2X2_54 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n297), .B(u_sdrc_core_u_bank_ctl__abc_21249_n310), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n311_1) );
  AND2X2 AND2X2_540 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n381), .B(\cfg_sdr_trcd_d[1] ), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n431_1) );
  AND2X2 AND2X2_541 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n434_1), .B(sdram_resetn_bF_buf17), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n435_1) );
  AND2X2 AND2X2_542 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n433), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n435_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_timer0_1__FF_INPUT) );
  AND2X2 AND2X2_543 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n424), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_timer0_2_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n439_1) );
  AND2X2 AND2X2_544 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n429), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n440_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n441) );
  AND2X2 AND2X2_545 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n381), .B(\cfg_sdr_trcd_d[2] ), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n442) );
  AND2X2 AND2X2_546 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n445_1), .B(sdram_resetn_bF_buf16), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n446_1) );
  AND2X2 AND2X2_547 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n444_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n446_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_timer0_2__FF_INPUT) );
  AND2X2 AND2X2_548 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n437_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_timer0_3_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n448_1) );
  AND2X2 AND2X2_549 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n449_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n450), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n451) );
  AND2X2 AND2X2_55 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n304), .B(u_sdrc_core_r2b_ba_1_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n312) );
  AND2X2 AND2X2_550 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n453_1), .B(sdram_resetn_bF_buf15), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n454) );
  AND2X2 AND2X2_551 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n452), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n454), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_timer0_3__FF_INPUT) );
  AND2X2 AND2X2_552 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n253_1), .B(u_sdrc_core_r2b_len_0_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n473) );
  AND2X2 AND2X2_553 ( .A(sdram_resetn_bF_buf14), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_0_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n474) );
  AND2X2 AND2X2_554 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf5), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n474), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n475) );
  AND2X2 AND2X2_555 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n253_1), .B(u_sdrc_core_r2b_len_1_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n477) );
  AND2X2 AND2X2_556 ( .A(sdram_resetn_bF_buf13), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_1_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n478) );
  AND2X2 AND2X2_557 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n478), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n479) );
  AND2X2 AND2X2_558 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n253_1), .B(u_sdrc_core_r2b_len_2_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n481) );
  AND2X2 AND2X2_559 ( .A(sdram_resetn_bF_buf12), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_2_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n482) );
  AND2X2 AND2X2_56 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n313_1), .B(sdram_resetn_bF_buf45), .Y(u_sdrc_core_u_bank_ctl_rank_ba_1__FF_INPUT) );
  AND2X2 AND2X2_560 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n482), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n483) );
  AND2X2 AND2X2_561 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n253_1), .B(u_sdrc_core_r2b_len_3_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n485) );
  AND2X2 AND2X2_562 ( .A(sdram_resetn_bF_buf11), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_3_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n486) );
  AND2X2 AND2X2_563 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n486), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n487) );
  AND2X2 AND2X2_564 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n253_1), .B(u_sdrc_core_r2b_len_4_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n489) );
  AND2X2 AND2X2_565 ( .A(sdram_resetn_bF_buf10), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_4_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n490) );
  AND2X2 AND2X2_566 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n490), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n491) );
  AND2X2 AND2X2_567 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n253_1), .B(u_sdrc_core_r2b_len_5_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n493) );
  AND2X2 AND2X2_568 ( .A(sdram_resetn_bF_buf9), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_5_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n494) );
  AND2X2 AND2X2_569 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n494), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n495) );
  AND2X2 AND2X2_57 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n253_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n216_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n315) );
  AND2X2 AND2X2_570 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n253_1), .B(u_sdrc_core_r2b_len_6_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n497) );
  AND2X2 AND2X2_571 ( .A(sdram_resetn_bF_buf8), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_6_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n498) );
  AND2X2 AND2X2_572 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf5), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n498), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n499) );
  AND2X2 AND2X2_573 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_0_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n501) );
  AND2X2 AND2X2_574 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf1), .B(u_sdrc_core_r2b_raddr_0_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n502) );
  AND2X2 AND2X2_575 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n503), .B(sdram_resetn_bF_buf7), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_0__FF_INPUT) );
  AND2X2 AND2X2_576 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_1_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n505) );
  AND2X2 AND2X2_577 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf0), .B(u_sdrc_core_r2b_raddr_1_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n506) );
  AND2X2 AND2X2_578 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n507), .B(sdram_resetn_bF_buf6), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_1__FF_INPUT) );
  AND2X2 AND2X2_579 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_2_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n509) );
  AND2X2 AND2X2_58 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n317_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n318), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n319) );
  AND2X2 AND2X2_580 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf4), .B(u_sdrc_core_r2b_raddr_2_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n510) );
  AND2X2 AND2X2_581 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n511), .B(sdram_resetn_bF_buf5), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_2__FF_INPUT) );
  AND2X2 AND2X2_582 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_3_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n513) );
  AND2X2 AND2X2_583 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf3), .B(u_sdrc_core_r2b_raddr_3_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n514) );
  AND2X2 AND2X2_584 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n515), .B(sdram_resetn_bF_buf4), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_3__FF_INPUT) );
  AND2X2 AND2X2_585 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_4_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n517) );
  AND2X2 AND2X2_586 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf2), .B(u_sdrc_core_r2b_raddr_4_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n518) );
  AND2X2 AND2X2_587 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n519), .B(sdram_resetn_bF_buf3), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_4__FF_INPUT) );
  AND2X2 AND2X2_588 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf5), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_5_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n521) );
  AND2X2 AND2X2_589 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf1), .B(u_sdrc_core_r2b_raddr_5_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n522) );
  AND2X2 AND2X2_59 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n241), .B(u_sdrc_core_u_bank_ctl_rank_ba_4_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n321) );
  AND2X2 AND2X2_590 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n523), .B(sdram_resetn_bF_buf2), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_5__FF_INPUT) );
  AND2X2 AND2X2_591 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_6_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n525) );
  AND2X2 AND2X2_592 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf0), .B(u_sdrc_core_r2b_raddr_6_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n526) );
  AND2X2 AND2X2_593 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n527), .B(sdram_resetn_bF_buf1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_6__FF_INPUT) );
  AND2X2 AND2X2_594 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_7_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n529) );
  AND2X2 AND2X2_595 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf4), .B(u_sdrc_core_r2b_raddr_7_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n530) );
  AND2X2 AND2X2_596 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n531), .B(sdram_resetn_bF_buf0), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_7__FF_INPUT) );
  AND2X2 AND2X2_597 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_8_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n533) );
  AND2X2 AND2X2_598 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf3), .B(u_sdrc_core_r2b_raddr_8_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n534) );
  AND2X2 AND2X2_599 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n535), .B(sdram_resetn_bF_buf49), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_8__FF_INPUT) );
  AND2X2 AND2X2_6 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n213), .B(u_sdrc_core_b2x_ba_0_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok) );
  AND2X2 AND2X2_60 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n294_1), .B(u_sdrc_core_u_bank_ctl_rank_ba_2_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n322_1) );
  AND2X2 AND2X2_600 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_9_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n537) );
  AND2X2 AND2X2_601 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf2), .B(u_sdrc_core_r2b_raddr_9_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n538) );
  AND2X2 AND2X2_602 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n539), .B(sdram_resetn_bF_buf48), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_9__FF_INPUT) );
  AND2X2 AND2X2_603 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_10_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n541) );
  AND2X2 AND2X2_604 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf1), .B(u_sdrc_core_r2b_raddr_10_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n542) );
  AND2X2 AND2X2_605 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n543), .B(sdram_resetn_bF_buf47), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_10__FF_INPUT) );
  AND2X2 AND2X2_606 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf5), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_11_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n545) );
  AND2X2 AND2X2_607 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf0), .B(u_sdrc_core_r2b_raddr_11_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n546) );
  AND2X2 AND2X2_608 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n547), .B(sdram_resetn_bF_buf46), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_11__FF_INPUT) );
  AND2X2 AND2X2_609 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_12_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n549) );
  AND2X2 AND2X2_61 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n325_1), .B(sdram_resetn_bF_buf44), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n326_1) );
  AND2X2 AND2X2_610 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf4), .B(u_sdrc_core_r2b_raddr_12_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n550) );
  AND2X2 AND2X2_611 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n551), .B(sdram_resetn_bF_buf45), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_12__FF_INPUT) );
  AND2X2 AND2X2_612 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_0_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n553) );
  AND2X2 AND2X2_613 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf3), .B(u_sdrc_core_r2b_caddr_0_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n554) );
  AND2X2 AND2X2_614 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n555), .B(sdram_resetn_bF_buf44), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_0__FF_INPUT) );
  AND2X2 AND2X2_615 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_1_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n557) );
  AND2X2 AND2X2_616 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf2), .B(u_sdrc_core_r2b_caddr_1_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n558) );
  AND2X2 AND2X2_617 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n559), .B(sdram_resetn_bF_buf43), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_1__FF_INPUT) );
  AND2X2 AND2X2_618 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_2_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n561) );
  AND2X2 AND2X2_619 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf1), .B(u_sdrc_core_r2b_caddr_2_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n562) );
  AND2X2 AND2X2_62 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n326_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n324_1), .Y(u_sdrc_core_u_bank_ctl_rank_ba_2__FF_INPUT) );
  AND2X2 AND2X2_620 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n563), .B(sdram_resetn_bF_buf42), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_2__FF_INPUT) );
  AND2X2 AND2X2_621 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_3_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n565) );
  AND2X2 AND2X2_622 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf0), .B(u_sdrc_core_r2b_caddr_3_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n566) );
  AND2X2 AND2X2_623 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n567), .B(sdram_resetn_bF_buf41), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_3__FF_INPUT) );
  AND2X2 AND2X2_624 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf5), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_4_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n569) );
  AND2X2 AND2X2_625 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf4), .B(u_sdrc_core_r2b_caddr_4_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n570) );
  AND2X2 AND2X2_626 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n571), .B(sdram_resetn_bF_buf40), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_4__FF_INPUT) );
  AND2X2 AND2X2_627 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_5_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n573) );
  AND2X2 AND2X2_628 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf3), .B(u_sdrc_core_r2b_caddr_5_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n574) );
  AND2X2 AND2X2_629 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n575), .B(sdram_resetn_bF_buf39), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_5__FF_INPUT) );
  AND2X2 AND2X2_63 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n241), .B(u_sdrc_core_u_bank_ctl_rank_ba_5_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n328_1) );
  AND2X2 AND2X2_630 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_6_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n577) );
  AND2X2 AND2X2_631 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf2), .B(u_sdrc_core_r2b_caddr_6_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n578) );
  AND2X2 AND2X2_632 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n579), .B(sdram_resetn_bF_buf38), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_6__FF_INPUT) );
  AND2X2 AND2X2_633 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_7_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n581) );
  AND2X2 AND2X2_634 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf1), .B(u_sdrc_core_r2b_caddr_7_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n582) );
  AND2X2 AND2X2_635 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n583), .B(sdram_resetn_bF_buf37), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_7__FF_INPUT) );
  AND2X2 AND2X2_636 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_8_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n585) );
  AND2X2 AND2X2_637 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf0), .B(u_sdrc_core_r2b_caddr_8_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n586) );
  AND2X2 AND2X2_638 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n587), .B(sdram_resetn_bF_buf36), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_8__FF_INPUT) );
  AND2X2 AND2X2_639 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_9_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n589) );
  AND2X2 AND2X2_64 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n294_1), .B(u_sdrc_core_u_bank_ctl_rank_ba_3_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n329) );
  AND2X2 AND2X2_640 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf4), .B(u_sdrc_core_r2b_caddr_9_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n590) );
  AND2X2 AND2X2_641 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n591), .B(sdram_resetn_bF_buf35), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_9__FF_INPUT) );
  AND2X2 AND2X2_642 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf5), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_10_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n593) );
  AND2X2 AND2X2_643 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf3), .B(u_sdrc_core_r2b_caddr_10_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n594) );
  AND2X2 AND2X2_644 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n595), .B(sdram_resetn_bF_buf34), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_10__FF_INPUT) );
  AND2X2 AND2X2_645 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_11_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n597) );
  AND2X2 AND2X2_646 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf2), .B(1'b0), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n598) );
  AND2X2 AND2X2_647 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n599), .B(sdram_resetn_bF_buf33), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_11__FF_INPUT) );
  AND2X2 AND2X2_648 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_12_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n601) );
  AND2X2 AND2X2_649 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf1), .B(1'b0), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n602) );
  AND2X2 AND2X2_65 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n332), .B(sdram_resetn_bF_buf43), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n333) );
  AND2X2 AND2X2_650 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n603), .B(sdram_resetn_bF_buf32), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_12__FF_INPUT) );
  AND2X2 AND2X2_651 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_4_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_0_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n605) );
  AND2X2 AND2X2_652 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_0_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n607) );
  AND2X2 AND2X2_653 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n609), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n610), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_0__FF_INPUT) );
  AND2X2 AND2X2_654 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_4_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_1_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n612) );
  AND2X2 AND2X2_655 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_1_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n613) );
  AND2X2 AND2X2_656 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n615), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n616), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_1__FF_INPUT) );
  AND2X2 AND2X2_657 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_4_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_2_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n618) );
  AND2X2 AND2X2_658 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_2_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n619) );
  AND2X2 AND2X2_659 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n621), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n622), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_2__FF_INPUT) );
  AND2X2 AND2X2_66 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n333), .B(u_sdrc_core_u_bank_ctl__abc_21249_n331), .Y(u_sdrc_core_u_bank_ctl_rank_ba_3__FF_INPUT) );
  AND2X2 AND2X2_660 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_4_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_3_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n624) );
  AND2X2 AND2X2_661 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_3_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n625) );
  AND2X2 AND2X2_662 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n627), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n628), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_3__FF_INPUT) );
  AND2X2 AND2X2_663 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_4_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_4_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n630) );
  AND2X2 AND2X2_664 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_4_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n631) );
  AND2X2 AND2X2_665 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n633), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n634), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_4__FF_INPUT) );
  AND2X2 AND2X2_666 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_4_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_5_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n636) );
  AND2X2 AND2X2_667 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_5_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n637) );
  AND2X2 AND2X2_668 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n639), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n640), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_5__FF_INPUT) );
  AND2X2 AND2X2_669 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_4_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_6_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n642) );
  AND2X2 AND2X2_67 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n336), .B(u_sdrc_core_u_bank_ctl__abc_21249_n337), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n338) );
  AND2X2 AND2X2_670 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_6_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n643) );
  AND2X2 AND2X2_671 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n645), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n646), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_6__FF_INPUT) );
  AND2X2 AND2X2_672 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_4_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_7_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n648) );
  AND2X2 AND2X2_673 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_7_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n649) );
  AND2X2 AND2X2_674 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n651), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n652), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_7__FF_INPUT) );
  AND2X2 AND2X2_675 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_4_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_8_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n654) );
  AND2X2 AND2X2_676 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_8_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n655) );
  AND2X2 AND2X2_677 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n657), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n658), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_8__FF_INPUT) );
  AND2X2 AND2X2_678 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_4_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_9_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n660) );
  AND2X2 AND2X2_679 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_9_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n661) );
  AND2X2 AND2X2_68 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n241), .B(u_sdrc_core_u_bank_ctl_rank_ba_6_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n340) );
  AND2X2 AND2X2_680 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n663), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n664), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_9__FF_INPUT) );
  AND2X2 AND2X2_681 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_4_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_10_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n666) );
  AND2X2 AND2X2_682 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n370), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_10_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n667) );
  AND2X2 AND2X2_683 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n669), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n670), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_10__FF_INPUT) );
  AND2X2 AND2X2_684 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_4_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_11_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n672) );
  AND2X2 AND2X2_685 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_11_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n673) );
  AND2X2 AND2X2_686 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n675), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n676), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_11__FF_INPUT) );
  AND2X2 AND2X2_687 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_4_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_12_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n678) );
  AND2X2 AND2X2_688 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n370), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_12_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n679) );
  AND2X2 AND2X2_689 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n681), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n682), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_12__FF_INPUT) );
  AND2X2 AND2X2_69 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n294_1), .B(u_sdrc_core_u_bank_ctl_rank_ba_4_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n341) );
  AND2X2 AND2X2_690 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n689), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n688), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_last) );
  AND2X2 AND2X2_691 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n704), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n703), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_len_0_) );
  AND2X2 AND2X2_692 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n707), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n706), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_len_1_) );
  AND2X2 AND2X2_693 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n710), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n709), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_len_2_) );
  AND2X2 AND2X2_694 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n713), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n712), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_len_3_) );
  AND2X2 AND2X2_695 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n716), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n715), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_len_4_) );
  AND2X2 AND2X2_696 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n719), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n718), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_len_5_) );
  AND2X2 AND2X2_697 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n722), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n721), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_len_6_) );
  AND2X2 AND2X2_698 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n725), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n724), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_wrap) );
  AND2X2 AND2X2_699 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_x2b_pre_ok_t), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_tras_ok), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n727) );
  AND2X2 AND2X2_7 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n213), .B(u_sdrc_core_u_bank_ctl__abc_21249_n211_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_xfr_ok) );
  AND2X2 AND2X2_70 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n344), .B(sdram_resetn_bF_buf42), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n345) );
  AND2X2 AND2X2_700 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n368_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n727), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n728) );
  AND2X2 AND2X2_701 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_2_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_x2b_act_ok_t), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n729) );
  AND2X2 AND2X2_702 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_4_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_r), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n733) );
  AND2X2 AND2X2_703 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n732), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n733), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n734) );
  AND2X2 AND2X2_704 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n734), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n731), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n735) );
  AND2X2 AND2X2_705 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n736), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_timer0_tc), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n737) );
  AND2X2 AND2X2_706 ( .A(sdram_resetn_bF_buf31), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_wrok), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_x2b_wrok_r_FF_INPUT) );
  AND2X2 AND2X2_707 ( .A(sdram_resetn_bF_buf30), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf2), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_r_FF_INPUT) );
  AND2X2 AND2X2_708 ( .A(sdram_resetn_bF_buf29), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_rdok), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_x2b_rdok_r_FF_INPUT) );
  AND2X2 AND2X2_709 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n380), .B(sdram_resetn_bF_buf28), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n743) );
  AND2X2 AND2X2_71 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n345), .B(u_sdrc_core_u_bank_ctl__abc_21249_n343), .Y(u_sdrc_core_u_bank_ctl_rank_ba_4__FF_INPUT) );
  AND2X2 AND2X2_710 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n742), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n743), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_timer0_tc_r_FF_INPUT) );
  AND2X2 AND2X2_711 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n745), .B(sdram_resetn_bF_buf27), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_tras_ok_r_FF_INPUT) );
  AND2X2 AND2X2_712 ( .A(sdram_resetn_bF_buf26), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_pre_ok), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_x2b_pre_ok_r_FF_INPUT) );
  AND2X2 AND2X2_713 ( .A(sdram_resetn_bF_buf25), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_act_ok), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_x2b_act_ok_r_FF_INPUT) );
  AND2X2 AND2X2_714 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n357), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n336), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n750) );
  AND2X2 AND2X2_715 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n749), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n750), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_valid_FF_INPUT) );
  AND2X2 AND2X2_716 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_last), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n756) );
  AND2X2 AND2X2_717 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf0), .B(u_sdrc_core_r2b_last), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n757) );
  AND2X2 AND2X2_718 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n758), .B(sdram_resetn_bF_buf24), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_l_last_FF_INPUT) );
  AND2X2 AND2X2_719 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_wrap), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n760) );
  AND2X2 AND2X2_72 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n241), .B(u_sdrc_core_u_bank_ctl_rank_ba_7_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n347) );
  AND2X2 AND2X2_720 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf4), .B(u_sdrc_core_r2b_wrap), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n761) );
  AND2X2 AND2X2_721 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n762), .B(sdram_resetn_bF_buf23), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_l_wrap_FF_INPUT) );
  AND2X2 AND2X2_722 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_write), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n764) );
  AND2X2 AND2X2_723 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf3), .B(u_sdrc_core_r2b_write), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n765) );
  AND2X2 AND2X2_724 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n766), .B(sdram_resetn_bF_buf22), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_l_write_FF_INPUT) );
  AND2X2 AND2X2_725 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf5), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_sdr_dma_last), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n768) );
  AND2X2 AND2X2_726 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf2), .B(1'b0), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n769) );
  AND2X2 AND2X2_727 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n770), .B(sdram_resetn_bF_buf21), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_l_sdr_dma_last_FF_INPUT) );
  AND2X2 AND2X2_728 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n249_1), .B(sdram_resetn_bF_buf20), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n250_1) );
  AND2X2 AND2X2_729 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n250_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_3_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n251) );
  AND2X2 AND2X2_73 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n294_1), .B(u_sdrc_core_u_bank_ctl_rank_ba_5_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n348) );
  AND2X2 AND2X2_730 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_r2b_req), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_0_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack) );
  AND2X2 AND2X2_731 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf3), .B(sdram_resetn_bF_buf19), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n253_1) );
  AND2X2 AND2X2_732 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n257), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n259_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n260) );
  AND2X2 AND2X2_733 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n260), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n255_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n261_1) );
  AND2X2 AND2X2_734 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n263), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n265_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n266) );
  AND2X2 AND2X2_735 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n268_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n270_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n271_1) );
  AND2X2 AND2X2_736 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n266), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n271_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n272) );
  AND2X2 AND2X2_737 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n272), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n261_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n273_1) );
  AND2X2 AND2X2_738 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n275), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n277_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n278) );
  AND2X2 AND2X2_739 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n280_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n282_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n283_1) );
  AND2X2 AND2X2_74 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n351), .B(sdram_resetn_bF_buf41), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n352) );
  AND2X2 AND2X2_740 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n278), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n283_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n284_1) );
  AND2X2 AND2X2_741 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n286_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n288_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n289) );
  AND2X2 AND2X2_742 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n291_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n293), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n294_1) );
  AND2X2 AND2X2_743 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n289), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n294_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n295_1) );
  AND2X2 AND2X2_744 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n284_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n295_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n296_1) );
  AND2X2 AND2X2_745 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n296_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n273_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n297) );
  AND2X2 AND2X2_746 ( .A(u_sdrc_core_r2b_raddr_10_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_10_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n298_1) );
  AND2X2 AND2X2_747 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n299_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n300_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n301) );
  AND2X2 AND2X2_748 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_8_), .B(u_sdrc_core_r2b_raddr_8_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n303_1) );
  AND2X2 AND2X2_749 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n304_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n305), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n306_1) );
  AND2X2 AND2X2_75 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n352), .B(u_sdrc_core_u_bank_ctl__abc_21249_n350), .Y(u_sdrc_core_u_bank_ctl_rank_ba_5__FF_INPUT) );
  AND2X2 AND2X2_750 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n302_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n307_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n308_1) );
  AND2X2 AND2X2_751 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n310_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n312_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n313) );
  AND2X2 AND2X2_752 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n315_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n317), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n318_1) );
  AND2X2 AND2X2_753 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n313), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n318_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n319_1) );
  AND2X2 AND2X2_754 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n321), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n323_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n324_1) );
  AND2X2 AND2X2_755 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n326_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_valid), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n327_1) );
  AND2X2 AND2X2_756 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n324_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n327_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n328_1) );
  AND2X2 AND2X2_757 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n319_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n328_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n329) );
  AND2X2 AND2X2_758 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n329), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n308_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n330_1) );
  AND2X2 AND2X2_759 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n297), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n330_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n331_1) );
  AND2X2 AND2X2_76 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n219_1), .B(u_sdrc_core_u_bank_ctl_rank_cnt_2_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n355) );
  AND2X2 AND2X2_760 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n332_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n253_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n333) );
  AND2X2 AND2X2_761 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n250_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_prech_page_closed), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n335) );
  AND2X2 AND2X2_762 ( .A(sdram_resetn_bF_buf18), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_4_bF_buf3), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n337) );
  AND2X2 AND2X2_763 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n337), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n336), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n338_1) );
  AND2X2 AND2X2_764 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n338_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_x2b_ack), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n339_1) );
  AND2X2 AND2X2_765 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n339_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_sdr_dma_last), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n340) );
  AND2X2 AND2X2_766 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n250_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_2_bF_buf3), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n342) );
  AND2X2 AND2X2_767 ( .A(sdram_resetn_bF_buf17), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_x2b_ack), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n343_1) );
  AND2X2 AND2X2_768 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n343_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_3_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n344_1) );
  AND2X2 AND2X2_769 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n337), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_refresh), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n345) );
  AND2X2 AND2X2_77 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n354), .B(u_sdrc_core_u_bank_ctl__abc_21249_n357), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n358) );
  AND2X2 AND2X2_770 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n343_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_2_bF_buf2), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n348_1) );
  AND2X2 AND2X2_771 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n338_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n249_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n349_1) );
  AND2X2 AND2X2_772 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n331_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n253_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n351) );
  AND2X2 AND2X2_773 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n339_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n353_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n354_1) );
  AND2X2 AND2X2_774 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n356), .B(sdram_resetn_bF_buf16), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n357) );
  AND2X2 AND2X2_775 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n355), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n358_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n359_1) );
  AND2X2 AND2X2_776 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n360), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_0_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n361) );
  AND2X2 AND2X2_777 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_4_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_write), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n364_1) );
  AND2X2 AND2X2_778 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n369_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n367), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n370) );
  AND2X2 AND2X2_779 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n370), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n371) );
  AND2X2 AND2X2_78 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n294_1), .B(u_sdrc_core_u_bank_ctl_rank_ba_6_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n360) );
  AND2X2 AND2X2_780 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n371), .B(u_sdrc_core_r2b_write), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n372) );
  AND2X2 AND2X2_781 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n331_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n372), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n373_1) );
  AND2X2 AND2X2_782 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n374_1), .B(sdram_resetn_bF_buf15), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_cmd_r_0__FF_INPUT) );
  AND2X2 AND2X2_783 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n371), .B(sdram_resetn_bF_buf14), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n376) );
  AND2X2 AND2X2_784 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n331_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n376), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n377) );
  AND2X2 AND2X2_785 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n381), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_cmd_0_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n382) );
  AND2X2 AND2X2_786 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n383_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n386_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n387_1) );
  AND2X2 AND2X2_787 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n387_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n379_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n388) );
  AND2X2 AND2X2_788 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n382), .B(\cfg_sdr_tras_d[0] ), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n389) );
  AND2X2 AND2X2_789 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n390), .B(sdram_resetn_bF_buf13), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_tras_cntr_0__FF_INPUT) );
  AND2X2 AND2X2_79 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n362), .B(sdram_resetn_bF_buf40), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n363) );
  AND2X2 AND2X2_790 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n382), .B(\cfg_sdr_tras_d[1] ), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n392_1) );
  AND2X2 AND2X2_791 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_tras_cntr_0_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_tras_cntr_1_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n394_1) );
  AND2X2 AND2X2_792 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n387_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n395_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n396_1) );
  AND2X2 AND2X2_793 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n397_1), .B(sdram_resetn_bF_buf12), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_tras_cntr_1__FF_INPUT) );
  AND2X2 AND2X2_794 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n382), .B(\cfg_sdr_tras_d[2] ), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n399_1) );
  AND2X2 AND2X2_795 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n384_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_tras_cntr_2_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n401_1) );
  AND2X2 AND2X2_796 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n387_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n402_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n403_1) );
  AND2X2 AND2X2_797 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n404_1), .B(sdram_resetn_bF_buf11), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_tras_cntr_2__FF_INPUT) );
  AND2X2 AND2X2_798 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n385), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_tras_cntr_3_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n406_1) );
  AND2X2 AND2X2_799 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n408_1), .B(sdram_resetn_bF_buf10), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n409_1) );
  AND2X2 AND2X2_8 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n217_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n218_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n219_1) );
  AND2X2 AND2X2_80 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n363), .B(u_sdrc_core_u_bank_ctl__abc_21249_n361), .Y(u_sdrc_core_u_bank_ctl_rank_ba_6__FF_INPUT) );
  AND2X2 AND2X2_800 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n409_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n407_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_tras_cntr_3__FF_INPUT) );
  AND2X2 AND2X2_801 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n415_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n413_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n416) );
  AND2X2 AND2X2_802 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n417_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n418), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n419_1) );
  AND2X2 AND2X2_803 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n421), .B(sdram_resetn_bF_buf9), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n422) );
  AND2X2 AND2X2_804 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n420_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n422), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_timer0_0__FF_INPUT) );
  AND2X2 AND2X2_805 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_timer0_1_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_timer0_0_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n426) );
  AND2X2 AND2X2_806 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n383_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n428_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n429) );
  AND2X2 AND2X2_807 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n429), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n427_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n430) );
  AND2X2 AND2X2_808 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n381), .B(\cfg_sdr_trcd_d[1] ), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n431_1) );
  AND2X2 AND2X2_809 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n434_1), .B(sdram_resetn_bF_buf8), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n435_1) );
  AND2X2 AND2X2_81 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n294_1), .B(u_sdrc_core_u_bank_ctl_rank_ba_7_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n365) );
  AND2X2 AND2X2_810 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n433), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n435_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_timer0_1__FF_INPUT) );
  AND2X2 AND2X2_811 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n424), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_timer0_2_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n439_1) );
  AND2X2 AND2X2_812 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n429), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n440_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n441) );
  AND2X2 AND2X2_813 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n381), .B(\cfg_sdr_trcd_d[2] ), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n442) );
  AND2X2 AND2X2_814 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n445_1), .B(sdram_resetn_bF_buf7), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n446_1) );
  AND2X2 AND2X2_815 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n444_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n446_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_timer0_2__FF_INPUT) );
  AND2X2 AND2X2_816 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n437_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_timer0_3_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n448_1) );
  AND2X2 AND2X2_817 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n449_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n450), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n451) );
  AND2X2 AND2X2_818 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n453_1), .B(sdram_resetn_bF_buf6), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n454) );
  AND2X2 AND2X2_819 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n452), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n454), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_timer0_3__FF_INPUT) );
  AND2X2 AND2X2_82 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n367), .B(sdram_resetn_bF_buf39), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n368) );
  AND2X2 AND2X2_820 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n253_1), .B(u_sdrc_core_r2b_len_0_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n473) );
  AND2X2 AND2X2_821 ( .A(sdram_resetn_bF_buf5), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_0_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n474) );
  AND2X2 AND2X2_822 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf5), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n474), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n475) );
  AND2X2 AND2X2_823 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n253_1), .B(u_sdrc_core_r2b_len_1_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n477) );
  AND2X2 AND2X2_824 ( .A(sdram_resetn_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_1_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n478) );
  AND2X2 AND2X2_825 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n478), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n479) );
  AND2X2 AND2X2_826 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n253_1), .B(u_sdrc_core_r2b_len_2_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n481) );
  AND2X2 AND2X2_827 ( .A(sdram_resetn_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_2_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n482) );
  AND2X2 AND2X2_828 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n482), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n483) );
  AND2X2 AND2X2_829 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n253_1), .B(u_sdrc_core_r2b_len_3_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n485) );
  AND2X2 AND2X2_83 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n368), .B(u_sdrc_core_u_bank_ctl__abc_21249_n366), .Y(u_sdrc_core_u_bank_ctl_rank_ba_7__FF_INPUT) );
  AND2X2 AND2X2_830 ( .A(sdram_resetn_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_3_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n486) );
  AND2X2 AND2X2_831 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n486), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n487) );
  AND2X2 AND2X2_832 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n253_1), .B(u_sdrc_core_r2b_len_4_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n489) );
  AND2X2 AND2X2_833 ( .A(sdram_resetn_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_4_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n490) );
  AND2X2 AND2X2_834 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n490), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n491) );
  AND2X2 AND2X2_835 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n253_1), .B(u_sdrc_core_r2b_len_5_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n493) );
  AND2X2 AND2X2_836 ( .A(sdram_resetn_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_5_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n494) );
  AND2X2 AND2X2_837 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n494), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n495) );
  AND2X2 AND2X2_838 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n253_1), .B(u_sdrc_core_r2b_len_6_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n497) );
  AND2X2 AND2X2_839 ( .A(sdram_resetn_bF_buf49), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_6_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n498) );
  AND2X2 AND2X2_84 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_0_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n370) );
  AND2X2 AND2X2_840 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf5), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n498), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n499) );
  AND2X2 AND2X2_841 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_0_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n501) );
  AND2X2 AND2X2_842 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf1), .B(u_sdrc_core_r2b_raddr_0_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n502) );
  AND2X2 AND2X2_843 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n503), .B(sdram_resetn_bF_buf48), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_0__FF_INPUT) );
  AND2X2 AND2X2_844 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_1_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n505) );
  AND2X2 AND2X2_845 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf0), .B(u_sdrc_core_r2b_raddr_1_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n506) );
  AND2X2 AND2X2_846 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n507), .B(sdram_resetn_bF_buf47), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_1__FF_INPUT) );
  AND2X2 AND2X2_847 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_2_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n509) );
  AND2X2 AND2X2_848 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf4), .B(u_sdrc_core_r2b_raddr_2_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n510) );
  AND2X2 AND2X2_849 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n511), .B(sdram_resetn_bF_buf46), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_2__FF_INPUT) );
  AND2X2 AND2X2_85 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n372), .B(u_sdrc_core_u_bank_ctl__abc_21249_n371), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n373) );
  AND2X2 AND2X2_850 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_3_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n513) );
  AND2X2 AND2X2_851 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf3), .B(u_sdrc_core_r2b_raddr_3_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n514) );
  AND2X2 AND2X2_852 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n515), .B(sdram_resetn_bF_buf45), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_3__FF_INPUT) );
  AND2X2 AND2X2_853 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_4_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n517) );
  AND2X2 AND2X2_854 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf2), .B(u_sdrc_core_r2b_raddr_4_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n518) );
  AND2X2 AND2X2_855 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n519), .B(sdram_resetn_bF_buf44), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_4__FF_INPUT) );
  AND2X2 AND2X2_856 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf5), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_5_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n521) );
  AND2X2 AND2X2_857 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf1), .B(u_sdrc_core_r2b_raddr_5_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n522) );
  AND2X2 AND2X2_858 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n523), .B(sdram_resetn_bF_buf43), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_5__FF_INPUT) );
  AND2X2 AND2X2_859 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_6_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n525) );
  AND2X2 AND2X2_86 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n374), .B(u_sdrc_core_u_bank_ctl__abc_21249_n375), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n376) );
  AND2X2 AND2X2_860 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf0), .B(u_sdrc_core_r2b_raddr_6_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n526) );
  AND2X2 AND2X2_861 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n527), .B(sdram_resetn_bF_buf42), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_6__FF_INPUT) );
  AND2X2 AND2X2_862 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_7_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n529) );
  AND2X2 AND2X2_863 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf4), .B(u_sdrc_core_r2b_raddr_7_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n530) );
  AND2X2 AND2X2_864 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n531), .B(sdram_resetn_bF_buf41), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_7__FF_INPUT) );
  AND2X2 AND2X2_865 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_8_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n533) );
  AND2X2 AND2X2_866 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf3), .B(u_sdrc_core_r2b_raddr_8_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n534) );
  AND2X2 AND2X2_867 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n535), .B(sdram_resetn_bF_buf40), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_8__FF_INPUT) );
  AND2X2 AND2X2_868 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_9_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n537) );
  AND2X2 AND2X2_869 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf2), .B(u_sdrc_core_r2b_raddr_9_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n538) );
  AND2X2 AND2X2_87 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n376), .B(u_sdrc_core_u_bank_ctl__abc_21249_n227_bF_buf2), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n377) );
  AND2X2 AND2X2_870 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n539), .B(sdram_resetn_bF_buf39), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_9__FF_INPUT) );
  AND2X2 AND2X2_871 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_10_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n541) );
  AND2X2 AND2X2_872 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf1), .B(u_sdrc_core_r2b_raddr_10_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n542) );
  AND2X2 AND2X2_873 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n543), .B(sdram_resetn_bF_buf38), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_10__FF_INPUT) );
  AND2X2 AND2X2_874 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf5), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_11_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n545) );
  AND2X2 AND2X2_875 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf0), .B(u_sdrc_core_r2b_raddr_11_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n546) );
  AND2X2 AND2X2_876 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n547), .B(sdram_resetn_bF_buf37), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_11__FF_INPUT) );
  AND2X2 AND2X2_877 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_12_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n549) );
  AND2X2 AND2X2_878 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf4), .B(u_sdrc_core_r2b_raddr_12_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n550) );
  AND2X2 AND2X2_879 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n551), .B(sdram_resetn_bF_buf36), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_12__FF_INPUT) );
  AND2X2 AND2X2_88 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_1_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n379) );
  AND2X2 AND2X2_880 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_0_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n553) );
  AND2X2 AND2X2_881 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf3), .B(u_sdrc_core_r2b_caddr_0_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n554) );
  AND2X2 AND2X2_882 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n555), .B(sdram_resetn_bF_buf35), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_0__FF_INPUT) );
  AND2X2 AND2X2_883 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_1_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n557) );
  AND2X2 AND2X2_884 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf2), .B(u_sdrc_core_r2b_caddr_1_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n558) );
  AND2X2 AND2X2_885 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n559), .B(sdram_resetn_bF_buf34), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_1__FF_INPUT) );
  AND2X2 AND2X2_886 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_2_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n561) );
  AND2X2 AND2X2_887 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf1), .B(u_sdrc_core_r2b_caddr_2_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n562) );
  AND2X2 AND2X2_888 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n563), .B(sdram_resetn_bF_buf33), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_2__FF_INPUT) );
  AND2X2 AND2X2_889 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_3_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n565) );
  AND2X2 AND2X2_89 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n381), .B(u_sdrc_core_u_bank_ctl__abc_21249_n380), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n382) );
  AND2X2 AND2X2_890 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf0), .B(u_sdrc_core_r2b_caddr_3_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n566) );
  AND2X2 AND2X2_891 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n567), .B(sdram_resetn_bF_buf32), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_3__FF_INPUT) );
  AND2X2 AND2X2_892 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf5), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_4_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n569) );
  AND2X2 AND2X2_893 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf4), .B(u_sdrc_core_r2b_caddr_4_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n570) );
  AND2X2 AND2X2_894 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n571), .B(sdram_resetn_bF_buf31), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_4__FF_INPUT) );
  AND2X2 AND2X2_895 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_5_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n573) );
  AND2X2 AND2X2_896 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf3), .B(u_sdrc_core_r2b_caddr_5_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n574) );
  AND2X2 AND2X2_897 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n575), .B(sdram_resetn_bF_buf30), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_5__FF_INPUT) );
  AND2X2 AND2X2_898 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_6_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n577) );
  AND2X2 AND2X2_899 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf2), .B(u_sdrc_core_r2b_caddr_6_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n578) );
  AND2X2 AND2X2_9 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n219_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n216_1), .Y(u_sdrc_core_b2x_idle) );
  AND2X2 AND2X2_90 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n383), .B(u_sdrc_core_u_bank_ctl__abc_21249_n384), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n385) );
  AND2X2 AND2X2_900 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n579), .B(sdram_resetn_bF_buf29), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_6__FF_INPUT) );
  AND2X2 AND2X2_901 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_7_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n581) );
  AND2X2 AND2X2_902 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf1), .B(u_sdrc_core_r2b_caddr_7_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n582) );
  AND2X2 AND2X2_903 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n583), .B(sdram_resetn_bF_buf28), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_7__FF_INPUT) );
  AND2X2 AND2X2_904 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_8_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n585) );
  AND2X2 AND2X2_905 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf0), .B(u_sdrc_core_r2b_caddr_8_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n586) );
  AND2X2 AND2X2_906 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n587), .B(sdram_resetn_bF_buf27), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_8__FF_INPUT) );
  AND2X2 AND2X2_907 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_9_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n589) );
  AND2X2 AND2X2_908 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf4), .B(u_sdrc_core_r2b_caddr_9_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n590) );
  AND2X2 AND2X2_909 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n591), .B(sdram_resetn_bF_buf26), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_9__FF_INPUT) );
  AND2X2 AND2X2_91 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n385), .B(u_sdrc_core_u_bank_ctl__abc_21249_n227_bF_buf1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n386) );
  AND2X2 AND2X2_910 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf5), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_10_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n593) );
  AND2X2 AND2X2_911 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf3), .B(u_sdrc_core_r2b_caddr_10_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n594) );
  AND2X2 AND2X2_912 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n595), .B(sdram_resetn_bF_buf25), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_10__FF_INPUT) );
  AND2X2 AND2X2_913 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_11_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n597) );
  AND2X2 AND2X2_914 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf2), .B(1'b0), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n598) );
  AND2X2 AND2X2_915 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n599), .B(sdram_resetn_bF_buf24), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_11__FF_INPUT) );
  AND2X2 AND2X2_916 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_12_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n601) );
  AND2X2 AND2X2_917 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf1), .B(1'b0), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n602) );
  AND2X2 AND2X2_918 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n603), .B(sdram_resetn_bF_buf23), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_12__FF_INPUT) );
  AND2X2 AND2X2_919 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_4_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_0_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n605) );
  AND2X2 AND2X2_92 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_2_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n388) );
  AND2X2 AND2X2_920 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_0_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n607) );
  AND2X2 AND2X2_921 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n609), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n610), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_0__FF_INPUT) );
  AND2X2 AND2X2_922 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_4_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_1_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n612) );
  AND2X2 AND2X2_923 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_1_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n613) );
  AND2X2 AND2X2_924 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n615), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n616), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_1__FF_INPUT) );
  AND2X2 AND2X2_925 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_4_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_2_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n618) );
  AND2X2 AND2X2_926 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_2_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n619) );
  AND2X2 AND2X2_927 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n621), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n622), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_2__FF_INPUT) );
  AND2X2 AND2X2_928 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_4_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_3_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n624) );
  AND2X2 AND2X2_929 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_3_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n625) );
  AND2X2 AND2X2_93 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n390), .B(u_sdrc_core_u_bank_ctl__abc_21249_n389), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n391) );
  AND2X2 AND2X2_930 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n627), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n628), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_3__FF_INPUT) );
  AND2X2 AND2X2_931 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_4_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_4_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n630) );
  AND2X2 AND2X2_932 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_4_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n631) );
  AND2X2 AND2X2_933 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n633), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n634), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_4__FF_INPUT) );
  AND2X2 AND2X2_934 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_4_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_5_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n636) );
  AND2X2 AND2X2_935 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_5_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n637) );
  AND2X2 AND2X2_936 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n639), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n640), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_5__FF_INPUT) );
  AND2X2 AND2X2_937 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_4_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_6_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n642) );
  AND2X2 AND2X2_938 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_6_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n643) );
  AND2X2 AND2X2_939 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n645), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n646), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_6__FF_INPUT) );
  AND2X2 AND2X2_94 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n392), .B(u_sdrc_core_u_bank_ctl__abc_21249_n393), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n394) );
  AND2X2 AND2X2_940 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_4_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_7_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n648) );
  AND2X2 AND2X2_941 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_7_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n649) );
  AND2X2 AND2X2_942 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n651), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n652), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_7__FF_INPUT) );
  AND2X2 AND2X2_943 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_4_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_8_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n654) );
  AND2X2 AND2X2_944 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_8_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n655) );
  AND2X2 AND2X2_945 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n657), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n658), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_8__FF_INPUT) );
  AND2X2 AND2X2_946 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_4_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_9_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n660) );
  AND2X2 AND2X2_947 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_9_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n661) );
  AND2X2 AND2X2_948 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n663), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n664), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_9__FF_INPUT) );
  AND2X2 AND2X2_949 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_4_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_10_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n666) );
  AND2X2 AND2X2_95 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n394), .B(u_sdrc_core_u_bank_ctl__abc_21249_n227_bF_buf0), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n395) );
  AND2X2 AND2X2_950 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n370), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_10_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n667) );
  AND2X2 AND2X2_951 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n669), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n670), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_10__FF_INPUT) );
  AND2X2 AND2X2_952 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_4_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_11_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n672) );
  AND2X2 AND2X2_953 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n606), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_11_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n673) );
  AND2X2 AND2X2_954 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n675), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n676), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_11__FF_INPUT) );
  AND2X2 AND2X2_955 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_4_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_12_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n678) );
  AND2X2 AND2X2_956 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n370), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_12_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n679) );
  AND2X2 AND2X2_957 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n681), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n682), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_12__FF_INPUT) );
  AND2X2 AND2X2_958 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n689), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n688), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_last) );
  AND2X2 AND2X2_959 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n704), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n703), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_len_0_) );
  AND2X2 AND2X2_96 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_3_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n397) );
  AND2X2 AND2X2_960 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n707), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n706), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_len_1_) );
  AND2X2 AND2X2_961 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n710), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n709), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_len_2_) );
  AND2X2 AND2X2_962 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n713), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n712), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_len_3_) );
  AND2X2 AND2X2_963 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n716), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n715), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_len_4_) );
  AND2X2 AND2X2_964 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n719), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n718), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_len_5_) );
  AND2X2 AND2X2_965 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n722), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n721), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_len_6_) );
  AND2X2 AND2X2_966 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n725), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n724), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_wrap) );
  AND2X2 AND2X2_967 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_x2b_pre_ok_t), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_tras_ok), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n727) );
  AND2X2 AND2X2_968 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n368_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n727), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n728) );
  AND2X2 AND2X2_969 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_2_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_x2b_act_ok_t), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n729) );
  AND2X2 AND2X2_97 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n399), .B(u_sdrc_core_u_bank_ctl__abc_21249_n398), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n400) );
  AND2X2 AND2X2_970 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_4_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_r), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n733) );
  AND2X2 AND2X2_971 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n732), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n733), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n734) );
  AND2X2 AND2X2_972 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n734), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n731), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n735) );
  AND2X2 AND2X2_973 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n736), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_timer0_tc), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n737) );
  AND2X2 AND2X2_974 ( .A(sdram_resetn_bF_buf22), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_wrok), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_x2b_wrok_r_FF_INPUT) );
  AND2X2 AND2X2_975 ( .A(sdram_resetn_bF_buf21), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf2), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_r_FF_INPUT) );
  AND2X2 AND2X2_976 ( .A(sdram_resetn_bF_buf20), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_rdok), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_x2b_rdok_r_FF_INPUT) );
  AND2X2 AND2X2_977 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n380), .B(sdram_resetn_bF_buf19), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n743) );
  AND2X2 AND2X2_978 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n742), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n743), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_timer0_tc_r_FF_INPUT) );
  AND2X2 AND2X2_979 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n745), .B(sdram_resetn_bF_buf18), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_tras_ok_r_FF_INPUT) );
  AND2X2 AND2X2_98 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n401), .B(u_sdrc_core_u_bank_ctl__abc_21249_n402), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n403) );
  AND2X2 AND2X2_980 ( .A(sdram_resetn_bF_buf17), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_pre_ok), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_x2b_pre_ok_r_FF_INPUT) );
  AND2X2 AND2X2_981 ( .A(sdram_resetn_bF_buf16), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_act_ok), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_x2b_act_ok_r_FF_INPUT) );
  AND2X2 AND2X2_982 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n357), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n336), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n750) );
  AND2X2 AND2X2_983 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n749), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n750), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_valid_FF_INPUT) );
  AND2X2 AND2X2_984 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_last), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n756) );
  AND2X2 AND2X2_985 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf0), .B(u_sdrc_core_r2b_last), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n757) );
  AND2X2 AND2X2_986 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n758), .B(sdram_resetn_bF_buf15), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_l_last_FF_INPUT) );
  AND2X2 AND2X2_987 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_wrap), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n760) );
  AND2X2 AND2X2_988 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf4), .B(u_sdrc_core_r2b_wrap), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n761) );
  AND2X2 AND2X2_989 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n762), .B(sdram_resetn_bF_buf14), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_l_wrap_FF_INPUT) );
  AND2X2 AND2X2_99 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n403), .B(u_sdrc_core_u_bank_ctl__abc_21249_n227_bF_buf3), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n404) );
  AND2X2 AND2X2_990 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_write), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n764) );
  AND2X2 AND2X2_991 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf3), .B(u_sdrc_core_r2b_write), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n765) );
  AND2X2 AND2X2_992 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n766), .B(sdram_resetn_bF_buf13), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_l_write_FF_INPUT) );
  AND2X2 AND2X2_993 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf5), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_sdr_dma_last), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n768) );
  AND2X2 AND2X2_994 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf2), .B(1'b0), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n769) );
  AND2X2 AND2X2_995 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n770), .B(sdram_resetn_bF_buf12), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_l_sdr_dma_last_FF_INPUT) );
  AND2X2 AND2X2_996 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n249_1), .B(sdram_resetn_bF_buf11), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n250_1) );
  AND2X2 AND2X2_997 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n250_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_3_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n251) );
  AND2X2 AND2X2_998 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_r2b_req), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_0_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack) );
  AND2X2 AND2X2_999 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf3), .B(sdram_resetn_bF_buf10), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n253_1) );
  BUFX2 BUFX2_1 ( .A(sdram_resetn), .Y(sdram_resetn_hier0_bF_buf6) );
  BUFX2 BUFX2_10 ( .A(wb_clk_i), .Y(wb_clk_i_hier0_bF_buf4) );
  BUFX2 BUFX2_100 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf0) );
  BUFX2 BUFX2_101 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf5) );
  BUFX2 BUFX2_102 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf4) );
  BUFX2 BUFX2_103 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf3) );
  BUFX2 BUFX2_104 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf2) );
  BUFX2 BUFX2_105 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf1) );
  BUFX2 BUFX2_106 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf0) );
  BUFX2 BUFX2_107 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf5) );
  BUFX2 BUFX2_108 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf4) );
  BUFX2 BUFX2_109 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf3) );
  BUFX2 BUFX2_11 ( .A(wb_clk_i), .Y(wb_clk_i_hier0_bF_buf3) );
  BUFX2 BUFX2_110 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf2) );
  BUFX2 BUFX2_111 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf1) );
  BUFX2 BUFX2_112 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf0) );
  BUFX2 BUFX2_113 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf5) );
  BUFX2 BUFX2_114 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf4) );
  BUFX2 BUFX2_115 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf3) );
  BUFX2 BUFX2_116 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf2) );
  BUFX2 BUFX2_117 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf1) );
  BUFX2 BUFX2_118 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf0) );
  BUFX2 BUFX2_119 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_2_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_2_bF_buf3) );
  BUFX2 BUFX2_12 ( .A(wb_clk_i), .Y(wb_clk_i_hier0_bF_buf2) );
  BUFX2 BUFX2_120 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_2_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_2_bF_buf2) );
  BUFX2 BUFX2_121 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_2_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_2_bF_buf1) );
  BUFX2 BUFX2_122 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_2_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_2_bF_buf0) );
  BUFX2 BUFX2_123 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf7) );
  BUFX2 BUFX2_124 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf6) );
  BUFX2 BUFX2_125 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf5) );
  BUFX2 BUFX2_126 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf4) );
  BUFX2 BUFX2_127 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf3) );
  BUFX2 BUFX2_128 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf2) );
  BUFX2 BUFX2_129 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf1) );
  BUFX2 BUFX2_13 ( .A(wb_clk_i), .Y(wb_clk_i_hier0_bF_buf1) );
  BUFX2 BUFX2_130 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf0) );
  BUFX2 BUFX2_131 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf5) );
  BUFX2 BUFX2_132 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf4) );
  BUFX2 BUFX2_133 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf3) );
  BUFX2 BUFX2_134 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf2) );
  BUFX2 BUFX2_135 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf1) );
  BUFX2 BUFX2_136 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf0) );
  BUFX2 BUFX2_137 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_4_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_4_bF_buf3) );
  BUFX2 BUFX2_138 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_4_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_4_bF_buf2) );
  BUFX2 BUFX2_139 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_4_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_4_bF_buf1) );
  BUFX2 BUFX2_14 ( .A(wb_clk_i), .Y(wb_clk_i_hier0_bF_buf0) );
  BUFX2 BUFX2_140 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_4_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_4_bF_buf0) );
  BUFX2 BUFX2_141 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf5) );
  BUFX2 BUFX2_142 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf4) );
  BUFX2 BUFX2_143 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf3) );
  BUFX2 BUFX2_144 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf2) );
  BUFX2 BUFX2_145 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf1) );
  BUFX2 BUFX2_146 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1_bF_buf0) );
  BUFX2 BUFX2_147 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf4) );
  BUFX2 BUFX2_148 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf3) );
  BUFX2 BUFX2_149 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf2) );
  BUFX2 BUFX2_15 ( .A(sdram_clk), .Y(sdram_clk_hier0_bF_buf8) );
  BUFX2 BUFX2_150 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf1) );
  BUFX2 BUFX2_151 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf0) );
  BUFX2 BUFX2_152 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n449), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf4) );
  BUFX2 BUFX2_153 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n449), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf3) );
  BUFX2 BUFX2_154 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n449), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf2) );
  BUFX2 BUFX2_155 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n449), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf1) );
  BUFX2 BUFX2_156 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n449), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n449_bF_buf0) );
  BUFX2 BUFX2_157 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_0_), .Y(u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf4) );
  BUFX2 BUFX2_158 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_0_), .Y(u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf3) );
  BUFX2 BUFX2_159 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_0_), .Y(u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf2) );
  BUFX2 BUFX2_16 ( .A(sdram_clk), .Y(sdram_clk_hier0_bF_buf7) );
  BUFX2 BUFX2_160 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_0_), .Y(u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf1) );
  BUFX2 BUFX2_161 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_0_), .Y(u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf0) );
  BUFX2 BUFX2_162 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n883), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n883_bF_buf3) );
  BUFX2 BUFX2_163 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n883), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n883_bF_buf2) );
  BUFX2 BUFX2_164 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n883), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n883_bF_buf1) );
  BUFX2 BUFX2_165 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n883), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n883_bF_buf0) );
  BUFX2 BUFX2_166 ( .A(u_sdrc_core_u_req_gen__abc_22171_n242), .Y(u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf4) );
  BUFX2 BUFX2_167 ( .A(u_sdrc_core_u_req_gen__abc_22171_n242), .Y(u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf3) );
  BUFX2 BUFX2_168 ( .A(u_sdrc_core_u_req_gen__abc_22171_n242), .Y(u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf2) );
  BUFX2 BUFX2_169 ( .A(u_sdrc_core_u_req_gen__abc_22171_n242), .Y(u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf1) );
  BUFX2 BUFX2_17 ( .A(sdram_clk), .Y(sdram_clk_hier0_bF_buf6) );
  BUFX2 BUFX2_170 ( .A(u_sdrc_core_u_req_gen__abc_22171_n242), .Y(u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf0) );
  BUFX2 BUFX2_171 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf5) );
  BUFX2 BUFX2_172 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf4) );
  BUFX2 BUFX2_173 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf3) );
  BUFX2 BUFX2_174 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf2) );
  BUFX2 BUFX2_175 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf1) );
  BUFX2 BUFX2_176 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf0) );
  BUFX2 BUFX2_177 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n523_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n523_1_bF_buf3) );
  BUFX2 BUFX2_178 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n523_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n523_1_bF_buf2) );
  BUFX2 BUFX2_179 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n523_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n523_1_bF_buf1) );
  BUFX2 BUFX2_18 ( .A(sdram_clk), .Y(sdram_clk_hier0_bF_buf5) );
  BUFX2 BUFX2_180 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n523_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n523_1_bF_buf0) );
  BUFX2 BUFX2_181 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf5) );
  BUFX2 BUFX2_182 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf4) );
  BUFX2 BUFX2_183 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf3) );
  BUFX2 BUFX2_184 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf2) );
  BUFX2 BUFX2_185 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf1) );
  BUFX2 BUFX2_186 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf0) );
  BUFX2 BUFX2_187 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf5) );
  BUFX2 BUFX2_188 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf4) );
  BUFX2 BUFX2_189 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf3) );
  BUFX2 BUFX2_19 ( .A(sdram_clk), .Y(sdram_clk_hier0_bF_buf4) );
  BUFX2 BUFX2_190 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf2) );
  BUFX2 BUFX2_191 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf1) );
  BUFX2 BUFX2_192 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf0) );
  BUFX2 BUFX2_193 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf5) );
  BUFX2 BUFX2_194 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf4) );
  BUFX2 BUFX2_195 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf3) );
  BUFX2 BUFX2_196 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf2) );
  BUFX2 BUFX2_197 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf1) );
  BUFX2 BUFX2_198 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n982), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n982_bF_buf0) );
  BUFX2 BUFX2_199 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf4) );
  BUFX2 BUFX2_2 ( .A(sdram_resetn), .Y(sdram_resetn_hier0_bF_buf5) );
  BUFX2 BUFX2_20 ( .A(sdram_clk), .Y(sdram_clk_hier0_bF_buf3) );
  BUFX2 BUFX2_200 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf3) );
  BUFX2 BUFX2_201 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf2) );
  BUFX2 BUFX2_202 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf1) );
  BUFX2 BUFX2_203 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf0) );
  BUFX2 BUFX2_204 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_2_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_2_bF_buf3) );
  BUFX2 BUFX2_205 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_2_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_2_bF_buf2) );
  BUFX2 BUFX2_206 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_2_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_2_bF_buf1) );
  BUFX2 BUFX2_207 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_2_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_2_bF_buf0) );
  BUFX2 BUFX2_208 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_), .Y(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf5) );
  BUFX2 BUFX2_209 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_), .Y(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf4) );
  BUFX2 BUFX2_21 ( .A(sdram_clk), .Y(sdram_clk_hier0_bF_buf2) );
  BUFX2 BUFX2_210 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_), .Y(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf3) );
  BUFX2 BUFX2_211 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_), .Y(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf2) );
  BUFX2 BUFX2_212 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_), .Y(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf1) );
  BUFX2 BUFX2_213 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_), .Y(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf0) );
  BUFX2 BUFX2_214 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf5) );
  BUFX2 BUFX2_215 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf4) );
  BUFX2 BUFX2_216 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf3) );
  BUFX2 BUFX2_217 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf2) );
  BUFX2 BUFX2_218 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf1) );
  BUFX2 BUFX2_219 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf0) );
  BUFX2 BUFX2_22 ( .A(sdram_clk), .Y(sdram_clk_hier0_bF_buf1) );
  BUFX2 BUFX2_220 ( .A(u_sdrc_core_u_req_gen__abc_22171_n335_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n335_1_bF_buf3) );
  BUFX2 BUFX2_221 ( .A(u_sdrc_core_u_req_gen__abc_22171_n335_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n335_1_bF_buf2) );
  BUFX2 BUFX2_222 ( .A(u_sdrc_core_u_req_gen__abc_22171_n335_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n335_1_bF_buf1) );
  BUFX2 BUFX2_223 ( .A(u_sdrc_core_u_req_gen__abc_22171_n335_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n335_1_bF_buf0) );
  BUFX2 BUFX2_224 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf5) );
  BUFX2 BUFX2_225 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf4) );
  BUFX2 BUFX2_226 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf3) );
  BUFX2 BUFX2_227 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf2) );
  BUFX2 BUFX2_228 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf1) );
  BUFX2 BUFX2_229 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf0) );
  BUFX2 BUFX2_23 ( .A(sdram_clk), .Y(sdram_clk_hier0_bF_buf0) );
  BUFX2 BUFX2_230 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1020), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf4) );
  BUFX2 BUFX2_231 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1020), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf3) );
  BUFX2 BUFX2_232 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1020), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf2) );
  BUFX2 BUFX2_233 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1020), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf1) );
  BUFX2 BUFX2_234 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1020), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf0) );
  BUFX2 BUFX2_235 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_), .Y(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf5) );
  BUFX2 BUFX2_236 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_), .Y(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf4) );
  BUFX2 BUFX2_237 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_), .Y(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf3) );
  BUFX2 BUFX2_238 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_), .Y(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf2) );
  BUFX2 BUFX2_239 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_), .Y(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf1) );
  BUFX2 BUFX2_24 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_), .Y(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf7) );
  BUFX2 BUFX2_240 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_), .Y(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf0) );
  BUFX2 BUFX2_241 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n171_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n171_1_bF_buf3) );
  BUFX2 BUFX2_242 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n171_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n171_1_bF_buf2) );
  BUFX2 BUFX2_243 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n171_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n171_1_bF_buf1) );
  BUFX2 BUFX2_244 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n171_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n171_1_bF_buf0) );
  BUFX2 BUFX2_245 ( .A(sdram_resetn_hier0_bF_buf6), .Y(sdram_resetn_bF_buf49) );
  BUFX2 BUFX2_246 ( .A(sdram_resetn_hier0_bF_buf5), .Y(sdram_resetn_bF_buf48) );
  BUFX2 BUFX2_247 ( .A(sdram_resetn_hier0_bF_buf4), .Y(sdram_resetn_bF_buf47) );
  BUFX2 BUFX2_248 ( .A(sdram_resetn_hier0_bF_buf3), .Y(sdram_resetn_bF_buf46) );
  BUFX2 BUFX2_249 ( .A(sdram_resetn_hier0_bF_buf2), .Y(sdram_resetn_bF_buf45) );
  BUFX2 BUFX2_25 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_), .Y(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf6) );
  BUFX2 BUFX2_250 ( .A(sdram_resetn_hier0_bF_buf1), .Y(sdram_resetn_bF_buf44) );
  BUFX2 BUFX2_251 ( .A(sdram_resetn_hier0_bF_buf0), .Y(sdram_resetn_bF_buf43) );
  BUFX2 BUFX2_252 ( .A(sdram_resetn_hier0_bF_buf6), .Y(sdram_resetn_bF_buf42) );
  BUFX2 BUFX2_253 ( .A(sdram_resetn_hier0_bF_buf5), .Y(sdram_resetn_bF_buf41) );
  BUFX2 BUFX2_254 ( .A(sdram_resetn_hier0_bF_buf4), .Y(sdram_resetn_bF_buf40) );
  BUFX2 BUFX2_255 ( .A(sdram_resetn_hier0_bF_buf3), .Y(sdram_resetn_bF_buf39) );
  BUFX2 BUFX2_256 ( .A(sdram_resetn_hier0_bF_buf2), .Y(sdram_resetn_bF_buf38) );
  BUFX2 BUFX2_257 ( .A(sdram_resetn_hier0_bF_buf1), .Y(sdram_resetn_bF_buf37) );
  BUFX2 BUFX2_258 ( .A(sdram_resetn_hier0_bF_buf0), .Y(sdram_resetn_bF_buf36) );
  BUFX2 BUFX2_259 ( .A(sdram_resetn_hier0_bF_buf6), .Y(sdram_resetn_bF_buf35) );
  BUFX2 BUFX2_26 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_), .Y(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf5) );
  BUFX2 BUFX2_260 ( .A(sdram_resetn_hier0_bF_buf5), .Y(sdram_resetn_bF_buf34) );
  BUFX2 BUFX2_261 ( .A(sdram_resetn_hier0_bF_buf4), .Y(sdram_resetn_bF_buf33) );
  BUFX2 BUFX2_262 ( .A(sdram_resetn_hier0_bF_buf3), .Y(sdram_resetn_bF_buf32) );
  BUFX2 BUFX2_263 ( .A(sdram_resetn_hier0_bF_buf2), .Y(sdram_resetn_bF_buf31) );
  BUFX2 BUFX2_264 ( .A(sdram_resetn_hier0_bF_buf1), .Y(sdram_resetn_bF_buf30) );
  BUFX2 BUFX2_265 ( .A(sdram_resetn_hier0_bF_buf0), .Y(sdram_resetn_bF_buf29) );
  BUFX2 BUFX2_266 ( .A(sdram_resetn_hier0_bF_buf6), .Y(sdram_resetn_bF_buf28) );
  BUFX2 BUFX2_267 ( .A(sdram_resetn_hier0_bF_buf5), .Y(sdram_resetn_bF_buf27) );
  BUFX2 BUFX2_268 ( .A(sdram_resetn_hier0_bF_buf4), .Y(sdram_resetn_bF_buf26) );
  BUFX2 BUFX2_269 ( .A(sdram_resetn_hier0_bF_buf3), .Y(sdram_resetn_bF_buf25) );
  BUFX2 BUFX2_27 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_), .Y(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf4) );
  BUFX2 BUFX2_270 ( .A(sdram_resetn_hier0_bF_buf2), .Y(sdram_resetn_bF_buf24) );
  BUFX2 BUFX2_271 ( .A(sdram_resetn_hier0_bF_buf1), .Y(sdram_resetn_bF_buf23) );
  BUFX2 BUFX2_272 ( .A(sdram_resetn_hier0_bF_buf0), .Y(sdram_resetn_bF_buf22) );
  BUFX2 BUFX2_273 ( .A(sdram_resetn_hier0_bF_buf6), .Y(sdram_resetn_bF_buf21) );
  BUFX2 BUFX2_274 ( .A(sdram_resetn_hier0_bF_buf5), .Y(sdram_resetn_bF_buf20) );
  BUFX2 BUFX2_275 ( .A(sdram_resetn_hier0_bF_buf4), .Y(sdram_resetn_bF_buf19) );
  BUFX2 BUFX2_276 ( .A(sdram_resetn_hier0_bF_buf3), .Y(sdram_resetn_bF_buf18) );
  BUFX2 BUFX2_277 ( .A(sdram_resetn_hier0_bF_buf2), .Y(sdram_resetn_bF_buf17) );
  BUFX2 BUFX2_278 ( .A(sdram_resetn_hier0_bF_buf1), .Y(sdram_resetn_bF_buf16) );
  BUFX2 BUFX2_279 ( .A(sdram_resetn_hier0_bF_buf0), .Y(sdram_resetn_bF_buf15) );
  BUFX2 BUFX2_28 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_), .Y(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf3) );
  BUFX2 BUFX2_280 ( .A(sdram_resetn_hier0_bF_buf6), .Y(sdram_resetn_bF_buf14) );
  BUFX2 BUFX2_281 ( .A(sdram_resetn_hier0_bF_buf5), .Y(sdram_resetn_bF_buf13) );
  BUFX2 BUFX2_282 ( .A(sdram_resetn_hier0_bF_buf4), .Y(sdram_resetn_bF_buf12) );
  BUFX2 BUFX2_283 ( .A(sdram_resetn_hier0_bF_buf3), .Y(sdram_resetn_bF_buf11) );
  BUFX2 BUFX2_284 ( .A(sdram_resetn_hier0_bF_buf2), .Y(sdram_resetn_bF_buf10) );
  BUFX2 BUFX2_285 ( .A(sdram_resetn_hier0_bF_buf1), .Y(sdram_resetn_bF_buf9) );
  BUFX2 BUFX2_286 ( .A(sdram_resetn_hier0_bF_buf0), .Y(sdram_resetn_bF_buf8) );
  BUFX2 BUFX2_287 ( .A(sdram_resetn_hier0_bF_buf6), .Y(sdram_resetn_bF_buf7) );
  BUFX2 BUFX2_288 ( .A(sdram_resetn_hier0_bF_buf5), .Y(sdram_resetn_bF_buf6) );
  BUFX2 BUFX2_289 ( .A(sdram_resetn_hier0_bF_buf4), .Y(sdram_resetn_bF_buf5) );
  BUFX2 BUFX2_29 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_), .Y(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf2) );
  BUFX2 BUFX2_290 ( .A(sdram_resetn_hier0_bF_buf3), .Y(sdram_resetn_bF_buf4) );
  BUFX2 BUFX2_291 ( .A(sdram_resetn_hier0_bF_buf2), .Y(sdram_resetn_bF_buf3) );
  BUFX2 BUFX2_292 ( .A(sdram_resetn_hier0_bF_buf1), .Y(sdram_resetn_bF_buf2) );
  BUFX2 BUFX2_293 ( .A(sdram_resetn_hier0_bF_buf0), .Y(sdram_resetn_bF_buf1) );
  BUFX2 BUFX2_294 ( .A(sdram_resetn_hier0_bF_buf6), .Y(sdram_resetn_bF_buf0) );
  BUFX2 BUFX2_295 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf5) );
  BUFX2 BUFX2_296 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf4) );
  BUFX2 BUFX2_297 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf3) );
  BUFX2 BUFX2_298 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf2) );
  BUFX2 BUFX2_299 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf1) );
  BUFX2 BUFX2_3 ( .A(sdram_resetn), .Y(sdram_resetn_hier0_bF_buf4) );
  BUFX2 BUFX2_30 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_), .Y(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf1) );
  BUFX2 BUFX2_300 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf0) );
  BUFX2 BUFX2_301 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf5) );
  BUFX2 BUFX2_302 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf4) );
  BUFX2 BUFX2_303 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf3) );
  BUFX2 BUFX2_304 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf2) );
  BUFX2 BUFX2_305 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf1) );
  BUFX2 BUFX2_306 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf0) );
  BUFX2 BUFX2_307 ( .A(wb_clk_i_hier0_bF_buf6), .Y(wb_clk_i_bF_buf59) );
  BUFX2 BUFX2_308 ( .A(wb_clk_i_hier0_bF_buf5), .Y(wb_clk_i_bF_buf58) );
  BUFX2 BUFX2_309 ( .A(wb_clk_i_hier0_bF_buf4), .Y(wb_clk_i_bF_buf57) );
  BUFX2 BUFX2_31 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_), .Y(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf0) );
  BUFX2 BUFX2_310 ( .A(wb_clk_i_hier0_bF_buf3), .Y(wb_clk_i_bF_buf56) );
  BUFX2 BUFX2_311 ( .A(wb_clk_i_hier0_bF_buf2), .Y(wb_clk_i_bF_buf55) );
  BUFX2 BUFX2_312 ( .A(wb_clk_i_hier0_bF_buf1), .Y(wb_clk_i_bF_buf54) );
  BUFX2 BUFX2_313 ( .A(wb_clk_i_hier0_bF_buf0), .Y(wb_clk_i_bF_buf53) );
  BUFX2 BUFX2_314 ( .A(wb_clk_i_hier0_bF_buf6), .Y(wb_clk_i_bF_buf52) );
  BUFX2 BUFX2_315 ( .A(wb_clk_i_hier0_bF_buf5), .Y(wb_clk_i_bF_buf51) );
  BUFX2 BUFX2_316 ( .A(wb_clk_i_hier0_bF_buf4), .Y(wb_clk_i_bF_buf50) );
  BUFX2 BUFX2_317 ( .A(wb_clk_i_hier0_bF_buf3), .Y(wb_clk_i_bF_buf49) );
  BUFX2 BUFX2_318 ( .A(wb_clk_i_hier0_bF_buf2), .Y(wb_clk_i_bF_buf48) );
  BUFX2 BUFX2_319 ( .A(wb_clk_i_hier0_bF_buf1), .Y(wb_clk_i_bF_buf47) );
  BUFX2 BUFX2_32 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf4) );
  BUFX2 BUFX2_320 ( .A(wb_clk_i_hier0_bF_buf0), .Y(wb_clk_i_bF_buf46) );
  BUFX2 BUFX2_321 ( .A(wb_clk_i_hier0_bF_buf6), .Y(wb_clk_i_bF_buf45) );
  BUFX2 BUFX2_322 ( .A(wb_clk_i_hier0_bF_buf5), .Y(wb_clk_i_bF_buf44) );
  BUFX2 BUFX2_323 ( .A(wb_clk_i_hier0_bF_buf4), .Y(wb_clk_i_bF_buf43) );
  BUFX2 BUFX2_324 ( .A(wb_clk_i_hier0_bF_buf3), .Y(wb_clk_i_bF_buf42) );
  BUFX2 BUFX2_325 ( .A(wb_clk_i_hier0_bF_buf2), .Y(wb_clk_i_bF_buf41) );
  BUFX2 BUFX2_326 ( .A(wb_clk_i_hier0_bF_buf1), .Y(wb_clk_i_bF_buf40) );
  BUFX2 BUFX2_327 ( .A(wb_clk_i_hier0_bF_buf0), .Y(wb_clk_i_bF_buf39) );
  BUFX2 BUFX2_328 ( .A(wb_clk_i_hier0_bF_buf6), .Y(wb_clk_i_bF_buf38) );
  BUFX2 BUFX2_329 ( .A(wb_clk_i_hier0_bF_buf5), .Y(wb_clk_i_bF_buf37) );
  BUFX2 BUFX2_33 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf3) );
  BUFX2 BUFX2_330 ( .A(wb_clk_i_hier0_bF_buf4), .Y(wb_clk_i_bF_buf36) );
  BUFX2 BUFX2_331 ( .A(wb_clk_i_hier0_bF_buf3), .Y(wb_clk_i_bF_buf35) );
  BUFX2 BUFX2_332 ( .A(wb_clk_i_hier0_bF_buf2), .Y(wb_clk_i_bF_buf34) );
  BUFX2 BUFX2_333 ( .A(wb_clk_i_hier0_bF_buf1), .Y(wb_clk_i_bF_buf33) );
  BUFX2 BUFX2_334 ( .A(wb_clk_i_hier0_bF_buf0), .Y(wb_clk_i_bF_buf32) );
  BUFX2 BUFX2_335 ( .A(wb_clk_i_hier0_bF_buf6), .Y(wb_clk_i_bF_buf31) );
  BUFX2 BUFX2_336 ( .A(wb_clk_i_hier0_bF_buf5), .Y(wb_clk_i_bF_buf30) );
  BUFX2 BUFX2_337 ( .A(wb_clk_i_hier0_bF_buf4), .Y(wb_clk_i_bF_buf29) );
  BUFX2 BUFX2_338 ( .A(wb_clk_i_hier0_bF_buf3), .Y(wb_clk_i_bF_buf28) );
  BUFX2 BUFX2_339 ( .A(wb_clk_i_hier0_bF_buf2), .Y(wb_clk_i_bF_buf27) );
  BUFX2 BUFX2_34 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf2) );
  BUFX2 BUFX2_340 ( .A(wb_clk_i_hier0_bF_buf1), .Y(wb_clk_i_bF_buf26) );
  BUFX2 BUFX2_341 ( .A(wb_clk_i_hier0_bF_buf0), .Y(wb_clk_i_bF_buf25) );
  BUFX2 BUFX2_342 ( .A(wb_clk_i_hier0_bF_buf6), .Y(wb_clk_i_bF_buf24) );
  BUFX2 BUFX2_343 ( .A(wb_clk_i_hier0_bF_buf5), .Y(wb_clk_i_bF_buf23) );
  BUFX2 BUFX2_344 ( .A(wb_clk_i_hier0_bF_buf4), .Y(wb_clk_i_bF_buf22) );
  BUFX2 BUFX2_345 ( .A(wb_clk_i_hier0_bF_buf3), .Y(wb_clk_i_bF_buf21) );
  BUFX2 BUFX2_346 ( .A(wb_clk_i_hier0_bF_buf2), .Y(wb_clk_i_bF_buf20) );
  BUFX2 BUFX2_347 ( .A(wb_clk_i_hier0_bF_buf1), .Y(wb_clk_i_bF_buf19) );
  BUFX2 BUFX2_348 ( .A(wb_clk_i_hier0_bF_buf0), .Y(wb_clk_i_bF_buf18) );
  BUFX2 BUFX2_349 ( .A(wb_clk_i_hier0_bF_buf6), .Y(wb_clk_i_bF_buf17) );
  BUFX2 BUFX2_35 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf1) );
  BUFX2 BUFX2_350 ( .A(wb_clk_i_hier0_bF_buf5), .Y(wb_clk_i_bF_buf16) );
  BUFX2 BUFX2_351 ( .A(wb_clk_i_hier0_bF_buf4), .Y(wb_clk_i_bF_buf15) );
  BUFX2 BUFX2_352 ( .A(wb_clk_i_hier0_bF_buf3), .Y(wb_clk_i_bF_buf14) );
  BUFX2 BUFX2_353 ( .A(wb_clk_i_hier0_bF_buf2), .Y(wb_clk_i_bF_buf13) );
  BUFX2 BUFX2_354 ( .A(wb_clk_i_hier0_bF_buf1), .Y(wb_clk_i_bF_buf12) );
  BUFX2 BUFX2_355 ( .A(wb_clk_i_hier0_bF_buf0), .Y(wb_clk_i_bF_buf11) );
  BUFX2 BUFX2_356 ( .A(wb_clk_i_hier0_bF_buf6), .Y(wb_clk_i_bF_buf10) );
  BUFX2 BUFX2_357 ( .A(wb_clk_i_hier0_bF_buf5), .Y(wb_clk_i_bF_buf9) );
  BUFX2 BUFX2_358 ( .A(wb_clk_i_hier0_bF_buf4), .Y(wb_clk_i_bF_buf8) );
  BUFX2 BUFX2_359 ( .A(wb_clk_i_hier0_bF_buf3), .Y(wb_clk_i_bF_buf7) );
  BUFX2 BUFX2_36 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf0) );
  BUFX2 BUFX2_360 ( .A(wb_clk_i_hier0_bF_buf2), .Y(wb_clk_i_bF_buf6) );
  BUFX2 BUFX2_361 ( .A(wb_clk_i_hier0_bF_buf1), .Y(wb_clk_i_bF_buf5) );
  BUFX2 BUFX2_362 ( .A(wb_clk_i_hier0_bF_buf0), .Y(wb_clk_i_bF_buf4) );
  BUFX2 BUFX2_363 ( .A(wb_clk_i_hier0_bF_buf6), .Y(wb_clk_i_bF_buf3) );
  BUFX2 BUFX2_364 ( .A(wb_clk_i_hier0_bF_buf5), .Y(wb_clk_i_bF_buf2) );
  BUFX2 BUFX2_365 ( .A(wb_clk_i_hier0_bF_buf4), .Y(wb_clk_i_bF_buf1) );
  BUFX2 BUFX2_366 ( .A(wb_clk_i_hier0_bF_buf3), .Y(wb_clk_i_bF_buf0) );
  BUFX2 BUFX2_367 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf5) );
  BUFX2 BUFX2_368 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf4) );
  BUFX2 BUFX2_369 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf3) );
  BUFX2 BUFX2_37 ( .A(u_sdrc_core_u_req_gen__abc_22171_n893), .Y(u_sdrc_core_u_req_gen__abc_22171_n893_bF_buf3) );
  BUFX2 BUFX2_370 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf2) );
  BUFX2 BUFX2_371 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf1) );
  BUFX2 BUFX2_372 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf0) );
  BUFX2 BUFX2_373 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n223_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n223_1_bF_buf3) );
  BUFX2 BUFX2_374 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n223_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n223_1_bF_buf2) );
  BUFX2 BUFX2_375 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n223_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n223_1_bF_buf1) );
  BUFX2 BUFX2_376 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n223_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n223_1_bF_buf0) );
  BUFX2 BUFX2_377 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf4) );
  BUFX2 BUFX2_378 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf3) );
  BUFX2 BUFX2_379 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf2) );
  BUFX2 BUFX2_38 ( .A(u_sdrc_core_u_req_gen__abc_22171_n893), .Y(u_sdrc_core_u_req_gen__abc_22171_n893_bF_buf2) );
  BUFX2 BUFX2_380 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf1) );
  BUFX2 BUFX2_381 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf0) );
  BUFX2 BUFX2_382 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n551), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf4) );
  BUFX2 BUFX2_383 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n551), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf3) );
  BUFX2 BUFX2_384 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n551), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf2) );
  BUFX2 BUFX2_385 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n551), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf1) );
  BUFX2 BUFX2_386 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n551), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf0) );
  BUFX2 BUFX2_387 ( .A(app_req_ack), .Y(app_req_ack_bF_buf6) );
  BUFX2 BUFX2_388 ( .A(app_req_ack), .Y(app_req_ack_bF_buf5) );
  BUFX2 BUFX2_389 ( .A(app_req_ack), .Y(app_req_ack_bF_buf4) );
  BUFX2 BUFX2_39 ( .A(u_sdrc_core_u_req_gen__abc_22171_n893), .Y(u_sdrc_core_u_req_gen__abc_22171_n893_bF_buf1) );
  BUFX2 BUFX2_390 ( .A(app_req_ack), .Y(app_req_ack_bF_buf3) );
  BUFX2 BUFX2_391 ( .A(app_req_ack), .Y(app_req_ack_bF_buf2) );
  BUFX2 BUFX2_392 ( .A(app_req_ack), .Y(app_req_ack_bF_buf1) );
  BUFX2 BUFX2_393 ( .A(app_req_ack), .Y(app_req_ack_bF_buf0) );
  BUFX2 BUFX2_394 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf5) );
  BUFX2 BUFX2_395 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf4) );
  BUFX2 BUFX2_396 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf3) );
  BUFX2 BUFX2_397 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf2) );
  BUFX2 BUFX2_398 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf1) );
  BUFX2 BUFX2_399 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf0) );
  BUFX2 BUFX2_4 ( .A(sdram_resetn), .Y(sdram_resetn_hier0_bF_buf3) );
  BUFX2 BUFX2_40 ( .A(u_sdrc_core_u_req_gen__abc_22171_n893), .Y(u_sdrc_core_u_req_gen__abc_22171_n893_bF_buf0) );
  BUFX2 BUFX2_400 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_4_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_4_bF_buf3) );
  BUFX2 BUFX2_401 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_4_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_4_bF_buf2) );
  BUFX2 BUFX2_402 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_4_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_4_bF_buf1) );
  BUFX2 BUFX2_403 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_4_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_4_bF_buf0) );
  BUFX2 BUFX2_404 ( .A(sdram_clk_hier0_bF_buf8), .Y(sdram_clk_bF_buf80) );
  BUFX2 BUFX2_405 ( .A(sdram_clk_hier0_bF_buf7), .Y(sdram_clk_bF_buf79) );
  BUFX2 BUFX2_406 ( .A(sdram_clk_hier0_bF_buf6), .Y(sdram_clk_bF_buf78) );
  BUFX2 BUFX2_407 ( .A(sdram_clk_hier0_bF_buf5), .Y(sdram_clk_bF_buf77) );
  BUFX2 BUFX2_408 ( .A(sdram_clk_hier0_bF_buf4), .Y(sdram_clk_bF_buf76) );
  BUFX2 BUFX2_409 ( .A(sdram_clk_hier0_bF_buf3), .Y(sdram_clk_bF_buf75) );
  BUFX2 BUFX2_41 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf4) );
  BUFX2 BUFX2_410 ( .A(sdram_clk_hier0_bF_buf2), .Y(sdram_clk_bF_buf74) );
  BUFX2 BUFX2_411 ( .A(sdram_clk_hier0_bF_buf1), .Y(sdram_clk_bF_buf73) );
  BUFX2 BUFX2_412 ( .A(sdram_clk_hier0_bF_buf0), .Y(sdram_clk_bF_buf72) );
  BUFX2 BUFX2_413 ( .A(sdram_clk_hier0_bF_buf8), .Y(sdram_clk_bF_buf71) );
  BUFX2 BUFX2_414 ( .A(sdram_clk_hier0_bF_buf7), .Y(sdram_clk_bF_buf70) );
  BUFX2 BUFX2_415 ( .A(sdram_clk_hier0_bF_buf6), .Y(sdram_clk_bF_buf69) );
  BUFX2 BUFX2_416 ( .A(sdram_clk_hier0_bF_buf5), .Y(sdram_clk_bF_buf68) );
  BUFX2 BUFX2_417 ( .A(sdram_clk_hier0_bF_buf4), .Y(sdram_clk_bF_buf67) );
  BUFX2 BUFX2_418 ( .A(sdram_clk_hier0_bF_buf3), .Y(sdram_clk_bF_buf66) );
  BUFX2 BUFX2_419 ( .A(sdram_clk_hier0_bF_buf2), .Y(sdram_clk_bF_buf65) );
  BUFX2 BUFX2_42 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf3) );
  BUFX2 BUFX2_420 ( .A(sdram_clk_hier0_bF_buf1), .Y(sdram_clk_bF_buf64) );
  BUFX2 BUFX2_421 ( .A(sdram_clk_hier0_bF_buf0), .Y(sdram_clk_bF_buf63) );
  BUFX2 BUFX2_422 ( .A(sdram_clk_hier0_bF_buf8), .Y(sdram_clk_bF_buf62) );
  BUFX2 BUFX2_423 ( .A(sdram_clk_hier0_bF_buf7), .Y(sdram_clk_bF_buf61) );
  BUFX2 BUFX2_424 ( .A(sdram_clk_hier0_bF_buf6), .Y(sdram_clk_bF_buf60) );
  BUFX2 BUFX2_425 ( .A(sdram_clk_hier0_bF_buf5), .Y(sdram_clk_bF_buf59) );
  BUFX2 BUFX2_426 ( .A(sdram_clk_hier0_bF_buf4), .Y(sdram_clk_bF_buf58) );
  BUFX2 BUFX2_427 ( .A(sdram_clk_hier0_bF_buf3), .Y(sdram_clk_bF_buf57) );
  BUFX2 BUFX2_428 ( .A(sdram_clk_hier0_bF_buf2), .Y(sdram_clk_bF_buf56) );
  BUFX2 BUFX2_429 ( .A(sdram_clk_hier0_bF_buf1), .Y(sdram_clk_bF_buf55) );
  BUFX2 BUFX2_43 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf2) );
  BUFX2 BUFX2_430 ( .A(sdram_clk_hier0_bF_buf0), .Y(sdram_clk_bF_buf54) );
  BUFX2 BUFX2_431 ( .A(sdram_clk_hier0_bF_buf8), .Y(sdram_clk_bF_buf53) );
  BUFX2 BUFX2_432 ( .A(sdram_clk_hier0_bF_buf7), .Y(sdram_clk_bF_buf52) );
  BUFX2 BUFX2_433 ( .A(sdram_clk_hier0_bF_buf6), .Y(sdram_clk_bF_buf51) );
  BUFX2 BUFX2_434 ( .A(sdram_clk_hier0_bF_buf5), .Y(sdram_clk_bF_buf50) );
  BUFX2 BUFX2_435 ( .A(sdram_clk_hier0_bF_buf4), .Y(sdram_clk_bF_buf49) );
  BUFX2 BUFX2_436 ( .A(sdram_clk_hier0_bF_buf3), .Y(sdram_clk_bF_buf48) );
  BUFX2 BUFX2_437 ( .A(sdram_clk_hier0_bF_buf2), .Y(sdram_clk_bF_buf47) );
  BUFX2 BUFX2_438 ( .A(sdram_clk_hier0_bF_buf1), .Y(sdram_clk_bF_buf46) );
  BUFX2 BUFX2_439 ( .A(sdram_clk_hier0_bF_buf0), .Y(sdram_clk_bF_buf45) );
  BUFX2 BUFX2_44 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf1) );
  BUFX2 BUFX2_440 ( .A(sdram_clk_hier0_bF_buf8), .Y(sdram_clk_bF_buf44) );
  BUFX2 BUFX2_441 ( .A(sdram_clk_hier0_bF_buf7), .Y(sdram_clk_bF_buf43) );
  BUFX2 BUFX2_442 ( .A(sdram_clk_hier0_bF_buf6), .Y(sdram_clk_bF_buf42) );
  BUFX2 BUFX2_443 ( .A(sdram_clk_hier0_bF_buf5), .Y(sdram_clk_bF_buf41) );
  BUFX2 BUFX2_444 ( .A(sdram_clk_hier0_bF_buf4), .Y(sdram_clk_bF_buf40) );
  BUFX2 BUFX2_445 ( .A(sdram_clk_hier0_bF_buf3), .Y(sdram_clk_bF_buf39) );
  BUFX2 BUFX2_446 ( .A(sdram_clk_hier0_bF_buf2), .Y(sdram_clk_bF_buf38) );
  BUFX2 BUFX2_447 ( .A(sdram_clk_hier0_bF_buf1), .Y(sdram_clk_bF_buf37) );
  BUFX2 BUFX2_448 ( .A(sdram_clk_hier0_bF_buf0), .Y(sdram_clk_bF_buf36) );
  BUFX2 BUFX2_449 ( .A(sdram_clk_hier0_bF_buf8), .Y(sdram_clk_bF_buf35) );
  BUFX2 BUFX2_45 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf0) );
  BUFX2 BUFX2_450 ( .A(sdram_clk_hier0_bF_buf7), .Y(sdram_clk_bF_buf34) );
  BUFX2 BUFX2_451 ( .A(sdram_clk_hier0_bF_buf6), .Y(sdram_clk_bF_buf33) );
  BUFX2 BUFX2_452 ( .A(sdram_clk_hier0_bF_buf5), .Y(sdram_clk_bF_buf32) );
  BUFX2 BUFX2_453 ( .A(sdram_clk_hier0_bF_buf4), .Y(sdram_clk_bF_buf31) );
  BUFX2 BUFX2_454 ( .A(sdram_clk_hier0_bF_buf3), .Y(sdram_clk_bF_buf30) );
  BUFX2 BUFX2_455 ( .A(sdram_clk_hier0_bF_buf2), .Y(sdram_clk_bF_buf29) );
  BUFX2 BUFX2_456 ( .A(sdram_clk_hier0_bF_buf1), .Y(sdram_clk_bF_buf28) );
  BUFX2 BUFX2_457 ( .A(sdram_clk_hier0_bF_buf0), .Y(sdram_clk_bF_buf27) );
  BUFX2 BUFX2_458 ( .A(sdram_clk_hier0_bF_buf8), .Y(sdram_clk_bF_buf26) );
  BUFX2 BUFX2_459 ( .A(sdram_clk_hier0_bF_buf7), .Y(sdram_clk_bF_buf25) );
  BUFX2 BUFX2_46 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n652), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf4) );
  BUFX2 BUFX2_460 ( .A(sdram_clk_hier0_bF_buf6), .Y(sdram_clk_bF_buf24) );
  BUFX2 BUFX2_461 ( .A(sdram_clk_hier0_bF_buf5), .Y(sdram_clk_bF_buf23) );
  BUFX2 BUFX2_462 ( .A(sdram_clk_hier0_bF_buf4), .Y(sdram_clk_bF_buf22) );
  BUFX2 BUFX2_463 ( .A(sdram_clk_hier0_bF_buf3), .Y(sdram_clk_bF_buf21) );
  BUFX2 BUFX2_464 ( .A(sdram_clk_hier0_bF_buf2), .Y(sdram_clk_bF_buf20) );
  BUFX2 BUFX2_465 ( .A(sdram_clk_hier0_bF_buf1), .Y(sdram_clk_bF_buf19) );
  BUFX2 BUFX2_466 ( .A(sdram_clk_hier0_bF_buf0), .Y(sdram_clk_bF_buf18) );
  BUFX2 BUFX2_467 ( .A(sdram_clk_hier0_bF_buf8), .Y(sdram_clk_bF_buf17) );
  BUFX2 BUFX2_468 ( .A(sdram_clk_hier0_bF_buf7), .Y(sdram_clk_bF_buf16) );
  BUFX2 BUFX2_469 ( .A(sdram_clk_hier0_bF_buf6), .Y(sdram_clk_bF_buf15) );
  BUFX2 BUFX2_47 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n652), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf3) );
  BUFX2 BUFX2_470 ( .A(sdram_clk_hier0_bF_buf5), .Y(sdram_clk_bF_buf14) );
  BUFX2 BUFX2_471 ( .A(sdram_clk_hier0_bF_buf4), .Y(sdram_clk_bF_buf13) );
  BUFX2 BUFX2_472 ( .A(sdram_clk_hier0_bF_buf3), .Y(sdram_clk_bF_buf12) );
  BUFX2 BUFX2_473 ( .A(sdram_clk_hier0_bF_buf2), .Y(sdram_clk_bF_buf11) );
  BUFX2 BUFX2_474 ( .A(sdram_clk_hier0_bF_buf1), .Y(sdram_clk_bF_buf10) );
  BUFX2 BUFX2_475 ( .A(sdram_clk_hier0_bF_buf0), .Y(sdram_clk_bF_buf9) );
  BUFX2 BUFX2_476 ( .A(sdram_clk_hier0_bF_buf8), .Y(sdram_clk_bF_buf8) );
  BUFX2 BUFX2_477 ( .A(sdram_clk_hier0_bF_buf7), .Y(sdram_clk_bF_buf7) );
  BUFX2 BUFX2_478 ( .A(sdram_clk_hier0_bF_buf6), .Y(sdram_clk_bF_buf6) );
  BUFX2 BUFX2_479 ( .A(sdram_clk_hier0_bF_buf5), .Y(sdram_clk_bF_buf5) );
  BUFX2 BUFX2_48 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n652), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf2) );
  BUFX2 BUFX2_480 ( .A(sdram_clk_hier0_bF_buf4), .Y(sdram_clk_bF_buf4) );
  BUFX2 BUFX2_481 ( .A(sdram_clk_hier0_bF_buf3), .Y(sdram_clk_bF_buf3) );
  BUFX2 BUFX2_482 ( .A(sdram_clk_hier0_bF_buf2), .Y(sdram_clk_bF_buf2) );
  BUFX2 BUFX2_483 ( .A(sdram_clk_hier0_bF_buf1), .Y(sdram_clk_bF_buf1) );
  BUFX2 BUFX2_484 ( .A(sdram_clk_hier0_bF_buf0), .Y(sdram_clk_bF_buf0) );
  BUFX2 BUFX2_485 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf5) );
  BUFX2 BUFX2_486 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf4) );
  BUFX2 BUFX2_487 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf3) );
  BUFX2 BUFX2_488 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf2) );
  BUFX2 BUFX2_489 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf1) );
  BUFX2 BUFX2_49 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n652), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf1) );
  BUFX2 BUFX2_490 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf0) );
  BUFX2 BUFX2_491 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n614), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n614_bF_buf3) );
  BUFX2 BUFX2_492 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n614), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n614_bF_buf2) );
  BUFX2 BUFX2_493 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n614), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n614_bF_buf1) );
  BUFX2 BUFX2_494 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n614), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n614_bF_buf0) );
  BUFX2 BUFX2_495 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_1_), .Y(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf5) );
  BUFX2 BUFX2_496 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_1_), .Y(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf4) );
  BUFX2 BUFX2_497 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_1_), .Y(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf3) );
  BUFX2 BUFX2_498 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_1_), .Y(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf2) );
  BUFX2 BUFX2_499 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_1_), .Y(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf1) );
  BUFX2 BUFX2_5 ( .A(sdram_resetn), .Y(sdram_resetn_hier0_bF_buf2) );
  BUFX2 BUFX2_50 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n652), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf0) );
  BUFX2 BUFX2_500 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_1_), .Y(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf0) );
  BUFX2 BUFX2_501 ( .A(u_sdrc_core_u_req_gen__abc_22171_n245_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf4) );
  BUFX2 BUFX2_502 ( .A(u_sdrc_core_u_req_gen__abc_22171_n245_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf3) );
  BUFX2 BUFX2_503 ( .A(u_sdrc_core_u_req_gen__abc_22171_n245_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf2) );
  BUFX2 BUFX2_504 ( .A(u_sdrc_core_u_req_gen__abc_22171_n245_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf1) );
  BUFX2 BUFX2_505 ( .A(u_sdrc_core_u_req_gen__abc_22171_n245_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf0) );
  BUFX2 BUFX2_506 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf5) );
  BUFX2 BUFX2_507 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf4) );
  BUFX2 BUFX2_508 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf3) );
  BUFX2 BUFX2_509 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf2) );
  BUFX2 BUFX2_51 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf5) );
  BUFX2 BUFX2_510 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf1) );
  BUFX2 BUFX2_511 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1_bF_buf0) );
  BUFX2 BUFX2_512 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n283), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n283_bF_buf3) );
  BUFX2 BUFX2_513 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n283), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n283_bF_buf2) );
  BUFX2 BUFX2_514 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n283), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n283_bF_buf1) );
  BUFX2 BUFX2_515 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n283), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n283_bF_buf0) );
  BUFX2 BUFX2_516 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n409), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf4) );
  BUFX2 BUFX2_517 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n409), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf3) );
  BUFX2 BUFX2_518 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n409), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf2) );
  BUFX2 BUFX2_519 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n409), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf1) );
  BUFX2 BUFX2_52 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf4) );
  BUFX2 BUFX2_520 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n409), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n409_bF_buf0) );
  BUFX2 BUFX2_521 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n227), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n227_bF_buf3) );
  BUFX2 BUFX2_522 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n227), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n227_bF_buf2) );
  BUFX2 BUFX2_523 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n227), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n227_bF_buf1) );
  BUFX2 BUFX2_524 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n227), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n227_bF_buf0) );
  BUFX2 BUFX2_525 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf5) );
  BUFX2 BUFX2_526 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf4) );
  BUFX2 BUFX2_527 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf3) );
  BUFX2 BUFX2_528 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf2) );
  BUFX2 BUFX2_529 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf1) );
  BUFX2 BUFX2_53 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf3) );
  BUFX2 BUFX2_530 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf0) );
  BUFX2 BUFX2_531 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf4) );
  BUFX2 BUFX2_532 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf3) );
  BUFX2 BUFX2_533 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf2) );
  BUFX2 BUFX2_534 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf1) );
  BUFX2 BUFX2_535 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf0) );
  BUFX2 BUFX2_536 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf4) );
  BUFX2 BUFX2_537 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf3) );
  BUFX2 BUFX2_538 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf2) );
  BUFX2 BUFX2_539 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf1) );
  BUFX2 BUFX2_54 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf2) );
  BUFX2 BUFX2_540 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf0) );
  BUFX2 BUFX2_541 ( .A(u_sdrc_core_u_bank_ctl_x2b_ack), .Y(u_sdrc_core_u_bank_ctl_x2b_ack_bF_buf3) );
  BUFX2 BUFX2_542 ( .A(u_sdrc_core_u_bank_ctl_x2b_ack), .Y(u_sdrc_core_u_bank_ctl_x2b_ack_bF_buf2) );
  BUFX2 BUFX2_543 ( .A(u_sdrc_core_u_bank_ctl_x2b_ack), .Y(u_sdrc_core_u_bank_ctl_x2b_ack_bF_buf1) );
  BUFX2 BUFX2_544 ( .A(u_sdrc_core_u_bank_ctl_x2b_ack), .Y(u_sdrc_core_u_bank_ctl_x2b_ack_bF_buf0) );
  BUFX2 BUFX2_545 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_4_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_4_bF_buf3) );
  BUFX2 BUFX2_546 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_4_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_4_bF_buf2) );
  BUFX2 BUFX2_547 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_4_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_4_bF_buf1) );
  BUFX2 BUFX2_548 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_4_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_4_bF_buf0) );
  BUFX2 BUFX2_549 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf4) );
  BUFX2 BUFX2_55 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf1) );
  BUFX2 BUFX2_550 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf3) );
  BUFX2 BUFX2_551 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf2) );
  BUFX2 BUFX2_552 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf1) );
  BUFX2 BUFX2_553 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf0) );
  BUFX2 BUFX2_554 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf4) );
  BUFX2 BUFX2_555 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf3) );
  BUFX2 BUFX2_556 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf2) );
  BUFX2 BUFX2_557 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf1) );
  BUFX2 BUFX2_558 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf0) );
  BUFX2 BUFX2_559 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf5) );
  BUFX2 BUFX2_56 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1_bF_buf0) );
  BUFX2 BUFX2_560 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf4) );
  BUFX2 BUFX2_561 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf3) );
  BUFX2 BUFX2_562 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf2) );
  BUFX2 BUFX2_563 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf1) );
  BUFX2 BUFX2_564 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf0) );
  BUFX2 BUFX2_565 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf4) );
  BUFX2 BUFX2_566 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf3) );
  BUFX2 BUFX2_567 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf2) );
  BUFX2 BUFX2_568 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf1) );
  BUFX2 BUFX2_569 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf0) );
  BUFX2 BUFX2_57 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_4_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_4_bF_buf3) );
  BUFX2 BUFX2_570 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n405_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n405_1_bF_buf3) );
  BUFX2 BUFX2_571 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n405_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n405_1_bF_buf2) );
  BUFX2 BUFX2_572 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n405_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n405_1_bF_buf1) );
  BUFX2 BUFX2_573 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n405_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n405_1_bF_buf0) );
  BUFX2 BUFX2_574 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf5) );
  BUFX2 BUFX2_575 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf4) );
  BUFX2 BUFX2_576 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf3) );
  BUFX2 BUFX2_577 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf2) );
  BUFX2 BUFX2_578 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf1) );
  BUFX2 BUFX2_579 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf0) );
  BUFX2 BUFX2_58 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_4_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_4_bF_buf2) );
  BUFX2 BUFX2_580 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf4) );
  BUFX2 BUFX2_581 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf3) );
  BUFX2 BUFX2_582 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf2) );
  BUFX2 BUFX2_583 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf1) );
  BUFX2 BUFX2_584 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf0) );
  BUFX2 BUFX2_585 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_2_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_2_bF_buf3) );
  BUFX2 BUFX2_586 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_2_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_2_bF_buf2) );
  BUFX2 BUFX2_587 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_2_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_2_bF_buf1) );
  BUFX2 BUFX2_588 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_2_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_2_bF_buf0) );
  BUFX2 BUFX2_589 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf5) );
  BUFX2 BUFX2_59 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_4_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_4_bF_buf1) );
  BUFX2 BUFX2_590 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf4) );
  BUFX2 BUFX2_591 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf3) );
  BUFX2 BUFX2_592 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf2) );
  BUFX2 BUFX2_593 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf1) );
  BUFX2 BUFX2_594 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf0) );
  BUFX2 BUFX2_595 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf5) );
  BUFX2 BUFX2_596 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf4) );
  BUFX2 BUFX2_597 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf3) );
  BUFX2 BUFX2_598 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf2) );
  BUFX2 BUFX2_599 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf1) );
  BUFX2 BUFX2_6 ( .A(sdram_resetn), .Y(sdram_resetn_hier0_bF_buf1) );
  BUFX2 BUFX2_60 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_4_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_4_bF_buf0) );
  BUFX2 BUFX2_600 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1_bF_buf0) );
  BUFX2 BUFX2_601 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf4) );
  BUFX2 BUFX2_602 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf3) );
  BUFX2 BUFX2_603 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf2) );
  BUFX2 BUFX2_604 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf1) );
  BUFX2 BUFX2_605 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf0) );
  BUFX2 BUFX2_606 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n170_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n170_1_bF_buf3) );
  BUFX2 BUFX2_607 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n170_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n170_1_bF_buf2) );
  BUFX2 BUFX2_608 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n170_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n170_1_bF_buf1) );
  BUFX2 BUFX2_609 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n170_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n170_1_bF_buf0) );
  BUFX2 BUFX2_61 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf5) );
  BUFX2 BUFX2_610 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf4) );
  BUFX2 BUFX2_611 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf3) );
  BUFX2 BUFX2_612 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf2) );
  BUFX2 BUFX2_613 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf1) );
  BUFX2 BUFX2_614 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf0) );
  BUFX2 BUFX2_615 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf5) );
  BUFX2 BUFX2_616 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf4) );
  BUFX2 BUFX2_617 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf3) );
  BUFX2 BUFX2_618 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf2) );
  BUFX2 BUFX2_619 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf1) );
  BUFX2 BUFX2_62 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf4) );
  BUFX2 BUFX2_620 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf0) );
  BUFX2 BUFX2_621 ( .A(u_sdrc_core_u_bs_convert_x2a_wrnext), .Y(u_sdrc_core_u_bs_convert_x2a_wrnext_bF_buf3) );
  BUFX2 BUFX2_622 ( .A(u_sdrc_core_u_bs_convert_x2a_wrnext), .Y(u_sdrc_core_u_bs_convert_x2a_wrnext_bF_buf2) );
  BUFX2 BUFX2_623 ( .A(u_sdrc_core_u_bs_convert_x2a_wrnext), .Y(u_sdrc_core_u_bs_convert_x2a_wrnext_bF_buf1) );
  BUFX2 BUFX2_624 ( .A(u_sdrc_core_u_bs_convert_x2a_wrnext), .Y(u_sdrc_core_u_bs_convert_x2a_wrnext_bF_buf0) );
  BUFX2 BUFX2_625 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n602), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n602_bF_buf3) );
  BUFX2 BUFX2_626 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n602), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n602_bF_buf2) );
  BUFX2 BUFX2_627 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n602), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n602_bF_buf1) );
  BUFX2 BUFX2_628 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n602), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n602_bF_buf0) );
  BUFX2 BUFX2_629 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_), .Y(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf7) );
  BUFX2 BUFX2_63 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf3) );
  BUFX2 BUFX2_630 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_), .Y(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf6) );
  BUFX2 BUFX2_631 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_), .Y(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf5) );
  BUFX2 BUFX2_632 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_), .Y(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf4) );
  BUFX2 BUFX2_633 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_), .Y(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf3) );
  BUFX2 BUFX2_634 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_), .Y(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf2) );
  BUFX2 BUFX2_635 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_), .Y(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf1) );
  BUFX2 BUFX2_636 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_), .Y(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf0) );
  BUFX2 BUFX2_637 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n782), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf7) );
  BUFX2 BUFX2_638 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n782), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf6) );
  BUFX2 BUFX2_639 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n782), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf5) );
  BUFX2 BUFX2_64 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf2) );
  BUFX2 BUFX2_640 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n782), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf4) );
  BUFX2 BUFX2_641 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n782), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf3) );
  BUFX2 BUFX2_642 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n782), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf2) );
  BUFX2 BUFX2_643 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n782), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf1) );
  BUFX2 BUFX2_644 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n782), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n782_bF_buf0) );
  BUFX2 BUFX2_645 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf4) );
  BUFX2 BUFX2_646 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf3) );
  BUFX2 BUFX2_647 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf2) );
  BUFX2 BUFX2_648 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf1) );
  BUFX2 BUFX2_649 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf0) );
  BUFX2 BUFX2_65 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf1) );
  BUFX2 BUFX2_650 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf5) );
  BUFX2 BUFX2_651 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf4) );
  BUFX2 BUFX2_652 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf3) );
  BUFX2 BUFX2_653 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf2) );
  BUFX2 BUFX2_654 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf1) );
  BUFX2 BUFX2_655 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf0) );
  BUFX2 BUFX2_656 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf5) );
  BUFX2 BUFX2_657 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf4) );
  BUFX2 BUFX2_658 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf3) );
  BUFX2 BUFX2_659 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf2) );
  BUFX2 BUFX2_66 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf0) );
  BUFX2 BUFX2_660 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf1) );
  BUFX2 BUFX2_661 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363_bF_buf0) );
  BUFX2 BUFX2_662 ( .A(u_sdrc_core_u_req_gen__abc_22171_n318), .Y(u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf4) );
  BUFX2 BUFX2_663 ( .A(u_sdrc_core_u_req_gen__abc_22171_n318), .Y(u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf3) );
  BUFX2 BUFX2_664 ( .A(u_sdrc_core_u_req_gen__abc_22171_n318), .Y(u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf2) );
  BUFX2 BUFX2_665 ( .A(u_sdrc_core_u_req_gen__abc_22171_n318), .Y(u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf1) );
  BUFX2 BUFX2_666 ( .A(u_sdrc_core_u_req_gen__abc_22171_n318), .Y(u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf0) );
  BUFX2 BUFX2_667 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf7) );
  BUFX2 BUFX2_668 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf6) );
  BUFX2 BUFX2_669 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf5) );
  BUFX2 BUFX2_67 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf5) );
  BUFX2 BUFX2_670 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf4) );
  BUFX2 BUFX2_671 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf3) );
  BUFX2 BUFX2_672 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf2) );
  BUFX2 BUFX2_673 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf1) );
  BUFX2 BUFX2_674 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1_bF_buf0) );
  BUFX2 BUFX2_675 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_2_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_2_bF_buf3) );
  BUFX2 BUFX2_676 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_2_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_2_bF_buf2) );
  BUFX2 BUFX2_677 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_2_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_2_bF_buf1) );
  BUFX2 BUFX2_678 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_2_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_2_bF_buf0) );
  BUFX2 BUFX2_679 ( .A(u_wb2sdrc_u_cmdfifo_wr_reset_n), .Y(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf5) );
  BUFX2 BUFX2_68 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf4) );
  BUFX2 BUFX2_680 ( .A(u_wb2sdrc_u_cmdfifo_wr_reset_n), .Y(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf4) );
  BUFX2 BUFX2_681 ( .A(u_wb2sdrc_u_cmdfifo_wr_reset_n), .Y(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf3) );
  BUFX2 BUFX2_682 ( .A(u_wb2sdrc_u_cmdfifo_wr_reset_n), .Y(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf2) );
  BUFX2 BUFX2_683 ( .A(u_wb2sdrc_u_cmdfifo_wr_reset_n), .Y(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf1) );
  BUFX2 BUFX2_684 ( .A(u_wb2sdrc_u_cmdfifo_wr_reset_n), .Y(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf0) );
  BUFX2 BUFX2_685 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf5) );
  BUFX2 BUFX2_686 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf4) );
  BUFX2 BUFX2_687 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf3) );
  BUFX2 BUFX2_688 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf2) );
  BUFX2 BUFX2_689 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf1) );
  BUFX2 BUFX2_69 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf3) );
  BUFX2 BUFX2_690 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf0) );
  BUFX2 BUFX2_691 ( .A(\cfg_sdr_width[1] ), .Y(cfg_sdr_width_1_bF_buf5) );
  BUFX2 BUFX2_692 ( .A(\cfg_sdr_width[1] ), .Y(cfg_sdr_width_1_bF_buf4) );
  BUFX2 BUFX2_693 ( .A(\cfg_sdr_width[1] ), .Y(cfg_sdr_width_1_bF_buf3) );
  BUFX2 BUFX2_694 ( .A(\cfg_sdr_width[1] ), .Y(cfg_sdr_width_1_bF_buf2) );
  BUFX2 BUFX2_695 ( .A(\cfg_sdr_width[1] ), .Y(cfg_sdr_width_1_bF_buf1) );
  BUFX2 BUFX2_696 ( .A(\cfg_sdr_width[1] ), .Y(cfg_sdr_width_1_bF_buf0) );
  BUFX2 BUFX2_697 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf5) );
  BUFX2 BUFX2_698 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf4) );
  BUFX2 BUFX2_699 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf3) );
  BUFX2 BUFX2_7 ( .A(sdram_resetn), .Y(sdram_resetn_hier0_bF_buf0) );
  BUFX2 BUFX2_70 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf2) );
  BUFX2 BUFX2_700 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf2) );
  BUFX2 BUFX2_701 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf1) );
  BUFX2 BUFX2_702 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1_bF_buf0) );
  BUFX2 BUFX2_703 ( .A(_auto_iopadmap_cc_313_execute_24675_0_), .Y(\sdr_addr[0] ) );
  BUFX2 BUFX2_704 ( .A(_auto_iopadmap_cc_313_execute_24675_1_), .Y(\sdr_addr[1] ) );
  BUFX2 BUFX2_705 ( .A(_auto_iopadmap_cc_313_execute_24675_2_), .Y(\sdr_addr[2] ) );
  BUFX2 BUFX2_706 ( .A(_auto_iopadmap_cc_313_execute_24675_3_), .Y(\sdr_addr[3] ) );
  BUFX2 BUFX2_707 ( .A(_auto_iopadmap_cc_313_execute_24675_4_), .Y(\sdr_addr[4] ) );
  BUFX2 BUFX2_708 ( .A(_auto_iopadmap_cc_313_execute_24675_5_), .Y(\sdr_addr[5] ) );
  BUFX2 BUFX2_709 ( .A(_auto_iopadmap_cc_313_execute_24675_6_), .Y(\sdr_addr[6] ) );
  BUFX2 BUFX2_71 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf1) );
  BUFX2 BUFX2_710 ( .A(_auto_iopadmap_cc_313_execute_24675_7_), .Y(\sdr_addr[7] ) );
  BUFX2 BUFX2_711 ( .A(_auto_iopadmap_cc_313_execute_24675_8_), .Y(\sdr_addr[8] ) );
  BUFX2 BUFX2_712 ( .A(_auto_iopadmap_cc_313_execute_24675_9_), .Y(\sdr_addr[9] ) );
  BUFX2 BUFX2_713 ( .A(_auto_iopadmap_cc_313_execute_24675_10_), .Y(\sdr_addr[10] ) );
  BUFX2 BUFX2_714 ( .A(_auto_iopadmap_cc_313_execute_24675_11_), .Y(\sdr_addr[11] ) );
  BUFX2 BUFX2_715 ( .A(_auto_iopadmap_cc_313_execute_24675_12_), .Y(\sdr_addr[12] ) );
  BUFX2 BUFX2_716 ( .A(_auto_iopadmap_cc_313_execute_24689_0_), .Y(\sdr_ba[0] ) );
  BUFX2 BUFX2_717 ( .A(_auto_iopadmap_cc_313_execute_24689_1_), .Y(\sdr_ba[1] ) );
  BUFX2 BUFX2_718 ( .A(_auto_iopadmap_cc_313_execute_24692), .Y(sdr_cas_n) );
  BUFX2 BUFX2_719 ( .A(_auto_iopadmap_cc_313_execute_24694), .Y(sdr_cke) );
  BUFX2 BUFX2_72 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf0) );
  BUFX2 BUFX2_720 ( .A(_auto_iopadmap_cc_313_execute_24696), .Y(sdr_cs_n) );
  BUFX2 BUFX2_721 ( .A(_auto_iopadmap_cc_313_execute_24698_0_), .Y(\sdr_dqm[0] ) );
  BUFX2 BUFX2_722 ( .A(_auto_iopadmap_cc_313_execute_24698_1_), .Y(\sdr_dqm[1] ) );
  BUFX2 BUFX2_723 ( .A(_auto_iopadmap_cc_313_execute_24701), .Y(sdr_init_done) );
  BUFX2 BUFX2_724 ( .A(_auto_iopadmap_cc_313_execute_24703), .Y(sdr_ras_n) );
  BUFX2 BUFX2_725 ( .A(_auto_iopadmap_cc_313_execute_24705), .Y(sdr_we_n) );
  BUFX2 BUFX2_726 ( .A(_auto_iopadmap_cc_313_execute_24707), .Y(wb_ack_o) );
  BUFX2 BUFX2_727 ( .A(_auto_iopadmap_cc_313_execute_24709_0_), .Y(\wb_dat_o[0] ) );
  BUFX2 BUFX2_728 ( .A(_auto_iopadmap_cc_313_execute_24709_1_), .Y(\wb_dat_o[1] ) );
  BUFX2 BUFX2_729 ( .A(_auto_iopadmap_cc_313_execute_24709_2_), .Y(\wb_dat_o[2] ) );
  BUFX2 BUFX2_73 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf5) );
  BUFX2 BUFX2_730 ( .A(_auto_iopadmap_cc_313_execute_24709_3_), .Y(\wb_dat_o[3] ) );
  BUFX2 BUFX2_731 ( .A(_auto_iopadmap_cc_313_execute_24709_4_), .Y(\wb_dat_o[4] ) );
  BUFX2 BUFX2_732 ( .A(_auto_iopadmap_cc_313_execute_24709_5_), .Y(\wb_dat_o[5] ) );
  BUFX2 BUFX2_733 ( .A(_auto_iopadmap_cc_313_execute_24709_6_), .Y(\wb_dat_o[6] ) );
  BUFX2 BUFX2_734 ( .A(_auto_iopadmap_cc_313_execute_24709_7_), .Y(\wb_dat_o[7] ) );
  BUFX2 BUFX2_735 ( .A(_auto_iopadmap_cc_313_execute_24709_8_), .Y(\wb_dat_o[8] ) );
  BUFX2 BUFX2_736 ( .A(_auto_iopadmap_cc_313_execute_24709_9_), .Y(\wb_dat_o[9] ) );
  BUFX2 BUFX2_737 ( .A(_auto_iopadmap_cc_313_execute_24709_10_), .Y(\wb_dat_o[10] ) );
  BUFX2 BUFX2_738 ( .A(_auto_iopadmap_cc_313_execute_24709_11_), .Y(\wb_dat_o[11] ) );
  BUFX2 BUFX2_739 ( .A(_auto_iopadmap_cc_313_execute_24709_12_), .Y(\wb_dat_o[12] ) );
  BUFX2 BUFX2_74 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf4) );
  BUFX2 BUFX2_740 ( .A(_auto_iopadmap_cc_313_execute_24709_13_), .Y(\wb_dat_o[13] ) );
  BUFX2 BUFX2_741 ( .A(_auto_iopadmap_cc_313_execute_24709_14_), .Y(\wb_dat_o[14] ) );
  BUFX2 BUFX2_742 ( .A(_auto_iopadmap_cc_313_execute_24709_15_), .Y(\wb_dat_o[15] ) );
  BUFX2 BUFX2_743 ( .A(_auto_iopadmap_cc_313_execute_24709_16_), .Y(\wb_dat_o[16] ) );
  BUFX2 BUFX2_744 ( .A(_auto_iopadmap_cc_313_execute_24709_17_), .Y(\wb_dat_o[17] ) );
  BUFX2 BUFX2_745 ( .A(_auto_iopadmap_cc_313_execute_24709_18_), .Y(\wb_dat_o[18] ) );
  BUFX2 BUFX2_746 ( .A(_auto_iopadmap_cc_313_execute_24709_19_), .Y(\wb_dat_o[19] ) );
  BUFX2 BUFX2_747 ( .A(_auto_iopadmap_cc_313_execute_24709_20_), .Y(\wb_dat_o[20] ) );
  BUFX2 BUFX2_748 ( .A(_auto_iopadmap_cc_313_execute_24709_21_), .Y(\wb_dat_o[21] ) );
  BUFX2 BUFX2_749 ( .A(_auto_iopadmap_cc_313_execute_24709_22_), .Y(\wb_dat_o[22] ) );
  BUFX2 BUFX2_75 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf3) );
  BUFX2 BUFX2_750 ( .A(_auto_iopadmap_cc_313_execute_24709_23_), .Y(\wb_dat_o[23] ) );
  BUFX2 BUFX2_751 ( .A(_auto_iopadmap_cc_313_execute_24709_24_), .Y(\wb_dat_o[24] ) );
  BUFX2 BUFX2_752 ( .A(_auto_iopadmap_cc_313_execute_24709_25_), .Y(\wb_dat_o[25] ) );
  BUFX2 BUFX2_753 ( .A(_auto_iopadmap_cc_313_execute_24709_26_), .Y(\wb_dat_o[26] ) );
  BUFX2 BUFX2_754 ( .A(_auto_iopadmap_cc_313_execute_24709_27_), .Y(\wb_dat_o[27] ) );
  BUFX2 BUFX2_755 ( .A(_auto_iopadmap_cc_313_execute_24709_28_), .Y(\wb_dat_o[28] ) );
  BUFX2 BUFX2_756 ( .A(_auto_iopadmap_cc_313_execute_24709_29_), .Y(\wb_dat_o[29] ) );
  BUFX2 BUFX2_757 ( .A(_auto_iopadmap_cc_313_execute_24709_30_), .Y(\wb_dat_o[30] ) );
  BUFX2 BUFX2_758 ( .A(_auto_iopadmap_cc_313_execute_24709_31_), .Y(\wb_dat_o[31] ) );
  BUFX2 BUFX2_76 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf2) );
  BUFX2 BUFX2_77 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf1) );
  BUFX2 BUFX2_78 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf0) );
  BUFX2 BUFX2_79 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf7) );
  BUFX2 BUFX2_8 ( .A(wb_clk_i), .Y(wb_clk_i_hier0_bF_buf6) );
  BUFX2 BUFX2_80 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf6) );
  BUFX2 BUFX2_81 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf5) );
  BUFX2 BUFX2_82 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf4) );
  BUFX2 BUFX2_83 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf3) );
  BUFX2 BUFX2_84 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf2) );
  BUFX2 BUFX2_85 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf1) );
  BUFX2 BUFX2_86 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf0) );
  BUFX2 BUFX2_87 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf7) );
  BUFX2 BUFX2_88 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf6) );
  BUFX2 BUFX2_89 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf5) );
  BUFX2 BUFX2_9 ( .A(wb_clk_i), .Y(wb_clk_i_hier0_bF_buf5) );
  BUFX2 BUFX2_90 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf4) );
  BUFX2 BUFX2_91 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf3) );
  BUFX2 BUFX2_92 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf2) );
  BUFX2 BUFX2_93 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf1) );
  BUFX2 BUFX2_94 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1158_bF_buf0) );
  BUFX2 BUFX2_95 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf5) );
  BUFX2 BUFX2_96 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf4) );
  BUFX2 BUFX2_97 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf3) );
  BUFX2 BUFX2_98 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf2) );
  BUFX2 BUFX2_99 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf1) );
  DFFPOSX1 DFFPOSX1_1 ( .CLK(sdram_clk_bF_buf80), .D(u_sdrc_core_pad_sdr_din1_0_), .Q(u_sdrc_core_pad_sdr_din2_0_) );
  DFFPOSX1 DFFPOSX1_10 ( .CLK(sdram_clk_bF_buf71), .D(u_sdrc_core_pad_sdr_din1_9_), .Q(u_sdrc_core_pad_sdr_din2_9_) );
  DFFPOSX1 DFFPOSX1_100 ( .CLK(sdram_clk_bF_buf62), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_tras_cntr_0__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_tras_cntr_0_) );
  DFFPOSX1 DFFPOSX1_1000 ( .CLK(wb_clk_i_bF_buf41), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n175), .Q(u_wb2sdrc_u_wrdatafifo_mem_0__7_) );
  DFFPOSX1 DFFPOSX1_1001 ( .CLK(wb_clk_i_bF_buf40), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n178), .Q(u_wb2sdrc_u_wrdatafifo_mem_0__8_) );
  DFFPOSX1 DFFPOSX1_1002 ( .CLK(wb_clk_i_bF_buf39), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n181), .Q(u_wb2sdrc_u_wrdatafifo_mem_0__9_) );
  DFFPOSX1 DFFPOSX1_1003 ( .CLK(wb_clk_i_bF_buf38), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n184), .Q(u_wb2sdrc_u_wrdatafifo_mem_0__10_) );
  DFFPOSX1 DFFPOSX1_1004 ( .CLK(wb_clk_i_bF_buf37), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n187), .Q(u_wb2sdrc_u_wrdatafifo_mem_0__11_) );
  DFFPOSX1 DFFPOSX1_1005 ( .CLK(wb_clk_i_bF_buf36), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n190), .Q(u_wb2sdrc_u_wrdatafifo_mem_0__12_) );
  DFFPOSX1 DFFPOSX1_1006 ( .CLK(wb_clk_i_bF_buf35), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n193), .Q(u_wb2sdrc_u_wrdatafifo_mem_0__13_) );
  DFFPOSX1 DFFPOSX1_1007 ( .CLK(wb_clk_i_bF_buf34), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n196), .Q(u_wb2sdrc_u_wrdatafifo_mem_0__14_) );
  DFFPOSX1 DFFPOSX1_1008 ( .CLK(wb_clk_i_bF_buf33), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n199), .Q(u_wb2sdrc_u_wrdatafifo_mem_0__15_) );
  DFFPOSX1 DFFPOSX1_1009 ( .CLK(wb_clk_i_bF_buf32), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n202), .Q(u_wb2sdrc_u_wrdatafifo_mem_0__16_) );
  DFFPOSX1 DFFPOSX1_101 ( .CLK(sdram_clk_bF_buf61), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_tras_cntr_1__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_tras_cntr_1_) );
  DFFPOSX1 DFFPOSX1_1010 ( .CLK(wb_clk_i_bF_buf31), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n205), .Q(u_wb2sdrc_u_wrdatafifo_mem_0__17_) );
  DFFPOSX1 DFFPOSX1_1011 ( .CLK(wb_clk_i_bF_buf30), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n208), .Q(u_wb2sdrc_u_wrdatafifo_mem_0__18_) );
  DFFPOSX1 DFFPOSX1_1012 ( .CLK(wb_clk_i_bF_buf29), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n211), .Q(u_wb2sdrc_u_wrdatafifo_mem_0__19_) );
  DFFPOSX1 DFFPOSX1_1013 ( .CLK(wb_clk_i_bF_buf28), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n214), .Q(u_wb2sdrc_u_wrdatafifo_mem_0__20_) );
  DFFPOSX1 DFFPOSX1_1014 ( .CLK(wb_clk_i_bF_buf27), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n217), .Q(u_wb2sdrc_u_wrdatafifo_mem_0__21_) );
  DFFPOSX1 DFFPOSX1_1015 ( .CLK(wb_clk_i_bF_buf26), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n220), .Q(u_wb2sdrc_u_wrdatafifo_mem_0__22_) );
  DFFPOSX1 DFFPOSX1_1016 ( .CLK(wb_clk_i_bF_buf25), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n223), .Q(u_wb2sdrc_u_wrdatafifo_mem_0__23_) );
  DFFPOSX1 DFFPOSX1_1017 ( .CLK(wb_clk_i_bF_buf24), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n226), .Q(u_wb2sdrc_u_wrdatafifo_mem_0__24_) );
  DFFPOSX1 DFFPOSX1_1018 ( .CLK(wb_clk_i_bF_buf23), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n229), .Q(u_wb2sdrc_u_wrdatafifo_mem_0__25_) );
  DFFPOSX1 DFFPOSX1_1019 ( .CLK(wb_clk_i_bF_buf22), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n232), .Q(u_wb2sdrc_u_wrdatafifo_mem_0__26_) );
  DFFPOSX1 DFFPOSX1_102 ( .CLK(sdram_clk_bF_buf60), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_tras_cntr_2__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_tras_cntr_2_) );
  DFFPOSX1 DFFPOSX1_1020 ( .CLK(wb_clk_i_bF_buf21), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n235), .Q(u_wb2sdrc_u_wrdatafifo_mem_0__27_) );
  DFFPOSX1 DFFPOSX1_1021 ( .CLK(wb_clk_i_bF_buf20), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n238), .Q(u_wb2sdrc_u_wrdatafifo_mem_0__28_) );
  DFFPOSX1 DFFPOSX1_1022 ( .CLK(wb_clk_i_bF_buf19), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n241), .Q(u_wb2sdrc_u_wrdatafifo_mem_0__29_) );
  DFFPOSX1 DFFPOSX1_1023 ( .CLK(wb_clk_i_bF_buf18), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n244), .Q(u_wb2sdrc_u_wrdatafifo_mem_0__30_) );
  DFFPOSX1 DFFPOSX1_1024 ( .CLK(wb_clk_i_bF_buf17), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n247), .Q(u_wb2sdrc_u_wrdatafifo_mem_0__31_) );
  DFFPOSX1 DFFPOSX1_1025 ( .CLK(wb_clk_i_bF_buf16), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n250), .Q(u_wb2sdrc_u_wrdatafifo_mem_0__32_) );
  DFFPOSX1 DFFPOSX1_1026 ( .CLK(wb_clk_i_bF_buf15), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n253), .Q(u_wb2sdrc_u_wrdatafifo_mem_0__33_) );
  DFFPOSX1 DFFPOSX1_1027 ( .CLK(wb_clk_i_bF_buf14), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n256), .Q(u_wb2sdrc_u_wrdatafifo_mem_0__34_) );
  DFFPOSX1 DFFPOSX1_1028 ( .CLK(wb_clk_i_bF_buf13), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n259), .Q(u_wb2sdrc_u_wrdatafifo_mem_0__35_) );
  DFFPOSX1 DFFPOSX1_1029 ( .CLK(wb_clk_i_bF_buf12), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1070), .Q(u_wb2sdrc_u_wrdatafifo_mem_7__0_) );
  DFFPOSX1 DFFPOSX1_103 ( .CLK(sdram_clk_bF_buf59), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_tras_cntr_3__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_tras_cntr_3_) );
  DFFPOSX1 DFFPOSX1_1030 ( .CLK(wb_clk_i_bF_buf11), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1071), .Q(u_wb2sdrc_u_wrdatafifo_mem_7__1_) );
  DFFPOSX1 DFFPOSX1_1031 ( .CLK(wb_clk_i_bF_buf10), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1072), .Q(u_wb2sdrc_u_wrdatafifo_mem_7__2_) );
  DFFPOSX1 DFFPOSX1_1032 ( .CLK(wb_clk_i_bF_buf9), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1073), .Q(u_wb2sdrc_u_wrdatafifo_mem_7__3_) );
  DFFPOSX1 DFFPOSX1_1033 ( .CLK(wb_clk_i_bF_buf8), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1074), .Q(u_wb2sdrc_u_wrdatafifo_mem_7__4_) );
  DFFPOSX1 DFFPOSX1_1034 ( .CLK(wb_clk_i_bF_buf7), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1075), .Q(u_wb2sdrc_u_wrdatafifo_mem_7__5_) );
  DFFPOSX1 DFFPOSX1_1035 ( .CLK(wb_clk_i_bF_buf6), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1076), .Q(u_wb2sdrc_u_wrdatafifo_mem_7__6_) );
  DFFPOSX1 DFFPOSX1_1036 ( .CLK(wb_clk_i_bF_buf5), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1077), .Q(u_wb2sdrc_u_wrdatafifo_mem_7__7_) );
  DFFPOSX1 DFFPOSX1_1037 ( .CLK(wb_clk_i_bF_buf4), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1078), .Q(u_wb2sdrc_u_wrdatafifo_mem_7__8_) );
  DFFPOSX1 DFFPOSX1_1038 ( .CLK(wb_clk_i_bF_buf3), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1079), .Q(u_wb2sdrc_u_wrdatafifo_mem_7__9_) );
  DFFPOSX1 DFFPOSX1_1039 ( .CLK(wb_clk_i_bF_buf2), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1080), .Q(u_wb2sdrc_u_wrdatafifo_mem_7__10_) );
  DFFPOSX1 DFFPOSX1_104 ( .CLK(sdram_clk_bF_buf58), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_timer0_0__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_timer0_0_) );
  DFFPOSX1 DFFPOSX1_1040 ( .CLK(wb_clk_i_bF_buf1), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1081), .Q(u_wb2sdrc_u_wrdatafifo_mem_7__11_) );
  DFFPOSX1 DFFPOSX1_1041 ( .CLK(wb_clk_i_bF_buf0), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1082), .Q(u_wb2sdrc_u_wrdatafifo_mem_7__12_) );
  DFFPOSX1 DFFPOSX1_1042 ( .CLK(wb_clk_i_bF_buf59), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1083), .Q(u_wb2sdrc_u_wrdatafifo_mem_7__13_) );
  DFFPOSX1 DFFPOSX1_1043 ( .CLK(wb_clk_i_bF_buf58), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1084), .Q(u_wb2sdrc_u_wrdatafifo_mem_7__14_) );
  DFFPOSX1 DFFPOSX1_1044 ( .CLK(wb_clk_i_bF_buf57), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1085), .Q(u_wb2sdrc_u_wrdatafifo_mem_7__15_) );
  DFFPOSX1 DFFPOSX1_1045 ( .CLK(wb_clk_i_bF_buf56), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1086), .Q(u_wb2sdrc_u_wrdatafifo_mem_7__16_) );
  DFFPOSX1 DFFPOSX1_1046 ( .CLK(wb_clk_i_bF_buf55), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1087), .Q(u_wb2sdrc_u_wrdatafifo_mem_7__17_) );
  DFFPOSX1 DFFPOSX1_1047 ( .CLK(wb_clk_i_bF_buf54), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1088), .Q(u_wb2sdrc_u_wrdatafifo_mem_7__18_) );
  DFFPOSX1 DFFPOSX1_1048 ( .CLK(wb_clk_i_bF_buf53), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1089), .Q(u_wb2sdrc_u_wrdatafifo_mem_7__19_) );
  DFFPOSX1 DFFPOSX1_1049 ( .CLK(wb_clk_i_bF_buf52), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1090), .Q(u_wb2sdrc_u_wrdatafifo_mem_7__20_) );
  DFFPOSX1 DFFPOSX1_105 ( .CLK(sdram_clk_bF_buf57), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_timer0_1__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_timer0_1_) );
  DFFPOSX1 DFFPOSX1_1050 ( .CLK(wb_clk_i_bF_buf51), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1091), .Q(u_wb2sdrc_u_wrdatafifo_mem_7__21_) );
  DFFPOSX1 DFFPOSX1_1051 ( .CLK(wb_clk_i_bF_buf50), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1092), .Q(u_wb2sdrc_u_wrdatafifo_mem_7__22_) );
  DFFPOSX1 DFFPOSX1_1052 ( .CLK(wb_clk_i_bF_buf49), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1093), .Q(u_wb2sdrc_u_wrdatafifo_mem_7__23_) );
  DFFPOSX1 DFFPOSX1_1053 ( .CLK(wb_clk_i_bF_buf48), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1094), .Q(u_wb2sdrc_u_wrdatafifo_mem_7__24_) );
  DFFPOSX1 DFFPOSX1_1054 ( .CLK(wb_clk_i_bF_buf47), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1095), .Q(u_wb2sdrc_u_wrdatafifo_mem_7__25_) );
  DFFPOSX1 DFFPOSX1_1055 ( .CLK(wb_clk_i_bF_buf46), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1096), .Q(u_wb2sdrc_u_wrdatafifo_mem_7__26_) );
  DFFPOSX1 DFFPOSX1_1056 ( .CLK(wb_clk_i_bF_buf45), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1097), .Q(u_wb2sdrc_u_wrdatafifo_mem_7__27_) );
  DFFPOSX1 DFFPOSX1_1057 ( .CLK(wb_clk_i_bF_buf44), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1098), .Q(u_wb2sdrc_u_wrdatafifo_mem_7__28_) );
  DFFPOSX1 DFFPOSX1_1058 ( .CLK(wb_clk_i_bF_buf43), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1099), .Q(u_wb2sdrc_u_wrdatafifo_mem_7__29_) );
  DFFPOSX1 DFFPOSX1_1059 ( .CLK(wb_clk_i_bF_buf42), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1100), .Q(u_wb2sdrc_u_wrdatafifo_mem_7__30_) );
  DFFPOSX1 DFFPOSX1_106 ( .CLK(sdram_clk_bF_buf56), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_timer0_2__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_timer0_2_) );
  DFFPOSX1 DFFPOSX1_1060 ( .CLK(wb_clk_i_bF_buf41), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1101), .Q(u_wb2sdrc_u_wrdatafifo_mem_7__31_) );
  DFFPOSX1 DFFPOSX1_1061 ( .CLK(wb_clk_i_bF_buf40), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1102), .Q(u_wb2sdrc_u_wrdatafifo_mem_7__32_) );
  DFFPOSX1 DFFPOSX1_1062 ( .CLK(wb_clk_i_bF_buf39), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1103), .Q(u_wb2sdrc_u_wrdatafifo_mem_7__33_) );
  DFFPOSX1 DFFPOSX1_1063 ( .CLK(wb_clk_i_bF_buf38), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1104), .Q(u_wb2sdrc_u_wrdatafifo_mem_7__34_) );
  DFFPOSX1 DFFPOSX1_1064 ( .CLK(wb_clk_i_bF_buf37), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1105), .Q(u_wb2sdrc_u_wrdatafifo_mem_7__35_) );
  DFFPOSX1 DFFPOSX1_1065 ( .CLK(wb_clk_i_bF_buf36), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n767), .Q(u_wb2sdrc_u_wrdatafifo_mem_6__0_) );
  DFFPOSX1 DFFPOSX1_1066 ( .CLK(wb_clk_i_bF_buf35), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n768), .Q(u_wb2sdrc_u_wrdatafifo_mem_6__1_) );
  DFFPOSX1 DFFPOSX1_1067 ( .CLK(wb_clk_i_bF_buf34), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n769), .Q(u_wb2sdrc_u_wrdatafifo_mem_6__2_) );
  DFFPOSX1 DFFPOSX1_1068 ( .CLK(wb_clk_i_bF_buf33), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n770), .Q(u_wb2sdrc_u_wrdatafifo_mem_6__3_) );
  DFFPOSX1 DFFPOSX1_1069 ( .CLK(wb_clk_i_bF_buf32), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n771), .Q(u_wb2sdrc_u_wrdatafifo_mem_6__4_) );
  DFFPOSX1 DFFPOSX1_107 ( .CLK(sdram_clk_bF_buf55), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_timer0_3__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_timer0_3_) );
  DFFPOSX1 DFFPOSX1_1070 ( .CLK(wb_clk_i_bF_buf31), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n772), .Q(u_wb2sdrc_u_wrdatafifo_mem_6__5_) );
  DFFPOSX1 DFFPOSX1_1071 ( .CLK(wb_clk_i_bF_buf30), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n773), .Q(u_wb2sdrc_u_wrdatafifo_mem_6__6_) );
  DFFPOSX1 DFFPOSX1_1072 ( .CLK(wb_clk_i_bF_buf29), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n774), .Q(u_wb2sdrc_u_wrdatafifo_mem_6__7_) );
  DFFPOSX1 DFFPOSX1_1073 ( .CLK(wb_clk_i_bF_buf28), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n775), .Q(u_wb2sdrc_u_wrdatafifo_mem_6__8_) );
  DFFPOSX1 DFFPOSX1_1074 ( .CLK(wb_clk_i_bF_buf27), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n776), .Q(u_wb2sdrc_u_wrdatafifo_mem_6__9_) );
  DFFPOSX1 DFFPOSX1_1075 ( .CLK(wb_clk_i_bF_buf26), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n777), .Q(u_wb2sdrc_u_wrdatafifo_mem_6__10_) );
  DFFPOSX1 DFFPOSX1_1076 ( .CLK(wb_clk_i_bF_buf25), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n778), .Q(u_wb2sdrc_u_wrdatafifo_mem_6__11_) );
  DFFPOSX1 DFFPOSX1_1077 ( .CLK(wb_clk_i_bF_buf24), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n779), .Q(u_wb2sdrc_u_wrdatafifo_mem_6__12_) );
  DFFPOSX1 DFFPOSX1_1078 ( .CLK(wb_clk_i_bF_buf23), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n780), .Q(u_wb2sdrc_u_wrdatafifo_mem_6__13_) );
  DFFPOSX1 DFFPOSX1_1079 ( .CLK(wb_clk_i_bF_buf22), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n781), .Q(u_wb2sdrc_u_wrdatafifo_mem_6__14_) );
  DFFPOSX1 DFFPOSX1_108 ( .CLK(sdram_clk_bF_buf54), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_wrok_r_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_wrok_r) );
  DFFPOSX1 DFFPOSX1_1080 ( .CLK(wb_clk_i_bF_buf21), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n782), .Q(u_wb2sdrc_u_wrdatafifo_mem_6__15_) );
  DFFPOSX1 DFFPOSX1_1081 ( .CLK(wb_clk_i_bF_buf20), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n783), .Q(u_wb2sdrc_u_wrdatafifo_mem_6__16_) );
  DFFPOSX1 DFFPOSX1_1082 ( .CLK(wb_clk_i_bF_buf19), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n784), .Q(u_wb2sdrc_u_wrdatafifo_mem_6__17_) );
  DFFPOSX1 DFFPOSX1_1083 ( .CLK(wb_clk_i_bF_buf18), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n785), .Q(u_wb2sdrc_u_wrdatafifo_mem_6__18_) );
  DFFPOSX1 DFFPOSX1_1084 ( .CLK(wb_clk_i_bF_buf17), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n786), .Q(u_wb2sdrc_u_wrdatafifo_mem_6__19_) );
  DFFPOSX1 DFFPOSX1_1085 ( .CLK(wb_clk_i_bF_buf16), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n787), .Q(u_wb2sdrc_u_wrdatafifo_mem_6__20_) );
  DFFPOSX1 DFFPOSX1_1086 ( .CLK(wb_clk_i_bF_buf15), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n788), .Q(u_wb2sdrc_u_wrdatafifo_mem_6__21_) );
  DFFPOSX1 DFFPOSX1_1087 ( .CLK(wb_clk_i_bF_buf14), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n789), .Q(u_wb2sdrc_u_wrdatafifo_mem_6__22_) );
  DFFPOSX1 DFFPOSX1_1088 ( .CLK(wb_clk_i_bF_buf13), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n790), .Q(u_wb2sdrc_u_wrdatafifo_mem_6__23_) );
  DFFPOSX1 DFFPOSX1_1089 ( .CLK(wb_clk_i_bF_buf12), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n791), .Q(u_wb2sdrc_u_wrdatafifo_mem_6__24_) );
  DFFPOSX1 DFFPOSX1_109 ( .CLK(sdram_clk_bF_buf53), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_xfr_ok_r_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_xfr_ok_r) );
  DFFPOSX1 DFFPOSX1_1090 ( .CLK(wb_clk_i_bF_buf11), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n792), .Q(u_wb2sdrc_u_wrdatafifo_mem_6__25_) );
  DFFPOSX1 DFFPOSX1_1091 ( .CLK(wb_clk_i_bF_buf10), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n793), .Q(u_wb2sdrc_u_wrdatafifo_mem_6__26_) );
  DFFPOSX1 DFFPOSX1_1092 ( .CLK(wb_clk_i_bF_buf9), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n794), .Q(u_wb2sdrc_u_wrdatafifo_mem_6__27_) );
  DFFPOSX1 DFFPOSX1_1093 ( .CLK(wb_clk_i_bF_buf8), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n795), .Q(u_wb2sdrc_u_wrdatafifo_mem_6__28_) );
  DFFPOSX1 DFFPOSX1_1094 ( .CLK(wb_clk_i_bF_buf7), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n796), .Q(u_wb2sdrc_u_wrdatafifo_mem_6__29_) );
  DFFPOSX1 DFFPOSX1_1095 ( .CLK(wb_clk_i_bF_buf6), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n797), .Q(u_wb2sdrc_u_wrdatafifo_mem_6__30_) );
  DFFPOSX1 DFFPOSX1_1096 ( .CLK(wb_clk_i_bF_buf5), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n798), .Q(u_wb2sdrc_u_wrdatafifo_mem_6__31_) );
  DFFPOSX1 DFFPOSX1_1097 ( .CLK(wb_clk_i_bF_buf4), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n799), .Q(u_wb2sdrc_u_wrdatafifo_mem_6__32_) );
  DFFPOSX1 DFFPOSX1_1098 ( .CLK(wb_clk_i_bF_buf3), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n800), .Q(u_wb2sdrc_u_wrdatafifo_mem_6__33_) );
  DFFPOSX1 DFFPOSX1_1099 ( .CLK(wb_clk_i_bF_buf2), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n801), .Q(u_wb2sdrc_u_wrdatafifo_mem_6__34_) );
  DFFPOSX1 DFFPOSX1_11 ( .CLK(sdram_clk_bF_buf70), .D(u_sdrc_core_pad_sdr_din1_10_), .Q(u_sdrc_core_pad_sdr_din2_10_) );
  DFFPOSX1 DFFPOSX1_110 ( .CLK(sdram_clk_bF_buf52), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_rdok_r_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_rdok_r) );
  DFFPOSX1 DFFPOSX1_1100 ( .CLK(wb_clk_i_bF_buf1), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n802), .Q(u_wb2sdrc_u_wrdatafifo_mem_6__35_) );
  DFFPOSX1 DFFPOSX1_1101 ( .CLK(wb_clk_i_bF_buf0), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n513), .Q(u_wb2sdrc_u_wrdatafifo_mem_4__0_) );
  DFFPOSX1 DFFPOSX1_1102 ( .CLK(wb_clk_i_bF_buf59), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n515), .Q(u_wb2sdrc_u_wrdatafifo_mem_4__1_) );
  DFFPOSX1 DFFPOSX1_1103 ( .CLK(wb_clk_i_bF_buf58), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n517), .Q(u_wb2sdrc_u_wrdatafifo_mem_4__2_) );
  DFFPOSX1 DFFPOSX1_1104 ( .CLK(wb_clk_i_bF_buf57), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n519), .Q(u_wb2sdrc_u_wrdatafifo_mem_4__3_) );
  DFFPOSX1 DFFPOSX1_1105 ( .CLK(wb_clk_i_bF_buf56), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n521), .Q(u_wb2sdrc_u_wrdatafifo_mem_4__4_) );
  DFFPOSX1 DFFPOSX1_1106 ( .CLK(wb_clk_i_bF_buf55), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n523), .Q(u_wb2sdrc_u_wrdatafifo_mem_4__5_) );
  DFFPOSX1 DFFPOSX1_1107 ( .CLK(wb_clk_i_bF_buf54), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n525), .Q(u_wb2sdrc_u_wrdatafifo_mem_4__6_) );
  DFFPOSX1 DFFPOSX1_1108 ( .CLK(wb_clk_i_bF_buf53), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n527), .Q(u_wb2sdrc_u_wrdatafifo_mem_4__7_) );
  DFFPOSX1 DFFPOSX1_1109 ( .CLK(wb_clk_i_bF_buf52), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n529), .Q(u_wb2sdrc_u_wrdatafifo_mem_4__8_) );
  DFFPOSX1 DFFPOSX1_111 ( .CLK(sdram_clk_bF_buf51), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_cmd_r_0__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_cmd_0_) );
  DFFPOSX1 DFFPOSX1_1110 ( .CLK(wb_clk_i_bF_buf51), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n531), .Q(u_wb2sdrc_u_wrdatafifo_mem_4__9_) );
  DFFPOSX1 DFFPOSX1_1111 ( .CLK(wb_clk_i_bF_buf50), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n533), .Q(u_wb2sdrc_u_wrdatafifo_mem_4__10_) );
  DFFPOSX1 DFFPOSX1_1112 ( .CLK(wb_clk_i_bF_buf49), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n535), .Q(u_wb2sdrc_u_wrdatafifo_mem_4__11_) );
  DFFPOSX1 DFFPOSX1_1113 ( .CLK(wb_clk_i_bF_buf48), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n537), .Q(u_wb2sdrc_u_wrdatafifo_mem_4__12_) );
  DFFPOSX1 DFFPOSX1_1114 ( .CLK(wb_clk_i_bF_buf47), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n539), .Q(u_wb2sdrc_u_wrdatafifo_mem_4__13_) );
  DFFPOSX1 DFFPOSX1_1115 ( .CLK(wb_clk_i_bF_buf46), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n541), .Q(u_wb2sdrc_u_wrdatafifo_mem_4__14_) );
  DFFPOSX1 DFFPOSX1_1116 ( .CLK(wb_clk_i_bF_buf45), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n543), .Q(u_wb2sdrc_u_wrdatafifo_mem_4__15_) );
  DFFPOSX1 DFFPOSX1_1117 ( .CLK(wb_clk_i_bF_buf44), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n545), .Q(u_wb2sdrc_u_wrdatafifo_mem_4__16_) );
  DFFPOSX1 DFFPOSX1_1118 ( .CLK(wb_clk_i_bF_buf43), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n547), .Q(u_wb2sdrc_u_wrdatafifo_mem_4__17_) );
  DFFPOSX1 DFFPOSX1_1119 ( .CLK(wb_clk_i_bF_buf42), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n549), .Q(u_wb2sdrc_u_wrdatafifo_mem_4__18_) );
  DFFPOSX1 DFFPOSX1_112 ( .CLK(sdram_clk_bF_buf50), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_cmd_r_1__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_cmd_1_) );
  DFFPOSX1 DFFPOSX1_1120 ( .CLK(wb_clk_i_bF_buf41), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n551), .Q(u_wb2sdrc_u_wrdatafifo_mem_4__19_) );
  DFFPOSX1 DFFPOSX1_1121 ( .CLK(wb_clk_i_bF_buf40), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n553), .Q(u_wb2sdrc_u_wrdatafifo_mem_4__20_) );
  DFFPOSX1 DFFPOSX1_1122 ( .CLK(wb_clk_i_bF_buf39), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n555), .Q(u_wb2sdrc_u_wrdatafifo_mem_4__21_) );
  DFFPOSX1 DFFPOSX1_1123 ( .CLK(wb_clk_i_bF_buf38), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n557), .Q(u_wb2sdrc_u_wrdatafifo_mem_4__22_) );
  DFFPOSX1 DFFPOSX1_1124 ( .CLK(wb_clk_i_bF_buf37), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n559), .Q(u_wb2sdrc_u_wrdatafifo_mem_4__23_) );
  DFFPOSX1 DFFPOSX1_1125 ( .CLK(wb_clk_i_bF_buf36), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n561), .Q(u_wb2sdrc_u_wrdatafifo_mem_4__24_) );
  DFFPOSX1 DFFPOSX1_1126 ( .CLK(wb_clk_i_bF_buf35), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n563), .Q(u_wb2sdrc_u_wrdatafifo_mem_4__25_) );
  DFFPOSX1 DFFPOSX1_1127 ( .CLK(wb_clk_i_bF_buf34), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n565), .Q(u_wb2sdrc_u_wrdatafifo_mem_4__26_) );
  DFFPOSX1 DFFPOSX1_1128 ( .CLK(wb_clk_i_bF_buf33), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n567), .Q(u_wb2sdrc_u_wrdatafifo_mem_4__27_) );
  DFFPOSX1 DFFPOSX1_1129 ( .CLK(wb_clk_i_bF_buf32), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n569), .Q(u_wb2sdrc_u_wrdatafifo_mem_4__28_) );
  DFFPOSX1 DFFPOSX1_113 ( .CLK(sdram_clk_bF_buf49), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_timer0_tc_r_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_timer0_tc) );
  DFFPOSX1 DFFPOSX1_1130 ( .CLK(wb_clk_i_bF_buf31), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n571), .Q(u_wb2sdrc_u_wrdatafifo_mem_4__29_) );
  DFFPOSX1 DFFPOSX1_1131 ( .CLK(wb_clk_i_bF_buf30), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n573), .Q(u_wb2sdrc_u_wrdatafifo_mem_4__30_) );
  DFFPOSX1 DFFPOSX1_1132 ( .CLK(wb_clk_i_bF_buf29), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n575), .Q(u_wb2sdrc_u_wrdatafifo_mem_4__31_) );
  DFFPOSX1 DFFPOSX1_1133 ( .CLK(wb_clk_i_bF_buf28), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n577), .Q(u_wb2sdrc_u_wrdatafifo_mem_4__32_) );
  DFFPOSX1 DFFPOSX1_1134 ( .CLK(wb_clk_i_bF_buf27), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n579), .Q(u_wb2sdrc_u_wrdatafifo_mem_4__33_) );
  DFFPOSX1 DFFPOSX1_1135 ( .CLK(wb_clk_i_bF_buf26), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n581), .Q(u_wb2sdrc_u_wrdatafifo_mem_4__34_) );
  DFFPOSX1 DFFPOSX1_1136 ( .CLK(wb_clk_i_bF_buf25), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n583), .Q(u_wb2sdrc_u_wrdatafifo_mem_4__35_) );
  DFFPOSX1 DFFPOSX1_114 ( .CLK(sdram_clk_bF_buf48), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_tras_ok_r_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_tras_ok) );
  DFFPOSX1 DFFPOSX1_115 ( .CLK(sdram_clk_bF_buf47), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_pre_ok_r_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_pre_ok_t) );
  DFFPOSX1 DFFPOSX1_116 ( .CLK(sdram_clk_bF_buf46), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_act_ok_r_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_act_ok_t) );
  DFFPOSX1 DFFPOSX1_117 ( .CLK(sdram_clk_bF_buf45), .D(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_17422_n90), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_0_) );
  DFFPOSX1 DFFPOSX1_118 ( .CLK(sdram_clk_bF_buf44), .D(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_17422_n61), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_prech_page_closed) );
  DFFPOSX1 DFFPOSX1_119 ( .CLK(sdram_clk_bF_buf43), .D(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_17422_n66), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_2_) );
  DFFPOSX1 DFFPOSX1_12 ( .CLK(sdram_clk_bF_buf69), .D(u_sdrc_core_pad_sdr_din1_11_), .Q(u_sdrc_core_pad_sdr_din2_11_) );
  DFFPOSX1 DFFPOSX1_120 ( .CLK(sdram_clk_bF_buf42), .D(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_17422_n55), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_3_) );
  DFFPOSX1 DFFPOSX1_121 ( .CLK(sdram_clk_bF_buf41), .D(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_17422_n82), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_4_) );
  DFFPOSX1 DFFPOSX1_122 ( .CLK(sdram_clk_bF_buf40), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_l_last_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_l_last) );
  DFFPOSX1 DFFPOSX1_123 ( .CLK(sdram_clk_bF_buf39), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_l_wrap_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_l_wrap) );
  DFFPOSX1 DFFPOSX1_124 ( .CLK(sdram_clk_bF_buf38), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_0__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_0_) );
  DFFPOSX1 DFFPOSX1_125 ( .CLK(sdram_clk_bF_buf37), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_1__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_1_) );
  DFFPOSX1 DFFPOSX1_126 ( .CLK(sdram_clk_bF_buf36), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_2__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_2_) );
  DFFPOSX1 DFFPOSX1_127 ( .CLK(sdram_clk_bF_buf35), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_3__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_3_) );
  DFFPOSX1 DFFPOSX1_128 ( .CLK(sdram_clk_bF_buf34), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_4__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_4_) );
  DFFPOSX1 DFFPOSX1_129 ( .CLK(sdram_clk_bF_buf33), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_5__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_5_) );
  DFFPOSX1 DFFPOSX1_13 ( .CLK(sdram_clk_bF_buf68), .D(u_sdrc_core_pad_sdr_din1_12_), .Q(u_sdrc_core_pad_sdr_din2_12_) );
  DFFPOSX1 DFFPOSX1_130 ( .CLK(sdram_clk_bF_buf32), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_6__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_6_) );
  DFFPOSX1 DFFPOSX1_131 ( .CLK(sdram_clk_bF_buf31), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_0__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_0_) );
  DFFPOSX1 DFFPOSX1_132 ( .CLK(sdram_clk_bF_buf30), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_1__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_1_) );
  DFFPOSX1 DFFPOSX1_133 ( .CLK(sdram_clk_bF_buf29), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_2__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_2_) );
  DFFPOSX1 DFFPOSX1_134 ( .CLK(sdram_clk_bF_buf28), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_3__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_3_) );
  DFFPOSX1 DFFPOSX1_135 ( .CLK(sdram_clk_bF_buf27), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_4__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_4_) );
  DFFPOSX1 DFFPOSX1_136 ( .CLK(sdram_clk_bF_buf26), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_5__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_5_) );
  DFFPOSX1 DFFPOSX1_137 ( .CLK(sdram_clk_bF_buf25), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_6__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_6_) );
  DFFPOSX1 DFFPOSX1_138 ( .CLK(sdram_clk_bF_buf24), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_7__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_7_) );
  DFFPOSX1 DFFPOSX1_139 ( .CLK(sdram_clk_bF_buf23), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_8__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_8_) );
  DFFPOSX1 DFFPOSX1_14 ( .CLK(sdram_clk_bF_buf67), .D(u_sdrc_core_pad_sdr_din1_13_), .Q(u_sdrc_core_pad_sdr_din2_13_) );
  DFFPOSX1 DFFPOSX1_140 ( .CLK(sdram_clk_bF_buf22), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_9__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_9_) );
  DFFPOSX1 DFFPOSX1_141 ( .CLK(sdram_clk_bF_buf21), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_10__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_10_) );
  DFFPOSX1 DFFPOSX1_142 ( .CLK(sdram_clk_bF_buf20), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_11__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_11_) );
  DFFPOSX1 DFFPOSX1_143 ( .CLK(sdram_clk_bF_buf19), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_12__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_12_) );
  DFFPOSX1 DFFPOSX1_144 ( .CLK(sdram_clk_bF_buf18), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_l_write_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_l_write) );
  DFFPOSX1 DFFPOSX1_145 ( .CLK(sdram_clk_bF_buf17), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_0__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_0_) );
  DFFPOSX1 DFFPOSX1_146 ( .CLK(sdram_clk_bF_buf16), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_1__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_1_) );
  DFFPOSX1 DFFPOSX1_147 ( .CLK(sdram_clk_bF_buf15), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_2__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_2_) );
  DFFPOSX1 DFFPOSX1_148 ( .CLK(sdram_clk_bF_buf14), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_3__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_3_) );
  DFFPOSX1 DFFPOSX1_149 ( .CLK(sdram_clk_bF_buf13), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_4__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_4_) );
  DFFPOSX1 DFFPOSX1_15 ( .CLK(sdram_clk_bF_buf66), .D(u_sdrc_core_pad_sdr_din1_14_), .Q(u_sdrc_core_pad_sdr_din2_14_) );
  DFFPOSX1 DFFPOSX1_150 ( .CLK(sdram_clk_bF_buf12), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_5__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_5_) );
  DFFPOSX1 DFFPOSX1_151 ( .CLK(sdram_clk_bF_buf11), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_6__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_6_) );
  DFFPOSX1 DFFPOSX1_152 ( .CLK(sdram_clk_bF_buf10), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_7__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_7_) );
  DFFPOSX1 DFFPOSX1_153 ( .CLK(sdram_clk_bF_buf9), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_8__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_8_) );
  DFFPOSX1 DFFPOSX1_154 ( .CLK(sdram_clk_bF_buf8), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_9__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_9_) );
  DFFPOSX1 DFFPOSX1_155 ( .CLK(sdram_clk_bF_buf7), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_10__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_10_) );
  DFFPOSX1 DFFPOSX1_156 ( .CLK(sdram_clk_bF_buf6), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_11__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_11_) );
  DFFPOSX1 DFFPOSX1_157 ( .CLK(sdram_clk_bF_buf5), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_12__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_l_raddr_12_) );
  DFFPOSX1 DFFPOSX1_158 ( .CLK(sdram_clk_bF_buf4), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_0__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_0_) );
  DFFPOSX1 DFFPOSX1_159 ( .CLK(sdram_clk_bF_buf3), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_1__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_1_) );
  DFFPOSX1 DFFPOSX1_16 ( .CLK(sdram_clk_bF_buf65), .D(u_sdrc_core_pad_sdr_din1_15_), .Q(u_sdrc_core_pad_sdr_din2_15_) );
  DFFPOSX1 DFFPOSX1_160 ( .CLK(sdram_clk_bF_buf2), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_2__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_2_) );
  DFFPOSX1 DFFPOSX1_161 ( .CLK(sdram_clk_bF_buf1), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_3__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_3_) );
  DFFPOSX1 DFFPOSX1_162 ( .CLK(sdram_clk_bF_buf0), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_4__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_4_) );
  DFFPOSX1 DFFPOSX1_163 ( .CLK(sdram_clk_bF_buf80), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_5__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_5_) );
  DFFPOSX1 DFFPOSX1_164 ( .CLK(sdram_clk_bF_buf79), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_6__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_6_) );
  DFFPOSX1 DFFPOSX1_165 ( .CLK(sdram_clk_bF_buf78), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_7__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_7_) );
  DFFPOSX1 DFFPOSX1_166 ( .CLK(sdram_clk_bF_buf77), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_8__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_8_) );
  DFFPOSX1 DFFPOSX1_167 ( .CLK(sdram_clk_bF_buf76), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_9__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_9_) );
  DFFPOSX1 DFFPOSX1_168 ( .CLK(sdram_clk_bF_buf75), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_10__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_10_) );
  DFFPOSX1 DFFPOSX1_169 ( .CLK(sdram_clk_bF_buf74), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_11__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_11_) );
  DFFPOSX1 DFFPOSX1_17 ( .CLK(sdram_clk_bF_buf64), .D(\sdr_dq[0] ), .Q(u_sdrc_core_pad_sdr_din1_0_) );
  DFFPOSX1 DFFPOSX1_170 ( .CLK(sdram_clk_bF_buf73), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_12__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_l_caddr_12_) );
  DFFPOSX1 DFFPOSX1_171 ( .CLK(sdram_clk_bF_buf72), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_l_sdr_dma_last_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_l_sdr_dma_last) );
  DFFPOSX1 DFFPOSX1_172 ( .CLK(sdram_clk_bF_buf71), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_valid_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_valid) );
  DFFPOSX1 DFFPOSX1_173 ( .CLK(sdram_clk_bF_buf70), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_tras_cntr_0__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_tras_cntr_0_) );
  DFFPOSX1 DFFPOSX1_174 ( .CLK(sdram_clk_bF_buf69), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_tras_cntr_1__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_tras_cntr_1_) );
  DFFPOSX1 DFFPOSX1_175 ( .CLK(sdram_clk_bF_buf68), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_tras_cntr_2__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_tras_cntr_2_) );
  DFFPOSX1 DFFPOSX1_176 ( .CLK(sdram_clk_bF_buf67), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_tras_cntr_3__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_tras_cntr_3_) );
  DFFPOSX1 DFFPOSX1_177 ( .CLK(sdram_clk_bF_buf66), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_timer0_0__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_timer0_0_) );
  DFFPOSX1 DFFPOSX1_178 ( .CLK(sdram_clk_bF_buf65), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_timer0_1__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_timer0_1_) );
  DFFPOSX1 DFFPOSX1_179 ( .CLK(sdram_clk_bF_buf64), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_timer0_2__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_timer0_2_) );
  DFFPOSX1 DFFPOSX1_18 ( .CLK(sdram_clk_bF_buf63), .D(\sdr_dq[1] ), .Q(u_sdrc_core_pad_sdr_din1_1_) );
  DFFPOSX1 DFFPOSX1_180 ( .CLK(sdram_clk_bF_buf63), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_timer0_3__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_timer0_3_) );
  DFFPOSX1 DFFPOSX1_181 ( .CLK(sdram_clk_bF_buf62), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_x2b_wrok_r_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_x2b_wrok_r) );
  DFFPOSX1 DFFPOSX1_182 ( .CLK(sdram_clk_bF_buf61), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_r_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_r) );
  DFFPOSX1 DFFPOSX1_183 ( .CLK(sdram_clk_bF_buf60), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_x2b_rdok_r_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_x2b_rdok_r) );
  DFFPOSX1 DFFPOSX1_184 ( .CLK(sdram_clk_bF_buf59), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_cmd_r_0__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_cmd_0_) );
  DFFPOSX1 DFFPOSX1_185 ( .CLK(sdram_clk_bF_buf58), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_cmd_r_1__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_cmd_1_) );
  DFFPOSX1 DFFPOSX1_186 ( .CLK(sdram_clk_bF_buf57), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_timer0_tc_r_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_timer0_tc) );
  DFFPOSX1 DFFPOSX1_187 ( .CLK(sdram_clk_bF_buf56), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_tras_ok_r_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_tras_ok) );
  DFFPOSX1 DFFPOSX1_188 ( .CLK(sdram_clk_bF_buf55), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_x2b_pre_ok_r_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_x2b_pre_ok_t) );
  DFFPOSX1 DFFPOSX1_189 ( .CLK(sdram_clk_bF_buf54), .D(u_sdrc_core_u_bank_ctl_bank1_fsm_x2b_act_ok_r_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank1_fsm_x2b_act_ok_t) );
  DFFPOSX1 DFFPOSX1_19 ( .CLK(sdram_clk_bF_buf62), .D(\sdr_dq[2] ), .Q(u_sdrc_core_pad_sdr_din1_2_) );
  DFFPOSX1 DFFPOSX1_190 ( .CLK(sdram_clk_bF_buf53), .D(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_17422_n90), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_0_) );
  DFFPOSX1 DFFPOSX1_191 ( .CLK(sdram_clk_bF_buf52), .D(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_17422_n61), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_prech_page_closed) );
  DFFPOSX1 DFFPOSX1_192 ( .CLK(sdram_clk_bF_buf51), .D(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_17422_n66), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_2_) );
  DFFPOSX1 DFFPOSX1_193 ( .CLK(sdram_clk_bF_buf50), .D(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_17422_n55), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_3_) );
  DFFPOSX1 DFFPOSX1_194 ( .CLK(sdram_clk_bF_buf49), .D(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_17422_n82), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_4_) );
  DFFPOSX1 DFFPOSX1_195 ( .CLK(sdram_clk_bF_buf48), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_l_last_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_l_last) );
  DFFPOSX1 DFFPOSX1_196 ( .CLK(sdram_clk_bF_buf47), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_l_wrap_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_l_wrap) );
  DFFPOSX1 DFFPOSX1_197 ( .CLK(sdram_clk_bF_buf46), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_0__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_0_) );
  DFFPOSX1 DFFPOSX1_198 ( .CLK(sdram_clk_bF_buf45), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_1__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_1_) );
  DFFPOSX1 DFFPOSX1_199 ( .CLK(sdram_clk_bF_buf44), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_2__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_2_) );
  DFFPOSX1 DFFPOSX1_2 ( .CLK(sdram_clk_bF_buf79), .D(u_sdrc_core_pad_sdr_din1_1_), .Q(u_sdrc_core_pad_sdr_din2_1_) );
  DFFPOSX1 DFFPOSX1_20 ( .CLK(sdram_clk_bF_buf61), .D(\sdr_dq[3] ), .Q(u_sdrc_core_pad_sdr_din1_3_) );
  DFFPOSX1 DFFPOSX1_200 ( .CLK(sdram_clk_bF_buf43), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_3__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_3_) );
  DFFPOSX1 DFFPOSX1_201 ( .CLK(sdram_clk_bF_buf42), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_4__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_4_) );
  DFFPOSX1 DFFPOSX1_202 ( .CLK(sdram_clk_bF_buf41), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_5__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_5_) );
  DFFPOSX1 DFFPOSX1_203 ( .CLK(sdram_clk_bF_buf40), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_6__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_6_) );
  DFFPOSX1 DFFPOSX1_204 ( .CLK(sdram_clk_bF_buf39), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_0__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_0_) );
  DFFPOSX1 DFFPOSX1_205 ( .CLK(sdram_clk_bF_buf38), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_1__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_1_) );
  DFFPOSX1 DFFPOSX1_206 ( .CLK(sdram_clk_bF_buf37), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_2__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_2_) );
  DFFPOSX1 DFFPOSX1_207 ( .CLK(sdram_clk_bF_buf36), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_3__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_3_) );
  DFFPOSX1 DFFPOSX1_208 ( .CLK(sdram_clk_bF_buf35), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_4__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_4_) );
  DFFPOSX1 DFFPOSX1_209 ( .CLK(sdram_clk_bF_buf34), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_5__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_5_) );
  DFFPOSX1 DFFPOSX1_21 ( .CLK(sdram_clk_bF_buf60), .D(\sdr_dq[4] ), .Q(u_sdrc_core_pad_sdr_din1_4_) );
  DFFPOSX1 DFFPOSX1_210 ( .CLK(sdram_clk_bF_buf33), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_6__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_6_) );
  DFFPOSX1 DFFPOSX1_211 ( .CLK(sdram_clk_bF_buf32), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_7__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_7_) );
  DFFPOSX1 DFFPOSX1_212 ( .CLK(sdram_clk_bF_buf31), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_8__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_8_) );
  DFFPOSX1 DFFPOSX1_213 ( .CLK(sdram_clk_bF_buf30), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_9__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_9_) );
  DFFPOSX1 DFFPOSX1_214 ( .CLK(sdram_clk_bF_buf29), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_10__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_10_) );
  DFFPOSX1 DFFPOSX1_215 ( .CLK(sdram_clk_bF_buf28), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_11__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_11_) );
  DFFPOSX1 DFFPOSX1_216 ( .CLK(sdram_clk_bF_buf27), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_12__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_12_) );
  DFFPOSX1 DFFPOSX1_217 ( .CLK(sdram_clk_bF_buf26), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_l_write_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_l_write) );
  DFFPOSX1 DFFPOSX1_218 ( .CLK(sdram_clk_bF_buf25), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_0__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_0_) );
  DFFPOSX1 DFFPOSX1_219 ( .CLK(sdram_clk_bF_buf24), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_1__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_1_) );
  DFFPOSX1 DFFPOSX1_22 ( .CLK(sdram_clk_bF_buf59), .D(\sdr_dq[5] ), .Q(u_sdrc_core_pad_sdr_din1_5_) );
  DFFPOSX1 DFFPOSX1_220 ( .CLK(sdram_clk_bF_buf23), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_2__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_2_) );
  DFFPOSX1 DFFPOSX1_221 ( .CLK(sdram_clk_bF_buf22), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_3__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_3_) );
  DFFPOSX1 DFFPOSX1_222 ( .CLK(sdram_clk_bF_buf21), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_4__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_4_) );
  DFFPOSX1 DFFPOSX1_223 ( .CLK(sdram_clk_bF_buf20), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_5__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_5_) );
  DFFPOSX1 DFFPOSX1_224 ( .CLK(sdram_clk_bF_buf19), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_6__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_6_) );
  DFFPOSX1 DFFPOSX1_225 ( .CLK(sdram_clk_bF_buf18), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_7__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_7_) );
  DFFPOSX1 DFFPOSX1_226 ( .CLK(sdram_clk_bF_buf17), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_8__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_8_) );
  DFFPOSX1 DFFPOSX1_227 ( .CLK(sdram_clk_bF_buf16), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_9__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_9_) );
  DFFPOSX1 DFFPOSX1_228 ( .CLK(sdram_clk_bF_buf15), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_10__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_10_) );
  DFFPOSX1 DFFPOSX1_229 ( .CLK(sdram_clk_bF_buf14), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_11__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_11_) );
  DFFPOSX1 DFFPOSX1_23 ( .CLK(sdram_clk_bF_buf58), .D(\sdr_dq[6] ), .Q(u_sdrc_core_pad_sdr_din1_6_) );
  DFFPOSX1 DFFPOSX1_230 ( .CLK(sdram_clk_bF_buf13), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_12__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_l_raddr_12_) );
  DFFPOSX1 DFFPOSX1_231 ( .CLK(sdram_clk_bF_buf12), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_0__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_0_) );
  DFFPOSX1 DFFPOSX1_232 ( .CLK(sdram_clk_bF_buf11), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_1__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_1_) );
  DFFPOSX1 DFFPOSX1_233 ( .CLK(sdram_clk_bF_buf10), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_2__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_2_) );
  DFFPOSX1 DFFPOSX1_234 ( .CLK(sdram_clk_bF_buf9), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_3__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_3_) );
  DFFPOSX1 DFFPOSX1_235 ( .CLK(sdram_clk_bF_buf8), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_4__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_4_) );
  DFFPOSX1 DFFPOSX1_236 ( .CLK(sdram_clk_bF_buf7), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_5__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_5_) );
  DFFPOSX1 DFFPOSX1_237 ( .CLK(sdram_clk_bF_buf6), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_6__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_6_) );
  DFFPOSX1 DFFPOSX1_238 ( .CLK(sdram_clk_bF_buf5), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_7__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_7_) );
  DFFPOSX1 DFFPOSX1_239 ( .CLK(sdram_clk_bF_buf4), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_8__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_8_) );
  DFFPOSX1 DFFPOSX1_24 ( .CLK(sdram_clk_bF_buf57), .D(\sdr_dq[7] ), .Q(u_sdrc_core_pad_sdr_din1_7_) );
  DFFPOSX1 DFFPOSX1_240 ( .CLK(sdram_clk_bF_buf3), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_9__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_9_) );
  DFFPOSX1 DFFPOSX1_241 ( .CLK(sdram_clk_bF_buf2), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_10__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_10_) );
  DFFPOSX1 DFFPOSX1_242 ( .CLK(sdram_clk_bF_buf1), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_11__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_11_) );
  DFFPOSX1 DFFPOSX1_243 ( .CLK(sdram_clk_bF_buf0), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_12__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_l_caddr_12_) );
  DFFPOSX1 DFFPOSX1_244 ( .CLK(sdram_clk_bF_buf80), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_l_sdr_dma_last_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_l_sdr_dma_last) );
  DFFPOSX1 DFFPOSX1_245 ( .CLK(sdram_clk_bF_buf79), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_valid_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_valid) );
  DFFPOSX1 DFFPOSX1_246 ( .CLK(sdram_clk_bF_buf78), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_tras_cntr_0__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_tras_cntr_0_) );
  DFFPOSX1 DFFPOSX1_247 ( .CLK(sdram_clk_bF_buf77), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_tras_cntr_1__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_tras_cntr_1_) );
  DFFPOSX1 DFFPOSX1_248 ( .CLK(sdram_clk_bF_buf76), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_tras_cntr_2__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_tras_cntr_2_) );
  DFFPOSX1 DFFPOSX1_249 ( .CLK(sdram_clk_bF_buf75), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_tras_cntr_3__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_tras_cntr_3_) );
  DFFPOSX1 DFFPOSX1_25 ( .CLK(sdram_clk_bF_buf56), .D(\sdr_dq[8] ), .Q(u_sdrc_core_pad_sdr_din1_8_) );
  DFFPOSX1 DFFPOSX1_250 ( .CLK(sdram_clk_bF_buf74), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_timer0_0__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_timer0_0_) );
  DFFPOSX1 DFFPOSX1_251 ( .CLK(sdram_clk_bF_buf73), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_timer0_1__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_timer0_1_) );
  DFFPOSX1 DFFPOSX1_252 ( .CLK(sdram_clk_bF_buf72), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_timer0_2__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_timer0_2_) );
  DFFPOSX1 DFFPOSX1_253 ( .CLK(sdram_clk_bF_buf71), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_timer0_3__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_timer0_3_) );
  DFFPOSX1 DFFPOSX1_254 ( .CLK(sdram_clk_bF_buf70), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_x2b_wrok_r_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_x2b_wrok_r) );
  DFFPOSX1 DFFPOSX1_255 ( .CLK(sdram_clk_bF_buf69), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_r_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_r) );
  DFFPOSX1 DFFPOSX1_256 ( .CLK(sdram_clk_bF_buf68), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_x2b_rdok_r_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_x2b_rdok_r) );
  DFFPOSX1 DFFPOSX1_257 ( .CLK(sdram_clk_bF_buf67), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_cmd_r_0__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_cmd_0_) );
  DFFPOSX1 DFFPOSX1_258 ( .CLK(sdram_clk_bF_buf66), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_cmd_r_1__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_cmd_1_) );
  DFFPOSX1 DFFPOSX1_259 ( .CLK(sdram_clk_bF_buf65), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_timer0_tc_r_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_timer0_tc) );
  DFFPOSX1 DFFPOSX1_26 ( .CLK(sdram_clk_bF_buf55), .D(\sdr_dq[9] ), .Q(u_sdrc_core_pad_sdr_din1_9_) );
  DFFPOSX1 DFFPOSX1_260 ( .CLK(sdram_clk_bF_buf64), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_tras_ok_r_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_tras_ok) );
  DFFPOSX1 DFFPOSX1_261 ( .CLK(sdram_clk_bF_buf63), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_x2b_pre_ok_r_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_x2b_pre_ok_t) );
  DFFPOSX1 DFFPOSX1_262 ( .CLK(sdram_clk_bF_buf62), .D(u_sdrc_core_u_bank_ctl_bank2_fsm_x2b_act_ok_r_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank2_fsm_x2b_act_ok_t) );
  DFFPOSX1 DFFPOSX1_263 ( .CLK(sdram_clk_bF_buf61), .D(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_17422_n90), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_0_) );
  DFFPOSX1 DFFPOSX1_264 ( .CLK(sdram_clk_bF_buf60), .D(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_17422_n61), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_prech_page_closed) );
  DFFPOSX1 DFFPOSX1_265 ( .CLK(sdram_clk_bF_buf59), .D(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_17422_n66), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_2_) );
  DFFPOSX1 DFFPOSX1_266 ( .CLK(sdram_clk_bF_buf58), .D(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_17422_n55), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_3_) );
  DFFPOSX1 DFFPOSX1_267 ( .CLK(sdram_clk_bF_buf57), .D(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_17422_n82), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_4_) );
  DFFPOSX1 DFFPOSX1_268 ( .CLK(sdram_clk_bF_buf56), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_l_last_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_l_last) );
  DFFPOSX1 DFFPOSX1_269 ( .CLK(sdram_clk_bF_buf55), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_l_wrap_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_l_wrap) );
  DFFPOSX1 DFFPOSX1_27 ( .CLK(sdram_clk_bF_buf54), .D(\sdr_dq[10] ), .Q(u_sdrc_core_pad_sdr_din1_10_) );
  DFFPOSX1 DFFPOSX1_270 ( .CLK(sdram_clk_bF_buf54), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_0__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_0_) );
  DFFPOSX1 DFFPOSX1_271 ( .CLK(sdram_clk_bF_buf53), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_1__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_1_) );
  DFFPOSX1 DFFPOSX1_272 ( .CLK(sdram_clk_bF_buf52), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_2__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_2_) );
  DFFPOSX1 DFFPOSX1_273 ( .CLK(sdram_clk_bF_buf51), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_3__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_3_) );
  DFFPOSX1 DFFPOSX1_274 ( .CLK(sdram_clk_bF_buf50), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_4__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_4_) );
  DFFPOSX1 DFFPOSX1_275 ( .CLK(sdram_clk_bF_buf49), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_5__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_5_) );
  DFFPOSX1 DFFPOSX1_276 ( .CLK(sdram_clk_bF_buf48), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_6__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_6_) );
  DFFPOSX1 DFFPOSX1_277 ( .CLK(sdram_clk_bF_buf47), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_0__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_0_) );
  DFFPOSX1 DFFPOSX1_278 ( .CLK(sdram_clk_bF_buf46), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_1__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_1_) );
  DFFPOSX1 DFFPOSX1_279 ( .CLK(sdram_clk_bF_buf45), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_2__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_2_) );
  DFFPOSX1 DFFPOSX1_28 ( .CLK(sdram_clk_bF_buf53), .D(\sdr_dq[11] ), .Q(u_sdrc_core_pad_sdr_din1_11_) );
  DFFPOSX1 DFFPOSX1_280 ( .CLK(sdram_clk_bF_buf44), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_3__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_3_) );
  DFFPOSX1 DFFPOSX1_281 ( .CLK(sdram_clk_bF_buf43), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_4__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_4_) );
  DFFPOSX1 DFFPOSX1_282 ( .CLK(sdram_clk_bF_buf42), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_5__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_5_) );
  DFFPOSX1 DFFPOSX1_283 ( .CLK(sdram_clk_bF_buf41), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_6__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_6_) );
  DFFPOSX1 DFFPOSX1_284 ( .CLK(sdram_clk_bF_buf40), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_7__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_7_) );
  DFFPOSX1 DFFPOSX1_285 ( .CLK(sdram_clk_bF_buf39), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_8__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_8_) );
  DFFPOSX1 DFFPOSX1_286 ( .CLK(sdram_clk_bF_buf38), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_9__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_9_) );
  DFFPOSX1 DFFPOSX1_287 ( .CLK(sdram_clk_bF_buf37), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_10__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_10_) );
  DFFPOSX1 DFFPOSX1_288 ( .CLK(sdram_clk_bF_buf36), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_11__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_11_) );
  DFFPOSX1 DFFPOSX1_289 ( .CLK(sdram_clk_bF_buf35), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_12__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_12_) );
  DFFPOSX1 DFFPOSX1_29 ( .CLK(sdram_clk_bF_buf52), .D(\sdr_dq[12] ), .Q(u_sdrc_core_pad_sdr_din1_12_) );
  DFFPOSX1 DFFPOSX1_290 ( .CLK(sdram_clk_bF_buf34), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_l_write_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_l_write) );
  DFFPOSX1 DFFPOSX1_291 ( .CLK(sdram_clk_bF_buf33), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_0__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_0_) );
  DFFPOSX1 DFFPOSX1_292 ( .CLK(sdram_clk_bF_buf32), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_1__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_1_) );
  DFFPOSX1 DFFPOSX1_293 ( .CLK(sdram_clk_bF_buf31), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_2__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_2_) );
  DFFPOSX1 DFFPOSX1_294 ( .CLK(sdram_clk_bF_buf30), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_3__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_3_) );
  DFFPOSX1 DFFPOSX1_295 ( .CLK(sdram_clk_bF_buf29), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_4__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_4_) );
  DFFPOSX1 DFFPOSX1_296 ( .CLK(sdram_clk_bF_buf28), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_5__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_5_) );
  DFFPOSX1 DFFPOSX1_297 ( .CLK(sdram_clk_bF_buf27), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_6__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_6_) );
  DFFPOSX1 DFFPOSX1_298 ( .CLK(sdram_clk_bF_buf26), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_7__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_7_) );
  DFFPOSX1 DFFPOSX1_299 ( .CLK(sdram_clk_bF_buf25), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_8__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_8_) );
  DFFPOSX1 DFFPOSX1_3 ( .CLK(sdram_clk_bF_buf78), .D(u_sdrc_core_pad_sdr_din1_2_), .Q(u_sdrc_core_pad_sdr_din2_2_) );
  DFFPOSX1 DFFPOSX1_30 ( .CLK(sdram_clk_bF_buf51), .D(\sdr_dq[13] ), .Q(u_sdrc_core_pad_sdr_din1_13_) );
  DFFPOSX1 DFFPOSX1_300 ( .CLK(sdram_clk_bF_buf24), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_9__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_9_) );
  DFFPOSX1 DFFPOSX1_301 ( .CLK(sdram_clk_bF_buf23), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_10__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_10_) );
  DFFPOSX1 DFFPOSX1_302 ( .CLK(sdram_clk_bF_buf22), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_11__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_11_) );
  DFFPOSX1 DFFPOSX1_303 ( .CLK(sdram_clk_bF_buf21), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_12__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_l_raddr_12_) );
  DFFPOSX1 DFFPOSX1_304 ( .CLK(sdram_clk_bF_buf20), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_0__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_0_) );
  DFFPOSX1 DFFPOSX1_305 ( .CLK(sdram_clk_bF_buf19), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_1__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_1_) );
  DFFPOSX1 DFFPOSX1_306 ( .CLK(sdram_clk_bF_buf18), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_2__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_2_) );
  DFFPOSX1 DFFPOSX1_307 ( .CLK(sdram_clk_bF_buf17), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_3__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_3_) );
  DFFPOSX1 DFFPOSX1_308 ( .CLK(sdram_clk_bF_buf16), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_4__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_4_) );
  DFFPOSX1 DFFPOSX1_309 ( .CLK(sdram_clk_bF_buf15), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_5__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_5_) );
  DFFPOSX1 DFFPOSX1_31 ( .CLK(sdram_clk_bF_buf50), .D(\sdr_dq[14] ), .Q(u_sdrc_core_pad_sdr_din1_14_) );
  DFFPOSX1 DFFPOSX1_310 ( .CLK(sdram_clk_bF_buf14), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_6__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_6_) );
  DFFPOSX1 DFFPOSX1_311 ( .CLK(sdram_clk_bF_buf13), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_7__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_7_) );
  DFFPOSX1 DFFPOSX1_312 ( .CLK(sdram_clk_bF_buf12), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_8__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_8_) );
  DFFPOSX1 DFFPOSX1_313 ( .CLK(sdram_clk_bF_buf11), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_9__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_9_) );
  DFFPOSX1 DFFPOSX1_314 ( .CLK(sdram_clk_bF_buf10), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_10__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_10_) );
  DFFPOSX1 DFFPOSX1_315 ( .CLK(sdram_clk_bF_buf9), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_11__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_11_) );
  DFFPOSX1 DFFPOSX1_316 ( .CLK(sdram_clk_bF_buf8), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_12__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_l_caddr_12_) );
  DFFPOSX1 DFFPOSX1_317 ( .CLK(sdram_clk_bF_buf7), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_l_sdr_dma_last_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_l_sdr_dma_last) );
  DFFPOSX1 DFFPOSX1_318 ( .CLK(sdram_clk_bF_buf6), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_valid_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_valid) );
  DFFPOSX1 DFFPOSX1_319 ( .CLK(sdram_clk_bF_buf5), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_tras_cntr_0__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_tras_cntr_0_) );
  DFFPOSX1 DFFPOSX1_32 ( .CLK(sdram_clk_bF_buf49), .D(\sdr_dq[15] ), .Q(u_sdrc_core_pad_sdr_din1_15_) );
  DFFPOSX1 DFFPOSX1_320 ( .CLK(sdram_clk_bF_buf4), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_tras_cntr_1__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_tras_cntr_1_) );
  DFFPOSX1 DFFPOSX1_321 ( .CLK(sdram_clk_bF_buf3), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_tras_cntr_2__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_tras_cntr_2_) );
  DFFPOSX1 DFFPOSX1_322 ( .CLK(sdram_clk_bF_buf2), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_tras_cntr_3__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_tras_cntr_3_) );
  DFFPOSX1 DFFPOSX1_323 ( .CLK(sdram_clk_bF_buf1), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_timer0_0__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_timer0_0_) );
  DFFPOSX1 DFFPOSX1_324 ( .CLK(sdram_clk_bF_buf0), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_timer0_1__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_timer0_1_) );
  DFFPOSX1 DFFPOSX1_325 ( .CLK(sdram_clk_bF_buf80), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_timer0_2__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_timer0_2_) );
  DFFPOSX1 DFFPOSX1_326 ( .CLK(sdram_clk_bF_buf79), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_timer0_3__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_timer0_3_) );
  DFFPOSX1 DFFPOSX1_327 ( .CLK(sdram_clk_bF_buf78), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_x2b_wrok_r_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_x2b_wrok_r) );
  DFFPOSX1 DFFPOSX1_328 ( .CLK(sdram_clk_bF_buf77), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_r_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_r) );
  DFFPOSX1 DFFPOSX1_329 ( .CLK(sdram_clk_bF_buf76), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_x2b_rdok_r_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_x2b_rdok_r) );
  DFFPOSX1 DFFPOSX1_33 ( .CLK(sdram_clk_bF_buf48), .D(u_sdrc_core_u_bank_ctl_rank_ba_0__FF_INPUT), .Q(u_sdrc_core_b2x_ba_0_) );
  DFFPOSX1 DFFPOSX1_330 ( .CLK(sdram_clk_bF_buf75), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_cmd_r_0__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_cmd_0_) );
  DFFPOSX1 DFFPOSX1_331 ( .CLK(sdram_clk_bF_buf74), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_cmd_r_1__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_cmd_1_) );
  DFFPOSX1 DFFPOSX1_332 ( .CLK(sdram_clk_bF_buf73), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_timer0_tc_r_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_timer0_tc) );
  DFFPOSX1 DFFPOSX1_333 ( .CLK(sdram_clk_bF_buf72), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_tras_ok_r_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_tras_ok) );
  DFFPOSX1 DFFPOSX1_334 ( .CLK(sdram_clk_bF_buf71), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_x2b_pre_ok_r_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_x2b_pre_ok_t) );
  DFFPOSX1 DFFPOSX1_335 ( .CLK(sdram_clk_bF_buf70), .D(u_sdrc_core_u_bank_ctl_bank3_fsm_x2b_act_ok_r_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank3_fsm_x2b_act_ok_t) );
  DFFPOSX1 DFFPOSX1_336 ( .CLK(sdram_clk_bF_buf69), .D(u_sdrc_core_u_bs_convert_saved_rd_data_0__FF_INPUT), .Q(u_sdrc_core_u_bs_convert_saved_rd_data_0_) );
  DFFPOSX1 DFFPOSX1_337 ( .CLK(sdram_clk_bF_buf68), .D(u_sdrc_core_u_bs_convert_saved_rd_data_1__FF_INPUT), .Q(u_sdrc_core_u_bs_convert_saved_rd_data_1_) );
  DFFPOSX1 DFFPOSX1_338 ( .CLK(sdram_clk_bF_buf67), .D(u_sdrc_core_u_bs_convert_saved_rd_data_2__FF_INPUT), .Q(u_sdrc_core_u_bs_convert_saved_rd_data_2_) );
  DFFPOSX1 DFFPOSX1_339 ( .CLK(sdram_clk_bF_buf66), .D(u_sdrc_core_u_bs_convert_saved_rd_data_3__FF_INPUT), .Q(u_sdrc_core_u_bs_convert_saved_rd_data_3_) );
  DFFPOSX1 DFFPOSX1_34 ( .CLK(sdram_clk_bF_buf47), .D(u_sdrc_core_u_bank_ctl_rank_ba_1__FF_INPUT), .Q(u_sdrc_core_b2x_ba_1_) );
  DFFPOSX1 DFFPOSX1_340 ( .CLK(sdram_clk_bF_buf65), .D(u_sdrc_core_u_bs_convert_saved_rd_data_4__FF_INPUT), .Q(u_sdrc_core_u_bs_convert_saved_rd_data_4_) );
  DFFPOSX1 DFFPOSX1_341 ( .CLK(sdram_clk_bF_buf64), .D(u_sdrc_core_u_bs_convert_saved_rd_data_5__FF_INPUT), .Q(u_sdrc_core_u_bs_convert_saved_rd_data_5_) );
  DFFPOSX1 DFFPOSX1_342 ( .CLK(sdram_clk_bF_buf63), .D(u_sdrc_core_u_bs_convert_saved_rd_data_6__FF_INPUT), .Q(u_sdrc_core_u_bs_convert_saved_rd_data_6_) );
  DFFPOSX1 DFFPOSX1_343 ( .CLK(sdram_clk_bF_buf62), .D(u_sdrc_core_u_bs_convert_saved_rd_data_7__FF_INPUT), .Q(u_sdrc_core_u_bs_convert_saved_rd_data_7_) );
  DFFPOSX1 DFFPOSX1_344 ( .CLK(sdram_clk_bF_buf61), .D(u_sdrc_core_u_bs_convert_saved_rd_data_8__FF_INPUT), .Q(u_sdrc_core_u_bs_convert_saved_rd_data_8_) );
  DFFPOSX1 DFFPOSX1_345 ( .CLK(sdram_clk_bF_buf60), .D(u_sdrc_core_u_bs_convert_saved_rd_data_9__FF_INPUT), .Q(u_sdrc_core_u_bs_convert_saved_rd_data_9_) );
  DFFPOSX1 DFFPOSX1_346 ( .CLK(sdram_clk_bF_buf59), .D(u_sdrc_core_u_bs_convert_saved_rd_data_10__FF_INPUT), .Q(u_sdrc_core_u_bs_convert_saved_rd_data_10_) );
  DFFPOSX1 DFFPOSX1_347 ( .CLK(sdram_clk_bF_buf58), .D(u_sdrc_core_u_bs_convert_saved_rd_data_11__FF_INPUT), .Q(u_sdrc_core_u_bs_convert_saved_rd_data_11_) );
  DFFPOSX1 DFFPOSX1_348 ( .CLK(sdram_clk_bF_buf57), .D(u_sdrc_core_u_bs_convert_saved_rd_data_12__FF_INPUT), .Q(u_sdrc_core_u_bs_convert_saved_rd_data_12_) );
  DFFPOSX1 DFFPOSX1_349 ( .CLK(sdram_clk_bF_buf56), .D(u_sdrc_core_u_bs_convert_saved_rd_data_13__FF_INPUT), .Q(u_sdrc_core_u_bs_convert_saved_rd_data_13_) );
  DFFPOSX1 DFFPOSX1_35 ( .CLK(sdram_clk_bF_buf46), .D(u_sdrc_core_u_bank_ctl_rank_ba_2__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_rank_ba_2_) );
  DFFPOSX1 DFFPOSX1_350 ( .CLK(sdram_clk_bF_buf55), .D(u_sdrc_core_u_bs_convert_saved_rd_data_14__FF_INPUT), .Q(u_sdrc_core_u_bs_convert_saved_rd_data_14_) );
  DFFPOSX1 DFFPOSX1_351 ( .CLK(sdram_clk_bF_buf54), .D(u_sdrc_core_u_bs_convert_saved_rd_data_15__FF_INPUT), .Q(u_sdrc_core_u_bs_convert_saved_rd_data_15_) );
  DFFPOSX1 DFFPOSX1_352 ( .CLK(sdram_clk_bF_buf53), .D(u_sdrc_core_u_bs_convert_saved_rd_data_16__FF_INPUT), .Q(u_sdrc_core_u_bs_convert_saved_rd_data_16_) );
  DFFPOSX1 DFFPOSX1_353 ( .CLK(sdram_clk_bF_buf52), .D(u_sdrc_core_u_bs_convert_saved_rd_data_17__FF_INPUT), .Q(u_sdrc_core_u_bs_convert_saved_rd_data_17_) );
  DFFPOSX1 DFFPOSX1_354 ( .CLK(sdram_clk_bF_buf51), .D(u_sdrc_core_u_bs_convert_saved_rd_data_18__FF_INPUT), .Q(u_sdrc_core_u_bs_convert_saved_rd_data_18_) );
  DFFPOSX1 DFFPOSX1_355 ( .CLK(sdram_clk_bF_buf50), .D(u_sdrc_core_u_bs_convert_saved_rd_data_19__FF_INPUT), .Q(u_sdrc_core_u_bs_convert_saved_rd_data_19_) );
  DFFPOSX1 DFFPOSX1_356 ( .CLK(sdram_clk_bF_buf49), .D(u_sdrc_core_u_bs_convert_saved_rd_data_20__FF_INPUT), .Q(u_sdrc_core_u_bs_convert_saved_rd_data_20_) );
  DFFPOSX1 DFFPOSX1_357 ( .CLK(sdram_clk_bF_buf48), .D(u_sdrc_core_u_bs_convert_saved_rd_data_21__FF_INPUT), .Q(u_sdrc_core_u_bs_convert_saved_rd_data_21_) );
  DFFPOSX1 DFFPOSX1_358 ( .CLK(sdram_clk_bF_buf47), .D(u_sdrc_core_u_bs_convert_saved_rd_data_22__FF_INPUT), .Q(u_sdrc_core_u_bs_convert_saved_rd_data_22_) );
  DFFPOSX1 DFFPOSX1_359 ( .CLK(sdram_clk_bF_buf46), .D(u_sdrc_core_u_bs_convert_saved_rd_data_23__FF_INPUT), .Q(u_sdrc_core_u_bs_convert_saved_rd_data_23_) );
  DFFPOSX1 DFFPOSX1_36 ( .CLK(sdram_clk_bF_buf45), .D(u_sdrc_core_u_bank_ctl_rank_ba_3__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_rank_ba_3_) );
  DFFPOSX1 DFFPOSX1_360 ( .CLK(sdram_clk_bF_buf45), .D(u_sdrc_core_u_bs_convert_rd_xfr_count_0__FF_INPUT), .Q(u_sdrc_core_u_bs_convert_rd_xfr_count_0_) );
  DFFPOSX1 DFFPOSX1_361 ( .CLK(sdram_clk_bF_buf44), .D(u_sdrc_core_u_bs_convert_rd_xfr_count_1__FF_INPUT), .Q(u_sdrc_core_u_bs_convert_rd_xfr_count_1_) );
  DFFPOSX1 DFFPOSX1_362 ( .CLK(sdram_clk_bF_buf43), .D(u_sdrc_core_u_bs_convert_wr_xfr_count_0__FF_INPUT), .Q(u_sdrc_core_u_bs_convert_wr_xfr_count_0_) );
  DFFPOSX1 DFFPOSX1_363 ( .CLK(sdram_clk_bF_buf42), .D(u_sdrc_core_u_bs_convert_wr_xfr_count_1__FF_INPUT), .Q(u_sdrc_core_u_bs_convert_wr_xfr_count_1_) );
  DFFPOSX1 DFFPOSX1_364 ( .CLK(sdram_clk_bF_buf41), .D(u_sdrc_core_u_req_gen__abc_16238_n57), .Q(u_sdrc_core_u_req_gen_req_st_0_) );
  DFFPOSX1 DFFPOSX1_365 ( .CLK(sdram_clk_bF_buf40), .D(u_sdrc_core_u_req_gen__abc_16238_n30), .Q(u_sdrc_core_u_req_gen_req_st_1_) );
  DFFPOSX1 DFFPOSX1_366 ( .CLK(sdram_clk_bF_buf39), .D(u_sdrc_core_u_req_gen__abc_16238_n38), .Q(u_sdrc_core_u_req_gen_req_st_2_) );
  DFFPOSX1 DFFPOSX1_367 ( .CLK(sdram_clk_bF_buf38), .D(u_sdrc_core_u_req_gen_r2b_ba_0__FF_INPUT), .Q(u_sdrc_core_r2b_ba_0_) );
  DFFPOSX1 DFFPOSX1_368 ( .CLK(sdram_clk_bF_buf37), .D(u_sdrc_core_u_req_gen_r2b_ba_1__FF_INPUT), .Q(u_sdrc_core_r2b_ba_1_) );
  DFFPOSX1 DFFPOSX1_369 ( .CLK(sdram_clk_bF_buf36), .D(u_sdrc_core_u_req_gen_r2b_raddr_0__FF_INPUT), .Q(u_sdrc_core_r2b_raddr_0_) );
  DFFPOSX1 DFFPOSX1_37 ( .CLK(sdram_clk_bF_buf44), .D(u_sdrc_core_u_bank_ctl_rank_ba_4__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_rank_ba_4_) );
  DFFPOSX1 DFFPOSX1_370 ( .CLK(sdram_clk_bF_buf35), .D(u_sdrc_core_u_req_gen_r2b_raddr_1__FF_INPUT), .Q(u_sdrc_core_r2b_raddr_1_) );
  DFFPOSX1 DFFPOSX1_371 ( .CLK(sdram_clk_bF_buf34), .D(u_sdrc_core_u_req_gen_r2b_raddr_2__FF_INPUT), .Q(u_sdrc_core_r2b_raddr_2_) );
  DFFPOSX1 DFFPOSX1_372 ( .CLK(sdram_clk_bF_buf33), .D(u_sdrc_core_u_req_gen_r2b_raddr_3__FF_INPUT), .Q(u_sdrc_core_r2b_raddr_3_) );
  DFFPOSX1 DFFPOSX1_373 ( .CLK(sdram_clk_bF_buf32), .D(u_sdrc_core_u_req_gen_r2b_raddr_4__FF_INPUT), .Q(u_sdrc_core_r2b_raddr_4_) );
  DFFPOSX1 DFFPOSX1_374 ( .CLK(sdram_clk_bF_buf31), .D(u_sdrc_core_u_req_gen_r2b_raddr_5__FF_INPUT), .Q(u_sdrc_core_r2b_raddr_5_) );
  DFFPOSX1 DFFPOSX1_375 ( .CLK(sdram_clk_bF_buf30), .D(u_sdrc_core_u_req_gen_r2b_raddr_6__FF_INPUT), .Q(u_sdrc_core_r2b_raddr_6_) );
  DFFPOSX1 DFFPOSX1_376 ( .CLK(sdram_clk_bF_buf29), .D(u_sdrc_core_u_req_gen_r2b_raddr_7__FF_INPUT), .Q(u_sdrc_core_r2b_raddr_7_) );
  DFFPOSX1 DFFPOSX1_377 ( .CLK(sdram_clk_bF_buf28), .D(u_sdrc_core_u_req_gen_r2b_raddr_8__FF_INPUT), .Q(u_sdrc_core_r2b_raddr_8_) );
  DFFPOSX1 DFFPOSX1_378 ( .CLK(sdram_clk_bF_buf27), .D(u_sdrc_core_u_req_gen_r2b_raddr_9__FF_INPUT), .Q(u_sdrc_core_r2b_raddr_9_) );
  DFFPOSX1 DFFPOSX1_379 ( .CLK(sdram_clk_bF_buf26), .D(u_sdrc_core_u_req_gen_r2b_raddr_10__FF_INPUT), .Q(u_sdrc_core_r2b_raddr_10_) );
  DFFPOSX1 DFFPOSX1_38 ( .CLK(sdram_clk_bF_buf43), .D(u_sdrc_core_u_bank_ctl_rank_ba_5__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_rank_ba_5_) );
  DFFPOSX1 DFFPOSX1_380 ( .CLK(sdram_clk_bF_buf25), .D(u_sdrc_core_u_req_gen_r2b_raddr_11__FF_INPUT), .Q(u_sdrc_core_r2b_raddr_11_) );
  DFFPOSX1 DFFPOSX1_381 ( .CLK(sdram_clk_bF_buf24), .D(u_sdrc_core_u_req_gen_r2b_raddr_12__FF_INPUT), .Q(u_sdrc_core_r2b_raddr_12_) );
  DFFPOSX1 DFFPOSX1_382 ( .CLK(sdram_clk_bF_buf23), .D(u_sdrc_core_u_req_gen_r2b_caddr_8__FF_INPUT), .Q(u_sdrc_core_r2b_caddr_8_) );
  DFFPOSX1 DFFPOSX1_383 ( .CLK(sdram_clk_bF_buf22), .D(u_sdrc_core_u_req_gen_r2b_caddr_9__FF_INPUT), .Q(u_sdrc_core_r2b_caddr_9_) );
  DFFPOSX1 DFFPOSX1_384 ( .CLK(sdram_clk_bF_buf21), .D(u_sdrc_core_u_req_gen_r2b_caddr_10__FF_INPUT), .Q(u_sdrc_core_r2b_caddr_10_) );
  DFFPOSX1 DFFPOSX1_385 ( .CLK(sdram_clk_bF_buf20), .D(u_sdrc_core_u_req_gen_r2b_start_FF_INPUT), .Q(u_sdrc_core_r2b_start) );
  DFFPOSX1 DFFPOSX1_386 ( .CLK(sdram_clk_bF_buf19), .D(u_sdrc_core_u_req_gen_r2b_write_FF_INPUT), .Q(u_sdrc_core_r2b_write) );
  DFFPOSX1 DFFPOSX1_387 ( .CLK(sdram_clk_bF_buf18), .D(u_sdrc_core_u_req_gen_lcl_wrap_FF_INPUT), .Q(u_sdrc_core_r2b_wrap) );
  DFFPOSX1 DFFPOSX1_388 ( .CLK(sdram_clk_bF_buf17), .D(u_sdrc_core_u_req_gen_lcl_req_len_0__FF_INPUT), .Q(u_sdrc_core_u_req_gen_lcl_req_len_0_) );
  DFFPOSX1 DFFPOSX1_389 ( .CLK(sdram_clk_bF_buf16), .D(u_sdrc_core_u_req_gen_lcl_req_len_1__FF_INPUT), .Q(u_sdrc_core_u_req_gen_lcl_req_len_1_) );
  DFFPOSX1 DFFPOSX1_39 ( .CLK(sdram_clk_bF_buf42), .D(u_sdrc_core_u_bank_ctl_rank_ba_6__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_rank_ba_6_) );
  DFFPOSX1 DFFPOSX1_390 ( .CLK(sdram_clk_bF_buf15), .D(u_sdrc_core_u_req_gen_lcl_req_len_2__FF_INPUT), .Q(u_sdrc_core_u_req_gen_lcl_req_len_2_) );
  DFFPOSX1 DFFPOSX1_391 ( .CLK(sdram_clk_bF_buf14), .D(u_sdrc_core_u_req_gen_lcl_req_len_3__FF_INPUT), .Q(u_sdrc_core_u_req_gen_lcl_req_len_3_) );
  DFFPOSX1 DFFPOSX1_392 ( .CLK(sdram_clk_bF_buf13), .D(u_sdrc_core_u_req_gen_lcl_req_len_4__FF_INPUT), .Q(u_sdrc_core_u_req_gen_lcl_req_len_4_) );
  DFFPOSX1 DFFPOSX1_393 ( .CLK(sdram_clk_bF_buf12), .D(u_sdrc_core_u_req_gen_lcl_req_len_5__FF_INPUT), .Q(u_sdrc_core_u_req_gen_lcl_req_len_5_) );
  DFFPOSX1 DFFPOSX1_394 ( .CLK(sdram_clk_bF_buf11), .D(u_sdrc_core_u_req_gen_lcl_req_len_6__FF_INPUT), .Q(u_sdrc_core_u_req_gen_lcl_req_len_6_) );
  DFFPOSX1 DFFPOSX1_395 ( .CLK(sdram_clk_bF_buf10), .D(u_sdrc_core_u_req_gen_page_ovflw_r_FF_INPUT), .Q(u_sdrc_core_u_req_gen_page_ovflw_r) );
  DFFPOSX1 DFFPOSX1_396 ( .CLK(sdram_clk_bF_buf9), .D(u_sdrc_core_u_req_gen_max_r2b_len_r_0__FF_INPUT), .Q(u_sdrc_core_u_req_gen_max_r2b_len_r_0_) );
  DFFPOSX1 DFFPOSX1_397 ( .CLK(sdram_clk_bF_buf8), .D(u_sdrc_core_u_req_gen_max_r2b_len_r_1__FF_INPUT), .Q(u_sdrc_core_u_req_gen_max_r2b_len_r_1_) );
  DFFPOSX1 DFFPOSX1_398 ( .CLK(sdram_clk_bF_buf7), .D(u_sdrc_core_u_req_gen_max_r2b_len_r_2__FF_INPUT), .Q(u_sdrc_core_u_req_gen_max_r2b_len_r_2_) );
  DFFPOSX1 DFFPOSX1_399 ( .CLK(sdram_clk_bF_buf6), .D(u_sdrc_core_u_req_gen_max_r2b_len_r_3__FF_INPUT), .Q(u_sdrc_core_u_req_gen_max_r2b_len_r_3_) );
  DFFPOSX1 DFFPOSX1_4 ( .CLK(sdram_clk_bF_buf77), .D(u_sdrc_core_pad_sdr_din1_3_), .Q(u_sdrc_core_pad_sdr_din2_3_) );
  DFFPOSX1 DFFPOSX1_40 ( .CLK(sdram_clk_bF_buf41), .D(u_sdrc_core_u_bank_ctl_rank_ba_7__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_rank_ba_7_) );
  DFFPOSX1 DFFPOSX1_400 ( .CLK(sdram_clk_bF_buf5), .D(u_sdrc_core_u_req_gen_max_r2b_len_r_4__FF_INPUT), .Q(u_sdrc_core_u_req_gen_max_r2b_len_r_4_) );
  DFFPOSX1 DFFPOSX1_401 ( .CLK(sdram_clk_bF_buf4), .D(u_sdrc_core_u_req_gen_max_r2b_len_r_5__FF_INPUT), .Q(u_sdrc_core_u_req_gen_max_r2b_len_r_5_) );
  DFFPOSX1 DFFPOSX1_402 ( .CLK(sdram_clk_bF_buf3), .D(u_sdrc_core_u_req_gen_max_r2b_len_r_6__FF_INPUT), .Q(u_sdrc_core_u_req_gen_max_r2b_len_r_6_) );
  DFFPOSX1 DFFPOSX1_403 ( .CLK(sdram_clk_bF_buf2), .D(u_sdrc_core_u_req_gen_map_address_0_), .Q(u_sdrc_core_r2b_caddr_0_) );
  DFFPOSX1 DFFPOSX1_404 ( .CLK(sdram_clk_bF_buf1), .D(u_sdrc_core_u_req_gen_map_address_1_), .Q(u_sdrc_core_r2b_caddr_1_) );
  DFFPOSX1 DFFPOSX1_405 ( .CLK(sdram_clk_bF_buf0), .D(u_sdrc_core_u_req_gen_map_address_2_), .Q(u_sdrc_core_r2b_caddr_2_) );
  DFFPOSX1 DFFPOSX1_406 ( .CLK(sdram_clk_bF_buf80), .D(u_sdrc_core_u_req_gen_map_address_3_), .Q(u_sdrc_core_r2b_caddr_3_) );
  DFFPOSX1 DFFPOSX1_407 ( .CLK(sdram_clk_bF_buf79), .D(u_sdrc_core_u_req_gen_map_address_4_), .Q(u_sdrc_core_r2b_caddr_4_) );
  DFFPOSX1 DFFPOSX1_408 ( .CLK(sdram_clk_bF_buf78), .D(u_sdrc_core_u_req_gen_map_address_5_), .Q(u_sdrc_core_r2b_caddr_5_) );
  DFFPOSX1 DFFPOSX1_409 ( .CLK(sdram_clk_bF_buf77), .D(u_sdrc_core_u_req_gen_map_address_6_), .Q(u_sdrc_core_r2b_caddr_6_) );
  DFFPOSX1 DFFPOSX1_41 ( .CLK(sdram_clk_bF_buf40), .D(u_sdrc_core_u_bank_ctl_rank_cnt_0__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_rank_cnt_0_) );
  DFFPOSX1 DFFPOSX1_410 ( .CLK(sdram_clk_bF_buf76), .D(u_sdrc_core_u_req_gen_map_address_7_), .Q(u_sdrc_core_r2b_caddr_7_) );
  DFFPOSX1 DFFPOSX1_411 ( .CLK(sdram_clk_bF_buf75), .D(u_sdrc_core_u_req_gen_map_address_8_), .Q(u_sdrc_core_u_req_gen_curr_sdr_addr_8_) );
  DFFPOSX1 DFFPOSX1_412 ( .CLK(sdram_clk_bF_buf74), .D(u_sdrc_core_u_req_gen_map_address_9_), .Q(u_sdrc_core_u_req_gen_curr_sdr_addr_9_) );
  DFFPOSX1 DFFPOSX1_413 ( .CLK(sdram_clk_bF_buf73), .D(u_sdrc_core_u_req_gen_map_address_10_), .Q(u_sdrc_core_u_req_gen_curr_sdr_addr_10_) );
  DFFPOSX1 DFFPOSX1_414 ( .CLK(sdram_clk_bF_buf72), .D(u_sdrc_core_u_req_gen_map_address_11_), .Q(u_sdrc_core_u_req_gen_curr_sdr_addr_11_) );
  DFFPOSX1 DFFPOSX1_415 ( .CLK(sdram_clk_bF_buf71), .D(u_sdrc_core_u_req_gen_map_address_12_), .Q(u_sdrc_core_u_req_gen_curr_sdr_addr_12_) );
  DFFPOSX1 DFFPOSX1_416 ( .CLK(sdram_clk_bF_buf70), .D(u_sdrc_core_u_req_gen_map_address_13_), .Q(u_sdrc_core_u_req_gen_curr_sdr_addr_13_) );
  DFFPOSX1 DFFPOSX1_417 ( .CLK(sdram_clk_bF_buf69), .D(u_sdrc_core_u_req_gen_map_address_14_), .Q(u_sdrc_core_u_req_gen_curr_sdr_addr_14_) );
  DFFPOSX1 DFFPOSX1_418 ( .CLK(sdram_clk_bF_buf68), .D(u_sdrc_core_u_req_gen_map_address_15_), .Q(u_sdrc_core_u_req_gen_curr_sdr_addr_15_) );
  DFFPOSX1 DFFPOSX1_419 ( .CLK(sdram_clk_bF_buf67), .D(u_sdrc_core_u_req_gen_map_address_16_), .Q(u_sdrc_core_u_req_gen_curr_sdr_addr_16_) );
  DFFPOSX1 DFFPOSX1_42 ( .CLK(sdram_clk_bF_buf39), .D(u_sdrc_core_u_bank_ctl_rank_cnt_1__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_rank_cnt_1_) );
  DFFPOSX1 DFFPOSX1_420 ( .CLK(sdram_clk_bF_buf66), .D(u_sdrc_core_u_req_gen_map_address_17_), .Q(u_sdrc_core_u_req_gen_curr_sdr_addr_17_) );
  DFFPOSX1 DFFPOSX1_421 ( .CLK(sdram_clk_bF_buf65), .D(u_sdrc_core_u_req_gen_map_address_18_), .Q(u_sdrc_core_u_req_gen_curr_sdr_addr_18_) );
  DFFPOSX1 DFFPOSX1_422 ( .CLK(sdram_clk_bF_buf64), .D(u_sdrc_core_u_req_gen_map_address_19_), .Q(u_sdrc_core_u_req_gen_curr_sdr_addr_19_) );
  DFFPOSX1 DFFPOSX1_423 ( .CLK(sdram_clk_bF_buf63), .D(u_sdrc_core_u_req_gen_map_address_20_), .Q(u_sdrc_core_u_req_gen_curr_sdr_addr_20_) );
  DFFPOSX1 DFFPOSX1_424 ( .CLK(sdram_clk_bF_buf62), .D(u_sdrc_core_u_req_gen_map_address_21_), .Q(u_sdrc_core_u_req_gen_curr_sdr_addr_21_) );
  DFFPOSX1 DFFPOSX1_425 ( .CLK(sdram_clk_bF_buf61), .D(u_sdrc_core_u_req_gen_map_address_22_), .Q(u_sdrc_core_u_req_gen_curr_sdr_addr_22_) );
  DFFPOSX1 DFFPOSX1_426 ( .CLK(sdram_clk_bF_buf60), .D(u_sdrc_core_u_req_gen_map_address_23_), .Q(u_sdrc_core_u_req_gen_curr_sdr_addr_23_) );
  DFFPOSX1 DFFPOSX1_427 ( .CLK(sdram_clk_bF_buf59), .D(u_sdrc_core_u_req_gen_map_address_24_), .Q(u_sdrc_core_u_req_gen_curr_sdr_addr_24_) );
  DFFPOSX1 DFFPOSX1_428 ( .CLK(sdram_clk_bF_buf58), .D(u_sdrc_core_u_req_gen_map_address_25_), .Q(u_sdrc_core_u_req_gen_curr_sdr_addr_25_) );
  DFFPOSX1 DFFPOSX1_429 ( .CLK(sdram_clk_bF_buf57), .D(u_sdrc_core_u_xfr_ctl__abc_16728_n178), .Q(u_sdrc_core_u_xfr_ctl_mgmt_st_0_) );
  DFFPOSX1 DFFPOSX1_43 ( .CLK(sdram_clk_bF_buf38), .D(u_sdrc_core_u_bank_ctl_rank_cnt_2__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_rank_cnt_2_) );
  DFFPOSX1 DFFPOSX1_430 ( .CLK(sdram_clk_bF_buf56), .D(u_sdrc_core_u_xfr_ctl__abc_16728_n181), .Q(u_sdrc_core_u_xfr_ctl_mgmt_st_1_) );
  DFFPOSX1 DFFPOSX1_431 ( .CLK(sdram_clk_bF_buf55), .D(u_sdrc_core_u_xfr_ctl__abc_16728_n270), .Q(u_sdrc_core_u_xfr_ctl_mgmt_st_2_) );
  DFFPOSX1 DFFPOSX1_432 ( .CLK(sdram_clk_bF_buf54), .D(u_sdrc_core_u_xfr_ctl__abc_16728_n258), .Q(u_sdrc_core_u_xfr_ctl_mgmt_st_3_) );
  DFFPOSX1 DFFPOSX1_433 ( .CLK(sdram_clk_bF_buf53), .D(u_sdrc_core_u_xfr_ctl__abc_16728_n189), .Q(u_sdrc_core_u_xfr_ctl_mgmt_st_4_) );
  DFFPOSX1 DFFPOSX1_434 ( .CLK(sdram_clk_bF_buf52), .D(u_sdrc_core_u_xfr_ctl__abc_16728_n184), .Q(u_sdrc_core_u_xfr_ctl_mgmt_st_5_) );
  DFFPOSX1 DFFPOSX1_435 ( .CLK(sdram_clk_bF_buf51), .D(u_sdrc_core_u_xfr_ctl__abc_16728_n43), .Q(u_sdrc_core_u_xfr_ctl_mgmt_st_6_) );
  DFFPOSX1 DFFPOSX1_436 ( .CLK(sdram_clk_bF_buf50), .D(u_sdrc_core_u_xfr_ctl__abc_16728_n35), .Q(u_sdrc_core_u_xfr_ctl_mgmt_st_7_) );
  DFFPOSX1 DFFPOSX1_437 ( .CLK(sdram_clk_bF_buf49), .D(u_sdrc_core_u_xfr_ctl_sdr_init_done_FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_24701) );
  DFFPOSX1 DFFPOSX1_438 ( .CLK(sdram_clk_bF_buf48), .D(u_sdrc_core_u_xfr_ctl_tmr0_0__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_tmr0_0_) );
  DFFPOSX1 DFFPOSX1_439 ( .CLK(sdram_clk_bF_buf47), .D(u_sdrc_core_u_xfr_ctl_tmr0_1__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_tmr0_1_) );
  DFFPOSX1 DFFPOSX1_44 ( .CLK(sdram_clk_bF_buf37), .D(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_17422_n90), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_0_) );
  DFFPOSX1 DFFPOSX1_440 ( .CLK(sdram_clk_bF_buf46), .D(u_sdrc_core_u_xfr_ctl_tmr0_2__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_tmr0_2_) );
  DFFPOSX1 DFFPOSX1_441 ( .CLK(sdram_clk_bF_buf45), .D(u_sdrc_core_u_xfr_ctl_tmr0_3__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_tmr0_3_) );
  DFFPOSX1 DFFPOSX1_442 ( .CLK(sdram_clk_bF_buf44), .D(u_sdrc_core_u_xfr_ctl_cntr1_0__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_cntr1_0_) );
  DFFPOSX1 DFFPOSX1_443 ( .CLK(sdram_clk_bF_buf43), .D(u_sdrc_core_u_xfr_ctl_cntr1_1__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_cntr1_1_) );
  DFFPOSX1 DFFPOSX1_444 ( .CLK(sdram_clk_bF_buf42), .D(u_sdrc_core_u_xfr_ctl_cntr1_2__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_cntr1_2_) );
  DFFPOSX1 DFFPOSX1_445 ( .CLK(sdram_clk_bF_buf41), .D(u_sdrc_core_u_xfr_ctl_cntr1_3__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_cntr1_3_) );
  DFFPOSX1 DFFPOSX1_446 ( .CLK(sdram_clk_bF_buf40), .D(u_sdrc_core_u_xfr_ctl_rfsh_timer_0__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_rfsh_timer_0_) );
  DFFPOSX1 DFFPOSX1_447 ( .CLK(sdram_clk_bF_buf39), .D(u_sdrc_core_u_xfr_ctl_rfsh_timer_1__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_rfsh_timer_1_) );
  DFFPOSX1 DFFPOSX1_448 ( .CLK(sdram_clk_bF_buf38), .D(u_sdrc_core_u_xfr_ctl_rfsh_timer_2__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_rfsh_timer_2_) );
  DFFPOSX1 DFFPOSX1_449 ( .CLK(sdram_clk_bF_buf37), .D(u_sdrc_core_u_xfr_ctl_rfsh_timer_3__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_rfsh_timer_3_) );
  DFFPOSX1 DFFPOSX1_45 ( .CLK(sdram_clk_bF_buf36), .D(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_17422_n61), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_prech_page_closed) );
  DFFPOSX1 DFFPOSX1_450 ( .CLK(sdram_clk_bF_buf36), .D(u_sdrc_core_u_xfr_ctl_rfsh_timer_4__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_rfsh_timer_4_) );
  DFFPOSX1 DFFPOSX1_451 ( .CLK(sdram_clk_bF_buf35), .D(u_sdrc_core_u_xfr_ctl_rfsh_timer_5__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_rfsh_timer_5_) );
  DFFPOSX1 DFFPOSX1_452 ( .CLK(sdram_clk_bF_buf34), .D(u_sdrc_core_u_xfr_ctl_rfsh_timer_6__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_rfsh_timer_6_) );
  DFFPOSX1 DFFPOSX1_453 ( .CLK(sdram_clk_bF_buf33), .D(u_sdrc_core_u_xfr_ctl_rfsh_timer_7__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_rfsh_timer_7_) );
  DFFPOSX1 DFFPOSX1_454 ( .CLK(sdram_clk_bF_buf32), .D(u_sdrc_core_u_xfr_ctl_rfsh_timer_8__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_rfsh_timer_8_) );
  DFFPOSX1 DFFPOSX1_455 ( .CLK(sdram_clk_bF_buf31), .D(u_sdrc_core_u_xfr_ctl_rfsh_timer_9__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_rfsh_timer_9_) );
  DFFPOSX1 DFFPOSX1_456 ( .CLK(sdram_clk_bF_buf30), .D(u_sdrc_core_u_xfr_ctl_rfsh_timer_10__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_rfsh_timer_10_) );
  DFFPOSX1 DFFPOSX1_457 ( .CLK(sdram_clk_bF_buf29), .D(u_sdrc_core_u_xfr_ctl_rfsh_timer_11__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_rfsh_timer_11_) );
  DFFPOSX1 DFFPOSX1_458 ( .CLK(sdram_clk_bF_buf28), .D(u_sdrc_core_u_xfr_ctl_rfsh_row_cnt_0__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_rfsh_row_cnt_0_) );
  DFFPOSX1 DFFPOSX1_459 ( .CLK(sdram_clk_bF_buf27), .D(u_sdrc_core_u_xfr_ctl_rfsh_row_cnt_1__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_rfsh_row_cnt_1_) );
  DFFPOSX1 DFFPOSX1_46 ( .CLK(sdram_clk_bF_buf35), .D(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_17422_n66), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_2_) );
  DFFPOSX1 DFFPOSX1_460 ( .CLK(sdram_clk_bF_buf26), .D(u_sdrc_core_u_xfr_ctl_rfsh_row_cnt_2__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_rfsh_row_cnt_2_) );
  DFFPOSX1 DFFPOSX1_461 ( .CLK(sdram_clk_bF_buf25), .D(u_sdrc_core_u_xfr_ctl_sdr_ba_0__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_24689_0_) );
  DFFPOSX1 DFFPOSX1_462 ( .CLK(sdram_clk_bF_buf24), .D(u_sdrc_core_u_xfr_ctl_sdr_ba_1__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_24689_1_) );
  DFFPOSX1 DFFPOSX1_463 ( .CLK(sdram_clk_bF_buf23), .D(u_sdrc_core_u_xfr_ctl_sdr_addr_0__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_24675_0_) );
  DFFPOSX1 DFFPOSX1_464 ( .CLK(sdram_clk_bF_buf22), .D(u_sdrc_core_u_xfr_ctl_sdr_addr_1__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_24675_1_) );
  DFFPOSX1 DFFPOSX1_465 ( .CLK(sdram_clk_bF_buf21), .D(u_sdrc_core_u_xfr_ctl_sdr_addr_2__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_24675_2_) );
  DFFPOSX1 DFFPOSX1_466 ( .CLK(sdram_clk_bF_buf20), .D(u_sdrc_core_u_xfr_ctl_sdr_addr_3__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_24675_3_) );
  DFFPOSX1 DFFPOSX1_467 ( .CLK(sdram_clk_bF_buf19), .D(u_sdrc_core_u_xfr_ctl_sdr_addr_4__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_24675_4_) );
  DFFPOSX1 DFFPOSX1_468 ( .CLK(sdram_clk_bF_buf18), .D(u_sdrc_core_u_xfr_ctl_sdr_addr_5__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_24675_5_) );
  DFFPOSX1 DFFPOSX1_469 ( .CLK(sdram_clk_bF_buf17), .D(u_sdrc_core_u_xfr_ctl_sdr_addr_6__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_24675_6_) );
  DFFPOSX1 DFFPOSX1_47 ( .CLK(sdram_clk_bF_buf34), .D(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_17422_n55), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_3_) );
  DFFPOSX1 DFFPOSX1_470 ( .CLK(sdram_clk_bF_buf16), .D(u_sdrc_core_u_xfr_ctl_sdr_addr_7__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_24675_7_) );
  DFFPOSX1 DFFPOSX1_471 ( .CLK(sdram_clk_bF_buf15), .D(u_sdrc_core_u_xfr_ctl_sdr_addr_8__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_24675_8_) );
  DFFPOSX1 DFFPOSX1_472 ( .CLK(sdram_clk_bF_buf14), .D(u_sdrc_core_u_xfr_ctl_sdr_addr_9__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_24675_9_) );
  DFFPOSX1 DFFPOSX1_473 ( .CLK(sdram_clk_bF_buf13), .D(u_sdrc_core_u_xfr_ctl_sdr_addr_10__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_24675_10_) );
  DFFPOSX1 DFFPOSX1_474 ( .CLK(sdram_clk_bF_buf12), .D(u_sdrc_core_u_xfr_ctl_sdr_addr_11__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_24675_11_) );
  DFFPOSX1 DFFPOSX1_475 ( .CLK(sdram_clk_bF_buf11), .D(u_sdrc_core_u_xfr_ctl_sdr_addr_12__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_24675_12_) );
  DFFPOSX1 DFFPOSX1_476 ( .CLK(sdram_clk_bF_buf10), .D(u_sdrc_core_u_xfr_ctl_sdr_dout_0__FF_INPUT), .Q(\sdr_dq[0] ) );
  DFFPOSX1 DFFPOSX1_477 ( .CLK(sdram_clk_bF_buf9), .D(u_sdrc_core_u_xfr_ctl_sdr_dout_1__FF_INPUT), .Q(\sdr_dq[1] ) );
  DFFPOSX1 DFFPOSX1_478 ( .CLK(sdram_clk_bF_buf8), .D(u_sdrc_core_u_xfr_ctl_sdr_dout_2__FF_INPUT), .Q(\sdr_dq[2] ) );
  DFFPOSX1 DFFPOSX1_479 ( .CLK(sdram_clk_bF_buf7), .D(u_sdrc_core_u_xfr_ctl_sdr_dout_3__FF_INPUT), .Q(\sdr_dq[3] ) );
  DFFPOSX1 DFFPOSX1_48 ( .CLK(sdram_clk_bF_buf33), .D(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_17422_n82), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_4_) );
  DFFPOSX1 DFFPOSX1_480 ( .CLK(sdram_clk_bF_buf6), .D(u_sdrc_core_u_xfr_ctl_sdr_dout_4__FF_INPUT), .Q(\sdr_dq[4] ) );
  DFFPOSX1 DFFPOSX1_481 ( .CLK(sdram_clk_bF_buf5), .D(u_sdrc_core_u_xfr_ctl_sdr_dout_5__FF_INPUT), .Q(\sdr_dq[5] ) );
  DFFPOSX1 DFFPOSX1_482 ( .CLK(sdram_clk_bF_buf4), .D(u_sdrc_core_u_xfr_ctl_sdr_dout_6__FF_INPUT), .Q(\sdr_dq[6] ) );
  DFFPOSX1 DFFPOSX1_483 ( .CLK(sdram_clk_bF_buf3), .D(u_sdrc_core_u_xfr_ctl_sdr_dout_7__FF_INPUT), .Q(\sdr_dq[7] ) );
  DFFPOSX1 DFFPOSX1_484 ( .CLK(sdram_clk_bF_buf2), .D(u_sdrc_core_u_xfr_ctl_sdr_dout_8__FF_INPUT), .Q(\sdr_dq[8] ) );
  DFFPOSX1 DFFPOSX1_485 ( .CLK(sdram_clk_bF_buf1), .D(u_sdrc_core_u_xfr_ctl_sdr_dout_9__FF_INPUT), .Q(\sdr_dq[9] ) );
  DFFPOSX1 DFFPOSX1_486 ( .CLK(sdram_clk_bF_buf0), .D(u_sdrc_core_u_xfr_ctl_sdr_dout_10__FF_INPUT), .Q(\sdr_dq[10] ) );
  DFFPOSX1 DFFPOSX1_487 ( .CLK(sdram_clk_bF_buf80), .D(u_sdrc_core_u_xfr_ctl_sdr_dout_11__FF_INPUT), .Q(\sdr_dq[11] ) );
  DFFPOSX1 DFFPOSX1_488 ( .CLK(sdram_clk_bF_buf79), .D(u_sdrc_core_u_xfr_ctl_sdr_dout_12__FF_INPUT), .Q(\sdr_dq[12] ) );
  DFFPOSX1 DFFPOSX1_489 ( .CLK(sdram_clk_bF_buf78), .D(u_sdrc_core_u_xfr_ctl_sdr_dout_13__FF_INPUT), .Q(\sdr_dq[13] ) );
  DFFPOSX1 DFFPOSX1_49 ( .CLK(sdram_clk_bF_buf32), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_l_last_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_l_last) );
  DFFPOSX1 DFFPOSX1_490 ( .CLK(sdram_clk_bF_buf77), .D(u_sdrc_core_u_xfr_ctl_sdr_dout_14__FF_INPUT), .Q(\sdr_dq[14] ) );
  DFFPOSX1 DFFPOSX1_491 ( .CLK(sdram_clk_bF_buf76), .D(u_sdrc_core_u_xfr_ctl_sdr_dout_15__FF_INPUT), .Q(\sdr_dq[15] ) );
  DFFPOSX1 DFFPOSX1_492 ( .CLK(sdram_clk_bF_buf75), .D(u_sdrc_core_u_xfr_ctl_sdr_cke_FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_24694) );
  DFFPOSX1 DFFPOSX1_493 ( .CLK(sdram_clk_bF_buf74), .D(u_sdrc_core_u_xfr_ctl_sdr_cs_n_FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_24696) );
  DFFPOSX1 DFFPOSX1_494 ( .CLK(sdram_clk_bF_buf73), .D(u_sdrc_core_u_xfr_ctl_sdr_ras_n_FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_24703) );
  DFFPOSX1 DFFPOSX1_495 ( .CLK(sdram_clk_bF_buf72), .D(u_sdrc_core_u_xfr_ctl_sdr_cas_n_FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_24692) );
  DFFPOSX1 DFFPOSX1_496 ( .CLK(sdram_clk_bF_buf71), .D(u_sdrc_core_u_xfr_ctl_sdr_we_n_FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_24705) );
  DFFPOSX1 DFFPOSX1_497 ( .CLK(sdram_clk_bF_buf70), .D(u_sdrc_core_u_xfr_ctl_sdr_dqm_0__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_24698_0_) );
  DFFPOSX1 DFFPOSX1_498 ( .CLK(sdram_clk_bF_buf69), .D(u_sdrc_core_u_xfr_ctl_sdr_dqm_1__FF_INPUT), .Q(_auto_iopadmap_cc_313_execute_24698_1_) );
  DFFPOSX1 DFFPOSX1_499 ( .CLK(sdram_clk_bF_buf68), .D(u_sdrc_core_u_xfr_ctl_xfr_st_0__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_xfr_st_0_) );
  DFFPOSX1 DFFPOSX1_5 ( .CLK(sdram_clk_bF_buf76), .D(u_sdrc_core_pad_sdr_din1_4_), .Q(u_sdrc_core_pad_sdr_din2_4_) );
  DFFPOSX1 DFFPOSX1_50 ( .CLK(sdram_clk_bF_buf31), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_l_wrap_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_l_wrap) );
  DFFPOSX1 DFFPOSX1_500 ( .CLK(sdram_clk_bF_buf67), .D(u_sdrc_core_u_xfr_ctl_xfr_st_1__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_xfr_st_1_) );
  DFFPOSX1 DFFPOSX1_501 ( .CLK(sdram_clk_bF_buf66), .D(u_sdrc_core_u_xfr_ctl_xfr_caddr_0__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_xfr_caddr_0_) );
  DFFPOSX1 DFFPOSX1_502 ( .CLK(sdram_clk_bF_buf65), .D(u_sdrc_core_u_xfr_ctl_xfr_caddr_1__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_xfr_caddr_1_) );
  DFFPOSX1 DFFPOSX1_503 ( .CLK(sdram_clk_bF_buf64), .D(u_sdrc_core_u_xfr_ctl_xfr_caddr_2__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_xfr_caddr_2_) );
  DFFPOSX1 DFFPOSX1_504 ( .CLK(sdram_clk_bF_buf63), .D(u_sdrc_core_u_xfr_ctl_xfr_caddr_3__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_xfr_caddr_3_) );
  DFFPOSX1 DFFPOSX1_505 ( .CLK(sdram_clk_bF_buf62), .D(u_sdrc_core_u_xfr_ctl_xfr_caddr_4__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_xfr_caddr_4_) );
  DFFPOSX1 DFFPOSX1_506 ( .CLK(sdram_clk_bF_buf61), .D(u_sdrc_core_u_xfr_ctl_xfr_caddr_5__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_xfr_caddr_5_) );
  DFFPOSX1 DFFPOSX1_507 ( .CLK(sdram_clk_bF_buf60), .D(u_sdrc_core_u_xfr_ctl_xfr_caddr_6__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_xfr_caddr_6_) );
  DFFPOSX1 DFFPOSX1_508 ( .CLK(sdram_clk_bF_buf59), .D(u_sdrc_core_u_xfr_ctl_xfr_caddr_7__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_xfr_caddr_7_) );
  DFFPOSX1 DFFPOSX1_509 ( .CLK(sdram_clk_bF_buf58), .D(u_sdrc_core_u_xfr_ctl_xfr_caddr_8__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_xfr_caddr_8_) );
  DFFPOSX1 DFFPOSX1_51 ( .CLK(sdram_clk_bF_buf30), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_0__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_0_) );
  DFFPOSX1 DFFPOSX1_510 ( .CLK(sdram_clk_bF_buf57), .D(u_sdrc_core_u_xfr_ctl_xfr_caddr_9__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_xfr_caddr_9_) );
  DFFPOSX1 DFFPOSX1_511 ( .CLK(sdram_clk_bF_buf56), .D(u_sdrc_core_u_xfr_ctl_xfr_caddr_10__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_xfr_caddr_10_) );
  DFFPOSX1 DFFPOSX1_512 ( .CLK(sdram_clk_bF_buf55), .D(u_sdrc_core_u_xfr_ctl_xfr_caddr_11__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_xfr_caddr_11_) );
  DFFPOSX1 DFFPOSX1_513 ( .CLK(sdram_clk_bF_buf54), .D(u_sdrc_core_u_xfr_ctl_xfr_caddr_12__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_xfr_caddr_12_) );
  DFFPOSX1 DFFPOSX1_514 ( .CLK(sdram_clk_bF_buf53), .D(u_sdrc_core_u_xfr_ctl_l_last_FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_l_last) );
  DFFPOSX1 DFFPOSX1_515 ( .CLK(sdram_clk_bF_buf52), .D(u_sdrc_core_u_xfr_ctl_l_wrap_FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_l_wrap) );
  DFFPOSX1 DFFPOSX1_516 ( .CLK(sdram_clk_bF_buf51), .D(u_sdrc_core_u_xfr_ctl_l_ba_0__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_xfr_bank_sel_0_) );
  DFFPOSX1 DFFPOSX1_517 ( .CLK(sdram_clk_bF_buf50), .D(u_sdrc_core_u_xfr_ctl_l_ba_1__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_xfr_bank_sel_1_) );
  DFFPOSX1 DFFPOSX1_518 ( .CLK(sdram_clk_bF_buf49), .D(u_sdrc_core_u_xfr_ctl_l_len_0__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_l_len_0_) );
  DFFPOSX1 DFFPOSX1_519 ( .CLK(sdram_clk_bF_buf48), .D(u_sdrc_core_u_xfr_ctl_l_len_1__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_l_len_1_) );
  DFFPOSX1 DFFPOSX1_52 ( .CLK(sdram_clk_bF_buf29), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_1__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_1_) );
  DFFPOSX1 DFFPOSX1_520 ( .CLK(sdram_clk_bF_buf47), .D(u_sdrc_core_u_xfr_ctl_l_len_2__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_l_len_2_) );
  DFFPOSX1 DFFPOSX1_521 ( .CLK(sdram_clk_bF_buf46), .D(u_sdrc_core_u_xfr_ctl_l_len_3__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_l_len_3_) );
  DFFPOSX1 DFFPOSX1_522 ( .CLK(sdram_clk_bF_buf45), .D(u_sdrc_core_u_xfr_ctl_l_len_4__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_l_len_4_) );
  DFFPOSX1 DFFPOSX1_523 ( .CLK(sdram_clk_bF_buf44), .D(u_sdrc_core_u_xfr_ctl_l_len_5__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_l_len_5_) );
  DFFPOSX1 DFFPOSX1_524 ( .CLK(sdram_clk_bF_buf43), .D(u_sdrc_core_u_xfr_ctl_l_len_6__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_l_len_6_) );
  DFFPOSX1 DFFPOSX1_525 ( .CLK(sdram_clk_bF_buf42), .D(u_sdrc_core_u_xfr_ctl_act_cmd_FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_act_cmd) );
  DFFPOSX1 DFFPOSX1_526 ( .CLK(sdram_clk_bF_buf41), .D(u_sdrc_core_u_xfr_ctl_d_act_cmd_FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_d_act_cmd) );
  DFFPOSX1 DFFPOSX1_527 ( .CLK(sdram_clk_bF_buf40), .D(u_sdrc_core_u_xfr_ctl_l_rd_next_0__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_l_rd_next_0_) );
  DFFPOSX1 DFFPOSX1_528 ( .CLK(sdram_clk_bF_buf39), .D(u_sdrc_core_u_xfr_ctl_l_rd_next_1__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_l_rd_next_1_) );
  DFFPOSX1 DFFPOSX1_529 ( .CLK(sdram_clk_bF_buf38), .D(u_sdrc_core_u_xfr_ctl_l_rd_next_2__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_l_rd_next_2_) );
  DFFPOSX1 DFFPOSX1_53 ( .CLK(sdram_clk_bF_buf28), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_2__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_2_) );
  DFFPOSX1 DFFPOSX1_530 ( .CLK(sdram_clk_bF_buf37), .D(u_sdrc_core_u_xfr_ctl_l_rd_next_3__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_l_rd_next_3_) );
  DFFPOSX1 DFFPOSX1_531 ( .CLK(sdram_clk_bF_buf36), .D(u_sdrc_core_u_xfr_ctl_l_rd_next_4__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_l_rd_next_4_) );
  DFFPOSX1 DFFPOSX1_532 ( .CLK(sdram_clk_bF_buf35), .D(u_sdrc_core_u_xfr_ctl_l_rd_next_5__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_l_rd_next_5_) );
  DFFPOSX1 DFFPOSX1_533 ( .CLK(sdram_clk_bF_buf34), .D(u_sdrc_core_u_xfr_ctl_l_rd_next_6__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_l_rd_next_6_) );
  DFFPOSX1 DFFPOSX1_534 ( .CLK(sdram_clk_bF_buf33), .D(u_sdrc_core_u_xfr_ctl_l_rd_last_0__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_l_rd_last_0_) );
  DFFPOSX1 DFFPOSX1_535 ( .CLK(sdram_clk_bF_buf32), .D(u_sdrc_core_u_xfr_ctl_l_rd_last_1__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_l_rd_last_1_) );
  DFFPOSX1 DFFPOSX1_536 ( .CLK(sdram_clk_bF_buf31), .D(u_sdrc_core_u_xfr_ctl_l_rd_last_2__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_l_rd_last_2_) );
  DFFPOSX1 DFFPOSX1_537 ( .CLK(sdram_clk_bF_buf30), .D(u_sdrc_core_u_xfr_ctl_l_rd_last_3__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_l_rd_last_3_) );
  DFFPOSX1 DFFPOSX1_538 ( .CLK(sdram_clk_bF_buf29), .D(u_sdrc_core_u_xfr_ctl_l_rd_last_4__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_l_rd_last_4_) );
  DFFPOSX1 DFFPOSX1_539 ( .CLK(sdram_clk_bF_buf28), .D(u_sdrc_core_u_xfr_ctl_l_rd_last_5__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_l_rd_last_5_) );
  DFFPOSX1 DFFPOSX1_54 ( .CLK(sdram_clk_bF_buf27), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_3__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_3_) );
  DFFPOSX1 DFFPOSX1_540 ( .CLK(sdram_clk_bF_buf27), .D(u_sdrc_core_u_xfr_ctl_l_rd_last_6__FF_INPUT), .Q(u_sdrc_core_u_xfr_ctl_l_rd_last_6_) );
  DFFPOSX1 DFFPOSX1_541 ( .CLK(wb_clk_i_bF_buf58), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n422), .Q(u_wb2sdrc_u_cmdfifo_mem_3__0_) );
  DFFPOSX1 DFFPOSX1_542 ( .CLK(wb_clk_i_bF_buf57), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n424), .Q(u_wb2sdrc_u_cmdfifo_mem_3__1_) );
  DFFPOSX1 DFFPOSX1_543 ( .CLK(wb_clk_i_bF_buf56), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n426), .Q(u_wb2sdrc_u_cmdfifo_mem_3__2_) );
  DFFPOSX1 DFFPOSX1_544 ( .CLK(wb_clk_i_bF_buf55), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n428), .Q(u_wb2sdrc_u_cmdfifo_mem_3__3_) );
  DFFPOSX1 DFFPOSX1_545 ( .CLK(wb_clk_i_bF_buf54), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n430), .Q(u_wb2sdrc_u_cmdfifo_mem_3__4_) );
  DFFPOSX1 DFFPOSX1_546 ( .CLK(wb_clk_i_bF_buf53), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n432), .Q(u_wb2sdrc_u_cmdfifo_mem_3__5_) );
  DFFPOSX1 DFFPOSX1_547 ( .CLK(wb_clk_i_bF_buf52), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n434), .Q(u_wb2sdrc_u_cmdfifo_mem_3__6_) );
  DFFPOSX1 DFFPOSX1_548 ( .CLK(wb_clk_i_bF_buf51), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n436), .Q(u_wb2sdrc_u_cmdfifo_mem_3__7_) );
  DFFPOSX1 DFFPOSX1_549 ( .CLK(wb_clk_i_bF_buf50), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n438), .Q(u_wb2sdrc_u_cmdfifo_mem_3__8_) );
  DFFPOSX1 DFFPOSX1_55 ( .CLK(sdram_clk_bF_buf26), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_4__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_4_) );
  DFFPOSX1 DFFPOSX1_550 ( .CLK(wb_clk_i_bF_buf49), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n440), .Q(u_wb2sdrc_u_cmdfifo_mem_3__9_) );
  DFFPOSX1 DFFPOSX1_551 ( .CLK(wb_clk_i_bF_buf48), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n442), .Q(u_wb2sdrc_u_cmdfifo_mem_3__10_) );
  DFFPOSX1 DFFPOSX1_552 ( .CLK(wb_clk_i_bF_buf47), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n444), .Q(u_wb2sdrc_u_cmdfifo_mem_3__11_) );
  DFFPOSX1 DFFPOSX1_553 ( .CLK(wb_clk_i_bF_buf46), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n446), .Q(u_wb2sdrc_u_cmdfifo_mem_3__12_) );
  DFFPOSX1 DFFPOSX1_554 ( .CLK(wb_clk_i_bF_buf45), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n448), .Q(u_wb2sdrc_u_cmdfifo_mem_3__13_) );
  DFFPOSX1 DFFPOSX1_555 ( .CLK(wb_clk_i_bF_buf44), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n450), .Q(u_wb2sdrc_u_cmdfifo_mem_3__14_) );
  DFFPOSX1 DFFPOSX1_556 ( .CLK(wb_clk_i_bF_buf43), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n452), .Q(u_wb2sdrc_u_cmdfifo_mem_3__15_) );
  DFFPOSX1 DFFPOSX1_557 ( .CLK(wb_clk_i_bF_buf42), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n454), .Q(u_wb2sdrc_u_cmdfifo_mem_3__16_) );
  DFFPOSX1 DFFPOSX1_558 ( .CLK(wb_clk_i_bF_buf41), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n456), .Q(u_wb2sdrc_u_cmdfifo_mem_3__17_) );
  DFFPOSX1 DFFPOSX1_559 ( .CLK(wb_clk_i_bF_buf40), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n458), .Q(u_wb2sdrc_u_cmdfifo_mem_3__18_) );
  DFFPOSX1 DFFPOSX1_56 ( .CLK(sdram_clk_bF_buf25), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_5__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_5_) );
  DFFPOSX1 DFFPOSX1_560 ( .CLK(wb_clk_i_bF_buf39), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n460), .Q(u_wb2sdrc_u_cmdfifo_mem_3__19_) );
  DFFPOSX1 DFFPOSX1_561 ( .CLK(wb_clk_i_bF_buf38), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n462), .Q(u_wb2sdrc_u_cmdfifo_mem_3__20_) );
  DFFPOSX1 DFFPOSX1_562 ( .CLK(wb_clk_i_bF_buf37), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n464), .Q(u_wb2sdrc_u_cmdfifo_mem_3__21_) );
  DFFPOSX1 DFFPOSX1_563 ( .CLK(wb_clk_i_bF_buf36), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n466), .Q(u_wb2sdrc_u_cmdfifo_mem_3__22_) );
  DFFPOSX1 DFFPOSX1_564 ( .CLK(wb_clk_i_bF_buf35), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n468), .Q(u_wb2sdrc_u_cmdfifo_mem_3__23_) );
  DFFPOSX1 DFFPOSX1_565 ( .CLK(wb_clk_i_bF_buf34), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n470), .Q(u_wb2sdrc_u_cmdfifo_mem_3__24_) );
  DFFPOSX1 DFFPOSX1_566 ( .CLK(wb_clk_i_bF_buf33), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n472), .Q(u_wb2sdrc_u_cmdfifo_mem_3__25_) );
  DFFPOSX1 DFFPOSX1_567 ( .CLK(wb_clk_i_bF_buf32), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n474), .Q(u_wb2sdrc_u_cmdfifo_mem_3__26_) );
  DFFPOSX1 DFFPOSX1_568 ( .CLK(wb_clk_i_bF_buf31), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n476), .Q(u_wb2sdrc_u_cmdfifo_mem_3__27_) );
  DFFPOSX1 DFFPOSX1_569 ( .CLK(wb_clk_i_bF_buf30), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n478), .Q(u_wb2sdrc_u_cmdfifo_mem_3__28_) );
  DFFPOSX1 DFFPOSX1_57 ( .CLK(sdram_clk_bF_buf24), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_6__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_6_) );
  DFFPOSX1 DFFPOSX1_570 ( .CLK(wb_clk_i_bF_buf29), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n480), .Q(u_wb2sdrc_u_cmdfifo_mem_3__29_) );
  DFFPOSX1 DFFPOSX1_571 ( .CLK(wb_clk_i_bF_buf28), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n482), .Q(u_wb2sdrc_u_cmdfifo_mem_3__30_) );
  DFFPOSX1 DFFPOSX1_572 ( .CLK(wb_clk_i_bF_buf27), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n484), .Q(u_wb2sdrc_u_cmdfifo_mem_3__31_) );
  DFFPOSX1 DFFPOSX1_573 ( .CLK(wb_clk_i_bF_buf26), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n486), .Q(u_wb2sdrc_u_cmdfifo_mem_3__32_) );
  DFFPOSX1 DFFPOSX1_574 ( .CLK(wb_clk_i_bF_buf25), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n488), .Q(u_wb2sdrc_u_cmdfifo_mem_3__33_) );
  DFFPOSX1 DFFPOSX1_575 ( .CLK(wb_clk_i_bF_buf24), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n490), .Q(u_wb2sdrc_u_cmdfifo_mem_3__34_) );
  DFFPOSX1 DFFPOSX1_576 ( .CLK(wb_clk_i_bF_buf23), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n492), .Q(u_wb2sdrc_u_cmdfifo_mem_3__35_) );
  DFFPOSX1 DFFPOSX1_577 ( .CLK(wb_clk_i_bF_buf22), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n532), .Q(u_wb2sdrc_u_cmdfifo_mem_2__0_) );
  DFFPOSX1 DFFPOSX1_578 ( .CLK(wb_clk_i_bF_buf21), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n534), .Q(u_wb2sdrc_u_cmdfifo_mem_2__1_) );
  DFFPOSX1 DFFPOSX1_579 ( .CLK(wb_clk_i_bF_buf20), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n536), .Q(u_wb2sdrc_u_cmdfifo_mem_2__2_) );
  DFFPOSX1 DFFPOSX1_58 ( .CLK(sdram_clk_bF_buf23), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_0__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_0_) );
  DFFPOSX1 DFFPOSX1_580 ( .CLK(wb_clk_i_bF_buf19), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n538), .Q(u_wb2sdrc_u_cmdfifo_mem_2__3_) );
  DFFPOSX1 DFFPOSX1_581 ( .CLK(wb_clk_i_bF_buf18), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n540), .Q(u_wb2sdrc_u_cmdfifo_mem_2__4_) );
  DFFPOSX1 DFFPOSX1_582 ( .CLK(wb_clk_i_bF_buf17), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n542), .Q(u_wb2sdrc_u_cmdfifo_mem_2__5_) );
  DFFPOSX1 DFFPOSX1_583 ( .CLK(wb_clk_i_bF_buf16), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n544), .Q(u_wb2sdrc_u_cmdfifo_mem_2__6_) );
  DFFPOSX1 DFFPOSX1_584 ( .CLK(wb_clk_i_bF_buf15), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n546), .Q(u_wb2sdrc_u_cmdfifo_mem_2__7_) );
  DFFPOSX1 DFFPOSX1_585 ( .CLK(wb_clk_i_bF_buf14), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n548), .Q(u_wb2sdrc_u_cmdfifo_mem_2__8_) );
  DFFPOSX1 DFFPOSX1_586 ( .CLK(wb_clk_i_bF_buf13), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n550), .Q(u_wb2sdrc_u_cmdfifo_mem_2__9_) );
  DFFPOSX1 DFFPOSX1_587 ( .CLK(wb_clk_i_bF_buf12), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n552), .Q(u_wb2sdrc_u_cmdfifo_mem_2__10_) );
  DFFPOSX1 DFFPOSX1_588 ( .CLK(wb_clk_i_bF_buf11), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n554), .Q(u_wb2sdrc_u_cmdfifo_mem_2__11_) );
  DFFPOSX1 DFFPOSX1_589 ( .CLK(wb_clk_i_bF_buf10), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n556), .Q(u_wb2sdrc_u_cmdfifo_mem_2__12_) );
  DFFPOSX1 DFFPOSX1_59 ( .CLK(sdram_clk_bF_buf22), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_1__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_1_) );
  DFFPOSX1 DFFPOSX1_590 ( .CLK(wb_clk_i_bF_buf9), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n558), .Q(u_wb2sdrc_u_cmdfifo_mem_2__13_) );
  DFFPOSX1 DFFPOSX1_591 ( .CLK(wb_clk_i_bF_buf8), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n560), .Q(u_wb2sdrc_u_cmdfifo_mem_2__14_) );
  DFFPOSX1 DFFPOSX1_592 ( .CLK(wb_clk_i_bF_buf7), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n562), .Q(u_wb2sdrc_u_cmdfifo_mem_2__15_) );
  DFFPOSX1 DFFPOSX1_593 ( .CLK(wb_clk_i_bF_buf6), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n564), .Q(u_wb2sdrc_u_cmdfifo_mem_2__16_) );
  DFFPOSX1 DFFPOSX1_594 ( .CLK(wb_clk_i_bF_buf5), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n566), .Q(u_wb2sdrc_u_cmdfifo_mem_2__17_) );
  DFFPOSX1 DFFPOSX1_595 ( .CLK(wb_clk_i_bF_buf4), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n568), .Q(u_wb2sdrc_u_cmdfifo_mem_2__18_) );
  DFFPOSX1 DFFPOSX1_596 ( .CLK(wb_clk_i_bF_buf3), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n570), .Q(u_wb2sdrc_u_cmdfifo_mem_2__19_) );
  DFFPOSX1 DFFPOSX1_597 ( .CLK(wb_clk_i_bF_buf2), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n572), .Q(u_wb2sdrc_u_cmdfifo_mem_2__20_) );
  DFFPOSX1 DFFPOSX1_598 ( .CLK(wb_clk_i_bF_buf1), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n574), .Q(u_wb2sdrc_u_cmdfifo_mem_2__21_) );
  DFFPOSX1 DFFPOSX1_599 ( .CLK(wb_clk_i_bF_buf0), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n576), .Q(u_wb2sdrc_u_cmdfifo_mem_2__22_) );
  DFFPOSX1 DFFPOSX1_6 ( .CLK(sdram_clk_bF_buf75), .D(u_sdrc_core_pad_sdr_din1_5_), .Q(u_sdrc_core_pad_sdr_din2_5_) );
  DFFPOSX1 DFFPOSX1_60 ( .CLK(sdram_clk_bF_buf21), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_2__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_2_) );
  DFFPOSX1 DFFPOSX1_600 ( .CLK(wb_clk_i_bF_buf59), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n578), .Q(u_wb2sdrc_u_cmdfifo_mem_2__23_) );
  DFFPOSX1 DFFPOSX1_601 ( .CLK(wb_clk_i_bF_buf58), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n580), .Q(u_wb2sdrc_u_cmdfifo_mem_2__24_) );
  DFFPOSX1 DFFPOSX1_602 ( .CLK(wb_clk_i_bF_buf57), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n582), .Q(u_wb2sdrc_u_cmdfifo_mem_2__25_) );
  DFFPOSX1 DFFPOSX1_603 ( .CLK(wb_clk_i_bF_buf56), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n584), .Q(u_wb2sdrc_u_cmdfifo_mem_2__26_) );
  DFFPOSX1 DFFPOSX1_604 ( .CLK(wb_clk_i_bF_buf55), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n586), .Q(u_wb2sdrc_u_cmdfifo_mem_2__27_) );
  DFFPOSX1 DFFPOSX1_605 ( .CLK(wb_clk_i_bF_buf54), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n588), .Q(u_wb2sdrc_u_cmdfifo_mem_2__28_) );
  DFFPOSX1 DFFPOSX1_606 ( .CLK(wb_clk_i_bF_buf53), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n590), .Q(u_wb2sdrc_u_cmdfifo_mem_2__29_) );
  DFFPOSX1 DFFPOSX1_607 ( .CLK(wb_clk_i_bF_buf52), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n592), .Q(u_wb2sdrc_u_cmdfifo_mem_2__30_) );
  DFFPOSX1 DFFPOSX1_608 ( .CLK(wb_clk_i_bF_buf51), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n594), .Q(u_wb2sdrc_u_cmdfifo_mem_2__31_) );
  DFFPOSX1 DFFPOSX1_609 ( .CLK(wb_clk_i_bF_buf50), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n596), .Q(u_wb2sdrc_u_cmdfifo_mem_2__32_) );
  DFFPOSX1 DFFPOSX1_61 ( .CLK(sdram_clk_bF_buf20), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_3__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_3_) );
  DFFPOSX1 DFFPOSX1_610 ( .CLK(wb_clk_i_bF_buf49), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n598), .Q(u_wb2sdrc_u_cmdfifo_mem_2__33_) );
  DFFPOSX1 DFFPOSX1_611 ( .CLK(wb_clk_i_bF_buf48), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n600), .Q(u_wb2sdrc_u_cmdfifo_mem_2__34_) );
  DFFPOSX1 DFFPOSX1_612 ( .CLK(wb_clk_i_bF_buf47), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n602), .Q(u_wb2sdrc_u_cmdfifo_mem_2__35_) );
  DFFPOSX1 DFFPOSX1_613 ( .CLK(wb_clk_i_bF_buf46), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n99), .Q(u_wb2sdrc_u_cmdfifo_mem_0__0_) );
  DFFPOSX1 DFFPOSX1_614 ( .CLK(wb_clk_i_bF_buf45), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n102), .Q(u_wb2sdrc_u_cmdfifo_mem_0__1_) );
  DFFPOSX1 DFFPOSX1_615 ( .CLK(wb_clk_i_bF_buf44), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n105), .Q(u_wb2sdrc_u_cmdfifo_mem_0__2_) );
  DFFPOSX1 DFFPOSX1_616 ( .CLK(wb_clk_i_bF_buf43), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n108), .Q(u_wb2sdrc_u_cmdfifo_mem_0__3_) );
  DFFPOSX1 DFFPOSX1_617 ( .CLK(wb_clk_i_bF_buf42), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n111), .Q(u_wb2sdrc_u_cmdfifo_mem_0__4_) );
  DFFPOSX1 DFFPOSX1_618 ( .CLK(wb_clk_i_bF_buf41), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n114), .Q(u_wb2sdrc_u_cmdfifo_mem_0__5_) );
  DFFPOSX1 DFFPOSX1_619 ( .CLK(wb_clk_i_bF_buf40), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n117), .Q(u_wb2sdrc_u_cmdfifo_mem_0__6_) );
  DFFPOSX1 DFFPOSX1_62 ( .CLK(sdram_clk_bF_buf19), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_4__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_4_) );
  DFFPOSX1 DFFPOSX1_620 ( .CLK(wb_clk_i_bF_buf39), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n120), .Q(u_wb2sdrc_u_cmdfifo_mem_0__7_) );
  DFFPOSX1 DFFPOSX1_621 ( .CLK(wb_clk_i_bF_buf38), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n123), .Q(u_wb2sdrc_u_cmdfifo_mem_0__8_) );
  DFFPOSX1 DFFPOSX1_622 ( .CLK(wb_clk_i_bF_buf37), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n126), .Q(u_wb2sdrc_u_cmdfifo_mem_0__9_) );
  DFFPOSX1 DFFPOSX1_623 ( .CLK(wb_clk_i_bF_buf36), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n129), .Q(u_wb2sdrc_u_cmdfifo_mem_0__10_) );
  DFFPOSX1 DFFPOSX1_624 ( .CLK(wb_clk_i_bF_buf35), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n132), .Q(u_wb2sdrc_u_cmdfifo_mem_0__11_) );
  DFFPOSX1 DFFPOSX1_625 ( .CLK(wb_clk_i_bF_buf34), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n135), .Q(u_wb2sdrc_u_cmdfifo_mem_0__12_) );
  DFFPOSX1 DFFPOSX1_626 ( .CLK(wb_clk_i_bF_buf33), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n138), .Q(u_wb2sdrc_u_cmdfifo_mem_0__13_) );
  DFFPOSX1 DFFPOSX1_627 ( .CLK(wb_clk_i_bF_buf32), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n141), .Q(u_wb2sdrc_u_cmdfifo_mem_0__14_) );
  DFFPOSX1 DFFPOSX1_628 ( .CLK(wb_clk_i_bF_buf31), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n144), .Q(u_wb2sdrc_u_cmdfifo_mem_0__15_) );
  DFFPOSX1 DFFPOSX1_629 ( .CLK(wb_clk_i_bF_buf30), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n147), .Q(u_wb2sdrc_u_cmdfifo_mem_0__16_) );
  DFFPOSX1 DFFPOSX1_63 ( .CLK(sdram_clk_bF_buf18), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_5__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_5_) );
  DFFPOSX1 DFFPOSX1_630 ( .CLK(wb_clk_i_bF_buf29), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n150), .Q(u_wb2sdrc_u_cmdfifo_mem_0__17_) );
  DFFPOSX1 DFFPOSX1_631 ( .CLK(wb_clk_i_bF_buf28), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n153), .Q(u_wb2sdrc_u_cmdfifo_mem_0__18_) );
  DFFPOSX1 DFFPOSX1_632 ( .CLK(wb_clk_i_bF_buf27), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n156), .Q(u_wb2sdrc_u_cmdfifo_mem_0__19_) );
  DFFPOSX1 DFFPOSX1_633 ( .CLK(wb_clk_i_bF_buf26), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n159), .Q(u_wb2sdrc_u_cmdfifo_mem_0__20_) );
  DFFPOSX1 DFFPOSX1_634 ( .CLK(wb_clk_i_bF_buf25), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n162), .Q(u_wb2sdrc_u_cmdfifo_mem_0__21_) );
  DFFPOSX1 DFFPOSX1_635 ( .CLK(wb_clk_i_bF_buf24), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n165), .Q(u_wb2sdrc_u_cmdfifo_mem_0__22_) );
  DFFPOSX1 DFFPOSX1_636 ( .CLK(wb_clk_i_bF_buf23), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n168), .Q(u_wb2sdrc_u_cmdfifo_mem_0__23_) );
  DFFPOSX1 DFFPOSX1_637 ( .CLK(wb_clk_i_bF_buf22), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n171), .Q(u_wb2sdrc_u_cmdfifo_mem_0__24_) );
  DFFPOSX1 DFFPOSX1_638 ( .CLK(wb_clk_i_bF_buf21), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n174), .Q(u_wb2sdrc_u_cmdfifo_mem_0__25_) );
  DFFPOSX1 DFFPOSX1_639 ( .CLK(wb_clk_i_bF_buf20), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n177), .Q(u_wb2sdrc_u_cmdfifo_mem_0__26_) );
  DFFPOSX1 DFFPOSX1_64 ( .CLK(sdram_clk_bF_buf17), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_6__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_6_) );
  DFFPOSX1 DFFPOSX1_640 ( .CLK(wb_clk_i_bF_buf19), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n180), .Q(u_wb2sdrc_u_cmdfifo_mem_0__27_) );
  DFFPOSX1 DFFPOSX1_641 ( .CLK(wb_clk_i_bF_buf18), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n183), .Q(u_wb2sdrc_u_cmdfifo_mem_0__28_) );
  DFFPOSX1 DFFPOSX1_642 ( .CLK(wb_clk_i_bF_buf17), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n186), .Q(u_wb2sdrc_u_cmdfifo_mem_0__29_) );
  DFFPOSX1 DFFPOSX1_643 ( .CLK(wb_clk_i_bF_buf16), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n189), .Q(u_wb2sdrc_u_cmdfifo_mem_0__30_) );
  DFFPOSX1 DFFPOSX1_644 ( .CLK(wb_clk_i_bF_buf15), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n192), .Q(u_wb2sdrc_u_cmdfifo_mem_0__31_) );
  DFFPOSX1 DFFPOSX1_645 ( .CLK(wb_clk_i_bF_buf14), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n195), .Q(u_wb2sdrc_u_cmdfifo_mem_0__32_) );
  DFFPOSX1 DFFPOSX1_646 ( .CLK(wb_clk_i_bF_buf13), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n198), .Q(u_wb2sdrc_u_cmdfifo_mem_0__33_) );
  DFFPOSX1 DFFPOSX1_647 ( .CLK(wb_clk_i_bF_buf12), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n201), .Q(u_wb2sdrc_u_cmdfifo_mem_0__34_) );
  DFFPOSX1 DFFPOSX1_648 ( .CLK(wb_clk_i_bF_buf11), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n204), .Q(u_wb2sdrc_u_cmdfifo_mem_0__35_) );
  DFFPOSX1 DFFPOSX1_649 ( .CLK(wb_clk_i_bF_buf10), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n494), .Q(u_wb2sdrc_u_cmdfifo_mem_1__0_) );
  DFFPOSX1 DFFPOSX1_65 ( .CLK(sdram_clk_bF_buf16), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_7__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_7_) );
  DFFPOSX1 DFFPOSX1_650 ( .CLK(wb_clk_i_bF_buf9), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n495), .Q(u_wb2sdrc_u_cmdfifo_mem_1__1_) );
  DFFPOSX1 DFFPOSX1_651 ( .CLK(wb_clk_i_bF_buf8), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n496), .Q(u_wb2sdrc_u_cmdfifo_mem_1__2_) );
  DFFPOSX1 DFFPOSX1_652 ( .CLK(wb_clk_i_bF_buf7), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n497), .Q(u_wb2sdrc_u_cmdfifo_mem_1__3_) );
  DFFPOSX1 DFFPOSX1_653 ( .CLK(wb_clk_i_bF_buf6), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n498), .Q(u_wb2sdrc_u_cmdfifo_mem_1__4_) );
  DFFPOSX1 DFFPOSX1_654 ( .CLK(wb_clk_i_bF_buf5), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n499), .Q(u_wb2sdrc_u_cmdfifo_mem_1__5_) );
  DFFPOSX1 DFFPOSX1_655 ( .CLK(wb_clk_i_bF_buf4), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n500), .Q(u_wb2sdrc_u_cmdfifo_mem_1__6_) );
  DFFPOSX1 DFFPOSX1_656 ( .CLK(wb_clk_i_bF_buf3), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n501), .Q(u_wb2sdrc_u_cmdfifo_mem_1__7_) );
  DFFPOSX1 DFFPOSX1_657 ( .CLK(wb_clk_i_bF_buf2), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n502), .Q(u_wb2sdrc_u_cmdfifo_mem_1__8_) );
  DFFPOSX1 DFFPOSX1_658 ( .CLK(wb_clk_i_bF_buf1), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n503), .Q(u_wb2sdrc_u_cmdfifo_mem_1__9_) );
  DFFPOSX1 DFFPOSX1_659 ( .CLK(wb_clk_i_bF_buf0), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n504), .Q(u_wb2sdrc_u_cmdfifo_mem_1__10_) );
  DFFPOSX1 DFFPOSX1_66 ( .CLK(sdram_clk_bF_buf15), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_8__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_8_) );
  DFFPOSX1 DFFPOSX1_660 ( .CLK(wb_clk_i_bF_buf59), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n505), .Q(u_wb2sdrc_u_cmdfifo_mem_1__11_) );
  DFFPOSX1 DFFPOSX1_661 ( .CLK(wb_clk_i_bF_buf58), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n506), .Q(u_wb2sdrc_u_cmdfifo_mem_1__12_) );
  DFFPOSX1 DFFPOSX1_662 ( .CLK(wb_clk_i_bF_buf57), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n507), .Q(u_wb2sdrc_u_cmdfifo_mem_1__13_) );
  DFFPOSX1 DFFPOSX1_663 ( .CLK(wb_clk_i_bF_buf56), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n508), .Q(u_wb2sdrc_u_cmdfifo_mem_1__14_) );
  DFFPOSX1 DFFPOSX1_664 ( .CLK(wb_clk_i_bF_buf55), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n509), .Q(u_wb2sdrc_u_cmdfifo_mem_1__15_) );
  DFFPOSX1 DFFPOSX1_665 ( .CLK(wb_clk_i_bF_buf54), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n510), .Q(u_wb2sdrc_u_cmdfifo_mem_1__16_) );
  DFFPOSX1 DFFPOSX1_666 ( .CLK(wb_clk_i_bF_buf53), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n511), .Q(u_wb2sdrc_u_cmdfifo_mem_1__17_) );
  DFFPOSX1 DFFPOSX1_667 ( .CLK(wb_clk_i_bF_buf52), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n512), .Q(u_wb2sdrc_u_cmdfifo_mem_1__18_) );
  DFFPOSX1 DFFPOSX1_668 ( .CLK(wb_clk_i_bF_buf51), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n513), .Q(u_wb2sdrc_u_cmdfifo_mem_1__19_) );
  DFFPOSX1 DFFPOSX1_669 ( .CLK(wb_clk_i_bF_buf50), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n514), .Q(u_wb2sdrc_u_cmdfifo_mem_1__20_) );
  DFFPOSX1 DFFPOSX1_67 ( .CLK(sdram_clk_bF_buf14), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_9__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_9_) );
  DFFPOSX1 DFFPOSX1_670 ( .CLK(wb_clk_i_bF_buf49), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n515), .Q(u_wb2sdrc_u_cmdfifo_mem_1__21_) );
  DFFPOSX1 DFFPOSX1_671 ( .CLK(wb_clk_i_bF_buf48), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n516), .Q(u_wb2sdrc_u_cmdfifo_mem_1__22_) );
  DFFPOSX1 DFFPOSX1_672 ( .CLK(wb_clk_i_bF_buf47), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n517), .Q(u_wb2sdrc_u_cmdfifo_mem_1__23_) );
  DFFPOSX1 DFFPOSX1_673 ( .CLK(wb_clk_i_bF_buf46), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n518), .Q(u_wb2sdrc_u_cmdfifo_mem_1__24_) );
  DFFPOSX1 DFFPOSX1_674 ( .CLK(wb_clk_i_bF_buf45), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n519), .Q(u_wb2sdrc_u_cmdfifo_mem_1__25_) );
  DFFPOSX1 DFFPOSX1_675 ( .CLK(wb_clk_i_bF_buf44), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n520), .Q(u_wb2sdrc_u_cmdfifo_mem_1__26_) );
  DFFPOSX1 DFFPOSX1_676 ( .CLK(wb_clk_i_bF_buf43), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n521), .Q(u_wb2sdrc_u_cmdfifo_mem_1__27_) );
  DFFPOSX1 DFFPOSX1_677 ( .CLK(wb_clk_i_bF_buf42), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n522), .Q(u_wb2sdrc_u_cmdfifo_mem_1__28_) );
  DFFPOSX1 DFFPOSX1_678 ( .CLK(wb_clk_i_bF_buf41), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n523), .Q(u_wb2sdrc_u_cmdfifo_mem_1__29_) );
  DFFPOSX1 DFFPOSX1_679 ( .CLK(wb_clk_i_bF_buf40), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n524), .Q(u_wb2sdrc_u_cmdfifo_mem_1__30_) );
  DFFPOSX1 DFFPOSX1_68 ( .CLK(sdram_clk_bF_buf13), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_10__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_10_) );
  DFFPOSX1 DFFPOSX1_680 ( .CLK(wb_clk_i_bF_buf39), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n525), .Q(u_wb2sdrc_u_cmdfifo_mem_1__31_) );
  DFFPOSX1 DFFPOSX1_681 ( .CLK(wb_clk_i_bF_buf38), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n526), .Q(u_wb2sdrc_u_cmdfifo_mem_1__32_) );
  DFFPOSX1 DFFPOSX1_682 ( .CLK(wb_clk_i_bF_buf37), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n527), .Q(u_wb2sdrc_u_cmdfifo_mem_1__33_) );
  DFFPOSX1 DFFPOSX1_683 ( .CLK(wb_clk_i_bF_buf36), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n528), .Q(u_wb2sdrc_u_cmdfifo_mem_1__34_) );
  DFFPOSX1 DFFPOSX1_684 ( .CLK(wb_clk_i_bF_buf35), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n529), .Q(u_wb2sdrc_u_cmdfifo_mem_1__35_) );
  DFFPOSX1 DFFPOSX1_685 ( .CLK(sdram_clk_bF_buf26), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n349), .Q(app_req_addr_0_) );
  DFFPOSX1 DFFPOSX1_686 ( .CLK(sdram_clk_bF_buf25), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n351), .Q(app_req_addr_1_) );
  DFFPOSX1 DFFPOSX1_687 ( .CLK(sdram_clk_bF_buf24), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n353), .Q(app_req_addr_2_) );
  DFFPOSX1 DFFPOSX1_688 ( .CLK(sdram_clk_bF_buf23), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n355), .Q(app_req_addr_3_) );
  DFFPOSX1 DFFPOSX1_689 ( .CLK(sdram_clk_bF_buf22), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n357), .Q(app_req_addr_4_) );
  DFFPOSX1 DFFPOSX1_69 ( .CLK(sdram_clk_bF_buf12), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_11__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_11_) );
  DFFPOSX1 DFFPOSX1_690 ( .CLK(sdram_clk_bF_buf21), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n359), .Q(app_req_addr_5_) );
  DFFPOSX1 DFFPOSX1_691 ( .CLK(sdram_clk_bF_buf20), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n361), .Q(app_req_addr_6_) );
  DFFPOSX1 DFFPOSX1_692 ( .CLK(sdram_clk_bF_buf19), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n363), .Q(app_req_addr_7_) );
  DFFPOSX1 DFFPOSX1_693 ( .CLK(sdram_clk_bF_buf18), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n365), .Q(app_req_addr_8_) );
  DFFPOSX1 DFFPOSX1_694 ( .CLK(sdram_clk_bF_buf17), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n367), .Q(app_req_addr_9_) );
  DFFPOSX1 DFFPOSX1_695 ( .CLK(sdram_clk_bF_buf16), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n369), .Q(app_req_addr_10_) );
  DFFPOSX1 DFFPOSX1_696 ( .CLK(sdram_clk_bF_buf15), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n371), .Q(app_req_addr_11_) );
  DFFPOSX1 DFFPOSX1_697 ( .CLK(sdram_clk_bF_buf14), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n373), .Q(app_req_addr_12_) );
  DFFPOSX1 DFFPOSX1_698 ( .CLK(sdram_clk_bF_buf13), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n375), .Q(app_req_addr_13_) );
  DFFPOSX1 DFFPOSX1_699 ( .CLK(sdram_clk_bF_buf12), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n377), .Q(app_req_addr_14_) );
  DFFPOSX1 DFFPOSX1_7 ( .CLK(sdram_clk_bF_buf74), .D(u_sdrc_core_pad_sdr_din1_6_), .Q(u_sdrc_core_pad_sdr_din2_6_) );
  DFFPOSX1 DFFPOSX1_70 ( .CLK(sdram_clk_bF_buf11), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_12__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_12_) );
  DFFPOSX1 DFFPOSX1_700 ( .CLK(sdram_clk_bF_buf11), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n379), .Q(app_req_addr_15_) );
  DFFPOSX1 DFFPOSX1_701 ( .CLK(sdram_clk_bF_buf10), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n381), .Q(app_req_addr_16_) );
  DFFPOSX1 DFFPOSX1_702 ( .CLK(sdram_clk_bF_buf9), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n383), .Q(app_req_addr_17_) );
  DFFPOSX1 DFFPOSX1_703 ( .CLK(sdram_clk_bF_buf8), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n385), .Q(app_req_addr_18_) );
  DFFPOSX1 DFFPOSX1_704 ( .CLK(sdram_clk_bF_buf7), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n387), .Q(app_req_addr_19_) );
  DFFPOSX1 DFFPOSX1_705 ( .CLK(sdram_clk_bF_buf6), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n389), .Q(app_req_addr_20_) );
  DFFPOSX1 DFFPOSX1_706 ( .CLK(sdram_clk_bF_buf5), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n391), .Q(app_req_addr_21_) );
  DFFPOSX1 DFFPOSX1_707 ( .CLK(sdram_clk_bF_buf4), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n393), .Q(app_req_addr_22_) );
  DFFPOSX1 DFFPOSX1_708 ( .CLK(sdram_clk_bF_buf3), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n395), .Q(app_req_addr_23_) );
  DFFPOSX1 DFFPOSX1_709 ( .CLK(sdram_clk_bF_buf2), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n397), .Q(app_req_addr_24_) );
  DFFPOSX1 DFFPOSX1_71 ( .CLK(sdram_clk_bF_buf10), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_l_write_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_l_write) );
  DFFPOSX1 DFFPOSX1_710 ( .CLK(sdram_clk_bF_buf1), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n399), .Q(app_req_addr_25_) );
  DFFPOSX1 DFFPOSX1_711 ( .CLK(sdram_clk_bF_buf0), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n401), .Q(app_req_wr_n) );
  DFFPOSX1 DFFPOSX1_712 ( .CLK(sdram_clk_bF_buf80), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n403), .Q(app_req_len_0_) );
  DFFPOSX1 DFFPOSX1_713 ( .CLK(sdram_clk_bF_buf79), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n405), .Q(app_req_len_1_) );
  DFFPOSX1 DFFPOSX1_714 ( .CLK(sdram_clk_bF_buf78), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n407), .Q(app_req_len_2_) );
  DFFPOSX1 DFFPOSX1_715 ( .CLK(sdram_clk_bF_buf77), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n409), .Q(app_req_len_3_) );
  DFFPOSX1 DFFPOSX1_716 ( .CLK(sdram_clk_bF_buf76), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n411), .Q(app_req_len_4_) );
  DFFPOSX1 DFFPOSX1_717 ( .CLK(sdram_clk_bF_buf75), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n413), .Q(app_req_len_5_) );
  DFFPOSX1 DFFPOSX1_718 ( .CLK(sdram_clk_bF_buf74), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n415), .Q(app_req_len_6_) );
  DFFPOSX1 DFFPOSX1_719 ( .CLK(sdram_clk_bF_buf73), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n417), .Q(app_req_len_7_) );
  DFFPOSX1 DFFPOSX1_72 ( .CLK(sdram_clk_bF_buf9), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_0__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_0_) );
  DFFPOSX1 DFFPOSX1_720 ( .CLK(sdram_clk_bF_buf72), .D(u_wb2sdrc_u_cmdfifo__abc_14585_n419), .Q(app_req_len_8_) );
  DFFPOSX1 DFFPOSX1_721 ( .CLK(sdram_clk_bF_buf58), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n464), .Q(u_wb2sdrc_u_rddatafifo_mem_1__0_) );
  DFFPOSX1 DFFPOSX1_722 ( .CLK(sdram_clk_bF_buf57), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n465), .Q(u_wb2sdrc_u_rddatafifo_mem_1__1_) );
  DFFPOSX1 DFFPOSX1_723 ( .CLK(sdram_clk_bF_buf56), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n466), .Q(u_wb2sdrc_u_rddatafifo_mem_1__2_) );
  DFFPOSX1 DFFPOSX1_724 ( .CLK(sdram_clk_bF_buf55), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n467), .Q(u_wb2sdrc_u_rddatafifo_mem_1__3_) );
  DFFPOSX1 DFFPOSX1_725 ( .CLK(sdram_clk_bF_buf54), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n468), .Q(u_wb2sdrc_u_rddatafifo_mem_1__4_) );
  DFFPOSX1 DFFPOSX1_726 ( .CLK(sdram_clk_bF_buf53), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n469), .Q(u_wb2sdrc_u_rddatafifo_mem_1__5_) );
  DFFPOSX1 DFFPOSX1_727 ( .CLK(sdram_clk_bF_buf52), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n470), .Q(u_wb2sdrc_u_rddatafifo_mem_1__6_) );
  DFFPOSX1 DFFPOSX1_728 ( .CLK(sdram_clk_bF_buf51), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n471), .Q(u_wb2sdrc_u_rddatafifo_mem_1__7_) );
  DFFPOSX1 DFFPOSX1_729 ( .CLK(sdram_clk_bF_buf50), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n472), .Q(u_wb2sdrc_u_rddatafifo_mem_1__8_) );
  DFFPOSX1 DFFPOSX1_73 ( .CLK(sdram_clk_bF_buf8), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_1__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_1_) );
  DFFPOSX1 DFFPOSX1_730 ( .CLK(sdram_clk_bF_buf49), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n473), .Q(u_wb2sdrc_u_rddatafifo_mem_1__9_) );
  DFFPOSX1 DFFPOSX1_731 ( .CLK(sdram_clk_bF_buf48), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n474), .Q(u_wb2sdrc_u_rddatafifo_mem_1__10_) );
  DFFPOSX1 DFFPOSX1_732 ( .CLK(sdram_clk_bF_buf47), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n475), .Q(u_wb2sdrc_u_rddatafifo_mem_1__11_) );
  DFFPOSX1 DFFPOSX1_733 ( .CLK(sdram_clk_bF_buf46), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n476), .Q(u_wb2sdrc_u_rddatafifo_mem_1__12_) );
  DFFPOSX1 DFFPOSX1_734 ( .CLK(sdram_clk_bF_buf45), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n477), .Q(u_wb2sdrc_u_rddatafifo_mem_1__13_) );
  DFFPOSX1 DFFPOSX1_735 ( .CLK(sdram_clk_bF_buf44), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n478), .Q(u_wb2sdrc_u_rddatafifo_mem_1__14_) );
  DFFPOSX1 DFFPOSX1_736 ( .CLK(sdram_clk_bF_buf43), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n479), .Q(u_wb2sdrc_u_rddatafifo_mem_1__15_) );
  DFFPOSX1 DFFPOSX1_737 ( .CLK(sdram_clk_bF_buf42), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n480), .Q(u_wb2sdrc_u_rddatafifo_mem_1__16_) );
  DFFPOSX1 DFFPOSX1_738 ( .CLK(sdram_clk_bF_buf41), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n481), .Q(u_wb2sdrc_u_rddatafifo_mem_1__17_) );
  DFFPOSX1 DFFPOSX1_739 ( .CLK(sdram_clk_bF_buf40), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n482), .Q(u_wb2sdrc_u_rddatafifo_mem_1__18_) );
  DFFPOSX1 DFFPOSX1_74 ( .CLK(sdram_clk_bF_buf7), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_2__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_2_) );
  DFFPOSX1 DFFPOSX1_740 ( .CLK(sdram_clk_bF_buf39), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n483), .Q(u_wb2sdrc_u_rddatafifo_mem_1__19_) );
  DFFPOSX1 DFFPOSX1_741 ( .CLK(sdram_clk_bF_buf38), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n484), .Q(u_wb2sdrc_u_rddatafifo_mem_1__20_) );
  DFFPOSX1 DFFPOSX1_742 ( .CLK(sdram_clk_bF_buf37), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n485), .Q(u_wb2sdrc_u_rddatafifo_mem_1__21_) );
  DFFPOSX1 DFFPOSX1_743 ( .CLK(sdram_clk_bF_buf36), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n486), .Q(u_wb2sdrc_u_rddatafifo_mem_1__22_) );
  DFFPOSX1 DFFPOSX1_744 ( .CLK(sdram_clk_bF_buf35), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n487), .Q(u_wb2sdrc_u_rddatafifo_mem_1__23_) );
  DFFPOSX1 DFFPOSX1_745 ( .CLK(sdram_clk_bF_buf34), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n488), .Q(u_wb2sdrc_u_rddatafifo_mem_1__24_) );
  DFFPOSX1 DFFPOSX1_746 ( .CLK(sdram_clk_bF_buf33), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n489), .Q(u_wb2sdrc_u_rddatafifo_mem_1__25_) );
  DFFPOSX1 DFFPOSX1_747 ( .CLK(sdram_clk_bF_buf32), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n490), .Q(u_wb2sdrc_u_rddatafifo_mem_1__26_) );
  DFFPOSX1 DFFPOSX1_748 ( .CLK(sdram_clk_bF_buf31), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n491), .Q(u_wb2sdrc_u_rddatafifo_mem_1__27_) );
  DFFPOSX1 DFFPOSX1_749 ( .CLK(sdram_clk_bF_buf30), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n492), .Q(u_wb2sdrc_u_rddatafifo_mem_1__28_) );
  DFFPOSX1 DFFPOSX1_75 ( .CLK(sdram_clk_bF_buf6), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_3__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_3_) );
  DFFPOSX1 DFFPOSX1_750 ( .CLK(sdram_clk_bF_buf29), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n493), .Q(u_wb2sdrc_u_rddatafifo_mem_1__29_) );
  DFFPOSX1 DFFPOSX1_751 ( .CLK(sdram_clk_bF_buf28), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n494), .Q(u_wb2sdrc_u_rddatafifo_mem_1__30_) );
  DFFPOSX1 DFFPOSX1_752 ( .CLK(sdram_clk_bF_buf27), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n495), .Q(u_wb2sdrc_u_rddatafifo_mem_1__31_) );
  DFFPOSX1 DFFPOSX1_753 ( .CLK(sdram_clk_bF_buf26), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n197), .Q(u_wb2sdrc_u_rddatafifo_mem_0__0_) );
  DFFPOSX1 DFFPOSX1_754 ( .CLK(sdram_clk_bF_buf25), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n199), .Q(u_wb2sdrc_u_rddatafifo_mem_0__1_) );
  DFFPOSX1 DFFPOSX1_755 ( .CLK(sdram_clk_bF_buf24), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n201), .Q(u_wb2sdrc_u_rddatafifo_mem_0__2_) );
  DFFPOSX1 DFFPOSX1_756 ( .CLK(sdram_clk_bF_buf23), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n203), .Q(u_wb2sdrc_u_rddatafifo_mem_0__3_) );
  DFFPOSX1 DFFPOSX1_757 ( .CLK(sdram_clk_bF_buf22), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n205), .Q(u_wb2sdrc_u_rddatafifo_mem_0__4_) );
  DFFPOSX1 DFFPOSX1_758 ( .CLK(sdram_clk_bF_buf21), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n207), .Q(u_wb2sdrc_u_rddatafifo_mem_0__5_) );
  DFFPOSX1 DFFPOSX1_759 ( .CLK(sdram_clk_bF_buf20), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n209), .Q(u_wb2sdrc_u_rddatafifo_mem_0__6_) );
  DFFPOSX1 DFFPOSX1_76 ( .CLK(sdram_clk_bF_buf5), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_4__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_4_) );
  DFFPOSX1 DFFPOSX1_760 ( .CLK(sdram_clk_bF_buf19), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n211), .Q(u_wb2sdrc_u_rddatafifo_mem_0__7_) );
  DFFPOSX1 DFFPOSX1_761 ( .CLK(sdram_clk_bF_buf18), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n213), .Q(u_wb2sdrc_u_rddatafifo_mem_0__8_) );
  DFFPOSX1 DFFPOSX1_762 ( .CLK(sdram_clk_bF_buf17), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n215), .Q(u_wb2sdrc_u_rddatafifo_mem_0__9_) );
  DFFPOSX1 DFFPOSX1_763 ( .CLK(sdram_clk_bF_buf16), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n217), .Q(u_wb2sdrc_u_rddatafifo_mem_0__10_) );
  DFFPOSX1 DFFPOSX1_764 ( .CLK(sdram_clk_bF_buf15), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n219), .Q(u_wb2sdrc_u_rddatafifo_mem_0__11_) );
  DFFPOSX1 DFFPOSX1_765 ( .CLK(sdram_clk_bF_buf14), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n221), .Q(u_wb2sdrc_u_rddatafifo_mem_0__12_) );
  DFFPOSX1 DFFPOSX1_766 ( .CLK(sdram_clk_bF_buf13), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n223), .Q(u_wb2sdrc_u_rddatafifo_mem_0__13_) );
  DFFPOSX1 DFFPOSX1_767 ( .CLK(sdram_clk_bF_buf12), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n225), .Q(u_wb2sdrc_u_rddatafifo_mem_0__14_) );
  DFFPOSX1 DFFPOSX1_768 ( .CLK(sdram_clk_bF_buf11), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n227), .Q(u_wb2sdrc_u_rddatafifo_mem_0__15_) );
  DFFPOSX1 DFFPOSX1_769 ( .CLK(sdram_clk_bF_buf10), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n229), .Q(u_wb2sdrc_u_rddatafifo_mem_0__16_) );
  DFFPOSX1 DFFPOSX1_77 ( .CLK(sdram_clk_bF_buf4), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_5__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_5_) );
  DFFPOSX1 DFFPOSX1_770 ( .CLK(sdram_clk_bF_buf9), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n231), .Q(u_wb2sdrc_u_rddatafifo_mem_0__17_) );
  DFFPOSX1 DFFPOSX1_771 ( .CLK(sdram_clk_bF_buf8), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n233), .Q(u_wb2sdrc_u_rddatafifo_mem_0__18_) );
  DFFPOSX1 DFFPOSX1_772 ( .CLK(sdram_clk_bF_buf7), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n235), .Q(u_wb2sdrc_u_rddatafifo_mem_0__19_) );
  DFFPOSX1 DFFPOSX1_773 ( .CLK(sdram_clk_bF_buf6), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n237), .Q(u_wb2sdrc_u_rddatafifo_mem_0__20_) );
  DFFPOSX1 DFFPOSX1_774 ( .CLK(sdram_clk_bF_buf5), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n239), .Q(u_wb2sdrc_u_rddatafifo_mem_0__21_) );
  DFFPOSX1 DFFPOSX1_775 ( .CLK(sdram_clk_bF_buf4), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n241), .Q(u_wb2sdrc_u_rddatafifo_mem_0__22_) );
  DFFPOSX1 DFFPOSX1_776 ( .CLK(sdram_clk_bF_buf3), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n243), .Q(u_wb2sdrc_u_rddatafifo_mem_0__23_) );
  DFFPOSX1 DFFPOSX1_777 ( .CLK(sdram_clk_bF_buf2), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n245), .Q(u_wb2sdrc_u_rddatafifo_mem_0__24_) );
  DFFPOSX1 DFFPOSX1_778 ( .CLK(sdram_clk_bF_buf1), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n247), .Q(u_wb2sdrc_u_rddatafifo_mem_0__25_) );
  DFFPOSX1 DFFPOSX1_779 ( .CLK(sdram_clk_bF_buf0), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n249), .Q(u_wb2sdrc_u_rddatafifo_mem_0__26_) );
  DFFPOSX1 DFFPOSX1_78 ( .CLK(sdram_clk_bF_buf3), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_6__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_6_) );
  DFFPOSX1 DFFPOSX1_780 ( .CLK(sdram_clk_bF_buf80), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n251), .Q(u_wb2sdrc_u_rddatafifo_mem_0__27_) );
  DFFPOSX1 DFFPOSX1_781 ( .CLK(sdram_clk_bF_buf79), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n253), .Q(u_wb2sdrc_u_rddatafifo_mem_0__28_) );
  DFFPOSX1 DFFPOSX1_782 ( .CLK(sdram_clk_bF_buf78), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n255), .Q(u_wb2sdrc_u_rddatafifo_mem_0__29_) );
  DFFPOSX1 DFFPOSX1_783 ( .CLK(sdram_clk_bF_buf77), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n257), .Q(u_wb2sdrc_u_rddatafifo_mem_0__30_) );
  DFFPOSX1 DFFPOSX1_784 ( .CLK(sdram_clk_bF_buf76), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n259), .Q(u_wb2sdrc_u_rddatafifo_mem_0__31_) );
  DFFPOSX1 DFFPOSX1_785 ( .CLK(sdram_clk_bF_buf75), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n98), .Q(u_wb2sdrc_u_rddatafifo_mem_3__0_) );
  DFFPOSX1 DFFPOSX1_786 ( .CLK(sdram_clk_bF_buf74), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n101), .Q(u_wb2sdrc_u_rddatafifo_mem_3__1_) );
  DFFPOSX1 DFFPOSX1_787 ( .CLK(sdram_clk_bF_buf73), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n104), .Q(u_wb2sdrc_u_rddatafifo_mem_3__2_) );
  DFFPOSX1 DFFPOSX1_788 ( .CLK(sdram_clk_bF_buf72), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n107), .Q(u_wb2sdrc_u_rddatafifo_mem_3__3_) );
  DFFPOSX1 DFFPOSX1_789 ( .CLK(sdram_clk_bF_buf71), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n110), .Q(u_wb2sdrc_u_rddatafifo_mem_3__4_) );
  DFFPOSX1 DFFPOSX1_79 ( .CLK(sdram_clk_bF_buf2), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_7__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_7_) );
  DFFPOSX1 DFFPOSX1_790 ( .CLK(sdram_clk_bF_buf70), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n113), .Q(u_wb2sdrc_u_rddatafifo_mem_3__5_) );
  DFFPOSX1 DFFPOSX1_791 ( .CLK(sdram_clk_bF_buf69), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n116), .Q(u_wb2sdrc_u_rddatafifo_mem_3__6_) );
  DFFPOSX1 DFFPOSX1_792 ( .CLK(sdram_clk_bF_buf68), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n119), .Q(u_wb2sdrc_u_rddatafifo_mem_3__7_) );
  DFFPOSX1 DFFPOSX1_793 ( .CLK(sdram_clk_bF_buf67), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n122), .Q(u_wb2sdrc_u_rddatafifo_mem_3__8_) );
  DFFPOSX1 DFFPOSX1_794 ( .CLK(sdram_clk_bF_buf66), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n125), .Q(u_wb2sdrc_u_rddatafifo_mem_3__9_) );
  DFFPOSX1 DFFPOSX1_795 ( .CLK(sdram_clk_bF_buf65), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n128), .Q(u_wb2sdrc_u_rddatafifo_mem_3__10_) );
  DFFPOSX1 DFFPOSX1_796 ( .CLK(sdram_clk_bF_buf64), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n131), .Q(u_wb2sdrc_u_rddatafifo_mem_3__11_) );
  DFFPOSX1 DFFPOSX1_797 ( .CLK(sdram_clk_bF_buf63), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n134), .Q(u_wb2sdrc_u_rddatafifo_mem_3__12_) );
  DFFPOSX1 DFFPOSX1_798 ( .CLK(sdram_clk_bF_buf62), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n137), .Q(u_wb2sdrc_u_rddatafifo_mem_3__13_) );
  DFFPOSX1 DFFPOSX1_799 ( .CLK(sdram_clk_bF_buf61), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n140), .Q(u_wb2sdrc_u_rddatafifo_mem_3__14_) );
  DFFPOSX1 DFFPOSX1_8 ( .CLK(sdram_clk_bF_buf73), .D(u_sdrc_core_pad_sdr_din1_7_), .Q(u_sdrc_core_pad_sdr_din2_7_) );
  DFFPOSX1 DFFPOSX1_80 ( .CLK(sdram_clk_bF_buf1), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_8__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_8_) );
  DFFPOSX1 DFFPOSX1_800 ( .CLK(sdram_clk_bF_buf60), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n143), .Q(u_wb2sdrc_u_rddatafifo_mem_3__15_) );
  DFFPOSX1 DFFPOSX1_801 ( .CLK(sdram_clk_bF_buf59), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n146), .Q(u_wb2sdrc_u_rddatafifo_mem_3__16_) );
  DFFPOSX1 DFFPOSX1_802 ( .CLK(sdram_clk_bF_buf58), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n149), .Q(u_wb2sdrc_u_rddatafifo_mem_3__17_) );
  DFFPOSX1 DFFPOSX1_803 ( .CLK(sdram_clk_bF_buf57), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n152), .Q(u_wb2sdrc_u_rddatafifo_mem_3__18_) );
  DFFPOSX1 DFFPOSX1_804 ( .CLK(sdram_clk_bF_buf56), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n155), .Q(u_wb2sdrc_u_rddatafifo_mem_3__19_) );
  DFFPOSX1 DFFPOSX1_805 ( .CLK(sdram_clk_bF_buf55), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n158), .Q(u_wb2sdrc_u_rddatafifo_mem_3__20_) );
  DFFPOSX1 DFFPOSX1_806 ( .CLK(sdram_clk_bF_buf54), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n161), .Q(u_wb2sdrc_u_rddatafifo_mem_3__21_) );
  DFFPOSX1 DFFPOSX1_807 ( .CLK(sdram_clk_bF_buf53), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n164), .Q(u_wb2sdrc_u_rddatafifo_mem_3__22_) );
  DFFPOSX1 DFFPOSX1_808 ( .CLK(sdram_clk_bF_buf52), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n167), .Q(u_wb2sdrc_u_rddatafifo_mem_3__23_) );
  DFFPOSX1 DFFPOSX1_809 ( .CLK(sdram_clk_bF_buf51), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n170), .Q(u_wb2sdrc_u_rddatafifo_mem_3__24_) );
  DFFPOSX1 DFFPOSX1_81 ( .CLK(sdram_clk_bF_buf0), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_9__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_9_) );
  DFFPOSX1 DFFPOSX1_810 ( .CLK(sdram_clk_bF_buf50), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n173), .Q(u_wb2sdrc_u_rddatafifo_mem_3__25_) );
  DFFPOSX1 DFFPOSX1_811 ( .CLK(sdram_clk_bF_buf49), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n176), .Q(u_wb2sdrc_u_rddatafifo_mem_3__26_) );
  DFFPOSX1 DFFPOSX1_812 ( .CLK(sdram_clk_bF_buf48), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n179), .Q(u_wb2sdrc_u_rddatafifo_mem_3__27_) );
  DFFPOSX1 DFFPOSX1_813 ( .CLK(sdram_clk_bF_buf47), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n182), .Q(u_wb2sdrc_u_rddatafifo_mem_3__28_) );
  DFFPOSX1 DFFPOSX1_814 ( .CLK(sdram_clk_bF_buf46), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n185), .Q(u_wb2sdrc_u_rddatafifo_mem_3__29_) );
  DFFPOSX1 DFFPOSX1_815 ( .CLK(sdram_clk_bF_buf45), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n188), .Q(u_wb2sdrc_u_rddatafifo_mem_3__30_) );
  DFFPOSX1 DFFPOSX1_816 ( .CLK(sdram_clk_bF_buf44), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n191), .Q(u_wb2sdrc_u_rddatafifo_mem_3__31_) );
  DFFPOSX1 DFFPOSX1_817 ( .CLK(sdram_clk_bF_buf43), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n264), .Q(u_wb2sdrc_u_rddatafifo_mem_2__0_) );
  DFFPOSX1 DFFPOSX1_818 ( .CLK(sdram_clk_bF_buf42), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n266), .Q(u_wb2sdrc_u_rddatafifo_mem_2__1_) );
  DFFPOSX1 DFFPOSX1_819 ( .CLK(sdram_clk_bF_buf41), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n268), .Q(u_wb2sdrc_u_rddatafifo_mem_2__2_) );
  DFFPOSX1 DFFPOSX1_82 ( .CLK(sdram_clk_bF_buf80), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_10__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_10_) );
  DFFPOSX1 DFFPOSX1_820 ( .CLK(sdram_clk_bF_buf40), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n270), .Q(u_wb2sdrc_u_rddatafifo_mem_2__3_) );
  DFFPOSX1 DFFPOSX1_821 ( .CLK(sdram_clk_bF_buf39), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n272), .Q(u_wb2sdrc_u_rddatafifo_mem_2__4_) );
  DFFPOSX1 DFFPOSX1_822 ( .CLK(sdram_clk_bF_buf38), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n274), .Q(u_wb2sdrc_u_rddatafifo_mem_2__5_) );
  DFFPOSX1 DFFPOSX1_823 ( .CLK(sdram_clk_bF_buf37), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n276), .Q(u_wb2sdrc_u_rddatafifo_mem_2__6_) );
  DFFPOSX1 DFFPOSX1_824 ( .CLK(sdram_clk_bF_buf36), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n278), .Q(u_wb2sdrc_u_rddatafifo_mem_2__7_) );
  DFFPOSX1 DFFPOSX1_825 ( .CLK(sdram_clk_bF_buf35), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n280), .Q(u_wb2sdrc_u_rddatafifo_mem_2__8_) );
  DFFPOSX1 DFFPOSX1_826 ( .CLK(sdram_clk_bF_buf34), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n282), .Q(u_wb2sdrc_u_rddatafifo_mem_2__9_) );
  DFFPOSX1 DFFPOSX1_827 ( .CLK(sdram_clk_bF_buf33), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n284), .Q(u_wb2sdrc_u_rddatafifo_mem_2__10_) );
  DFFPOSX1 DFFPOSX1_828 ( .CLK(sdram_clk_bF_buf32), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n286), .Q(u_wb2sdrc_u_rddatafifo_mem_2__11_) );
  DFFPOSX1 DFFPOSX1_829 ( .CLK(sdram_clk_bF_buf31), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n288), .Q(u_wb2sdrc_u_rddatafifo_mem_2__12_) );
  DFFPOSX1 DFFPOSX1_83 ( .CLK(sdram_clk_bF_buf79), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_11__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_11_) );
  DFFPOSX1 DFFPOSX1_830 ( .CLK(sdram_clk_bF_buf30), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n290), .Q(u_wb2sdrc_u_rddatafifo_mem_2__13_) );
  DFFPOSX1 DFFPOSX1_831 ( .CLK(sdram_clk_bF_buf29), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n292), .Q(u_wb2sdrc_u_rddatafifo_mem_2__14_) );
  DFFPOSX1 DFFPOSX1_832 ( .CLK(sdram_clk_bF_buf28), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n294), .Q(u_wb2sdrc_u_rddatafifo_mem_2__15_) );
  DFFPOSX1 DFFPOSX1_833 ( .CLK(sdram_clk_bF_buf27), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n296), .Q(u_wb2sdrc_u_rddatafifo_mem_2__16_) );
  DFFPOSX1 DFFPOSX1_834 ( .CLK(sdram_clk_bF_buf26), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n298), .Q(u_wb2sdrc_u_rddatafifo_mem_2__17_) );
  DFFPOSX1 DFFPOSX1_835 ( .CLK(sdram_clk_bF_buf25), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n300), .Q(u_wb2sdrc_u_rddatafifo_mem_2__18_) );
  DFFPOSX1 DFFPOSX1_836 ( .CLK(sdram_clk_bF_buf24), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n302), .Q(u_wb2sdrc_u_rddatafifo_mem_2__19_) );
  DFFPOSX1 DFFPOSX1_837 ( .CLK(sdram_clk_bF_buf23), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n304), .Q(u_wb2sdrc_u_rddatafifo_mem_2__20_) );
  DFFPOSX1 DFFPOSX1_838 ( .CLK(sdram_clk_bF_buf22), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n306), .Q(u_wb2sdrc_u_rddatafifo_mem_2__21_) );
  DFFPOSX1 DFFPOSX1_839 ( .CLK(sdram_clk_bF_buf21), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n308), .Q(u_wb2sdrc_u_rddatafifo_mem_2__22_) );
  DFFPOSX1 DFFPOSX1_84 ( .CLK(sdram_clk_bF_buf78), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_12__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_l_raddr_12_) );
  DFFPOSX1 DFFPOSX1_840 ( .CLK(sdram_clk_bF_buf20), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n310), .Q(u_wb2sdrc_u_rddatafifo_mem_2__23_) );
  DFFPOSX1 DFFPOSX1_841 ( .CLK(sdram_clk_bF_buf19), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n312), .Q(u_wb2sdrc_u_rddatafifo_mem_2__24_) );
  DFFPOSX1 DFFPOSX1_842 ( .CLK(sdram_clk_bF_buf18), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n314), .Q(u_wb2sdrc_u_rddatafifo_mem_2__25_) );
  DFFPOSX1 DFFPOSX1_843 ( .CLK(sdram_clk_bF_buf17), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n316), .Q(u_wb2sdrc_u_rddatafifo_mem_2__26_) );
  DFFPOSX1 DFFPOSX1_844 ( .CLK(sdram_clk_bF_buf16), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n318), .Q(u_wb2sdrc_u_rddatafifo_mem_2__27_) );
  DFFPOSX1 DFFPOSX1_845 ( .CLK(sdram_clk_bF_buf15), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n320), .Q(u_wb2sdrc_u_rddatafifo_mem_2__28_) );
  DFFPOSX1 DFFPOSX1_846 ( .CLK(sdram_clk_bF_buf14), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n322), .Q(u_wb2sdrc_u_rddatafifo_mem_2__29_) );
  DFFPOSX1 DFFPOSX1_847 ( .CLK(sdram_clk_bF_buf13), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n324), .Q(u_wb2sdrc_u_rddatafifo_mem_2__30_) );
  DFFPOSX1 DFFPOSX1_848 ( .CLK(sdram_clk_bF_buf12), .D(u_wb2sdrc_u_rddatafifo__abc_14216_n326), .Q(u_wb2sdrc_u_rddatafifo_mem_2__31_) );
  DFFPOSX1 DFFPOSX1_849 ( .CLK(wb_clk_i_bF_buf12), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n586), .Q(u_wb2sdrc_u_wrdatafifo_mem_3__0_) );
  DFFPOSX1 DFFPOSX1_85 ( .CLK(sdram_clk_bF_buf77), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_0__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_0_) );
  DFFPOSX1 DFFPOSX1_850 ( .CLK(wb_clk_i_bF_buf11), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n588), .Q(u_wb2sdrc_u_wrdatafifo_mem_3__1_) );
  DFFPOSX1 DFFPOSX1_851 ( .CLK(wb_clk_i_bF_buf10), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n590), .Q(u_wb2sdrc_u_wrdatafifo_mem_3__2_) );
  DFFPOSX1 DFFPOSX1_852 ( .CLK(wb_clk_i_bF_buf9), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n592), .Q(u_wb2sdrc_u_wrdatafifo_mem_3__3_) );
  DFFPOSX1 DFFPOSX1_853 ( .CLK(wb_clk_i_bF_buf8), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n594), .Q(u_wb2sdrc_u_wrdatafifo_mem_3__4_) );
  DFFPOSX1 DFFPOSX1_854 ( .CLK(wb_clk_i_bF_buf7), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n596), .Q(u_wb2sdrc_u_wrdatafifo_mem_3__5_) );
  DFFPOSX1 DFFPOSX1_855 ( .CLK(wb_clk_i_bF_buf6), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n598), .Q(u_wb2sdrc_u_wrdatafifo_mem_3__6_) );
  DFFPOSX1 DFFPOSX1_856 ( .CLK(wb_clk_i_bF_buf5), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n600), .Q(u_wb2sdrc_u_wrdatafifo_mem_3__7_) );
  DFFPOSX1 DFFPOSX1_857 ( .CLK(wb_clk_i_bF_buf4), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n602), .Q(u_wb2sdrc_u_wrdatafifo_mem_3__8_) );
  DFFPOSX1 DFFPOSX1_858 ( .CLK(wb_clk_i_bF_buf3), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n604), .Q(u_wb2sdrc_u_wrdatafifo_mem_3__9_) );
  DFFPOSX1 DFFPOSX1_859 ( .CLK(wb_clk_i_bF_buf2), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n606), .Q(u_wb2sdrc_u_wrdatafifo_mem_3__10_) );
  DFFPOSX1 DFFPOSX1_86 ( .CLK(sdram_clk_bF_buf76), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_1__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_1_) );
  DFFPOSX1 DFFPOSX1_860 ( .CLK(wb_clk_i_bF_buf1), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n608), .Q(u_wb2sdrc_u_wrdatafifo_mem_3__11_) );
  DFFPOSX1 DFFPOSX1_861 ( .CLK(wb_clk_i_bF_buf0), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n610), .Q(u_wb2sdrc_u_wrdatafifo_mem_3__12_) );
  DFFPOSX1 DFFPOSX1_862 ( .CLK(wb_clk_i_bF_buf59), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n612), .Q(u_wb2sdrc_u_wrdatafifo_mem_3__13_) );
  DFFPOSX1 DFFPOSX1_863 ( .CLK(wb_clk_i_bF_buf58), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n614), .Q(u_wb2sdrc_u_wrdatafifo_mem_3__14_) );
  DFFPOSX1 DFFPOSX1_864 ( .CLK(wb_clk_i_bF_buf57), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n616), .Q(u_wb2sdrc_u_wrdatafifo_mem_3__15_) );
  DFFPOSX1 DFFPOSX1_865 ( .CLK(wb_clk_i_bF_buf56), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n618), .Q(u_wb2sdrc_u_wrdatafifo_mem_3__16_) );
  DFFPOSX1 DFFPOSX1_866 ( .CLK(wb_clk_i_bF_buf55), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n620), .Q(u_wb2sdrc_u_wrdatafifo_mem_3__17_) );
  DFFPOSX1 DFFPOSX1_867 ( .CLK(wb_clk_i_bF_buf54), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n622), .Q(u_wb2sdrc_u_wrdatafifo_mem_3__18_) );
  DFFPOSX1 DFFPOSX1_868 ( .CLK(wb_clk_i_bF_buf53), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n624), .Q(u_wb2sdrc_u_wrdatafifo_mem_3__19_) );
  DFFPOSX1 DFFPOSX1_869 ( .CLK(wb_clk_i_bF_buf52), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n626), .Q(u_wb2sdrc_u_wrdatafifo_mem_3__20_) );
  DFFPOSX1 DFFPOSX1_87 ( .CLK(sdram_clk_bF_buf75), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_2__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_2_) );
  DFFPOSX1 DFFPOSX1_870 ( .CLK(wb_clk_i_bF_buf51), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n628), .Q(u_wb2sdrc_u_wrdatafifo_mem_3__21_) );
  DFFPOSX1 DFFPOSX1_871 ( .CLK(wb_clk_i_bF_buf50), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n630), .Q(u_wb2sdrc_u_wrdatafifo_mem_3__22_) );
  DFFPOSX1 DFFPOSX1_872 ( .CLK(wb_clk_i_bF_buf49), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n632), .Q(u_wb2sdrc_u_wrdatafifo_mem_3__23_) );
  DFFPOSX1 DFFPOSX1_873 ( .CLK(wb_clk_i_bF_buf48), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n634), .Q(u_wb2sdrc_u_wrdatafifo_mem_3__24_) );
  DFFPOSX1 DFFPOSX1_874 ( .CLK(wb_clk_i_bF_buf47), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n636), .Q(u_wb2sdrc_u_wrdatafifo_mem_3__25_) );
  DFFPOSX1 DFFPOSX1_875 ( .CLK(wb_clk_i_bF_buf46), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n638), .Q(u_wb2sdrc_u_wrdatafifo_mem_3__26_) );
  DFFPOSX1 DFFPOSX1_876 ( .CLK(wb_clk_i_bF_buf45), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n640), .Q(u_wb2sdrc_u_wrdatafifo_mem_3__27_) );
  DFFPOSX1 DFFPOSX1_877 ( .CLK(wb_clk_i_bF_buf44), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n642), .Q(u_wb2sdrc_u_wrdatafifo_mem_3__28_) );
  DFFPOSX1 DFFPOSX1_878 ( .CLK(wb_clk_i_bF_buf43), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n644), .Q(u_wb2sdrc_u_wrdatafifo_mem_3__29_) );
  DFFPOSX1 DFFPOSX1_879 ( .CLK(wb_clk_i_bF_buf42), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n646), .Q(u_wb2sdrc_u_wrdatafifo_mem_3__30_) );
  DFFPOSX1 DFFPOSX1_88 ( .CLK(sdram_clk_bF_buf74), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_3__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_3_) );
  DFFPOSX1 DFFPOSX1_880 ( .CLK(wb_clk_i_bF_buf41), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n648), .Q(u_wb2sdrc_u_wrdatafifo_mem_3__31_) );
  DFFPOSX1 DFFPOSX1_881 ( .CLK(wb_clk_i_bF_buf40), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n650), .Q(u_wb2sdrc_u_wrdatafifo_mem_3__32_) );
  DFFPOSX1 DFFPOSX1_882 ( .CLK(wb_clk_i_bF_buf39), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n652), .Q(u_wb2sdrc_u_wrdatafifo_mem_3__33_) );
  DFFPOSX1 DFFPOSX1_883 ( .CLK(wb_clk_i_bF_buf38), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n654), .Q(u_wb2sdrc_u_wrdatafifo_mem_3__34_) );
  DFFPOSX1 DFFPOSX1_884 ( .CLK(wb_clk_i_bF_buf37), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n656), .Q(u_wb2sdrc_u_wrdatafifo_mem_3__35_) );
  DFFPOSX1 DFFPOSX1_885 ( .CLK(wb_clk_i_bF_buf36), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n914), .Q(u_wb2sdrc_u_wrdatafifo_mem_2__0_) );
  DFFPOSX1 DFFPOSX1_886 ( .CLK(wb_clk_i_bF_buf35), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n916), .Q(u_wb2sdrc_u_wrdatafifo_mem_2__1_) );
  DFFPOSX1 DFFPOSX1_887 ( .CLK(wb_clk_i_bF_buf34), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n918), .Q(u_wb2sdrc_u_wrdatafifo_mem_2__2_) );
  DFFPOSX1 DFFPOSX1_888 ( .CLK(wb_clk_i_bF_buf33), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n920), .Q(u_wb2sdrc_u_wrdatafifo_mem_2__3_) );
  DFFPOSX1 DFFPOSX1_889 ( .CLK(wb_clk_i_bF_buf32), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n922), .Q(u_wb2sdrc_u_wrdatafifo_mem_2__4_) );
  DFFPOSX1 DFFPOSX1_89 ( .CLK(sdram_clk_bF_buf73), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_4__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_4_) );
  DFFPOSX1 DFFPOSX1_890 ( .CLK(wb_clk_i_bF_buf31), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n924), .Q(u_wb2sdrc_u_wrdatafifo_mem_2__5_) );
  DFFPOSX1 DFFPOSX1_891 ( .CLK(wb_clk_i_bF_buf30), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n926), .Q(u_wb2sdrc_u_wrdatafifo_mem_2__6_) );
  DFFPOSX1 DFFPOSX1_892 ( .CLK(wb_clk_i_bF_buf29), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n928), .Q(u_wb2sdrc_u_wrdatafifo_mem_2__7_) );
  DFFPOSX1 DFFPOSX1_893 ( .CLK(wb_clk_i_bF_buf28), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n930), .Q(u_wb2sdrc_u_wrdatafifo_mem_2__8_) );
  DFFPOSX1 DFFPOSX1_894 ( .CLK(wb_clk_i_bF_buf27), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n932), .Q(u_wb2sdrc_u_wrdatafifo_mem_2__9_) );
  DFFPOSX1 DFFPOSX1_895 ( .CLK(wb_clk_i_bF_buf26), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n934), .Q(u_wb2sdrc_u_wrdatafifo_mem_2__10_) );
  DFFPOSX1 DFFPOSX1_896 ( .CLK(wb_clk_i_bF_buf25), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n936), .Q(u_wb2sdrc_u_wrdatafifo_mem_2__11_) );
  DFFPOSX1 DFFPOSX1_897 ( .CLK(wb_clk_i_bF_buf24), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n938), .Q(u_wb2sdrc_u_wrdatafifo_mem_2__12_) );
  DFFPOSX1 DFFPOSX1_898 ( .CLK(wb_clk_i_bF_buf23), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n940), .Q(u_wb2sdrc_u_wrdatafifo_mem_2__13_) );
  DFFPOSX1 DFFPOSX1_899 ( .CLK(wb_clk_i_bF_buf22), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n942), .Q(u_wb2sdrc_u_wrdatafifo_mem_2__14_) );
  DFFPOSX1 DFFPOSX1_9 ( .CLK(sdram_clk_bF_buf72), .D(u_sdrc_core_pad_sdr_din1_8_), .Q(u_sdrc_core_pad_sdr_din2_8_) );
  DFFPOSX1 DFFPOSX1_90 ( .CLK(sdram_clk_bF_buf72), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_5__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_5_) );
  DFFPOSX1 DFFPOSX1_900 ( .CLK(wb_clk_i_bF_buf21), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n944), .Q(u_wb2sdrc_u_wrdatafifo_mem_2__15_) );
  DFFPOSX1 DFFPOSX1_901 ( .CLK(wb_clk_i_bF_buf20), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n946), .Q(u_wb2sdrc_u_wrdatafifo_mem_2__16_) );
  DFFPOSX1 DFFPOSX1_902 ( .CLK(wb_clk_i_bF_buf19), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n948), .Q(u_wb2sdrc_u_wrdatafifo_mem_2__17_) );
  DFFPOSX1 DFFPOSX1_903 ( .CLK(wb_clk_i_bF_buf18), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n950), .Q(u_wb2sdrc_u_wrdatafifo_mem_2__18_) );
  DFFPOSX1 DFFPOSX1_904 ( .CLK(wb_clk_i_bF_buf17), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n952), .Q(u_wb2sdrc_u_wrdatafifo_mem_2__19_) );
  DFFPOSX1 DFFPOSX1_905 ( .CLK(wb_clk_i_bF_buf16), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n954), .Q(u_wb2sdrc_u_wrdatafifo_mem_2__20_) );
  DFFPOSX1 DFFPOSX1_906 ( .CLK(wb_clk_i_bF_buf15), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n956), .Q(u_wb2sdrc_u_wrdatafifo_mem_2__21_) );
  DFFPOSX1 DFFPOSX1_907 ( .CLK(wb_clk_i_bF_buf14), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n958), .Q(u_wb2sdrc_u_wrdatafifo_mem_2__22_) );
  DFFPOSX1 DFFPOSX1_908 ( .CLK(wb_clk_i_bF_buf13), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n960), .Q(u_wb2sdrc_u_wrdatafifo_mem_2__23_) );
  DFFPOSX1 DFFPOSX1_909 ( .CLK(wb_clk_i_bF_buf12), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n962), .Q(u_wb2sdrc_u_wrdatafifo_mem_2__24_) );
  DFFPOSX1 DFFPOSX1_91 ( .CLK(sdram_clk_bF_buf71), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_6__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_6_) );
  DFFPOSX1 DFFPOSX1_910 ( .CLK(wb_clk_i_bF_buf11), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n964), .Q(u_wb2sdrc_u_wrdatafifo_mem_2__25_) );
  DFFPOSX1 DFFPOSX1_911 ( .CLK(wb_clk_i_bF_buf10), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n966), .Q(u_wb2sdrc_u_wrdatafifo_mem_2__26_) );
  DFFPOSX1 DFFPOSX1_912 ( .CLK(wb_clk_i_bF_buf9), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n968), .Q(u_wb2sdrc_u_wrdatafifo_mem_2__27_) );
  DFFPOSX1 DFFPOSX1_913 ( .CLK(wb_clk_i_bF_buf8), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n970), .Q(u_wb2sdrc_u_wrdatafifo_mem_2__28_) );
  DFFPOSX1 DFFPOSX1_914 ( .CLK(wb_clk_i_bF_buf7), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n972), .Q(u_wb2sdrc_u_wrdatafifo_mem_2__29_) );
  DFFPOSX1 DFFPOSX1_915 ( .CLK(wb_clk_i_bF_buf6), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n974), .Q(u_wb2sdrc_u_wrdatafifo_mem_2__30_) );
  DFFPOSX1 DFFPOSX1_916 ( .CLK(wb_clk_i_bF_buf5), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n976), .Q(u_wb2sdrc_u_wrdatafifo_mem_2__31_) );
  DFFPOSX1 DFFPOSX1_917 ( .CLK(wb_clk_i_bF_buf4), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n978), .Q(u_wb2sdrc_u_wrdatafifo_mem_2__32_) );
  DFFPOSX1 DFFPOSX1_918 ( .CLK(wb_clk_i_bF_buf3), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n980), .Q(u_wb2sdrc_u_wrdatafifo_mem_2__33_) );
  DFFPOSX1 DFFPOSX1_919 ( .CLK(wb_clk_i_bF_buf2), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n982), .Q(u_wb2sdrc_u_wrdatafifo_mem_2__34_) );
  DFFPOSX1 DFFPOSX1_92 ( .CLK(sdram_clk_bF_buf70), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_7__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_7_) );
  DFFPOSX1 DFFPOSX1_920 ( .CLK(wb_clk_i_bF_buf1), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n984), .Q(u_wb2sdrc_u_wrdatafifo_mem_2__35_) );
  DFFPOSX1 DFFPOSX1_921 ( .CLK(wb_clk_i_bF_buf0), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n876), .Q(u_wb2sdrc_u_wrdatafifo_mem_1__0_) );
  DFFPOSX1 DFFPOSX1_922 ( .CLK(wb_clk_i_bF_buf59), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n877), .Q(u_wb2sdrc_u_wrdatafifo_mem_1__1_) );
  DFFPOSX1 DFFPOSX1_923 ( .CLK(wb_clk_i_bF_buf58), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n878), .Q(u_wb2sdrc_u_wrdatafifo_mem_1__2_) );
  DFFPOSX1 DFFPOSX1_924 ( .CLK(wb_clk_i_bF_buf57), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n879), .Q(u_wb2sdrc_u_wrdatafifo_mem_1__3_) );
  DFFPOSX1 DFFPOSX1_925 ( .CLK(wb_clk_i_bF_buf56), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n880), .Q(u_wb2sdrc_u_wrdatafifo_mem_1__4_) );
  DFFPOSX1 DFFPOSX1_926 ( .CLK(wb_clk_i_bF_buf55), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n881), .Q(u_wb2sdrc_u_wrdatafifo_mem_1__5_) );
  DFFPOSX1 DFFPOSX1_927 ( .CLK(wb_clk_i_bF_buf54), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n882), .Q(u_wb2sdrc_u_wrdatafifo_mem_1__6_) );
  DFFPOSX1 DFFPOSX1_928 ( .CLK(wb_clk_i_bF_buf53), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n883), .Q(u_wb2sdrc_u_wrdatafifo_mem_1__7_) );
  DFFPOSX1 DFFPOSX1_929 ( .CLK(wb_clk_i_bF_buf52), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n884), .Q(u_wb2sdrc_u_wrdatafifo_mem_1__8_) );
  DFFPOSX1 DFFPOSX1_93 ( .CLK(sdram_clk_bF_buf69), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_8__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_8_) );
  DFFPOSX1 DFFPOSX1_930 ( .CLK(wb_clk_i_bF_buf51), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n885), .Q(u_wb2sdrc_u_wrdatafifo_mem_1__9_) );
  DFFPOSX1 DFFPOSX1_931 ( .CLK(wb_clk_i_bF_buf50), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n886), .Q(u_wb2sdrc_u_wrdatafifo_mem_1__10_) );
  DFFPOSX1 DFFPOSX1_932 ( .CLK(wb_clk_i_bF_buf49), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n887), .Q(u_wb2sdrc_u_wrdatafifo_mem_1__11_) );
  DFFPOSX1 DFFPOSX1_933 ( .CLK(wb_clk_i_bF_buf48), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n888), .Q(u_wb2sdrc_u_wrdatafifo_mem_1__12_) );
  DFFPOSX1 DFFPOSX1_934 ( .CLK(wb_clk_i_bF_buf47), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n889), .Q(u_wb2sdrc_u_wrdatafifo_mem_1__13_) );
  DFFPOSX1 DFFPOSX1_935 ( .CLK(wb_clk_i_bF_buf46), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n890), .Q(u_wb2sdrc_u_wrdatafifo_mem_1__14_) );
  DFFPOSX1 DFFPOSX1_936 ( .CLK(wb_clk_i_bF_buf45), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n891), .Q(u_wb2sdrc_u_wrdatafifo_mem_1__15_) );
  DFFPOSX1 DFFPOSX1_937 ( .CLK(wb_clk_i_bF_buf44), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n892), .Q(u_wb2sdrc_u_wrdatafifo_mem_1__16_) );
  DFFPOSX1 DFFPOSX1_938 ( .CLK(wb_clk_i_bF_buf43), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n893), .Q(u_wb2sdrc_u_wrdatafifo_mem_1__17_) );
  DFFPOSX1 DFFPOSX1_939 ( .CLK(wb_clk_i_bF_buf42), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n894), .Q(u_wb2sdrc_u_wrdatafifo_mem_1__18_) );
  DFFPOSX1 DFFPOSX1_94 ( .CLK(sdram_clk_bF_buf68), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_9__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_9_) );
  DFFPOSX1 DFFPOSX1_940 ( .CLK(wb_clk_i_bF_buf41), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n895), .Q(u_wb2sdrc_u_wrdatafifo_mem_1__19_) );
  DFFPOSX1 DFFPOSX1_941 ( .CLK(wb_clk_i_bF_buf40), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n896), .Q(u_wb2sdrc_u_wrdatafifo_mem_1__20_) );
  DFFPOSX1 DFFPOSX1_942 ( .CLK(wb_clk_i_bF_buf39), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n897), .Q(u_wb2sdrc_u_wrdatafifo_mem_1__21_) );
  DFFPOSX1 DFFPOSX1_943 ( .CLK(wb_clk_i_bF_buf38), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n898), .Q(u_wb2sdrc_u_wrdatafifo_mem_1__22_) );
  DFFPOSX1 DFFPOSX1_944 ( .CLK(wb_clk_i_bF_buf37), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n899), .Q(u_wb2sdrc_u_wrdatafifo_mem_1__23_) );
  DFFPOSX1 DFFPOSX1_945 ( .CLK(wb_clk_i_bF_buf36), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n900), .Q(u_wb2sdrc_u_wrdatafifo_mem_1__24_) );
  DFFPOSX1 DFFPOSX1_946 ( .CLK(wb_clk_i_bF_buf35), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n901), .Q(u_wb2sdrc_u_wrdatafifo_mem_1__25_) );
  DFFPOSX1 DFFPOSX1_947 ( .CLK(wb_clk_i_bF_buf34), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n902), .Q(u_wb2sdrc_u_wrdatafifo_mem_1__26_) );
  DFFPOSX1 DFFPOSX1_948 ( .CLK(wb_clk_i_bF_buf33), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n903), .Q(u_wb2sdrc_u_wrdatafifo_mem_1__27_) );
  DFFPOSX1 DFFPOSX1_949 ( .CLK(wb_clk_i_bF_buf32), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n904), .Q(u_wb2sdrc_u_wrdatafifo_mem_1__28_) );
  DFFPOSX1 DFFPOSX1_95 ( .CLK(sdram_clk_bF_buf67), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_10__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_10_) );
  DFFPOSX1 DFFPOSX1_950 ( .CLK(wb_clk_i_bF_buf31), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n905), .Q(u_wb2sdrc_u_wrdatafifo_mem_1__29_) );
  DFFPOSX1 DFFPOSX1_951 ( .CLK(wb_clk_i_bF_buf30), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n906), .Q(u_wb2sdrc_u_wrdatafifo_mem_1__30_) );
  DFFPOSX1 DFFPOSX1_952 ( .CLK(wb_clk_i_bF_buf29), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n907), .Q(u_wb2sdrc_u_wrdatafifo_mem_1__31_) );
  DFFPOSX1 DFFPOSX1_953 ( .CLK(wb_clk_i_bF_buf28), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n908), .Q(u_wb2sdrc_u_wrdatafifo_mem_1__32_) );
  DFFPOSX1 DFFPOSX1_954 ( .CLK(wb_clk_i_bF_buf27), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n909), .Q(u_wb2sdrc_u_wrdatafifo_mem_1__33_) );
  DFFPOSX1 DFFPOSX1_955 ( .CLK(wb_clk_i_bF_buf26), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n910), .Q(u_wb2sdrc_u_wrdatafifo_mem_1__34_) );
  DFFPOSX1 DFFPOSX1_956 ( .CLK(wb_clk_i_bF_buf25), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n911), .Q(u_wb2sdrc_u_wrdatafifo_mem_1__35_) );
  DFFPOSX1 DFFPOSX1_957 ( .CLK(wb_clk_i_bF_buf24), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n986), .Q(u_wb2sdrc_u_wrdatafifo_mem_5__0_) );
  DFFPOSX1 DFFPOSX1_958 ( .CLK(wb_clk_i_bF_buf23), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n987), .Q(u_wb2sdrc_u_wrdatafifo_mem_5__1_) );
  DFFPOSX1 DFFPOSX1_959 ( .CLK(wb_clk_i_bF_buf22), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n988), .Q(u_wb2sdrc_u_wrdatafifo_mem_5__2_) );
  DFFPOSX1 DFFPOSX1_96 ( .CLK(sdram_clk_bF_buf66), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_11__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_11_) );
  DFFPOSX1 DFFPOSX1_960 ( .CLK(wb_clk_i_bF_buf21), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n989), .Q(u_wb2sdrc_u_wrdatafifo_mem_5__3_) );
  DFFPOSX1 DFFPOSX1_961 ( .CLK(wb_clk_i_bF_buf20), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n990), .Q(u_wb2sdrc_u_wrdatafifo_mem_5__4_) );
  DFFPOSX1 DFFPOSX1_962 ( .CLK(wb_clk_i_bF_buf19), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n991), .Q(u_wb2sdrc_u_wrdatafifo_mem_5__5_) );
  DFFPOSX1 DFFPOSX1_963 ( .CLK(wb_clk_i_bF_buf18), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n992), .Q(u_wb2sdrc_u_wrdatafifo_mem_5__6_) );
  DFFPOSX1 DFFPOSX1_964 ( .CLK(wb_clk_i_bF_buf17), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n993), .Q(u_wb2sdrc_u_wrdatafifo_mem_5__7_) );
  DFFPOSX1 DFFPOSX1_965 ( .CLK(wb_clk_i_bF_buf16), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n994), .Q(u_wb2sdrc_u_wrdatafifo_mem_5__8_) );
  DFFPOSX1 DFFPOSX1_966 ( .CLK(wb_clk_i_bF_buf15), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n995), .Q(u_wb2sdrc_u_wrdatafifo_mem_5__9_) );
  DFFPOSX1 DFFPOSX1_967 ( .CLK(wb_clk_i_bF_buf14), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n996), .Q(u_wb2sdrc_u_wrdatafifo_mem_5__10_) );
  DFFPOSX1 DFFPOSX1_968 ( .CLK(wb_clk_i_bF_buf13), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n997), .Q(u_wb2sdrc_u_wrdatafifo_mem_5__11_) );
  DFFPOSX1 DFFPOSX1_969 ( .CLK(wb_clk_i_bF_buf12), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n998), .Q(u_wb2sdrc_u_wrdatafifo_mem_5__12_) );
  DFFPOSX1 DFFPOSX1_97 ( .CLK(sdram_clk_bF_buf65), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_12__FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_l_caddr_12_) );
  DFFPOSX1 DFFPOSX1_970 ( .CLK(wb_clk_i_bF_buf11), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n999), .Q(u_wb2sdrc_u_wrdatafifo_mem_5__13_) );
  DFFPOSX1 DFFPOSX1_971 ( .CLK(wb_clk_i_bF_buf10), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1000), .Q(u_wb2sdrc_u_wrdatafifo_mem_5__14_) );
  DFFPOSX1 DFFPOSX1_972 ( .CLK(wb_clk_i_bF_buf9), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1001), .Q(u_wb2sdrc_u_wrdatafifo_mem_5__15_) );
  DFFPOSX1 DFFPOSX1_973 ( .CLK(wb_clk_i_bF_buf8), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1002), .Q(u_wb2sdrc_u_wrdatafifo_mem_5__16_) );
  DFFPOSX1 DFFPOSX1_974 ( .CLK(wb_clk_i_bF_buf7), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1003), .Q(u_wb2sdrc_u_wrdatafifo_mem_5__17_) );
  DFFPOSX1 DFFPOSX1_975 ( .CLK(wb_clk_i_bF_buf6), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1004), .Q(u_wb2sdrc_u_wrdatafifo_mem_5__18_) );
  DFFPOSX1 DFFPOSX1_976 ( .CLK(wb_clk_i_bF_buf5), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1005), .Q(u_wb2sdrc_u_wrdatafifo_mem_5__19_) );
  DFFPOSX1 DFFPOSX1_977 ( .CLK(wb_clk_i_bF_buf4), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1006), .Q(u_wb2sdrc_u_wrdatafifo_mem_5__20_) );
  DFFPOSX1 DFFPOSX1_978 ( .CLK(wb_clk_i_bF_buf3), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1007), .Q(u_wb2sdrc_u_wrdatafifo_mem_5__21_) );
  DFFPOSX1 DFFPOSX1_979 ( .CLK(wb_clk_i_bF_buf2), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1008), .Q(u_wb2sdrc_u_wrdatafifo_mem_5__22_) );
  DFFPOSX1 DFFPOSX1_98 ( .CLK(sdram_clk_bF_buf64), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_l_sdr_dma_last_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_l_sdr_dma_last) );
  DFFPOSX1 DFFPOSX1_980 ( .CLK(wb_clk_i_bF_buf1), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1009), .Q(u_wb2sdrc_u_wrdatafifo_mem_5__23_) );
  DFFPOSX1 DFFPOSX1_981 ( .CLK(wb_clk_i_bF_buf0), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1010), .Q(u_wb2sdrc_u_wrdatafifo_mem_5__24_) );
  DFFPOSX1 DFFPOSX1_982 ( .CLK(wb_clk_i_bF_buf59), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1011), .Q(u_wb2sdrc_u_wrdatafifo_mem_5__25_) );
  DFFPOSX1 DFFPOSX1_983 ( .CLK(wb_clk_i_bF_buf58), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1012), .Q(u_wb2sdrc_u_wrdatafifo_mem_5__26_) );
  DFFPOSX1 DFFPOSX1_984 ( .CLK(wb_clk_i_bF_buf57), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1013), .Q(u_wb2sdrc_u_wrdatafifo_mem_5__27_) );
  DFFPOSX1 DFFPOSX1_985 ( .CLK(wb_clk_i_bF_buf56), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1014), .Q(u_wb2sdrc_u_wrdatafifo_mem_5__28_) );
  DFFPOSX1 DFFPOSX1_986 ( .CLK(wb_clk_i_bF_buf55), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1015), .Q(u_wb2sdrc_u_wrdatafifo_mem_5__29_) );
  DFFPOSX1 DFFPOSX1_987 ( .CLK(wb_clk_i_bF_buf54), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1016), .Q(u_wb2sdrc_u_wrdatafifo_mem_5__30_) );
  DFFPOSX1 DFFPOSX1_988 ( .CLK(wb_clk_i_bF_buf53), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1017), .Q(u_wb2sdrc_u_wrdatafifo_mem_5__31_) );
  DFFPOSX1 DFFPOSX1_989 ( .CLK(wb_clk_i_bF_buf52), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1018), .Q(u_wb2sdrc_u_wrdatafifo_mem_5__32_) );
  DFFPOSX1 DFFPOSX1_99 ( .CLK(sdram_clk_bF_buf63), .D(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_valid_FF_INPUT), .Q(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_valid) );
  DFFPOSX1 DFFPOSX1_990 ( .CLK(wb_clk_i_bF_buf51), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1019), .Q(u_wb2sdrc_u_wrdatafifo_mem_5__33_) );
  DFFPOSX1 DFFPOSX1_991 ( .CLK(wb_clk_i_bF_buf50), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1020), .Q(u_wb2sdrc_u_wrdatafifo_mem_5__34_) );
  DFFPOSX1 DFFPOSX1_992 ( .CLK(wb_clk_i_bF_buf49), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n1021), .Q(u_wb2sdrc_u_wrdatafifo_mem_5__35_) );
  DFFPOSX1 DFFPOSX1_993 ( .CLK(wb_clk_i_bF_buf48), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n154), .Q(u_wb2sdrc_u_wrdatafifo_mem_0__0_) );
  DFFPOSX1 DFFPOSX1_994 ( .CLK(wb_clk_i_bF_buf47), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n157), .Q(u_wb2sdrc_u_wrdatafifo_mem_0__1_) );
  DFFPOSX1 DFFPOSX1_995 ( .CLK(wb_clk_i_bF_buf46), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n160), .Q(u_wb2sdrc_u_wrdatafifo_mem_0__2_) );
  DFFPOSX1 DFFPOSX1_996 ( .CLK(wb_clk_i_bF_buf45), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n163), .Q(u_wb2sdrc_u_wrdatafifo_mem_0__3_) );
  DFFPOSX1 DFFPOSX1_997 ( .CLK(wb_clk_i_bF_buf44), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n166), .Q(u_wb2sdrc_u_wrdatafifo_mem_0__4_) );
  DFFPOSX1 DFFPOSX1_998 ( .CLK(wb_clk_i_bF_buf43), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n169), .Q(u_wb2sdrc_u_wrdatafifo_mem_0__5_) );
  DFFPOSX1 DFFPOSX1_999 ( .CLK(wb_clk_i_bF_buf42), .D(u_wb2sdrc_u_wrdatafifo__abc_14975_n172), .Q(u_wb2sdrc_u_wrdatafifo_mem_0__6_) );
  DFFSR DFFSR_1 ( .CLK(wb_clk_i_bF_buf59), .D(u_wb2sdrc_pending_read_FF_INPUT), .Q(u_wb2sdrc_pending_read), .R(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_10 ( .CLK(sdram_clk_bF_buf63), .D(u_wb2sdrc_u_cmdfifo_grey_rd_ptr_2__FF_INPUT), .Q(u_wb2sdrc_u_cmdfifo_grey_rd_ptr_2_), .R(sdram_resetn_bF_buf8), .S(1'b1) );
  DFFSR DFFSR_11 ( .CLK(sdram_clk_bF_buf62), .D(u_wb2sdrc_u_cmdfifo_rd_ptr_0__FF_INPUT), .Q(u_wb2sdrc_u_cmdfifo_rd_ptr_0_), .R(sdram_resetn_bF_buf7), .S(1'b1) );
  DFFSR DFFSR_12 ( .CLK(sdram_clk_bF_buf61), .D(u_wb2sdrc_u_cmdfifo_rd_ptr_1__FF_INPUT), .Q(u_wb2sdrc_u_cmdfifo_rd_ptr_1_), .R(sdram_resetn_bF_buf6), .S(1'b1) );
  DFFSR DFFSR_13 ( .CLK(sdram_clk_bF_buf60), .D(u_wb2sdrc_u_cmdfifo_rd_ptr_2__FF_INPUT), .Q(u_wb2sdrc_u_cmdfifo_rd_ptr_2_), .R(sdram_resetn_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_14 ( .CLK(sdram_clk_bF_buf59), .D(u_wb2sdrc_u_cmdfifo_empty_q_FF_INPUT), .Q(u_wb2sdrc_cmdfifo_empty), .R(1'b1), .S(sdram_resetn_bF_buf4) );
  DFFSR DFFSR_15 ( .CLK(wb_clk_i_bF_buf34), .D(u_wb2sdrc_u_cmdfifo_grey_rd_ptr_0_), .Q(u_wb2sdrc_u_cmdfifo_sync_rd_ptr_0_0_), .R(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_16 ( .CLK(wb_clk_i_bF_buf33), .D(u_wb2sdrc_u_cmdfifo_grey_rd_ptr_1_), .Q(u_wb2sdrc_u_cmdfifo_sync_rd_ptr_0_1_), .R(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_17 ( .CLK(wb_clk_i_bF_buf32), .D(u_wb2sdrc_u_cmdfifo_grey_rd_ptr_2_), .Q(u_wb2sdrc_u_cmdfifo_sync_rd_ptr_0_2_), .R(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_18 ( .CLK(wb_clk_i_bF_buf31), .D(u_wb2sdrc_u_cmdfifo_sync_rd_ptr_0_0_), .Q(u_wb2sdrc_u_cmdfifo_sync_rd_ptr_1_0_), .R(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_19 ( .CLK(wb_clk_i_bF_buf30), .D(u_wb2sdrc_u_cmdfifo_sync_rd_ptr_0_1_), .Q(u_wb2sdrc_u_cmdfifo_sync_rd_ptr_1_1_), .R(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_2 ( .CLK(sdram_clk_bF_buf71), .D(u_wb2sdrc_u_cmdfifo_grey_wr_ptr_0_), .Q(u_wb2sdrc_u_cmdfifo_sync_wr_ptr_0_0_), .R(sdram_resetn_bF_buf16), .S(1'b1) );
  DFFSR DFFSR_20 ( .CLK(wb_clk_i_bF_buf29), .D(u_wb2sdrc_u_cmdfifo_sync_rd_ptr_0_2_), .Q(u_wb2sdrc_u_cmdfifo_sync_rd_ptr_2_), .R(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_21 ( .CLK(wb_clk_i_bF_buf28), .D(u_wb2sdrc_u_cmdfifo_wr_ptr_0__FF_INPUT), .Q(u_wb2sdrc_u_cmdfifo_wr_ptr_0_), .R(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_22 ( .CLK(wb_clk_i_bF_buf27), .D(u_wb2sdrc_u_cmdfifo_wr_ptr_1__FF_INPUT), .Q(u_wb2sdrc_u_cmdfifo_wr_ptr_1_), .R(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_23 ( .CLK(wb_clk_i_bF_buf26), .D(u_wb2sdrc_u_cmdfifo_wr_ptr_2__FF_INPUT), .Q(u_wb2sdrc_u_cmdfifo_wr_ptr_2_), .R(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_24 ( .CLK(wb_clk_i_bF_buf25), .D(u_wb2sdrc_u_cmdfifo_grey_wr_ptr_0__FF_INPUT), .Q(u_wb2sdrc_u_cmdfifo_grey_wr_ptr_0_), .R(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_25 ( .CLK(wb_clk_i_bF_buf24), .D(u_wb2sdrc_u_cmdfifo_grey_wr_ptr_1__FF_INPUT), .Q(u_wb2sdrc_u_cmdfifo_grey_wr_ptr_1_), .R(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_26 ( .CLK(wb_clk_i_bF_buf23), .D(u_wb2sdrc_u_cmdfifo_grey_wr_ptr_2__FF_INPUT), .Q(u_wb2sdrc_u_cmdfifo_grey_wr_ptr_2_), .R(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_27 ( .CLK(wb_clk_i_bF_buf22), .D(u_wb2sdrc_u_cmdfifo_full_q_FF_INPUT), .Q(u_wb2sdrc_cmdfifo_full), .R(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_28 ( .CLK(wb_clk_i_bF_buf21), .D(u_wb2sdrc_u_rddatafifo_grey_wr_ptr_0_), .Q(u_wb2sdrc_u_rddatafifo_sync_wr_ptr_0_0_), .R(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_29 ( .CLK(wb_clk_i_bF_buf20), .D(u_wb2sdrc_u_rddatafifo_grey_wr_ptr_1_), .Q(u_wb2sdrc_u_rddatafifo_sync_wr_ptr_0_1_), .R(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_3 ( .CLK(sdram_clk_bF_buf70), .D(u_wb2sdrc_u_cmdfifo_grey_wr_ptr_1_), .Q(u_wb2sdrc_u_cmdfifo_sync_wr_ptr_0_1_), .R(sdram_resetn_bF_buf15), .S(1'b1) );
  DFFSR DFFSR_30 ( .CLK(wb_clk_i_bF_buf19), .D(u_wb2sdrc_u_rddatafifo_grey_wr_ptr_2_), .Q(u_wb2sdrc_u_rddatafifo_sync_wr_ptr_0_2_), .R(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_31 ( .CLK(wb_clk_i_bF_buf18), .D(u_wb2sdrc_u_rddatafifo_sync_wr_ptr_0_0_), .Q(u_wb2sdrc_u_rddatafifo_sync_wr_ptr_1_0_), .R(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_32 ( .CLK(wb_clk_i_bF_buf17), .D(u_wb2sdrc_u_rddatafifo_sync_wr_ptr_0_1_), .Q(u_wb2sdrc_u_rddatafifo_sync_wr_ptr_1_1_), .R(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_33 ( .CLK(wb_clk_i_bF_buf16), .D(u_wb2sdrc_u_rddatafifo_sync_wr_ptr_0_2_), .Q(u_wb2sdrc_u_rddatafifo_sync_wr_ptr_2_), .R(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_34 ( .CLK(wb_clk_i_bF_buf15), .D(u_wb2sdrc_u_rddatafifo_rd_ptr_0__FF_INPUT), .Q(u_wb2sdrc_u_rddatafifo_rd_ptr_0_), .R(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_35 ( .CLK(wb_clk_i_bF_buf14), .D(u_wb2sdrc_u_rddatafifo_rd_ptr_1__FF_INPUT), .Q(u_wb2sdrc_u_rddatafifo_rd_ptr_1_), .R(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_36 ( .CLK(wb_clk_i_bF_buf13), .D(u_wb2sdrc_u_rddatafifo_rd_ptr_2__FF_INPUT), .Q(u_wb2sdrc_u_rddatafifo_rd_ptr_2_), .R(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_37 ( .CLK(sdram_clk_bF_buf11), .D(u_wb2sdrc_u_rddatafifo_wr_ptr_0__FF_INPUT), .Q(u_wb2sdrc_u_rddatafifo_wr_ptr_0_), .R(sdram_resetn_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_38 ( .CLK(sdram_clk_bF_buf10), .D(u_wb2sdrc_u_rddatafifo_wr_ptr_1__FF_INPUT), .Q(u_wb2sdrc_u_rddatafifo_wr_ptr_1_), .R(sdram_resetn_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_39 ( .CLK(sdram_clk_bF_buf9), .D(u_wb2sdrc_u_rddatafifo_wr_ptr_2__FF_INPUT), .Q(u_wb2sdrc_u_rddatafifo_wr_ptr_2_), .R(sdram_resetn_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_4 ( .CLK(sdram_clk_bF_buf69), .D(u_wb2sdrc_u_cmdfifo_grey_wr_ptr_2_), .Q(u_wb2sdrc_u_cmdfifo_sync_wr_ptr_0_2_), .R(sdram_resetn_bF_buf14), .S(1'b1) );
  DFFSR DFFSR_40 ( .CLK(sdram_clk_bF_buf8), .D(u_wb2sdrc_u_rddatafifo_grey_wr_ptr_0__FF_INPUT), .Q(u_wb2sdrc_u_rddatafifo_grey_wr_ptr_0_), .R(sdram_resetn_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_41 ( .CLK(sdram_clk_bF_buf7), .D(u_wb2sdrc_u_rddatafifo_grey_wr_ptr_1__FF_INPUT), .Q(u_wb2sdrc_u_rddatafifo_grey_wr_ptr_1_), .R(sdram_resetn_bF_buf49), .S(1'b1) );
  DFFSR DFFSR_42 ( .CLK(sdram_clk_bF_buf6), .D(u_wb2sdrc_u_rddatafifo_grey_wr_ptr_2__FF_INPUT), .Q(u_wb2sdrc_u_rddatafifo_grey_wr_ptr_2_), .R(sdram_resetn_bF_buf48), .S(1'b1) );
  DFFSR DFFSR_43 ( .CLK(sdram_clk_bF_buf5), .D(u_wb2sdrc_u_wrdatafifo_grey_rd_ptr_0__FF_INPUT), .Q(u_wb2sdrc_u_wrdatafifo_grey_rd_ptr_0_), .R(sdram_resetn_bF_buf47), .S(1'b1) );
  DFFSR DFFSR_44 ( .CLK(sdram_clk_bF_buf4), .D(u_wb2sdrc_u_wrdatafifo_grey_rd_ptr_1__FF_INPUT), .Q(u_wb2sdrc_u_wrdatafifo_grey_rd_ptr_1_), .R(sdram_resetn_bF_buf46), .S(1'b1) );
  DFFSR DFFSR_45 ( .CLK(sdram_clk_bF_buf3), .D(u_wb2sdrc_u_wrdatafifo_grey_rd_ptr_2__FF_INPUT), .Q(u_wb2sdrc_u_wrdatafifo_grey_rd_ptr_2_), .R(sdram_resetn_bF_buf45), .S(1'b1) );
  DFFSR DFFSR_46 ( .CLK(sdram_clk_bF_buf2), .D(u_wb2sdrc_u_wrdatafifo_grey_rd_ptr_3__FF_INPUT), .Q(u_wb2sdrc_u_wrdatafifo_grey_rd_ptr_3_), .R(sdram_resetn_bF_buf44), .S(1'b1) );
  DFFSR DFFSR_47 ( .CLK(sdram_clk_bF_buf1), .D(u_wb2sdrc_u_wrdatafifo_rd_ptr_0__FF_INPUT), .Q(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_), .R(sdram_resetn_bF_buf43), .S(1'b1) );
  DFFSR DFFSR_48 ( .CLK(sdram_clk_bF_buf0), .D(u_wb2sdrc_u_wrdatafifo_rd_ptr_1__FF_INPUT), .Q(u_wb2sdrc_u_wrdatafifo_rd_ptr_1_), .R(sdram_resetn_bF_buf42), .S(1'b1) );
  DFFSR DFFSR_49 ( .CLK(sdram_clk_bF_buf80), .D(u_wb2sdrc_u_wrdatafifo_rd_ptr_2__FF_INPUT), .Q(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_), .R(sdram_resetn_bF_buf41), .S(1'b1) );
  DFFSR DFFSR_5 ( .CLK(sdram_clk_bF_buf68), .D(u_wb2sdrc_u_cmdfifo_sync_wr_ptr_0_0_), .Q(u_wb2sdrc_u_cmdfifo_sync_wr_ptr_1_0_), .R(sdram_resetn_bF_buf13), .S(1'b1) );
  DFFSR DFFSR_50 ( .CLK(sdram_clk_bF_buf79), .D(u_wb2sdrc_u_wrdatafifo_rd_ptr_3__FF_INPUT), .Q(u_wb2sdrc_u_wrdatafifo_rd_ptr_3_), .R(sdram_resetn_bF_buf40), .S(1'b1) );
  DFFSR DFFSR_51 ( .CLK(wb_clk_i_bF_buf24), .D(u_wb2sdrc_u_wrdatafifo_grey_rd_ptr_0_), .Q(u_wb2sdrc_u_wrdatafifo_sync_rd_ptr_0_0_), .R(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_52 ( .CLK(wb_clk_i_bF_buf23), .D(u_wb2sdrc_u_wrdatafifo_grey_rd_ptr_1_), .Q(u_wb2sdrc_u_wrdatafifo_sync_rd_ptr_0_1_), .R(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_53 ( .CLK(wb_clk_i_bF_buf22), .D(u_wb2sdrc_u_wrdatafifo_grey_rd_ptr_2_), .Q(u_wb2sdrc_u_wrdatafifo_sync_rd_ptr_0_2_), .R(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_54 ( .CLK(wb_clk_i_bF_buf21), .D(u_wb2sdrc_u_wrdatafifo_grey_rd_ptr_3_), .Q(u_wb2sdrc_u_wrdatafifo_sync_rd_ptr_0_3_), .R(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_55 ( .CLK(wb_clk_i_bF_buf20), .D(u_wb2sdrc_u_wrdatafifo_sync_rd_ptr_0_0_), .Q(u_wb2sdrc_u_wrdatafifo_sync_rd_ptr_1_0_), .R(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_56 ( .CLK(wb_clk_i_bF_buf19), .D(u_wb2sdrc_u_wrdatafifo_sync_rd_ptr_0_1_), .Q(u_wb2sdrc_u_wrdatafifo_sync_rd_ptr_1_1_), .R(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_57 ( .CLK(wb_clk_i_bF_buf18), .D(u_wb2sdrc_u_wrdatafifo_sync_rd_ptr_0_2_), .Q(u_wb2sdrc_u_wrdatafifo_sync_rd_ptr_1_2_), .R(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_58 ( .CLK(wb_clk_i_bF_buf17), .D(u_wb2sdrc_u_wrdatafifo_sync_rd_ptr_0_3_), .Q(u_wb2sdrc_u_wrdatafifo_sync_rd_ptr_1_3_), .R(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf5), .S(1'b1) );
  DFFSR DFFSR_59 ( .CLK(wb_clk_i_bF_buf16), .D(u_wb2sdrc_u_wrdatafifo_wr_ptr_0__FF_INPUT), .Q(u_wb2sdrc_u_wrdatafifo_wr_ptr_0_), .R(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf4), .S(1'b1) );
  DFFSR DFFSR_6 ( .CLK(sdram_clk_bF_buf67), .D(u_wb2sdrc_u_cmdfifo_sync_wr_ptr_0_1_), .Q(u_wb2sdrc_u_cmdfifo_sync_wr_ptr_1_1_), .R(sdram_resetn_bF_buf12), .S(1'b1) );
  DFFSR DFFSR_60 ( .CLK(wb_clk_i_bF_buf15), .D(u_wb2sdrc_u_wrdatafifo_wr_ptr_1__FF_INPUT), .Q(u_wb2sdrc_u_wrdatafifo_wr_ptr_1_), .R(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf3), .S(1'b1) );
  DFFSR DFFSR_61 ( .CLK(wb_clk_i_bF_buf14), .D(u_wb2sdrc_u_wrdatafifo_wr_ptr_2__FF_INPUT), .Q(u_wb2sdrc_u_wrdatafifo_wr_ptr_2_), .R(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf2), .S(1'b1) );
  DFFSR DFFSR_62 ( .CLK(wb_clk_i_bF_buf13), .D(u_wb2sdrc_u_wrdatafifo_wr_ptr_3__FF_INPUT), .Q(u_wb2sdrc_u_wrdatafifo_wr_ptr_3_), .R(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf1), .S(1'b1) );
  DFFSR DFFSR_63 ( .CLK(wb_clk_i_bF_buf12), .D(u_wb2sdrc_u_wrdatafifo_full_q_FF_INPUT), .Q(u_wb2sdrc_u_wrdatafifo_full), .R(u_wb2sdrc_u_cmdfifo_wr_reset_n_bF_buf0), .S(1'b1) );
  DFFSR DFFSR_7 ( .CLK(sdram_clk_bF_buf66), .D(u_wb2sdrc_u_cmdfifo_sync_wr_ptr_0_2_), .Q(u_wb2sdrc_u_cmdfifo_sync_wr_ptr_2_), .R(sdram_resetn_bF_buf11), .S(1'b1) );
  DFFSR DFFSR_8 ( .CLK(sdram_clk_bF_buf65), .D(u_wb2sdrc_u_cmdfifo_grey_rd_ptr_0__FF_INPUT), .Q(u_wb2sdrc_u_cmdfifo_grey_rd_ptr_0_), .R(sdram_resetn_bF_buf10), .S(1'b1) );
  DFFSR DFFSR_9 ( .CLK(sdram_clk_bF_buf64), .D(u_wb2sdrc_u_cmdfifo_grey_rd_ptr_1__FF_INPUT), .Q(u_wb2sdrc_u_cmdfifo_grey_rd_ptr_1_), .R(sdram_resetn_bF_buf9), .S(1'b1) );
  INVX1 INVX1_1 ( .A(u_sdrc_core_b2x_ba_0_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n211_1) );
  INVX1 INVX1_10 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n255), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n256_1) );
  INVX1 INVX1_100 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_2_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n314_1) );
  INVX1 INVX1_101 ( .A(u_sdrc_core_r2b_raddr_1_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n316_1) );
  INVX1 INVX1_102 ( .A(u_sdrc_core_r2b_raddr_4_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n320_1) );
  INVX1 INVX1_103 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_4_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n322_1) );
  INVX1 INVX1_104 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_5_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n325) );
  INVX1 INVX1_105 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n331_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n332_1) );
  INVX1 INVX1_106 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_refresh), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n336) );
  INVX1 INVX1_107 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_l_sdr_dma_last), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n353_1) );
  INVX1 INVX1_108 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n250_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n355) );
  INVX1 INVX1_109 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_prech_page_closed), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n356) );
  INVX1 INVX1_11 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n257), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n259_1) );
  INVX1 INVX1_110 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n357), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n358_1) );
  INVX1 INVX1_111 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_r2b_req), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n360) );
  INVX1 INVX1_112 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_4_bF_buf1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n367) );
  INVX1 INVX1_113 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n368_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n369_1) );
  INVX1 INVX1_114 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_tras_cntr_0_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n379_1) );
  INVX1 INVX1_115 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n380), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n381) );
  INVX1 INVX1_116 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n382), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n383_1) );
  INVX1 INVX1_117 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n384_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n393) );
  INVX1 INVX1_118 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n385), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n400_1) );
  INVX1 INVX1_119 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_timer0_0_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n413_1) );
  INVX1 INVX1_12 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n219_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n264) );
  INVX1 INVX1_120 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n424), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n425) );
  INVX1 INVX1_121 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n437_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n438_1) );
  INVX1 INVX1_122 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_l_write), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n730) );
  INVX1 INVX1_123 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n428_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n742) );
  INVX1 INVX1_124 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n386_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n745) );
  INVX1 INVX1_125 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_x2b_ack), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n249_1) );
  INVX1 INVX1_126 ( .A(u_sdrc_core_r2b_raddr_12_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n254) );
  INVX1 INVX1_127 ( .A(u_sdrc_core_r2b_raddr_11_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n256_1) );
  INVX1 INVX1_128 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_12_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n258_1) );
  INVX1 INVX1_129 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_11_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n262_1) );
  INVX1 INVX1_13 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n268_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n270_1) );
  INVX1 INVX1_130 ( .A(u_sdrc_core_r2b_raddr_9_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n264_1) );
  INVX1 INVX1_131 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_9_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n267_1) );
  INVX1 INVX1_132 ( .A(u_sdrc_core_r2b_raddr_7_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n269) );
  INVX1 INVX1_133 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_7_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n274_1) );
  INVX1 INVX1_134 ( .A(u_sdrc_core_r2b_raddr_3_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n276_1) );
  INVX1 INVX1_135 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_6_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n279_1) );
  INVX1 INVX1_136 ( .A(u_sdrc_core_r2b_raddr_6_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n281) );
  INVX1 INVX1_137 ( .A(u_sdrc_core_r2b_raddr_5_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n285) );
  INVX1 INVX1_138 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_1_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n287_1) );
  INVX1 INVX1_139 ( .A(u_sdrc_core_r2b_raddr_0_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n290_1) );
  INVX1 INVX1_14 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n278), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n279_1) );
  INVX1 INVX1_140 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_0_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n292_1) );
  INVX1 INVX1_141 ( .A(u_sdrc_core_r2b_raddr_10_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n299_1) );
  INVX1 INVX1_142 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_10_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n300_1) );
  INVX1 INVX1_143 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_8_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n304_1) );
  INVX1 INVX1_144 ( .A(u_sdrc_core_r2b_raddr_8_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n305) );
  INVX1 INVX1_145 ( .A(u_sdrc_core_r2b_raddr_2_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n309) );
  INVX1 INVX1_146 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_3_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n311_1) );
  INVX1 INVX1_147 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_2_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n314_1) );
  INVX1 INVX1_148 ( .A(u_sdrc_core_r2b_raddr_1_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n316_1) );
  INVX1 INVX1_149 ( .A(u_sdrc_core_r2b_raddr_4_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n320_1) );
  INVX1 INVX1_15 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n280_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n281_1) );
  INVX1 INVX1_150 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_4_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n322_1) );
  INVX1 INVX1_151 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_5_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n325) );
  INVX1 INVX1_152 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n331_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n332_1) );
  INVX1 INVX1_153 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_refresh), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n336) );
  INVX1 INVX1_154 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_l_sdr_dma_last), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n353_1) );
  INVX1 INVX1_155 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n250_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n355) );
  INVX1 INVX1_156 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_prech_page_closed), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n356) );
  INVX1 INVX1_157 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n357), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n358_1) );
  INVX1 INVX1_158 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_r2b_req), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n360) );
  INVX1 INVX1_159 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_4_bF_buf1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n367) );
  INVX1 INVX1_16 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n221_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n282_1) );
  INVX1 INVX1_160 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n368_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n369_1) );
  INVX1 INVX1_161 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_tras_cntr_0_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n379_1) );
  INVX1 INVX1_162 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n380), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n381) );
  INVX1 INVX1_163 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n382), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n383_1) );
  INVX1 INVX1_164 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n384_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n393) );
  INVX1 INVX1_165 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n385), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n400_1) );
  INVX1 INVX1_166 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_timer0_0_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n413_1) );
  INVX1 INVX1_167 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n424), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n425) );
  INVX1 INVX1_168 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n437_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n438_1) );
  INVX1 INVX1_169 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_l_write), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n730) );
  INVX1 INVX1_17 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_cmd_1_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n284_1) );
  INVX1 INVX1_170 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n428_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n742) );
  INVX1 INVX1_171 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n386_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n745) );
  INVX1 INVX1_172 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_x2b_ack), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n249_1) );
  INVX1 INVX1_173 ( .A(u_sdrc_core_r2b_raddr_12_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n254) );
  INVX1 INVX1_174 ( .A(u_sdrc_core_r2b_raddr_11_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n256_1) );
  INVX1 INVX1_175 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_12_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n258_1) );
  INVX1 INVX1_176 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_11_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n262_1) );
  INVX1 INVX1_177 ( .A(u_sdrc_core_r2b_raddr_9_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n264_1) );
  INVX1 INVX1_178 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_9_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n267_1) );
  INVX1 INVX1_179 ( .A(u_sdrc_core_r2b_raddr_7_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n269) );
  INVX1 INVX1_18 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_cmd_1_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n286_1) );
  INVX1 INVX1_180 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_7_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n274_1) );
  INVX1 INVX1_181 ( .A(u_sdrc_core_r2b_raddr_3_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n276_1) );
  INVX1 INVX1_182 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_6_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n279_1) );
  INVX1 INVX1_183 ( .A(u_sdrc_core_r2b_raddr_6_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n281) );
  INVX1 INVX1_184 ( .A(u_sdrc_core_r2b_raddr_5_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n285) );
  INVX1 INVX1_185 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_1_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n287_1) );
  INVX1 INVX1_186 ( .A(u_sdrc_core_r2b_raddr_0_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n290_1) );
  INVX1 INVX1_187 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_0_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n292_1) );
  INVX1 INVX1_188 ( .A(u_sdrc_core_r2b_raddr_10_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n299_1) );
  INVX1 INVX1_189 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_10_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n300_1) );
  INVX1 INVX1_19 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n229), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n290) );
  INVX1 INVX1_190 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_8_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n304_1) );
  INVX1 INVX1_191 ( .A(u_sdrc_core_r2b_raddr_8_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n305) );
  INVX1 INVX1_192 ( .A(u_sdrc_core_r2b_raddr_2_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n309) );
  INVX1 INVX1_193 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_3_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n311_1) );
  INVX1 INVX1_194 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_2_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n314_1) );
  INVX1 INVX1_195 ( .A(u_sdrc_core_r2b_raddr_1_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n316_1) );
  INVX1 INVX1_196 ( .A(u_sdrc_core_r2b_raddr_4_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n320_1) );
  INVX1 INVX1_197 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_4_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n322_1) );
  INVX1 INVX1_198 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_5_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n325) );
  INVX1 INVX1_199 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n331_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n332_1) );
  INVX1 INVX1_2 ( .A(u_sdrc_core_b2x_ba_1_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n213) );
  INVX1 INVX1_20 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n240_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n293) );
  INVX1 INVX1_200 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_refresh), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n336) );
  INVX1 INVX1_201 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_l_sdr_dma_last), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n353_1) );
  INVX1 INVX1_202 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n250_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n355) );
  INVX1 INVX1_203 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_prech_page_closed), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n356) );
  INVX1 INVX1_204 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n357), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n358_1) );
  INVX1 INVX1_205 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_r2b_req), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n360) );
  INVX1 INVX1_206 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_4_bF_buf1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n367) );
  INVX1 INVX1_207 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n368_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n369_1) );
  INVX1 INVX1_208 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_tras_cntr_0_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n379_1) );
  INVX1 INVX1_209 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n380), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n381) );
  INVX1 INVX1_21 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n315), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n316) );
  INVX1 INVX1_210 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n382), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n383_1) );
  INVX1 INVX1_211 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n384_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n393) );
  INVX1 INVX1_212 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n385), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n400_1) );
  INVX1 INVX1_213 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_timer0_0_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n413_1) );
  INVX1 INVX1_214 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n424), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n425) );
  INVX1 INVX1_215 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n437_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n438_1) );
  INVX1 INVX1_216 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_l_write), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n730) );
  INVX1 INVX1_217 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n428_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n742) );
  INVX1 INVX1_218 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n386_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n745) );
  INVX1 INVX1_219 ( .A(\cfg_sdr_width[0] ), .Y(u_sdrc_core_u_bs_convert__abc_21684_n168_1) );
  INVX1 INVX1_22 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n319), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n320_1) );
  INVX1 INVX1_220 ( .A(cfg_sdr_width_1_bF_buf5), .Y(u_sdrc_core_u_bs_convert__abc_21684_n169_1) );
  INVX1 INVX1_221 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_1_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n173_1) );
  INVX1 INVX1_222 ( .A(app_wr_data_24_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n186_1) );
  INVX1 INVX1_223 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n188_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n189_1) );
  INVX1 INVX1_224 ( .A(app_wr_data_25_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n205) );
  INVX1 INVX1_225 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n206_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n207_1) );
  INVX1 INVX1_226 ( .A(app_wr_data_26_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n223) );
  INVX1 INVX1_227 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n224_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n225) );
  INVX1 INVX1_228 ( .A(app_wr_data_27_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n239) );
  INVX1 INVX1_229 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n240), .Y(u_sdrc_core_u_bs_convert__abc_21684_n241) );
  INVX1 INVX1_23 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n269), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n335) );
  INVX1 INVX1_230 ( .A(app_wr_data_28_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n256) );
  INVX1 INVX1_231 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n257), .Y(u_sdrc_core_u_bs_convert__abc_21684_n258_1) );
  INVX1 INVX1_232 ( .A(app_wr_data_29_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n274) );
  INVX1 INVX1_233 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n275), .Y(u_sdrc_core_u_bs_convert__abc_21684_n276) );
  INVX1 INVX1_234 ( .A(app_wr_data_30_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n293) );
  INVX1 INVX1_235 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n294), .Y(u_sdrc_core_u_bs_convert__abc_21684_n295) );
  INVX1 INVX1_236 ( .A(app_wr_data_31_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n309) );
  INVX1 INVX1_237 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n310), .Y(u_sdrc_core_u_bs_convert__abc_21684_n311) );
  INVX1 INVX1_238 ( .A(app_wr_en_n_3_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n360) );
  INVX1 INVX1_239 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n361_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n362) );
  INVX1 INVX1_24 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n338), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n339) );
  INVX1 INVX1_240 ( .A(app_last_wr), .Y(u_sdrc_core_u_bs_convert__abc_21684_n481) );
  INVX1 INVX1_241 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n483), .Y(u_sdrc_core_u_bs_convert__abc_21684_n484) );
  INVX1 INVX1_242 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n488), .Y(u_sdrc_core_u_bs_convert__abc_21684_n489) );
  INVX1 INVX1_243 ( .A(app_last_rd), .Y(u_sdrc_core_u_bs_convert__abc_21684_n493) );
  INVX1 INVX1_244 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n495), .Y(u_sdrc_core_u_bs_convert__abc_21684_n496) );
  INVX1 INVX1_245 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n500), .Y(u_sdrc_core_u_bs_convert__abc_21684_n501) );
  INVX1 INVX1_246 ( .A(u_sdrc_core_u_bs_convert_rd_xfr_count_0_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n505) );
  INVX1 INVX1_247 ( .A(u_sdrc_core_b2r_ack), .Y(u_sdrc_core_u_req_gen__abc_22171_n181) );
  INVX1 INVX1_248 ( .A(u_sdrc_core_u_req_gen__abc_22171_n190), .Y(u_sdrc_core_u_req_gen__abc_22171_n193) );
  INVX1 INVX1_249 ( .A(u_sdrc_core_u_req_gen_page_ovflw_r), .Y(u_sdrc_core_u_req_gen__abc_22171_n195_1) );
  INVX1 INVX1_25 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n355), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n356) );
  INVX1 INVX1_250 ( .A(sdram_resetn_bF_buf23), .Y(u_sdrc_core_u_req_gen__abc_22171_n197) );
  INVX1 INVX1_251 ( .A(u_sdrc_core_u_req_gen__abc_22171_n202), .Y(u_sdrc_core_u_req_gen__abc_22171_n204) );
  INVX1 INVX1_252 ( .A(u_sdrc_core_u_req_gen_max_r2b_len_r_1_), .Y(u_sdrc_core_u_req_gen__abc_22171_n208) );
  INVX1 INVX1_253 ( .A(u_sdrc_core_u_req_gen__abc_22171_n209), .Y(u_sdrc_core_u_req_gen__abc_22171_n210_1) );
  INVX1 INVX1_254 ( .A(u_sdrc_core_u_req_gen_lcl_req_len_2_), .Y(u_sdrc_core_u_req_gen__abc_22171_n212) );
  INVX1 INVX1_255 ( .A(u_sdrc_core_u_req_gen_max_r2b_len_r_2_), .Y(u_sdrc_core_u_req_gen__abc_22171_n214) );
  INVX1 INVX1_256 ( .A(u_sdrc_core_u_req_gen_lcl_req_len_3_), .Y(u_sdrc_core_u_req_gen__abc_22171_n218) );
  INVX1 INVX1_257 ( .A(u_sdrc_core_u_req_gen_max_r2b_len_r_3_), .Y(u_sdrc_core_u_req_gen__abc_22171_n220) );
  INVX1 INVX1_258 ( .A(u_sdrc_core_u_req_gen_max_r2b_len_r_4_), .Y(u_sdrc_core_u_req_gen__abc_22171_n225) );
  INVX1 INVX1_259 ( .A(u_sdrc_core_u_req_gen__abc_22171_n226_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n227) );
  INVX1 INVX1_26 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n358), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n359) );
  INVX1 INVX1_260 ( .A(u_sdrc_core_u_req_gen_max_r2b_len_r_5_), .Y(u_sdrc_core_u_req_gen__abc_22171_n230) );
  INVX1 INVX1_261 ( .A(u_sdrc_core_u_req_gen__abc_22171_n231), .Y(u_sdrc_core_u_req_gen__abc_22171_n232) );
  INVX1 INVX1_262 ( .A(u_sdrc_core_u_req_gen_max_r2b_len_r_6_), .Y(u_sdrc_core_u_req_gen__abc_22171_n235) );
  INVX1 INVX1_263 ( .A(u_sdrc_core_u_req_gen__abc_22171_n236_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n237) );
  INVX1 INVX1_264 ( .A(\cfg_sdr_width[0] ), .Y(u_sdrc_core_u_req_gen__abc_22171_n240) );
  INVX1 INVX1_265 ( .A(u_sdrc_core_u_req_gen__abc_22171_n249), .Y(u_sdrc_core_u_req_gen__abc_22171_n250) );
  INVX1 INVX1_266 ( .A(u_sdrc_core_u_req_gen__abc_22171_n252), .Y(u_sdrc_core_u_req_gen__abc_22171_n253) );
  INVX1 INVX1_267 ( .A(app_req_addr_2_), .Y(u_sdrc_core_u_req_gen__abc_22171_n255) );
  INVX1 INVX1_268 ( .A(app_req_addr_0_), .Y(u_sdrc_core_u_req_gen__abc_22171_n257) );
  INVX1 INVX1_269 ( .A(app_req_addr_1_), .Y(u_sdrc_core_u_req_gen__abc_22171_n259) );
  INVX1 INVX1_27 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n615), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n616) );
  INVX1 INVX1_270 ( .A(u_sdrc_core_u_req_gen__abc_22171_n262_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n264) );
  INVX1 INVX1_271 ( .A(u_sdrc_core_u_req_gen__abc_22171_n266), .Y(u_sdrc_core_u_req_gen__abc_22171_n267) );
  INVX1 INVX1_272 ( .A(app_req_addr_3_), .Y(u_sdrc_core_u_req_gen__abc_22171_n269) );
  INVX1 INVX1_273 ( .A(u_sdrc_core_u_req_gen__abc_22171_n275), .Y(u_sdrc_core_u_req_gen__abc_22171_n276) );
  INVX1 INVX1_274 ( .A(app_req_addr_4_), .Y(u_sdrc_core_u_req_gen__abc_22171_n280) );
  INVX1 INVX1_275 ( .A(u_sdrc_core_u_req_gen__abc_22171_n285), .Y(u_sdrc_core_u_req_gen__abc_22171_n287) );
  INVX1 INVX1_276 ( .A(u_sdrc_core_u_req_gen__abc_22171_n289), .Y(u_sdrc_core_u_req_gen__abc_22171_n290_1) );
  INVX1 INVX1_277 ( .A(app_req_addr_5_), .Y(u_sdrc_core_u_req_gen__abc_22171_n292) );
  INVX1 INVX1_278 ( .A(u_sdrc_core_u_req_gen__abc_22171_n298_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n299) );
  INVX1 INVX1_279 ( .A(u_sdrc_core_u_req_gen__abc_22171_n307_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n308) );
  INVX1 INVX1_28 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n619), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n620) );
  INVX1 INVX1_280 ( .A(u_sdrc_core_u_req_gen__abc_22171_n311), .Y(u_sdrc_core_u_req_gen__abc_22171_n312) );
  INVX1 INVX1_281 ( .A(u_sdrc_core_u_req_gen__abc_22171_n314), .Y(u_sdrc_core_u_req_gen__abc_22171_n315) );
  INVX1 INVX1_282 ( .A(u_sdrc_core_u_req_gen_req_st_0_), .Y(u_sdrc_core_r2b_req) );
  INVX1 INVX1_283 ( .A(u_sdrc_core_u_req_gen__abc_22171_n336), .Y(u_sdrc_core_u_req_gen__abc_22171_n337_1) );
  INVX1 INVX1_284 ( .A(u_sdrc_core_u_req_gen_lcl_req_len_0_), .Y(u_sdrc_core_u_req_gen__abc_22171_n339) );
  INVX1 INVX1_285 ( .A(u_sdrc_core_u_req_gen_lcl_req_len_1_), .Y(u_sdrc_core_u_req_gen__abc_22171_n349) );
  INVX1 INVX1_286 ( .A(u_sdrc_core_u_req_gen__abc_22171_n347), .Y(u_sdrc_core_u_req_gen__abc_22171_n353) );
  INVX1 INVX1_287 ( .A(u_sdrc_core_u_req_gen__abc_22171_n351), .Y(u_sdrc_core_u_req_gen__abc_22171_n354_1) );
  INVX1 INVX1_288 ( .A(u_sdrc_core_u_req_gen__abc_22171_n348), .Y(u_sdrc_core_u_req_gen__abc_22171_n366) );
  INVX1 INVX1_289 ( .A(u_sdrc_core_u_req_gen__abc_22171_n367), .Y(u_sdrc_core_u_req_gen__abc_22171_n372) );
  INVX1 INVX1_29 ( .A(u_sdrc_core_r2b_ba_0_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n625) );
  INVX1 INVX1_290 ( .A(u_sdrc_core_u_req_gen__abc_22171_n370), .Y(u_sdrc_core_u_req_gen__abc_22171_n373_1) );
  INVX1 INVX1_291 ( .A(app_req_len_2_), .Y(u_sdrc_core_u_req_gen__abc_22171_n380) );
  INVX1 INVX1_292 ( .A(app_req_len_0_), .Y(u_sdrc_core_u_req_gen__abc_22171_n382_1) );
  INVX1 INVX1_293 ( .A(app_req_len_1_), .Y(u_sdrc_core_u_req_gen__abc_22171_n384) );
  INVX1 INVX1_294 ( .A(u_sdrc_core_u_req_gen__abc_22171_n387), .Y(u_sdrc_core_u_req_gen__abc_22171_n388_1) );
  INVX1 INVX1_295 ( .A(u_sdrc_core_u_req_gen__abc_22171_n395), .Y(u_sdrc_core_u_req_gen__abc_22171_n396_1) );
  INVX1 INVX1_296 ( .A(u_sdrc_core_u_req_gen__abc_22171_n368), .Y(u_sdrc_core_u_req_gen__abc_22171_n400_1) );
  INVX1 INVX1_297 ( .A(u_sdrc_core_u_req_gen__abc_22171_n401), .Y(u_sdrc_core_u_req_gen__abc_22171_n402) );
  INVX1 INVX1_298 ( .A(u_sdrc_core_u_req_gen__abc_22171_n405), .Y(u_sdrc_core_u_req_gen__abc_22171_n406_1) );
  INVX1 INVX1_299 ( .A(u_sdrc_core_u_req_gen__abc_22171_n403), .Y(u_sdrc_core_u_req_gen__abc_22171_n422) );
  INVX1 INVX1_3 ( .A(u_sdrc_core_u_bank_ctl_rank_cnt_0_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n217_1) );
  INVX1 INVX1_30 ( .A(u_sdrc_core_r2b_ba_1_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n626) );
  INVX1 INVX1_300 ( .A(u_sdrc_core_u_req_gen__abc_22171_n423_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n424) );
  INVX1 INVX1_301 ( .A(u_sdrc_core_u_req_gen__abc_22171_n425_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n426) );
  INVX1 INVX1_302 ( .A(u_sdrc_core_r2b_len_4_), .Y(u_sdrc_core_u_req_gen__abc_22171_n427) );
  INVX1 INVX1_303 ( .A(u_sdrc_core_u_req_gen__abc_22171_n429_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n431_1) );
  INVX1 INVX1_304 ( .A(u_sdrc_core_u_req_gen__abc_22171_n445), .Y(u_sdrc_core_u_req_gen__abc_22171_n446) );
  INVX1 INVX1_305 ( .A(u_sdrc_core_u_req_gen__abc_22171_n447), .Y(u_sdrc_core_u_req_gen__abc_22171_n448_1) );
  INVX1 INVX1_306 ( .A(u_sdrc_core_r2b_len_5_), .Y(u_sdrc_core_u_req_gen__abc_22171_n449) );
  INVX1 INVX1_307 ( .A(u_sdrc_core_u_req_gen__abc_22171_n451_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n453) );
  INVX1 INVX1_308 ( .A(u_sdrc_core_u_req_gen_lcl_req_len_6_), .Y(u_sdrc_core_u_req_gen__abc_22171_n466_1) );
  INVX1 INVX1_309 ( .A(u_sdrc_core_u_req_gen__abc_22171_n468_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n469) );
  INVX1 INVX1_31 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_ack), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n249_1) );
  INVX1 INVX1_310 ( .A(u_sdrc_core_u_req_gen__abc_22171_n472), .Y(u_sdrc_core_u_req_gen__abc_22171_n473) );
  INVX1 INVX1_311 ( .A(u_sdrc_core_u_req_gen__abc_22171_n479), .Y(u_sdrc_core_u_req_gen__abc_22171_n480_1) );
  INVX1 INVX1_312 ( .A(u_sdrc_core_r2b_caddr_1_), .Y(u_sdrc_core_u_req_gen__abc_22171_n486_1) );
  INVX1 INVX1_313 ( .A(u_sdrc_core_u_req_gen__abc_22171_n492_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n493) );
  INVX1 INVX1_314 ( .A(u_sdrc_core_u_req_gen__abc_22171_n504_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n505) );
  INVX1 INVX1_315 ( .A(u_sdrc_core_u_req_gen__abc_22171_n508_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n509_1) );
  INVX1 INVX1_316 ( .A(u_sdrc_core_u_req_gen__abc_22171_n519), .Y(u_sdrc_core_u_req_gen__abc_22171_n520) );
  INVX1 INVX1_317 ( .A(u_sdrc_core_r2b_caddr_3_), .Y(u_sdrc_core_u_req_gen__abc_22171_n521) );
  INVX1 INVX1_318 ( .A(u_sdrc_core_u_req_gen__abc_22171_n523), .Y(u_sdrc_core_u_req_gen__abc_22171_n524) );
  INVX1 INVX1_319 ( .A(u_sdrc_core_u_req_gen__abc_22171_n525), .Y(u_sdrc_core_u_req_gen__abc_22171_n527_1) );
  INVX1 INVX1_32 ( .A(u_sdrc_core_r2b_raddr_12_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n254) );
  INVX1 INVX1_320 ( .A(u_sdrc_core_u_req_gen__abc_22171_n274), .Y(u_sdrc_core_u_req_gen__abc_22171_n533) );
  INVX1 INVX1_321 ( .A(u_sdrc_core_u_req_gen__abc_22171_n538), .Y(u_sdrc_core_u_req_gen__abc_22171_n539) );
  INVX1 INVX1_322 ( .A(u_sdrc_core_u_req_gen__abc_22171_n522), .Y(u_sdrc_core_u_req_gen__abc_22171_n542) );
  INVX1 INVX1_323 ( .A(u_sdrc_core_u_req_gen__abc_22171_n549), .Y(u_sdrc_core_u_req_gen__abc_22171_n550) );
  INVX1 INVX1_324 ( .A(u_sdrc_core_u_req_gen__abc_22171_n557), .Y(u_sdrc_core_u_req_gen__abc_22171_n558) );
  INVX1 INVX1_325 ( .A(u_sdrc_core_u_req_gen__abc_22171_n559), .Y(u_sdrc_core_u_req_gen__abc_22171_n560) );
  INVX1 INVX1_326 ( .A(u_sdrc_core_u_req_gen__abc_22171_n562), .Y(u_sdrc_core_u_req_gen__abc_22171_n564) );
  INVX1 INVX1_327 ( .A(u_sdrc_core_u_req_gen__abc_22171_n297), .Y(u_sdrc_core_u_req_gen__abc_22171_n570) );
  INVX1 INVX1_328 ( .A(u_sdrc_core_u_req_gen__abc_22171_n580), .Y(u_sdrc_core_u_req_gen__abc_22171_n581) );
  INVX1 INVX1_329 ( .A(u_sdrc_core_u_req_gen__abc_22171_n585), .Y(u_sdrc_core_u_req_gen__abc_22171_n586) );
  INVX1 INVX1_33 ( .A(u_sdrc_core_r2b_raddr_11_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n256_1) );
  INVX1 INVX1_330 ( .A(u_sdrc_core_r2b_caddr_7_), .Y(u_sdrc_core_u_req_gen__abc_22171_n598) );
  INVX1 INVX1_331 ( .A(u_sdrc_core_u_req_gen__abc_22171_n600), .Y(u_sdrc_core_u_req_gen__abc_22171_n601) );
  INVX1 INVX1_332 ( .A(u_sdrc_core_u_req_gen__abc_22171_n622), .Y(u_sdrc_core_u_req_gen__abc_22171_n623) );
  INVX1 INVX1_333 ( .A(u_sdrc_core_u_req_gen__abc_22171_n635), .Y(u_sdrc_core_u_req_gen__abc_22171_n636) );
  INVX1 INVX1_334 ( .A(u_sdrc_core_u_req_gen__abc_22171_n646), .Y(u_sdrc_core_u_req_gen__abc_22171_n647) );
  INVX1 INVX1_335 ( .A(u_sdrc_core_u_req_gen__abc_22171_n660), .Y(u_sdrc_core_u_req_gen__abc_22171_n661) );
  INVX1 INVX1_336 ( .A(u_sdrc_core_u_req_gen__abc_22171_n672), .Y(u_sdrc_core_u_req_gen__abc_22171_n673) );
  INVX1 INVX1_337 ( .A(u_sdrc_core_u_req_gen__abc_22171_n681), .Y(u_sdrc_core_u_req_gen__abc_22171_n682) );
  INVX1 INVX1_338 ( .A(u_sdrc_core_u_req_gen__abc_22171_n693), .Y(u_sdrc_core_u_req_gen__abc_22171_n694) );
  INVX1 INVX1_339 ( .A(u_sdrc_core_u_req_gen__abc_22171_n714), .Y(u_sdrc_core_u_req_gen__abc_22171_n715) );
  INVX1 INVX1_34 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_12_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n258_1) );
  INVX1 INVX1_340 ( .A(u_sdrc_core_u_req_gen__abc_22171_n725), .Y(u_sdrc_core_u_req_gen__abc_22171_n726) );
  INVX1 INVX1_341 ( .A(u_sdrc_core_u_req_gen__abc_22171_n738), .Y(u_sdrc_core_u_req_gen__abc_22171_n739) );
  INVX1 INVX1_342 ( .A(u_sdrc_core_u_req_gen_curr_sdr_addr_18_), .Y(u_sdrc_core_u_req_gen__abc_22171_n751) );
  INVX1 INVX1_343 ( .A(u_sdrc_core_u_req_gen__abc_22171_n761), .Y(u_sdrc_core_u_req_gen__abc_22171_n762) );
  INVX1 INVX1_344 ( .A(u_sdrc_core_u_req_gen__abc_22171_n780), .Y(u_sdrc_core_u_req_gen__abc_22171_n781) );
  INVX1 INVX1_345 ( .A(u_sdrc_core_u_req_gen__abc_22171_n785), .Y(u_sdrc_core_u_req_gen__abc_22171_n786) );
  INVX1 INVX1_346 ( .A(u_sdrc_core_u_req_gen__abc_22171_n790), .Y(u_sdrc_core_u_req_gen__abc_22171_n791) );
  INVX1 INVX1_347 ( .A(u_sdrc_core_u_req_gen__abc_22171_n793), .Y(u_sdrc_core_u_req_gen__abc_22171_n794) );
  INVX1 INVX1_348 ( .A(u_sdrc_core_u_req_gen__abc_22171_n798), .Y(u_sdrc_core_u_req_gen_map_address_21_) );
  INVX1 INVX1_349 ( .A(u_sdrc_core_u_req_gen__abc_22171_n804), .Y(u_sdrc_core_u_req_gen__abc_22171_n805) );
  INVX1 INVX1_35 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_11_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n262_1) );
  INVX1 INVX1_350 ( .A(u_sdrc_core_u_req_gen_curr_sdr_addr_22_), .Y(u_sdrc_core_u_req_gen__abc_22171_n807) );
  INVX1 INVX1_351 ( .A(u_sdrc_core_u_req_gen__abc_22171_n808), .Y(u_sdrc_core_u_req_gen__abc_22171_n809) );
  INVX1 INVX1_352 ( .A(u_sdrc_core_u_req_gen__abc_22171_n813), .Y(u_sdrc_core_u_req_gen_map_address_22_) );
  INVX1 INVX1_353 ( .A(u_sdrc_core_u_req_gen__abc_22171_n820), .Y(u_sdrc_core_u_req_gen__abc_22171_n821) );
  INVX1 INVX1_354 ( .A(u_sdrc_core_u_req_gen_curr_sdr_addr_23_), .Y(u_sdrc_core_u_req_gen__abc_22171_n822) );
  INVX1 INVX1_355 ( .A(u_sdrc_core_u_req_gen__abc_22171_n825), .Y(u_sdrc_core_u_req_gen__abc_22171_n826) );
  INVX1 INVX1_356 ( .A(u_sdrc_core_u_req_gen__abc_22171_n831), .Y(u_sdrc_core_u_req_gen_map_address_23_) );
  INVX1 INVX1_357 ( .A(u_sdrc_core_u_req_gen__abc_22171_n838), .Y(u_sdrc_core_u_req_gen__abc_22171_n839) );
  INVX1 INVX1_358 ( .A(u_sdrc_core_u_req_gen_curr_sdr_addr_24_), .Y(u_sdrc_core_u_req_gen__abc_22171_n840) );
  INVX1 INVX1_359 ( .A(u_sdrc_core_u_req_gen__abc_22171_n844), .Y(u_sdrc_core_u_req_gen__abc_22171_n845) );
  INVX1 INVX1_36 ( .A(u_sdrc_core_r2b_raddr_9_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n264_1) );
  INVX1 INVX1_360 ( .A(u_sdrc_core_u_req_gen__abc_22171_n850), .Y(u_sdrc_core_u_req_gen_map_address_24_) );
  INVX1 INVX1_361 ( .A(u_sdrc_core_u_req_gen__abc_22171_n857), .Y(u_sdrc_core_u_req_gen__abc_22171_n858) );
  INVX1 INVX1_362 ( .A(u_sdrc_core_u_req_gen_curr_sdr_addr_25_), .Y(u_sdrc_core_u_req_gen__abc_22171_n859) );
  INVX1 INVX1_363 ( .A(u_sdrc_core_u_req_gen__abc_22171_n863), .Y(u_sdrc_core_u_req_gen__abc_22171_n865) );
  INVX1 INVX1_364 ( .A(u_sdrc_core_u_req_gen__abc_22171_n869), .Y(u_sdrc_core_u_req_gen_map_address_25_) );
  INVX1 INVX1_365 ( .A(\cfg_colbits[0] ), .Y(u_sdrc_core_u_req_gen__abc_22171_n873) );
  INVX1 INVX1_366 ( .A(u_sdrc_core_u_req_gen__abc_22171_n874), .Y(u_sdrc_core_u_req_gen__abc_22171_n886) );
  INVX1 INVX1_367 ( .A(u_sdrc_core_u_req_gen__abc_22171_n879), .Y(u_sdrc_core_u_req_gen__abc_22171_n887) );
  INVX1 INVX1_368 ( .A(u_sdrc_core_u_req_gen__abc_22171_n888), .Y(u_sdrc_core_u_req_gen__abc_22171_n980) );
  INVX1 INVX1_369 ( .A(u_sdrc_core_u_req_gen__abc_22171_n983), .Y(u_sdrc_core_u_req_gen__abc_22171_n984) );
  INVX1 INVX1_37 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_9_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n267_1) );
  INVX1 INVX1_370 ( .A(u_sdrc_core_u_req_gen__abc_22171_n993), .Y(u_sdrc_core_u_req_gen__abc_22171_n994) );
  INVX1 INVX1_371 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1001), .Y(u_sdrc_core_u_req_gen__abc_22171_n1002) );
  INVX1 INVX1_372 ( .A(app_req), .Y(u_sdrc_core_u_req_gen__abc_22171_n1005) );
  INVX1 INVX1_373 ( .A(u_sdrc_core_u_req_gen__abc_22171_n596), .Y(u_sdrc_core_u_req_gen__abc_22171_n1009) );
  INVX1 INVX1_374 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1010), .Y(u_sdrc_core_u_req_gen__abc_22171_n1011) );
  INVX1 INVX1_375 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1018), .Y(u_sdrc_core_u_req_gen__abc_22171_n1019) );
  INVX1 INVX1_376 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1020), .Y(u_sdrc_core_u_req_gen__abc_22171_n1021) );
  INVX1 INVX1_377 ( .A(u_sdrc_core_u_req_gen__abc_22171_n397), .Y(u_sdrc_core_u_req_gen__abc_22171_n1023) );
  INVX1 INVX1_378 ( .A(u_sdrc_core_u_req_gen__abc_22171_n363), .Y(u_sdrc_core_u_req_gen__abc_22171_n1029) );
  INVX1 INVX1_379 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1035), .Y(u_sdrc_core_u_req_gen__abc_22171_n1036) );
  INVX1 INVX1_38 ( .A(u_sdrc_core_r2b_raddr_7_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n269) );
  INVX1 INVX1_380 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1024), .Y(u_sdrc_core_u_req_gen__abc_22171_n1042) );
  INVX1 INVX1_381 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1026), .Y(u_sdrc_core_u_req_gen__abc_22171_n1044) );
  INVX1 INVX1_382 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1033), .Y(u_sdrc_core_u_req_gen__abc_22171_n1045) );
  INVX1 INVX1_383 ( .A(u_sdrc_core_u_req_gen__abc_22171_n301), .Y(u_sdrc_core_u_req_gen__abc_22171_n1052) );
  INVX1 INVX1_384 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1013), .Y(u_sdrc_core_u_req_gen__abc_22171_n1062) );
  INVX1 INVX1_385 ( .A(u_sdrc_core_u_req_gen__abc_22171_n611), .Y(u_sdrc_core_u_req_gen__abc_22171_n1064) );
  INVX1 INVX1_386 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1065), .Y(u_sdrc_core_u_req_gen__abc_22171_n1067) );
  INVX1 INVX1_387 ( .A(u_sdrc_core_u_req_gen__abc_22171_n631), .Y(u_sdrc_core_u_req_gen__abc_22171_n1078) );
  INVX1 INVX1_388 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1082), .Y(u_sdrc_core_u_req_gen__abc_22171_n1083) );
  INVX1 INVX1_389 ( .A(u_sdrc_core_r2b_wrap), .Y(u_sdrc_core_u_req_gen__abc_22171_n1087) );
  INVX1 INVX1_39 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_7_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n274_1) );
  INVX1 INVX1_390 ( .A(u_sdrc_core_u_req_gen__abc_22171_n644), .Y(u_sdrc_core_u_req_gen__abc_22171_n1089) );
  INVX1 INVX1_391 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1091), .Y(u_sdrc_core_u_req_gen__abc_22171_n1092) );
  INVX1 INVX1_392 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1066), .Y(u_sdrc_core_u_req_gen__abc_22171_n1094) );
  INVX1 INVX1_393 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1095), .Y(u_sdrc_core_u_req_gen__abc_22171_n1096) );
  INVX1 INVX1_394 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n353_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n354) );
  INVX1 INVX1_395 ( .A(u_sdrc_core_u_xfr_ctl_cntr1_3_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n355) );
  INVX1 INVX1_396 ( .A(u_sdrc_core_u_xfr_ctl_cntr1_2_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n356_1) );
  INVX1 INVX1_397 ( .A(u_sdrc_core_u_xfr_ctl_cntr1_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n357) );
  INVX1 INVX1_398 ( .A(u_sdrc_core_u_xfr_ctl_cntr1_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n358_1) );
  INVX1 INVX1_399 ( .A(u_sdrc_core_u_xfr_ctl_rfsh_row_cnt_2_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n366) );
  INVX1 INVX1_4 ( .A(u_sdrc_core_u_bank_ctl_rank_cnt_1_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n218_1) );
  INVX1 INVX1_40 ( .A(u_sdrc_core_r2b_raddr_3_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n276_1) );
  INVX1 INVX1_400 ( .A(u_sdrc_core_u_xfr_ctl_rfsh_row_cnt_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n368) );
  INVX1 INVX1_401 ( .A(u_sdrc_core_u_xfr_ctl_rfsh_row_cnt_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n370) );
  INVX1 INVX1_402 ( .A(u_sdrc_core_u_xfr_ctl_xfr_st_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n385) );
  INVX1 INVX1_403 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n386), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n387_1) );
  INVX1 INVX1_404 ( .A(u_sdrc_core_u_xfr_ctl_xfr_st_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n388) );
  INVX1 INVX1_405 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n389_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n390) );
  INVX1 INVX1_406 ( .A(u_sdrc_core_u_xfr_ctl_mgmt_st_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n392) );
  INVX1 INVX1_407 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n394), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n395) );
  INVX1 INVX1_408 ( .A(u_sdrc_core_u_xfr_ctl_mgmt_st_4_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n396_1) );
  INVX1 INVX1_409 ( .A(u_sdrc_core_u_xfr_ctl_mgmt_st_6_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n397) );
  INVX1 INVX1_41 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_6_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n279_1) );
  INVX1 INVX1_410 ( .A(u_sdrc_core_u_xfr_ctl_mgmt_st_5_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n398_1) );
  INVX1 INVX1_411 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n400_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n401_1) );
  INVX1 INVX1_412 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n361), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n408_1) );
  INVX1 INVX1_413 ( .A(cfg_sdr_en), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n414_1) );
  INVX1 INVX1_414 ( .A(_auto_iopadmap_cc_313_execute_24701), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n424) );
  INVX1 INVX1_415 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n430), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n431) );
  INVX1 INVX1_416 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n377_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n433) );
  INVX1 INVX1_417 ( .A(u_sdrc_core_u_xfr_ctl_l_len_4_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n447) );
  INVX1 INVX1_418 ( .A(u_sdrc_core_u_xfr_ctl_l_len_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n448_1) );
  INVX1 INVX1_419 ( .A(u_sdrc_core_u_xfr_ctl_l_len_3_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n450_1) );
  INVX1 INVX1_42 ( .A(u_sdrc_core_r2b_raddr_6_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n281) );
  INVX1 INVX1_420 ( .A(u_sdrc_core_u_xfr_ctl_l_len_2_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n451_1) );
  INVX1 INVX1_421 ( .A(u_sdrc_core_u_xfr_ctl_l_len_6_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n454_1) );
  INVX1 INVX1_422 ( .A(u_sdrc_core_u_xfr_ctl_l_len_5_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n455_1) );
  INVX1 INVX1_423 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n459_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n460_1) );
  INVX1 INVX1_424 ( .A(u_sdrc_core_b2x_cmd_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n461_1) );
  INVX1 INVX1_425 ( .A(u_sdrc_core_u_xfr_ctl_l_wrap), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n462_1) );
  INVX1 INVX1_426 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n463_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n464_1) );
  INVX1 INVX1_427 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n467_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n468_1) );
  INVX1 INVX1_428 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n469_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n470_1) );
  INVX1 INVX1_429 ( .A(u_sdrc_core_b2x_cmd_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n471_1) );
  INVX1 INVX1_43 ( .A(u_sdrc_core_r2b_raddr_5_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n285) );
  INVX1 INVX1_430 ( .A(u_sdrc_core_u_bank_ctl_xfr_bank_sel_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n473) );
  INVX1 INVX1_431 ( .A(u_sdrc_core_b2x_ba_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n474) );
  INVX1 INVX1_432 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n483), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n484_1) );
  INVX1 INVX1_433 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n458), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n491_1) );
  INVX1 INVX1_434 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n493_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n494_1) );
  INVX1 INVX1_435 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n445), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n505_1) );
  INVX1 INVX1_436 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n446_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n506_1) );
  INVX1 INVX1_437 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n465_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n507) );
  INVX1 INVX1_438 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n472), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n508) );
  INVX1 INVX1_439 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n476), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n510) );
  INVX1 INVX1_44 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_1_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n287_1) );
  INVX1 INVX1_440 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n486), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n517_1) );
  INVX1 INVX1_441 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n503), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n522) );
  INVX1 INVX1_442 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n524_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n525) );
  INVX1 INVX1_443 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n537), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n538) );
  INVX1 INVX1_444 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n543), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n544) );
  INVX1 INVX1_445 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n501_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n547) );
  INVX1 INVX1_446 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n548_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n549) );
  INVX1 INVX1_447 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n554_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n555) );
  INVX1 INVX1_448 ( .A(\cfg_sdr_cas[2] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n557_1) );
  INVX1 INVX1_449 ( .A(\cfg_sdr_cas[1] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n558_1) );
  INVX1 INVX1_45 ( .A(u_sdrc_core_r2b_raddr_0_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n290_1) );
  INVX1 INVX1_450 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n560_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n561) );
  INVX1 INVX1_451 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n562), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n563_1) );
  INVX1 INVX1_452 ( .A(\cfg_sdr_cas[0] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n564_1) );
  INVX1 INVX1_453 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n566_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n567) );
  INVX1 INVX1_454 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n571), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n572_1) );
  INVX1 INVX1_455 ( .A(u_sdrc_core_u_xfr_ctl_xfr_caddr_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n597) );
  INVX1 INVX1_456 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n552_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n598) );
  INVX1 INVX1_457 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n550), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n599_1) );
  INVX1 INVX1_458 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n593_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n603_1) );
  INVX1 INVX1_459 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n492_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n619) );
  INVX1 INVX1_46 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_0_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n292_1) );
  INVX1 INVX1_460 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n629), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n630_1) );
  INVX1 INVX1_461 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n640), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n641_1) );
  INVX1 INVX1_462 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n651), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n652_1) );
  INVX1 INVX1_463 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n662), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n663) );
  INVX1 INVX1_464 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n673), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n674) );
  INVX1 INVX1_465 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n684_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n685_1) );
  INVX1 INVX1_466 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n695_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n696_1) );
  INVX1 INVX1_467 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n706), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n707_1) );
  INVX1 INVX1_468 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n717), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n718_1) );
  INVX1 INVX1_469 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n728), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n729) );
  INVX1 INVX1_47 ( .A(u_sdrc_core_r2b_raddr_10_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n299_1) );
  INVX1 INVX1_470 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n740_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n741) );
  INVX1 INVX1_471 ( .A(u_sdrc_core_u_xfr_ctl_l_len_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n773) );
  INVX1 INVX1_472 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n780), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n787) );
  INVX1 INVX1_473 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n786), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n795) );
  INVX1 INVX1_474 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n794_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n803_1) );
  INVX1 INVX1_475 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n802), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n811_1) );
  INVX1 INVX1_476 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n810_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n819_1) );
  INVX1 INVX1_477 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n606_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n826_1) );
  INVX1 INVX1_478 ( .A(u_sdrc_core_b2x_len_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n846_1) );
  INVX1 INVX1_479 ( .A(u_sdrc_core_b2x_len_2_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n847_1) );
  INVX1 INVX1_48 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_10_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n300_1) );
  INVX1 INVX1_480 ( .A(u_sdrc_core_b2x_len_3_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n852_1) );
  INVX1 INVX1_481 ( .A(u_sdrc_core_b2x_len_4_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n853) );
  INVX1 INVX1_482 ( .A(u_sdrc_core_b2x_len_5_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n856_1) );
  INVX1 INVX1_483 ( .A(u_sdrc_core_b2x_len_6_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n857_1) );
  INVX1 INVX1_484 ( .A(u_sdrc_core_u_xfr_ctl_mgmt_st_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n871_1) );
  INVX1 INVX1_485 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n873), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n874) );
  INVX1 INVX1_486 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n500_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n875) );
  INVX1 INVX1_487 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n876), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n877) );
  INVX1 INVX1_488 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n888), .Y(u_sdrc_core_u_xfr_ctl_sdr_ras_n_FF_INPUT) );
  INVX1 INVX1_489 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n577), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n895) );
  INVX1 INVX1_49 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_8_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n304_1) );
  INVX1 INVX1_490 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n527), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n905) );
  INVX1 INVX1_491 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n912), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1013) );
  INVX1 INVX1_492 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1041), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1045) );
  INVX1 INVX1_493 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1042), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1047) );
  INVX1 INVX1_494 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1040), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1052) );
  INVX1 INVX1_495 ( .A(u_sdrc_core_u_xfr_ctl_tmr0_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1053) );
  INVX1 INVX1_496 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n351_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1058) );
  INVX1 INVX1_497 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n352), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1071) );
  INVX1 INVX1_498 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1091), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1092) );
  INVX1 INVX1_499 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n539_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1093) );
  INVX1 INVX1_5 ( .A(u_sdrc_core_b2r_ack), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n239_1) );
  INVX1 INVX1_50 ( .A(u_sdrc_core_r2b_raddr_8_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n305) );
  INVX1 INVX1_500 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1095), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1105) );
  INVX1 INVX1_501 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1107), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1115) );
  INVX1 INVX1_502 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1117), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1125) );
  INVX1 INVX1_503 ( .A(u_sdrc_core_u_xfr_ctl_rfsh_timer_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1132) );
  INVX1 INVX1_504 ( .A(\cfg_sdr_rfsh[5] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1133) );
  INVX1 INVX1_505 ( .A(u_sdrc_core_u_xfr_ctl_rfsh_timer_5_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1135) );
  INVX1 INVX1_506 ( .A(\cfg_sdr_rfsh[4] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1138) );
  INVX1 INVX1_507 ( .A(u_sdrc_core_u_xfr_ctl_rfsh_timer_4_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1140) );
  INVX1 INVX1_508 ( .A(\cfg_sdr_rfsh[7] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1144) );
  INVX1 INVX1_509 ( .A(u_sdrc_core_u_xfr_ctl_rfsh_timer_7_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1146) );
  INVX1 INVX1_51 ( .A(u_sdrc_core_r2b_raddr_2_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n309) );
  INVX1 INVX1_510 ( .A(\cfg_sdr_rfsh[11] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1150) );
  INVX1 INVX1_511 ( .A(u_sdrc_core_u_xfr_ctl_rfsh_timer_11_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1152) );
  INVX1 INVX1_512 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1156), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1157) );
  INVX1 INVX1_513 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1158), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1159) );
  INVX1 INVX1_514 ( .A(\cfg_sdr_rfsh[8] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1161) );
  INVX1 INVX1_515 ( .A(u_sdrc_core_u_xfr_ctl_rfsh_timer_8_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1162) );
  INVX1 INVX1_516 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1169), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1170) );
  INVX1 INVX1_517 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1171), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1172) );
  INVX1 INVX1_518 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1174), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1175) );
  INVX1 INVX1_519 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1176), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1177) );
  INVX1 INVX1_52 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_3_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n311_1) );
  INVX1 INVX1_520 ( .A(\cfg_sdr_rfsh[0] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1179) );
  INVX1 INVX1_521 ( .A(\cfg_sdr_rfsh[2] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1184) );
  INVX1 INVX1_522 ( .A(u_sdrc_core_u_xfr_ctl_rfsh_timer_2_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1186) );
  INVX1 INVX1_523 ( .A(\cfg_sdr_rfsh[10] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1190) );
  INVX1 INVX1_524 ( .A(u_sdrc_core_u_xfr_ctl_rfsh_timer_10_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1191) );
  INVX1 INVX1_525 ( .A(\cfg_sdr_rfsh[6] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1195) );
  INVX1 INVX1_526 ( .A(u_sdrc_core_u_xfr_ctl_rfsh_timer_6_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1196) );
  INVX1 INVX1_527 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1202), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1203) );
  INVX1 INVX1_528 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1207), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1208) );
  INVX1 INVX1_529 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1212), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1213) );
  INVX1 INVX1_53 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_2_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n314_1) );
  INVX1 INVX1_530 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1217), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1218) );
  INVX1 INVX1_531 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1222), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1223) );
  INVX1 INVX1_532 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1227), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1228) );
  INVX1 INVX1_533 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1232), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1233) );
  INVX1 INVX1_534 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1236), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1237) );
  INVX1 INVX1_535 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1241), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1242) );
  INVX1 INVX1_536 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1246), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1247) );
  INVX1 INVX1_537 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1251), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1252) );
  INVX1 INVX1_538 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1260), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1261) );
  INVX1 INVX1_539 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1265), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1266) );
  INVX1 INVX1_54 ( .A(u_sdrc_core_r2b_raddr_1_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n316_1) );
  INVX1 INVX1_540 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1270), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1271) );
  INVX1 INVX1_541 ( .A(u_sdrc_core_u_xfr_ctl_act_cmd), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1374) );
  INVX1 INVX1_542 ( .A(u_sdrc_core_u_xfr_ctl_d_act_cmd), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1375) );
  INVX1 INVX1_543 ( .A(u_wb2sdrc_cmdfifo_empty), .Y(app_req) );
  INVX1 INVX1_544 ( .A(u_wb2sdrc_cmdfifo_full), .Y(u_wb2sdrc__abc_24125_n28_1) );
  INVX1 INVX1_545 ( .A(u_wb2sdrc_u_wrdatafifo_full), .Y(u_wb2sdrc__abc_24125_n31) );
  INVX1 INVX1_546 ( .A(u_wb2sdrc__abc_24125_n29_1), .Y(u_wb2sdrc__abc_24125_n34) );
  INVX1 INVX1_547 ( .A(u_wb2sdrc_pending_read), .Y(u_wb2sdrc__abc_24125_n39_1) );
  INVX1 INVX1_548 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n400_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n401_1) );
  INVX1 INVX1_549 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n402), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n403_1) );
  INVX1 INVX1_55 ( .A(u_sdrc_core_r2b_raddr_4_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n320_1) );
  INVX1 INVX1_550 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n404_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n405) );
  INVX1 INVX1_551 ( .A(u_wb2sdrc_u_cmdfifo_wr_ptr_0_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n406_1) );
  INVX1 INVX1_552 ( .A(u_wb2sdrc_u_cmdfifo_sync_rd_ptr_1_0_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n408) );
  INVX1 INVX1_553 ( .A(u_wb2sdrc_u_cmdfifo_wr_ptr_1_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n412_1) );
  INVX1 INVX1_554 ( .A(u_wb2sdrc_u_cmdfifo_sync_rd_ptr_2_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n417) );
  INVX1 INVX1_555 ( .A(u_wb2sdrc_u_cmdfifo_wr_ptr_2_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n418_1) );
  INVX1 INVX1_556 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n421_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n422_1) );
  INVX1 INVX1_557 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n416_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n424_1) );
  INVX1 INVX1_558 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n407_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n427_1) );
  INVX1 INVX1_559 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n409_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n428_1) );
  INVX1 INVX1_56 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_4_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n322_1) );
  INVX1 INVX1_560 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n414), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n430_1) );
  INVX1 INVX1_561 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n438), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n439_1) );
  INVX1 INVX1_562 ( .A(u_wb2sdrc_u_cmdfifo_sync_wr_ptr_1_1_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n443_1) );
  INVX1 INVX1_563 ( .A(u_wb2sdrc_u_cmdfifo_sync_wr_ptr_2_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n444) );
  INVX1 INVX1_564 ( .A(u_wb2sdrc_u_cmdfifo_sync_wr_ptr_1_0_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n448_1) );
  INVX1 INVX1_565 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n453), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n454_1) );
  INVX1 INVX1_566 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_2_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n458_1) );
  INVX1 INVX1_567 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n441), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n462_1) );
  INVX1 INVX1_568 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n460_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n469_1) );
  INVX1 INVX1_569 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n596), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n597) );
  INVX1 INVX1_57 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_5_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n325) );
  INVX1 INVX1_570 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n595), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n603) );
  INVX1 INVX1_571 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n475_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n619) );
  INVX1 INVX1_572 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n635), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n636) );
  INVX1 INVX1_573 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n644), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n645) );
  INVX1 INVX1_574 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n426), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n654) );
  INVX1 INVX1_575 ( .A(u_wb2sdrc_u_rddatafifo_wr_ptr_0_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n375_1) );
  INVX1 INVX1_576 ( .A(u_wb2sdrc_u_rddatafifo_wr_ptr_1_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n384_1) );
  INVX1 INVX1_577 ( .A(u_wb2sdrc_u_rddatafifo_wr_ptr_2_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n389) );
  INVX1 INVX1_578 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n411_1), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n412_1) );
  INVX1 INVX1_579 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n413), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n415_1) );
  INVX1 INVX1_58 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n331_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n332_1) );
  INVX1 INVX1_580 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n417), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n418) );
  INVX1 INVX1_581 ( .A(u_wb2sdrc_u_rddatafifo_sync_wr_ptr_1_0_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n421) );
  INVX1 INVX1_582 ( .A(u_wb2sdrc_u_rddatafifo_sync_wr_ptr_2_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n426) );
  INVX1 INVX1_583 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_2_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n428_1) );
  INVX1 INVX1_584 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n431_1), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n432_1) );
  INVX1 INVX1_585 ( .A(u_wb2sdrc_rddatafifo_rd), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1119) );
  INVX1 INVX1_586 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1130), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1131) );
  INVX1 INVX1_587 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1156), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1157) );
  INVX1 INVX1_588 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1155), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1163) );
  INVX1 INVX1_589 ( .A(u_wb2sdrc_u_wrdatafifo_sync_rd_ptr_1_2_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n696_1) );
  INVX1 INVX1_59 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_refresh), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n336) );
  INVX1 INVX1_590 ( .A(u_wb2sdrc_u_wrdatafifo_sync_rd_ptr_1_3_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n697_1) );
  INVX1 INVX1_591 ( .A(u_wb2sdrc_u_wrdatafifo_sync_rd_ptr_1_1_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n702_1) );
  INVX1 INVX1_592 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n699_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n704_1) );
  INVX1 INVX1_593 ( .A(u_wb2sdrc_u_wrdatafifo_sync_rd_ptr_1_0_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n710) );
  INVX1 INVX1_594 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n712), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n716_1) );
  INVX1 INVX1_595 ( .A(u_wb2sdrc_u_wrdatafifo_wr_ptr_2_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n724) );
  INVX1 INVX1_596 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n726_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n727) );
  INVX1 INVX1_597 ( .A(u_wb2sdrc_u_wrdatafifo_wr_ptr_3_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n731) );
  INVX1 INVX1_598 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n733_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n734) );
  INVX1 INVX1_599 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n701), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n736) );
  INVX1 INVX1_6 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n243), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n244_1) );
  INVX1 INVX1_60 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_l_sdr_dma_last), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n353_1) );
  INVX1 INVX1_600 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n709_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n737) );
  INVX1 INVX1_601 ( .A(u_wb2sdrc_u_wrdatafifo_wr_ptr_0_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n738_1) );
  INVX1 INVX1_602 ( .A(u_wb2sdrc_u_wrdatafifo_wr_ptr_1_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n743) );
  INVX1 INVX1_603 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n754), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n757_1) );
  INVX1 INVX1_604 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_3_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n792_1) );
  INVX1 INVX1_605 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2286), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2287) );
  INVX1 INVX1_606 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2290), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2291) );
  INVX1 INVX1_607 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2294), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2310) );
  INVX1 INVX1_608 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n753_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2319) );
  INVX1 INVX1_609 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2328), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2329) );
  INVX1 INVX1_61 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n250_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n355) );
  INVX1 INVX1_610 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2334), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2335) );
  INVX1 INVX1_611 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2342), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2343) );
  INVX1 INVX1_62 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_prech_page_closed), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n356) );
  INVX1 INVX1_63 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n357), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n358_1) );
  INVX1 INVX1_64 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_r2b_req), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n360) );
  INVX1 INVX1_65 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_4_bF_buf1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n367) );
  INVX1 INVX1_66 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n368_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n369_1) );
  INVX1 INVX1_67 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_tras_cntr_0_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n379_1) );
  INVX1 INVX1_68 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n380), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n381) );
  INVX1 INVX1_69 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n382), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n383_1) );
  INVX1 INVX1_7 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n245_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n246_1) );
  INVX1 INVX1_70 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n384_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n393) );
  INVX1 INVX1_71 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n385), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n400_1) );
  INVX1 INVX1_72 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_timer0_0_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n413_1) );
  INVX1 INVX1_73 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n424), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n425) );
  INVX1 INVX1_74 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n437_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n438_1) );
  INVX1 INVX1_75 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_l_write), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n730) );
  INVX1 INVX1_76 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n428_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n742) );
  INVX1 INVX1_77 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n386_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n745) );
  INVX1 INVX1_78 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_x2b_ack), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n249_1) );
  INVX1 INVX1_79 ( .A(u_sdrc_core_r2b_raddr_12_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n254) );
  INVX1 INVX1_8 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n242_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n252_1) );
  INVX1 INVX1_80 ( .A(u_sdrc_core_r2b_raddr_11_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n256_1) );
  INVX1 INVX1_81 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_12_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n258_1) );
  INVX1 INVX1_82 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_11_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n262_1) );
  INVX1 INVX1_83 ( .A(u_sdrc_core_r2b_raddr_9_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n264_1) );
  INVX1 INVX1_84 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_9_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n267_1) );
  INVX1 INVX1_85 ( .A(u_sdrc_core_r2b_raddr_7_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n269) );
  INVX1 INVX1_86 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_7_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n274_1) );
  INVX1 INVX1_87 ( .A(u_sdrc_core_r2b_raddr_3_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n276_1) );
  INVX1 INVX1_88 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_6_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n279_1) );
  INVX1 INVX1_89 ( .A(u_sdrc_core_r2b_raddr_6_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n281) );
  INVX1 INVX1_9 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n253_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n254_1) );
  INVX1 INVX1_90 ( .A(u_sdrc_core_r2b_raddr_5_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n285) );
  INVX1 INVX1_91 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_1_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n287_1) );
  INVX1 INVX1_92 ( .A(u_sdrc_core_r2b_raddr_0_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n290_1) );
  INVX1 INVX1_93 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_0_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n292_1) );
  INVX1 INVX1_94 ( .A(u_sdrc_core_r2b_raddr_10_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n299_1) );
  INVX1 INVX1_95 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_10_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n300_1) );
  INVX1 INVX1_96 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_8_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n304_1) );
  INVX1 INVX1_97 ( .A(u_sdrc_core_r2b_raddr_8_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n305) );
  INVX1 INVX1_98 ( .A(u_sdrc_core_r2b_raddr_2_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n309) );
  INVX1 INVX1_99 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_3_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n311_1) );
  INVX2 INVX2_1 ( .A(u_sdrc_core_u_bank_ctl_rank_cnt_2_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n216_1) );
  INVX2 INVX2_10 ( .A(u_sdrc_core_u_req_gen__abc_22171_n242_bF_buf4), .Y(u_sdrc_core_u_req_gen__abc_22171_n391) );
  INVX2 INVX2_11 ( .A(u_sdrc_core_u_req_gen__abc_22171_n245_1_bF_buf0), .Y(u_sdrc_core_u_req_gen__abc_22171_n416) );
  INVX2 INVX2_12 ( .A(u_sdrc_core_u_xfr_ctl_mgmt_st_2_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n393_1) );
  INVX2 INVX2_13 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n403_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n444_1) );
  INVX2 INVX2_14 ( .A(wb_we_i), .Y(u_wb2sdrc_u_cmdfifo_wr_data_26_) );
  INVX2 INVX2_15 ( .A(u_wb2sdrc__abc_24125_n36_1), .Y(u_wb2sdrc_rddatafifo_rd) );
  INVX2 INVX2_16 ( .A(\wb_sel_i[0] ), .Y(u_wb2sdrc_u_wrdatafifo_wr_data_32_) );
  INVX2 INVX2_17 ( .A(\wb_sel_i[1] ), .Y(u_wb2sdrc_u_wrdatafifo_wr_data_33_) );
  INVX2 INVX2_18 ( .A(\wb_sel_i[2] ), .Y(u_wb2sdrc_u_wrdatafifo_wr_data_34_) );
  INVX2 INVX2_19 ( .A(\wb_sel_i[3] ), .Y(u_wb2sdrc_u_wrdatafifo_wr_data_35_) );
  INVX2 INVX2_2 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n411_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n412_1) );
  INVX2 INVX2_20 ( .A(app_req_ack_bF_buf6), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n590) );
  INVX2 INVX2_21 ( .A(u_wb2sdrc_cmdfifo_wr), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n624) );
  INVX2 INVX2_22 ( .A(app_rd_valid), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1151) );
  INVX2 INVX2_23 ( .A(app_wr_next_req), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2279) );
  INVX2 INVX2_24 ( .A(u_wb2sdrc_u_wrdatafifo_wr_en), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2323) );
  INVX2 INVX2_3 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n411_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n412_1) );
  INVX2 INVX2_4 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n411_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n412_1) );
  INVX2 INVX2_5 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n411_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n412_1) );
  INVX2 INVX2_6 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf3), .Y(u_sdrc_core_u_bs_convert__abc_21684_n175_1) );
  INVX2 INVX2_7 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n508), .Y(u_sdrc_core_u_bs_convert__abc_21684_n510) );
  INVX2 INVX2_8 ( .A(u_sdrc_core_u_req_gen__abc_22171_n222), .Y(u_sdrc_core_r2b_len_3_) );
  INVX2 INVX2_9 ( .A(cfg_sdr_width_1_bF_buf1), .Y(u_sdrc_core_u_req_gen__abc_22171_n241) );
  INVX4 INVX4_1 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_xfr_ok_bF_buf3), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n227) );
  INVX4 INVX4_10 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n184_1_bF_buf5), .Y(u_sdrc_core_u_bs_convert__abc_21684_n185_1) );
  INVX4 INVX4_11 ( .A(u_sdrc_core_u_bs_convert_x2a_rdok), .Y(u_sdrc_core_u_bs_convert__abc_21684_n542) );
  INVX4 INVX4_12 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n545), .Y(u_sdrc_core_u_bs_convert__abc_21684_n546) );
  INVX4 INVX4_13 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n579), .Y(u_sdrc_core_u_bs_convert__abc_21684_n580) );
  INVX4 INVX4_14 ( .A(u_sdrc_core_u_req_gen__abc_22171_n216_1), .Y(u_sdrc_core_r2b_len_2_) );
  INVX4 INVX4_15 ( .A(u_sdrc_core_u_req_gen__abc_22171_n335_1_bF_buf2), .Y(u_sdrc_core_u_req_gen__abc_22171_n346_1) );
  INVX4 INVX4_16 ( .A(\cfg_colbits[1] ), .Y(u_sdrc_core_u_req_gen__abc_22171_n876) );
  INVX4 INVX4_17 ( .A(u_sdrc_core_u_req_gen__abc_22171_n877), .Y(u_sdrc_core_u_req_gen__abc_22171_n893) );
  INVX4 INVX4_18 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n404_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n405_1) );
  INVX4 INVX4_19 ( .A(sdram_resetn_bF_buf18), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n413_1) );
  INVX4 INVX4_2 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_2_bF_buf0), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n366) );
  INVX4 INVX4_20 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n607), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n610_1) );
  INVX4 INVX4_21 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n883_bF_buf1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n911) );
  INVX4 INVX4_3 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_0_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n685) );
  INVX4 INVX4_4 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_2_bF_buf0), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n366) );
  INVX4 INVX4_5 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_0_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n685) );
  INVX4 INVX4_6 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_2_bF_buf0), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n366) );
  INVX4 INVX4_7 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_0_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n685) );
  INVX4 INVX4_8 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_2_bF_buf0), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n366) );
  INVX4 INVX4_9 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_0_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n685) );
  INVX8 INVX8_1 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf2), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n283) );
  INVX8 INVX8_10 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf7), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1) );
  INVX8 INVX8_11 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf4), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1) );
  INVX8 INVX8_12 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n981_bF_buf5), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n982) );
  INVX8 INVX8_13 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf3), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1092) );
  INVX8 INVX8_14 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf3), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1201) );
  INVX8 INVX8_15 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_1_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n409) );
  INVX8 INVX8_16 ( .A(u_wb2sdrc_u_rddatafifo_rd_ptr_0_bF_buf5), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1) );
  INVX8 INVX8_17 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n447_1_bF_buf3), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n449) );
  INVX8 INVX8_18 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf3), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n551) );
  INVX8 INVX8_19 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf3), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n652) );
  INVX8 INVX8_2 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf2), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n457_1) );
  INVX8 INVX8_20 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf3), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1020) );
  INVX8 INVX8_21 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_0_bF_buf7), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n764_1) );
  INVX8 INVX8_22 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_1_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n782) );
  INVX8 INVX8_23 ( .A(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf5), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1) );
  INVX8 INVX8_24 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf4), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1) );
  INVX8 INVX8_25 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf4), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1) );
  INVX8 INVX8_26 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf4), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1) );
  INVX8 INVX8_27 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf4), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841) );
  INVX8 INVX8_28 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf4), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951) );
  INVX8 INVX8_29 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf4), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061) );
  INVX8 INVX8_3 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf2), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n457_1) );
  INVX8 INVX8_30 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf4), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171) );
  INVX8 INVX8_31 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2362_bF_buf5), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2363) );
  INVX8 INVX8_4 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf2), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n457_1) );
  INVX8 INVX8_5 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf2), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n457_1) );
  INVX8 INVX8_6 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n170_1_bF_buf3), .Y(u_sdrc_core_u_bs_convert__abc_21684_n171_1) );
  INVX8 INVX8_7 ( .A(app_req_ack_bF_buf4), .Y(u_sdrc_core_u_req_gen__abc_22171_n318) );
  INVX8 INVX8_8 ( .A(wb_rst_i), .Y(u_wb2sdrc_u_cmdfifo_wr_reset_n) );
  INVX8 INVX8_9 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_1_bF_buf5), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n436_1) );
  OR2X2 OR2X2_1 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2r_ack_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_b2r_ack_bF_buf4), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n207_1) );
  OR2X2 OR2X2_10 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n232_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n233_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n234) );
  OR2X2 OR2X2_100 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_9_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n452) );
  OR2X2 OR2X2_1000 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n579), .B(u_sdrc_core_pad_sdr_din2_0_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n582) );
  OR2X2 OR2X2_1001 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n453), .B(u_sdrc_core_u_bs_convert__abc_21684_n542), .Y(u_sdrc_core_u_bs_convert__abc_21684_n585) );
  OR2X2 OR2X2_1002 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n584), .B(u_sdrc_core_u_bs_convert__abc_21684_n585), .Y(u_sdrc_core_u_bs_convert__abc_21684_n586) );
  OR2X2 OR2X2_1003 ( .A(u_sdrc_core_u_bs_convert_saved_rd_data_8_), .B(u_sdrc_core_u_bs_convert_x2a_rdok), .Y(u_sdrc_core_u_bs_convert__abc_21684_n587) );
  OR2X2 OR2X2_1004 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n580), .B(u_sdrc_core_u_bs_convert_saved_rd_data_9_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n590) );
  OR2X2 OR2X2_1005 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n579), .B(u_sdrc_core_pad_sdr_din2_1_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n591) );
  OR2X2 OR2X2_1006 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n456), .B(u_sdrc_core_u_bs_convert__abc_21684_n542), .Y(u_sdrc_core_u_bs_convert__abc_21684_n594) );
  OR2X2 OR2X2_1007 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n593), .B(u_sdrc_core_u_bs_convert__abc_21684_n594), .Y(u_sdrc_core_u_bs_convert__abc_21684_n595) );
  OR2X2 OR2X2_1008 ( .A(u_sdrc_core_u_bs_convert_saved_rd_data_9_), .B(u_sdrc_core_u_bs_convert_x2a_rdok), .Y(u_sdrc_core_u_bs_convert__abc_21684_n596) );
  OR2X2 OR2X2_1009 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n580), .B(u_sdrc_core_u_bs_convert_saved_rd_data_10_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n599) );
  OR2X2 OR2X2_101 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n223_1_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_9_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n453) );
  OR2X2 OR2X2_1010 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n579), .B(u_sdrc_core_pad_sdr_din2_2_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n600) );
  OR2X2 OR2X2_1011 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n459), .B(u_sdrc_core_u_bs_convert__abc_21684_n542), .Y(u_sdrc_core_u_bs_convert__abc_21684_n603) );
  OR2X2 OR2X2_1012 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n602), .B(u_sdrc_core_u_bs_convert__abc_21684_n603), .Y(u_sdrc_core_u_bs_convert__abc_21684_n604) );
  OR2X2 OR2X2_1013 ( .A(u_sdrc_core_u_bs_convert_saved_rd_data_10_), .B(u_sdrc_core_u_bs_convert_x2a_rdok), .Y(u_sdrc_core_u_bs_convert__abc_21684_n605) );
  OR2X2 OR2X2_1014 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n580), .B(u_sdrc_core_u_bs_convert_saved_rd_data_11_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n608) );
  OR2X2 OR2X2_1015 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n579), .B(u_sdrc_core_pad_sdr_din2_3_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n609) );
  OR2X2 OR2X2_1016 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n462), .B(u_sdrc_core_u_bs_convert__abc_21684_n542), .Y(u_sdrc_core_u_bs_convert__abc_21684_n612) );
  OR2X2 OR2X2_1017 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n611), .B(u_sdrc_core_u_bs_convert__abc_21684_n612), .Y(u_sdrc_core_u_bs_convert__abc_21684_n613) );
  OR2X2 OR2X2_1018 ( .A(u_sdrc_core_u_bs_convert_saved_rd_data_11_), .B(u_sdrc_core_u_bs_convert_x2a_rdok), .Y(u_sdrc_core_u_bs_convert__abc_21684_n614) );
  OR2X2 OR2X2_1019 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n580), .B(u_sdrc_core_u_bs_convert_saved_rd_data_12_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n617) );
  OR2X2 OR2X2_102 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n454), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf2), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n455) );
  OR2X2 OR2X2_1020 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n579), .B(u_sdrc_core_pad_sdr_din2_4_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n618) );
  OR2X2 OR2X2_1021 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n465), .B(u_sdrc_core_u_bs_convert__abc_21684_n542), .Y(u_sdrc_core_u_bs_convert__abc_21684_n621) );
  OR2X2 OR2X2_1022 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n620), .B(u_sdrc_core_u_bs_convert__abc_21684_n621), .Y(u_sdrc_core_u_bs_convert__abc_21684_n622) );
  OR2X2 OR2X2_1023 ( .A(u_sdrc_core_u_bs_convert_saved_rd_data_12_), .B(u_sdrc_core_u_bs_convert_x2a_rdok), .Y(u_sdrc_core_u_bs_convert__abc_21684_n623) );
  OR2X2 OR2X2_1024 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n580), .B(u_sdrc_core_u_bs_convert_saved_rd_data_13_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n626) );
  OR2X2 OR2X2_1025 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n579), .B(u_sdrc_core_pad_sdr_din2_5_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n627) );
  OR2X2 OR2X2_1026 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n468), .B(u_sdrc_core_u_bs_convert__abc_21684_n542), .Y(u_sdrc_core_u_bs_convert__abc_21684_n630) );
  OR2X2 OR2X2_1027 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n629), .B(u_sdrc_core_u_bs_convert__abc_21684_n630), .Y(u_sdrc_core_u_bs_convert__abc_21684_n631) );
  OR2X2 OR2X2_1028 ( .A(u_sdrc_core_u_bs_convert_saved_rd_data_13_), .B(u_sdrc_core_u_bs_convert_x2a_rdok), .Y(u_sdrc_core_u_bs_convert__abc_21684_n632) );
  OR2X2 OR2X2_1029 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n580), .B(u_sdrc_core_u_bs_convert_saved_rd_data_14_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n635) );
  OR2X2 OR2X2_103 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n283_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_9_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n456) );
  OR2X2 OR2X2_1030 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n579), .B(u_sdrc_core_pad_sdr_din2_6_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n636) );
  OR2X2 OR2X2_1031 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n471), .B(u_sdrc_core_u_bs_convert__abc_21684_n542), .Y(u_sdrc_core_u_bs_convert__abc_21684_n639) );
  OR2X2 OR2X2_1032 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n638), .B(u_sdrc_core_u_bs_convert__abc_21684_n639), .Y(u_sdrc_core_u_bs_convert__abc_21684_n640) );
  OR2X2 OR2X2_1033 ( .A(u_sdrc_core_u_bs_convert_saved_rd_data_14_), .B(u_sdrc_core_u_bs_convert_x2a_rdok), .Y(u_sdrc_core_u_bs_convert__abc_21684_n641) );
  OR2X2 OR2X2_1034 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n580), .B(u_sdrc_core_u_bs_convert_saved_rd_data_15_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n644) );
  OR2X2 OR2X2_1035 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n579), .B(u_sdrc_core_pad_sdr_din2_7_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n645) );
  OR2X2 OR2X2_1036 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n474), .B(u_sdrc_core_u_bs_convert__abc_21684_n542), .Y(u_sdrc_core_u_bs_convert__abc_21684_n648) );
  OR2X2 OR2X2_1037 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n647), .B(u_sdrc_core_u_bs_convert__abc_21684_n648), .Y(u_sdrc_core_u_bs_convert__abc_21684_n649) );
  OR2X2 OR2X2_1038 ( .A(u_sdrc_core_u_bs_convert_saved_rd_data_15_), .B(u_sdrc_core_u_bs_convert_x2a_rdok), .Y(u_sdrc_core_u_bs_convert__abc_21684_n650) );
  OR2X2 OR2X2_1039 ( .A(u_sdrc_core_u_req_gen__abc_22171_n183), .B(u_sdrc_core_u_req_gen__abc_22171_n186), .Y(u_sdrc_core_u_req_gen__abc_16238_n30) );
  OR2X2 OR2X2_104 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n458), .B(u_sdrc_core_u_bank_ctl__abc_21249_n451), .Y(u_sdrc_core_b2x_addr_9_) );
  OR2X2 OR2X2_1040 ( .A(u_sdrc_core_u_req_gen__abc_22171_n188), .B(u_sdrc_core_u_req_gen__abc_22171_n191), .Y(u_sdrc_core_u_req_gen__abc_16238_n38) );
  OR2X2 OR2X2_1041 ( .A(u_sdrc_core_u_req_gen__abc_22171_n198), .B(u_sdrc_core_u_req_gen__abc_22171_n197), .Y(u_sdrc_core_u_req_gen__abc_22171_n199) );
  OR2X2 OR2X2_1042 ( .A(u_sdrc_core_u_req_gen__abc_22171_n199), .B(u_sdrc_core_u_req_gen__abc_22171_n196), .Y(u_sdrc_core_u_req_gen__abc_22171_n200_1) );
  OR2X2 OR2X2_1043 ( .A(u_sdrc_core_u_req_gen__abc_22171_n200_1), .B(u_sdrc_core_u_req_gen__abc_22171_n194), .Y(u_sdrc_core_u_req_gen__abc_16238_n57) );
  OR2X2 OR2X2_1044 ( .A(u_sdrc_core_u_req_gen__abc_22171_n205), .B(u_sdrc_core_u_req_gen__abc_22171_n203), .Y(u_sdrc_core_r2b_len_0_) );
  OR2X2 OR2X2_1045 ( .A(u_sdrc_core_u_req_gen__abc_22171_n202), .B(u_sdrc_core_u_req_gen_lcl_req_len_1_), .Y(u_sdrc_core_u_req_gen__abc_22171_n207) );
  OR2X2 OR2X2_1046 ( .A(u_sdrc_core_u_req_gen__abc_22171_n213), .B(u_sdrc_core_u_req_gen__abc_22171_n215_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n216_1) );
  OR2X2 OR2X2_1047 ( .A(u_sdrc_core_u_req_gen__abc_22171_n219_1), .B(u_sdrc_core_u_req_gen__abc_22171_n221_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n222) );
  OR2X2 OR2X2_1048 ( .A(u_sdrc_core_u_req_gen__abc_22171_n202), .B(u_sdrc_core_u_req_gen_lcl_req_len_4_), .Y(u_sdrc_core_u_req_gen__abc_22171_n224) );
  OR2X2 OR2X2_1049 ( .A(u_sdrc_core_u_req_gen__abc_22171_n202), .B(u_sdrc_core_u_req_gen_lcl_req_len_5_), .Y(u_sdrc_core_u_req_gen__abc_22171_n229) );
  OR2X2 OR2X2_105 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_10_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n461) );
  OR2X2 OR2X2_1050 ( .A(u_sdrc_core_u_req_gen__abc_22171_n202), .B(u_sdrc_core_u_req_gen_lcl_req_len_6_), .Y(u_sdrc_core_u_req_gen__abc_22171_n234_1) );
  OR2X2 OR2X2_1051 ( .A(u_sdrc_core_u_req_gen__abc_22171_n247), .B(u_sdrc_core_u_req_gen__abc_22171_n246), .Y(u_sdrc_core_u_req_gen__abc_22171_n248) );
  OR2X2 OR2X2_1052 ( .A(u_sdrc_core_u_req_gen__abc_22171_n248), .B(u_sdrc_core_u_req_gen__abc_22171_n243_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n249) );
  OR2X2 OR2X2_1053 ( .A(u_sdrc_core_u_req_gen__abc_22171_n250), .B(u_sdrc_core_u_req_gen__abc_22171_n251), .Y(u_sdrc_core_u_req_gen__abc_22171_n252) );
  OR2X2 OR2X2_1054 ( .A(u_sdrc_core_u_req_gen__abc_22171_n260), .B(u_sdrc_core_u_req_gen__abc_22171_n258), .Y(u_sdrc_core_u_req_gen__abc_22171_n261) );
  OR2X2 OR2X2_1055 ( .A(u_sdrc_core_u_req_gen__abc_22171_n261), .B(u_sdrc_core_u_req_gen__abc_22171_n256_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n262_1) );
  OR2X2 OR2X2_1056 ( .A(u_sdrc_core_u_req_gen__abc_22171_n263_1), .B(u_sdrc_core_u_req_gen__abc_22171_n265), .Y(u_sdrc_core_u_req_gen__abc_22171_n266) );
  OR2X2 OR2X2_1057 ( .A(u_sdrc_core_u_req_gen__abc_22171_n272), .B(u_sdrc_core_u_req_gen__abc_22171_n271), .Y(u_sdrc_core_u_req_gen__abc_22171_n273_1) );
  OR2X2 OR2X2_1058 ( .A(u_sdrc_core_u_req_gen__abc_22171_n273_1), .B(u_sdrc_core_u_req_gen__abc_22171_n270), .Y(u_sdrc_core_u_req_gen__abc_22171_n274) );
  OR2X2 OR2X2_1059 ( .A(u_sdrc_core_u_req_gen__abc_22171_n263_1), .B(u_sdrc_core_u_req_gen__abc_22171_n274), .Y(u_sdrc_core_u_req_gen__abc_22171_n277_1) );
  OR2X2 OR2X2_106 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n223_1_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_10_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n462) );
  OR2X2 OR2X2_1060 ( .A(u_sdrc_core_u_req_gen__abc_22171_n283_1), .B(u_sdrc_core_u_req_gen__abc_22171_n282), .Y(u_sdrc_core_u_req_gen__abc_22171_n284) );
  OR2X2 OR2X2_1061 ( .A(u_sdrc_core_u_req_gen__abc_22171_n284), .B(u_sdrc_core_u_req_gen__abc_22171_n281_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n285) );
  OR2X2 OR2X2_1062 ( .A(u_sdrc_core_u_req_gen__abc_22171_n288), .B(u_sdrc_core_u_req_gen__abc_22171_n286), .Y(u_sdrc_core_u_req_gen__abc_22171_n289) );
  OR2X2 OR2X2_1063 ( .A(u_sdrc_core_u_req_gen__abc_22171_n295), .B(u_sdrc_core_u_req_gen__abc_22171_n294_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n296_1) );
  OR2X2 OR2X2_1064 ( .A(u_sdrc_core_u_req_gen__abc_22171_n296_1), .B(u_sdrc_core_u_req_gen__abc_22171_n293), .Y(u_sdrc_core_u_req_gen__abc_22171_n297) );
  OR2X2 OR2X2_1065 ( .A(u_sdrc_core_u_req_gen__abc_22171_n286), .B(u_sdrc_core_u_req_gen__abc_22171_n297), .Y(u_sdrc_core_u_req_gen__abc_22171_n300) );
  OR2X2 OR2X2_1066 ( .A(u_sdrc_core_u_req_gen__abc_22171_n305), .B(u_sdrc_core_u_req_gen__abc_22171_n304_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n306) );
  OR2X2 OR2X2_1067 ( .A(u_sdrc_core_u_req_gen__abc_22171_n306), .B(u_sdrc_core_u_req_gen__abc_22171_n303), .Y(u_sdrc_core_u_req_gen__abc_22171_n307_1) );
  OR2X2 OR2X2_1068 ( .A(u_sdrc_core_u_req_gen__abc_22171_n310_1), .B(u_sdrc_core_u_req_gen__abc_22171_n309), .Y(u_sdrc_core_u_req_gen__abc_22171_n311) );
  OR2X2 OR2X2_1069 ( .A(app_req_ack_bF_buf5), .B(u_sdrc_core_r2b_write), .Y(u_sdrc_core_u_req_gen__abc_22171_n316) );
  OR2X2 OR2X2_107 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n463), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n464) );
  OR2X2 OR2X2_1070 ( .A(u_sdrc_core_u_req_gen__abc_22171_n331), .B(u_sdrc_core_u_req_gen__abc_22171_n332), .Y(u_sdrc_core_u_req_gen_lcl_wrap_FF_INPUT) );
  OR2X2 OR2X2_1071 ( .A(u_sdrc_core_u_req_gen__abc_22171_n338), .B(u_sdrc_core_u_req_gen__abc_22171_n340), .Y(u_sdrc_core_u_req_gen__abc_22171_n341_1) );
  OR2X2 OR2X2_1072 ( .A(u_sdrc_core_u_req_gen__abc_22171_n342), .B(u_sdrc_core_u_req_gen__abc_22171_n344), .Y(u_sdrc_core_u_req_gen_lcl_req_len_0__FF_INPUT) );
  OR2X2 OR2X2_1073 ( .A(u_sdrc_core_u_req_gen__abc_22171_n350_1), .B(u_sdrc_core_u_req_gen__abc_22171_n348), .Y(u_sdrc_core_u_req_gen__abc_22171_n351) );
  OR2X2 OR2X2_1074 ( .A(u_sdrc_core_u_req_gen__abc_22171_n351), .B(u_sdrc_core_u_req_gen__abc_22171_n347), .Y(u_sdrc_core_u_req_gen__abc_22171_n352_1) );
  OR2X2 OR2X2_1075 ( .A(u_sdrc_core_u_req_gen__abc_22171_n354_1), .B(u_sdrc_core_u_req_gen__abc_22171_n353), .Y(u_sdrc_core_u_req_gen__abc_22171_n355) );
  OR2X2 OR2X2_1076 ( .A(u_sdrc_core_u_req_gen__abc_22171_n356), .B(u_sdrc_core_u_req_gen__abc_22171_n346_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n357) );
  OR2X2 OR2X2_1077 ( .A(u_sdrc_core_u_req_gen__abc_22171_n335_1_bF_buf1), .B(u_sdrc_core_u_req_gen_lcl_req_len_1_), .Y(u_sdrc_core_u_req_gen__abc_22171_n358_1) );
  OR2X2 OR2X2_1078 ( .A(u_sdrc_core_u_req_gen__abc_22171_n359), .B(app_req_ack_bF_buf1), .Y(u_sdrc_core_u_req_gen__abc_22171_n360_1) );
  OR2X2 OR2X2_1079 ( .A(u_sdrc_core_u_req_gen__abc_22171_n362), .B(u_sdrc_core_u_req_gen__abc_22171_n361), .Y(u_sdrc_core_u_req_gen__abc_22171_n363) );
  OR2X2 OR2X2_108 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n283_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_10_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n465) );
  OR2X2 OR2X2_1080 ( .A(u_sdrc_core_u_req_gen__abc_22171_n363), .B(u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf2), .Y(u_sdrc_core_u_req_gen__abc_22171_n364) );
  OR2X2 OR2X2_1081 ( .A(u_sdrc_core_u_req_gen__abc_22171_n369_1), .B(u_sdrc_core_u_req_gen__abc_22171_n368), .Y(u_sdrc_core_u_req_gen__abc_22171_n370) );
  OR2X2 OR2X2_1082 ( .A(u_sdrc_core_u_req_gen__abc_22171_n367), .B(u_sdrc_core_u_req_gen__abc_22171_n370), .Y(u_sdrc_core_u_req_gen__abc_22171_n371_1) );
  OR2X2 OR2X2_1083 ( .A(u_sdrc_core_u_req_gen__abc_22171_n372), .B(u_sdrc_core_u_req_gen__abc_22171_n373_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n374) );
  OR2X2 OR2X2_1084 ( .A(u_sdrc_core_u_req_gen__abc_22171_n375), .B(u_sdrc_core_u_req_gen__abc_22171_n346_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n376) );
  OR2X2 OR2X2_1085 ( .A(u_sdrc_core_u_req_gen__abc_22171_n335_1_bF_buf0), .B(u_sdrc_core_u_req_gen_lcl_req_len_2_), .Y(u_sdrc_core_u_req_gen__abc_22171_n377_1) );
  OR2X2 OR2X2_1086 ( .A(u_sdrc_core_u_req_gen__abc_22171_n378), .B(app_req_ack_bF_buf0), .Y(u_sdrc_core_u_req_gen__abc_22171_n379_1) );
  OR2X2 OR2X2_1087 ( .A(u_sdrc_core_u_req_gen__abc_22171_n385), .B(u_sdrc_core_u_req_gen__abc_22171_n383), .Y(u_sdrc_core_u_req_gen__abc_22171_n386_1) );
  OR2X2 OR2X2_1088 ( .A(u_sdrc_core_u_req_gen__abc_22171_n386_1), .B(u_sdrc_core_u_req_gen__abc_22171_n381), .Y(u_sdrc_core_u_req_gen__abc_22171_n387) );
  OR2X2 OR2X2_1089 ( .A(u_sdrc_core_u_req_gen__abc_22171_n388_1), .B(u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf1), .Y(u_sdrc_core_u_req_gen__abc_22171_n389) );
  OR2X2 OR2X2_109 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n467), .B(u_sdrc_core_u_bank_ctl__abc_21249_n460), .Y(u_sdrc_core_b2x_addr_10_) );
  OR2X2 OR2X2_1090 ( .A(u_sdrc_core_u_req_gen__abc_22171_n391), .B(app_req_len_3_), .Y(u_sdrc_core_u_req_gen__abc_22171_n392) );
  OR2X2 OR2X2_1091 ( .A(u_sdrc_core_u_req_gen__abc_22171_n394_1), .B(u_sdrc_core_u_req_gen__abc_22171_n393), .Y(u_sdrc_core_u_req_gen__abc_22171_n395) );
  OR2X2 OR2X2_1092 ( .A(u_sdrc_core_u_req_gen__abc_22171_n404_1), .B(u_sdrc_core_u_req_gen__abc_22171_n403), .Y(u_sdrc_core_u_req_gen__abc_22171_n405) );
  OR2X2 OR2X2_1093 ( .A(u_sdrc_core_u_req_gen__abc_22171_n402), .B(u_sdrc_core_u_req_gen__abc_22171_n406_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n407) );
  OR2X2 OR2X2_1094 ( .A(u_sdrc_core_u_req_gen__abc_22171_n401), .B(u_sdrc_core_u_req_gen__abc_22171_n405), .Y(u_sdrc_core_u_req_gen__abc_22171_n408_1) );
  OR2X2 OR2X2_1095 ( .A(u_sdrc_core_u_req_gen__abc_22171_n410), .B(u_sdrc_core_u_req_gen__abc_22171_n399), .Y(u_sdrc_core_u_req_gen__abc_22171_n411) );
  OR2X2 OR2X2_1096 ( .A(u_sdrc_core_u_req_gen__abc_22171_n412_1), .B(u_sdrc_core_u_req_gen__abc_22171_n398), .Y(u_sdrc_core_u_req_gen_lcl_req_len_3__FF_INPUT) );
  OR2X2 OR2X2_1097 ( .A(u_sdrc_core_u_req_gen__abc_22171_n391), .B(app_req_len_4_), .Y(u_sdrc_core_u_req_gen__abc_22171_n414_1) );
  OR2X2 OR2X2_1098 ( .A(u_sdrc_core_u_req_gen__abc_22171_n241), .B(app_req_len_2_), .Y(u_sdrc_core_u_req_gen__abc_22171_n415) );
  OR2X2 OR2X2_1099 ( .A(u_sdrc_core_u_req_gen__abc_22171_n416), .B(app_req_len_3_), .Y(u_sdrc_core_u_req_gen__abc_22171_n417_1) );
  OR2X2 OR2X2_11 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n235_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n236), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n237_1) );
  OR2X2 OR2X2_110 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_11_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n470) );
  OR2X2 OR2X2_1100 ( .A(u_sdrc_core_u_req_gen__abc_22171_n427), .B(u_sdrc_core_u_req_gen_lcl_req_len_4_), .Y(u_sdrc_core_u_req_gen__abc_22171_n428) );
  OR2X2 OR2X2_1101 ( .A(u_sdrc_core_u_req_gen__abc_22171_n424), .B(u_sdrc_core_u_req_gen__abc_22171_n429_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n430) );
  OR2X2 OR2X2_1102 ( .A(u_sdrc_core_u_req_gen__abc_22171_n423_1), .B(u_sdrc_core_u_req_gen__abc_22171_n431_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n432) );
  OR2X2 OR2X2_1103 ( .A(u_sdrc_core_u_req_gen__abc_22171_n434), .B(u_sdrc_core_u_req_gen__abc_22171_n421_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n435) );
  OR2X2 OR2X2_1104 ( .A(u_sdrc_core_u_req_gen__abc_22171_n436_1), .B(u_sdrc_core_u_req_gen__abc_22171_n420), .Y(u_sdrc_core_u_req_gen_lcl_req_len_4__FF_INPUT) );
  OR2X2 OR2X2_1105 ( .A(u_sdrc_core_u_req_gen__abc_22171_n391), .B(app_req_len_5_), .Y(u_sdrc_core_u_req_gen__abc_22171_n438) );
  OR2X2 OR2X2_1106 ( .A(u_sdrc_core_u_req_gen__abc_22171_n241), .B(app_req_len_3_), .Y(u_sdrc_core_u_req_gen__abc_22171_n439) );
  OR2X2 OR2X2_1107 ( .A(u_sdrc_core_u_req_gen__abc_22171_n416), .B(app_req_len_4_), .Y(u_sdrc_core_u_req_gen__abc_22171_n440_1) );
  OR2X2 OR2X2_1108 ( .A(u_sdrc_core_u_req_gen__abc_22171_n449), .B(u_sdrc_core_u_req_gen_lcl_req_len_5_), .Y(u_sdrc_core_u_req_gen__abc_22171_n450_1) );
  OR2X2 OR2X2_1109 ( .A(u_sdrc_core_u_req_gen__abc_22171_n446), .B(u_sdrc_core_u_req_gen__abc_22171_n451_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n452_1) );
  OR2X2 OR2X2_111 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n223_1_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_11_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n471) );
  OR2X2 OR2X2_1110 ( .A(u_sdrc_core_u_req_gen__abc_22171_n445), .B(u_sdrc_core_u_req_gen__abc_22171_n453), .Y(u_sdrc_core_u_req_gen__abc_22171_n454) );
  OR2X2 OR2X2_1111 ( .A(u_sdrc_core_u_req_gen__abc_22171_n456), .B(u_sdrc_core_u_req_gen__abc_22171_n444_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n457) );
  OR2X2 OR2X2_1112 ( .A(u_sdrc_core_u_req_gen__abc_22171_n458), .B(u_sdrc_core_u_req_gen__abc_22171_n443), .Y(u_sdrc_core_u_req_gen_lcl_req_len_5__FF_INPUT) );
  OR2X2 OR2X2_1113 ( .A(u_sdrc_core_u_req_gen__abc_22171_n391), .B(app_req_len_6_), .Y(u_sdrc_core_u_req_gen__abc_22171_n460) );
  OR2X2 OR2X2_1114 ( .A(u_sdrc_core_u_req_gen__abc_22171_n241), .B(app_req_len_4_), .Y(u_sdrc_core_u_req_gen__abc_22171_n461) );
  OR2X2 OR2X2_1115 ( .A(u_sdrc_core_u_req_gen__abc_22171_n416), .B(app_req_len_5_), .Y(u_sdrc_core_u_req_gen__abc_22171_n462_1) );
  OR2X2 OR2X2_1116 ( .A(u_sdrc_core_u_req_gen__abc_22171_n464_1), .B(u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf2), .Y(u_sdrc_core_u_req_gen__abc_22171_n465) );
  OR2X2 OR2X2_1117 ( .A(u_sdrc_core_u_req_gen__abc_22171_n467), .B(u_sdrc_core_r2b_len_6_), .Y(u_sdrc_core_u_req_gen__abc_22171_n470) );
  OR2X2 OR2X2_1118 ( .A(u_sdrc_core_u_req_gen__abc_22171_n473), .B(u_sdrc_core_u_req_gen__abc_22171_n466_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n474_1) );
  OR2X2 OR2X2_1119 ( .A(u_sdrc_core_u_req_gen__abc_22171_n472), .B(u_sdrc_core_u_req_gen_lcl_req_len_6_), .Y(u_sdrc_core_u_req_gen__abc_22171_n475) );
  OR2X2 OR2X2_112 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n472), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf0), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n473) );
  OR2X2 OR2X2_1120 ( .A(u_sdrc_core_u_req_gen__abc_22171_n476), .B(app_req_ack_bF_buf3), .Y(u_sdrc_core_u_req_gen__abc_22171_n477_1) );
  OR2X2 OR2X2_1121 ( .A(u_sdrc_core_u_req_gen__abc_22171_n480_1), .B(u_sdrc_core_u_req_gen__abc_22171_n346_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n481) );
  OR2X2 OR2X2_1122 ( .A(u_sdrc_core_u_req_gen__abc_22171_n336), .B(u_sdrc_core_r2b_caddr_0_), .Y(u_sdrc_core_u_req_gen__abc_22171_n482) );
  OR2X2 OR2X2_1123 ( .A(u_sdrc_core_u_req_gen__abc_22171_n484), .B(u_sdrc_core_u_req_gen_max_r2b_len_r_0__FF_INPUT), .Y(u_sdrc_core_u_req_gen_map_address_0_) );
  OR2X2 OR2X2_1124 ( .A(u_sdrc_core_u_req_gen__abc_22171_n487), .B(u_sdrc_core_u_req_gen__abc_22171_n209), .Y(u_sdrc_core_u_req_gen__abc_22171_n488) );
  OR2X2 OR2X2_1125 ( .A(u_sdrc_core_u_req_gen__abc_22171_n488), .B(u_sdrc_core_u_req_gen__abc_22171_n486_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n489_1) );
  OR2X2 OR2X2_1126 ( .A(u_sdrc_core_r2b_len_1_), .B(u_sdrc_core_r2b_caddr_1_), .Y(u_sdrc_core_u_req_gen__abc_22171_n490) );
  OR2X2 OR2X2_1127 ( .A(u_sdrc_core_u_req_gen__abc_22171_n491), .B(u_sdrc_core_u_req_gen__abc_22171_n479), .Y(u_sdrc_core_u_req_gen__abc_22171_n494) );
  OR2X2 OR2X2_1128 ( .A(u_sdrc_core_u_req_gen__abc_22171_n495_1), .B(u_sdrc_core_u_req_gen__abc_22171_n346_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n496) );
  OR2X2 OR2X2_1129 ( .A(u_sdrc_core_u_req_gen__abc_22171_n335_1_bF_buf3), .B(u_sdrc_core_r2b_caddr_1_), .Y(u_sdrc_core_u_req_gen__abc_22171_n497) );
  OR2X2 OR2X2_113 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n283_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_11_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n474) );
  OR2X2 OR2X2_1130 ( .A(u_sdrc_core_u_req_gen__abc_22171_n498_1), .B(app_req_ack_bF_buf2), .Y(u_sdrc_core_u_req_gen__abc_22171_n499) );
  OR2X2 OR2X2_1131 ( .A(u_sdrc_core_u_req_gen__abc_22171_n248), .B(u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf0), .Y(u_sdrc_core_u_req_gen__abc_22171_n500) );
  OR2X2 OR2X2_1132 ( .A(u_sdrc_core_u_req_gen__abc_22171_n492_1), .B(u_sdrc_core_u_req_gen__abc_22171_n502), .Y(u_sdrc_core_u_req_gen__abc_22171_n503) );
  OR2X2 OR2X2_1133 ( .A(u_sdrc_core_r2b_len_2_), .B(u_sdrc_core_r2b_caddr_2_), .Y(u_sdrc_core_u_req_gen__abc_22171_n506) );
  OR2X2 OR2X2_1134 ( .A(u_sdrc_core_u_req_gen__abc_22171_n503), .B(u_sdrc_core_u_req_gen__abc_22171_n507_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n510_1) );
  OR2X2 OR2X2_1135 ( .A(u_sdrc_core_u_req_gen__abc_22171_n511), .B(u_sdrc_core_u_req_gen__abc_22171_n346_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n512) );
  OR2X2 OR2X2_1136 ( .A(u_sdrc_core_u_req_gen__abc_22171_n335_1_bF_buf2), .B(u_sdrc_core_r2b_caddr_2_), .Y(u_sdrc_core_u_req_gen__abc_22171_n513) );
  OR2X2 OR2X2_1137 ( .A(u_sdrc_core_u_req_gen__abc_22171_n514), .B(app_req_ack_bF_buf1), .Y(u_sdrc_core_u_req_gen__abc_22171_n515) );
  OR2X2 OR2X2_1138 ( .A(u_sdrc_core_u_req_gen__abc_22171_n264), .B(u_sdrc_core_u_req_gen__abc_22171_n318_bF_buf4), .Y(u_sdrc_core_u_req_gen__abc_22171_n516) );
  OR2X2 OR2X2_1139 ( .A(u_sdrc_core_u_req_gen__abc_22171_n222), .B(u_sdrc_core_u_req_gen__abc_22171_n521), .Y(u_sdrc_core_u_req_gen__abc_22171_n522) );
  OR2X2 OR2X2_114 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n476), .B(u_sdrc_core_u_bank_ctl__abc_21249_n469), .Y(u_sdrc_core_b2x_addr_11_) );
  OR2X2 OR2X2_1140 ( .A(u_sdrc_core_u_req_gen__abc_22171_n520), .B(u_sdrc_core_u_req_gen__abc_22171_n525), .Y(u_sdrc_core_u_req_gen__abc_22171_n526) );
  OR2X2 OR2X2_1141 ( .A(u_sdrc_core_u_req_gen__abc_22171_n519), .B(u_sdrc_core_u_req_gen__abc_22171_n527_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n528) );
  OR2X2 OR2X2_1142 ( .A(u_sdrc_core_u_req_gen__abc_22171_n530), .B(u_sdrc_core_u_req_gen__abc_22171_n518), .Y(u_sdrc_core_u_req_gen__abc_22171_n531) );
  OR2X2 OR2X2_1143 ( .A(u_sdrc_core_u_req_gen__abc_22171_n532), .B(u_sdrc_core_u_req_gen__abc_22171_n534), .Y(u_sdrc_core_u_req_gen_map_address_3_) );
  OR2X2 OR2X2_1144 ( .A(u_sdrc_core_r2b_len_4_), .B(u_sdrc_core_r2b_caddr_4_), .Y(u_sdrc_core_u_req_gen__abc_22171_n540) );
  OR2X2 OR2X2_1145 ( .A(u_sdrc_core_u_req_gen__abc_22171_n543), .B(u_sdrc_core_u_req_gen__abc_22171_n542), .Y(u_sdrc_core_u_req_gen__abc_22171_n544) );
  OR2X2 OR2X2_1146 ( .A(u_sdrc_core_u_req_gen__abc_22171_n546), .B(u_sdrc_core_u_req_gen__abc_22171_n544), .Y(u_sdrc_core_u_req_gen__abc_22171_n547) );
  OR2X2 OR2X2_1147 ( .A(u_sdrc_core_u_req_gen__abc_22171_n547), .B(u_sdrc_core_u_req_gen__abc_22171_n541), .Y(u_sdrc_core_u_req_gen__abc_22171_n548) );
  OR2X2 OR2X2_1148 ( .A(u_sdrc_core_u_req_gen__abc_22171_n552), .B(u_sdrc_core_u_req_gen__abc_22171_n537), .Y(u_sdrc_core_u_req_gen__abc_22171_n553) );
  OR2X2 OR2X2_1149 ( .A(u_sdrc_core_u_req_gen__abc_22171_n554), .B(u_sdrc_core_u_req_gen__abc_22171_n536), .Y(u_sdrc_core_u_req_gen_map_address_4_) );
  OR2X2 OR2X2_115 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_12_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n479) );
  OR2X2 OR2X2_1150 ( .A(u_sdrc_core_r2b_len_5_), .B(u_sdrc_core_r2b_caddr_5_), .Y(u_sdrc_core_u_req_gen__abc_22171_n561) );
  OR2X2 OR2X2_1151 ( .A(u_sdrc_core_u_req_gen__abc_22171_n558), .B(u_sdrc_core_u_req_gen__abc_22171_n562), .Y(u_sdrc_core_u_req_gen__abc_22171_n563) );
  OR2X2 OR2X2_1152 ( .A(u_sdrc_core_u_req_gen__abc_22171_n557), .B(u_sdrc_core_u_req_gen__abc_22171_n564), .Y(u_sdrc_core_u_req_gen__abc_22171_n565) );
  OR2X2 OR2X2_1153 ( .A(u_sdrc_core_u_req_gen__abc_22171_n567), .B(u_sdrc_core_u_req_gen__abc_22171_n556), .Y(u_sdrc_core_u_req_gen__abc_22171_n568) );
  OR2X2 OR2X2_1154 ( .A(u_sdrc_core_u_req_gen__abc_22171_n569), .B(u_sdrc_core_u_req_gen__abc_22171_n571), .Y(u_sdrc_core_u_req_gen_map_address_5_) );
  OR2X2 OR2X2_1155 ( .A(u_sdrc_core_u_req_gen__abc_22171_n538), .B(u_sdrc_core_u_req_gen__abc_22171_n559), .Y(u_sdrc_core_u_req_gen__abc_22171_n575) );
  OR2X2 OR2X2_1156 ( .A(u_sdrc_core_u_req_gen__abc_22171_n578), .B(u_sdrc_core_u_req_gen__abc_22171_n576), .Y(u_sdrc_core_u_req_gen__abc_22171_n579) );
  OR2X2 OR2X2_1157 ( .A(u_sdrc_core_r2b_len_6_), .B(u_sdrc_core_r2b_caddr_6_), .Y(u_sdrc_core_u_req_gen__abc_22171_n582) );
  OR2X2 OR2X2_1158 ( .A(u_sdrc_core_u_req_gen__abc_22171_n579), .B(u_sdrc_core_u_req_gen__abc_22171_n583), .Y(u_sdrc_core_u_req_gen__abc_22171_n584) );
  OR2X2 OR2X2_1159 ( .A(u_sdrc_core_u_req_gen__abc_22171_n588_1), .B(u_sdrc_core_u_req_gen__abc_22171_n574), .Y(u_sdrc_core_u_req_gen__abc_22171_n589) );
  OR2X2 OR2X2_116 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n223_1_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_12_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n480) );
  OR2X2 OR2X2_1160 ( .A(u_sdrc_core_u_req_gen__abc_22171_n590), .B(u_sdrc_core_u_req_gen__abc_22171_n573), .Y(u_sdrc_core_u_req_gen_map_address_6_) );
  OR2X2 OR2X2_1161 ( .A(u_sdrc_core_u_req_gen__abc_22171_n594), .B(u_sdrc_core_u_req_gen__abc_22171_n593), .Y(u_sdrc_core_u_req_gen__abc_22171_n595) );
  OR2X2 OR2X2_1162 ( .A(u_sdrc_core_u_req_gen__abc_22171_n595), .B(u_sdrc_core_u_req_gen__abc_22171_n592), .Y(u_sdrc_core_u_req_gen__abc_22171_n596) );
  OR2X2 OR2X2_1163 ( .A(u_sdrc_core_u_req_gen__abc_22171_n599), .B(u_sdrc_core_u_req_gen__abc_22171_n346_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n600) );
  OR2X2 OR2X2_1164 ( .A(u_sdrc_core_u_req_gen__abc_22171_n602), .B(u_sdrc_core_u_req_gen__abc_22171_n603), .Y(u_sdrc_core_u_req_gen__abc_22171_n604) );
  OR2X2 OR2X2_1165 ( .A(u_sdrc_core_u_req_gen__abc_22171_n605), .B(u_sdrc_core_u_req_gen__abc_22171_n597), .Y(u_sdrc_core_u_req_gen_map_address_7_) );
  OR2X2 OR2X2_1166 ( .A(u_sdrc_core_u_req_gen__abc_22171_n609), .B(u_sdrc_core_u_req_gen__abc_22171_n608), .Y(u_sdrc_core_u_req_gen__abc_22171_n610) );
  OR2X2 OR2X2_1167 ( .A(u_sdrc_core_u_req_gen__abc_22171_n610), .B(u_sdrc_core_u_req_gen__abc_22171_n607), .Y(u_sdrc_core_u_req_gen__abc_22171_n611) );
  OR2X2 OR2X2_1168 ( .A(u_sdrc_core_u_req_gen__abc_22171_n576), .B(u_sdrc_core_u_req_gen__abc_22171_n580), .Y(u_sdrc_core_u_req_gen__abc_22171_n616) );
  OR2X2 OR2X2_1169 ( .A(u_sdrc_core_u_req_gen__abc_22171_n615), .B(u_sdrc_core_u_req_gen__abc_22171_n618), .Y(u_sdrc_core_u_req_gen__abc_22171_n619) );
  OR2X2 OR2X2_117 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n481), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf4), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n482) );
  OR2X2 OR2X2_1170 ( .A(u_sdrc_core_u_req_gen__abc_22171_n620), .B(u_sdrc_core_u_req_gen_curr_sdr_addr_8_), .Y(u_sdrc_core_u_req_gen__abc_22171_n621) );
  OR2X2 OR2X2_1171 ( .A(u_sdrc_core_u_req_gen__abc_22171_n625), .B(u_sdrc_core_u_req_gen__abc_22171_n612), .Y(u_sdrc_core_u_req_gen_map_address_8_) );
  OR2X2 OR2X2_1172 ( .A(u_sdrc_core_u_req_gen__abc_22171_n629), .B(u_sdrc_core_u_req_gen__abc_22171_n628), .Y(u_sdrc_core_u_req_gen__abc_22171_n630) );
  OR2X2 OR2X2_1173 ( .A(u_sdrc_core_u_req_gen__abc_22171_n630), .B(u_sdrc_core_u_req_gen__abc_22171_n627), .Y(u_sdrc_core_u_req_gen__abc_22171_n631) );
  OR2X2 OR2X2_1174 ( .A(u_sdrc_core_u_req_gen__abc_22171_n622), .B(u_sdrc_core_u_req_gen_curr_sdr_addr_9_), .Y(u_sdrc_core_u_req_gen__abc_22171_n633) );
  OR2X2 OR2X2_1175 ( .A(u_sdrc_core_u_req_gen__abc_22171_n638), .B(u_sdrc_core_u_req_gen__abc_22171_n632), .Y(u_sdrc_core_u_req_gen_map_address_9_) );
  OR2X2 OR2X2_1176 ( .A(u_sdrc_core_u_req_gen__abc_22171_n391), .B(app_req_addr_10_), .Y(u_sdrc_core_u_req_gen__abc_22171_n640) );
  OR2X2 OR2X2_1177 ( .A(u_sdrc_core_u_req_gen__abc_22171_n241), .B(app_req_addr_8_), .Y(u_sdrc_core_u_req_gen__abc_22171_n641) );
  OR2X2 OR2X2_1178 ( .A(u_sdrc_core_u_req_gen__abc_22171_n416), .B(app_req_addr_9_), .Y(u_sdrc_core_u_req_gen__abc_22171_n642) );
  OR2X2 OR2X2_1179 ( .A(u_sdrc_core_u_req_gen__abc_22171_n635), .B(u_sdrc_core_u_req_gen_curr_sdr_addr_10_), .Y(u_sdrc_core_u_req_gen__abc_22171_n648) );
  OR2X2 OR2X2_118 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n283_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_12_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n483) );
  OR2X2 OR2X2_1180 ( .A(u_sdrc_core_u_req_gen__abc_22171_n650), .B(u_sdrc_core_u_req_gen__abc_22171_n645), .Y(u_sdrc_core_u_req_gen_map_address_10_) );
  OR2X2 OR2X2_1181 ( .A(u_sdrc_core_u_req_gen__abc_22171_n653), .B(u_sdrc_core_u_req_gen__abc_22171_n654), .Y(u_sdrc_core_u_req_gen__abc_22171_n655) );
  OR2X2 OR2X2_1182 ( .A(u_sdrc_core_u_req_gen__abc_22171_n655), .B(u_sdrc_core_u_req_gen__abc_22171_n652), .Y(u_sdrc_core_u_req_gen__abc_22171_n656) );
  OR2X2 OR2X2_1183 ( .A(u_sdrc_core_u_req_gen__abc_22171_n646), .B(u_sdrc_core_u_req_gen_curr_sdr_addr_11_), .Y(u_sdrc_core_u_req_gen__abc_22171_n662) );
  OR2X2 OR2X2_1184 ( .A(u_sdrc_core_u_req_gen__abc_22171_n664), .B(u_sdrc_core_u_req_gen__abc_22171_n657), .Y(u_sdrc_core_u_req_gen_map_address_11_) );
  OR2X2 OR2X2_1185 ( .A(u_sdrc_core_u_req_gen__abc_22171_n668), .B(u_sdrc_core_u_req_gen__abc_22171_n667), .Y(u_sdrc_core_u_req_gen__abc_22171_n669) );
  OR2X2 OR2X2_1186 ( .A(u_sdrc_core_u_req_gen__abc_22171_n669), .B(u_sdrc_core_u_req_gen__abc_22171_n666), .Y(u_sdrc_core_u_req_gen__abc_22171_n670) );
  OR2X2 OR2X2_1187 ( .A(u_sdrc_core_u_req_gen__abc_22171_n660), .B(u_sdrc_core_u_req_gen_curr_sdr_addr_12_), .Y(u_sdrc_core_u_req_gen__abc_22171_n674) );
  OR2X2 OR2X2_1188 ( .A(u_sdrc_core_u_req_gen__abc_22171_n676), .B(u_sdrc_core_u_req_gen__abc_22171_n671), .Y(u_sdrc_core_u_req_gen_map_address_12_) );
  OR2X2 OR2X2_1189 ( .A(u_sdrc_core_u_req_gen__abc_22171_n672), .B(u_sdrc_core_u_req_gen_curr_sdr_addr_13_), .Y(u_sdrc_core_u_req_gen__abc_22171_n678) );
  OR2X2 OR2X2_119 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n485), .B(u_sdrc_core_u_bank_ctl__abc_21249_n478), .Y(u_sdrc_core_b2x_addr_12_) );
  OR2X2 OR2X2_1190 ( .A(u_sdrc_core_u_req_gen__abc_22171_n687), .B(u_sdrc_core_u_req_gen__abc_22171_n686), .Y(u_sdrc_core_u_req_gen__abc_22171_n688) );
  OR2X2 OR2X2_1191 ( .A(u_sdrc_core_u_req_gen__abc_22171_n688), .B(u_sdrc_core_u_req_gen__abc_22171_n685), .Y(u_sdrc_core_u_req_gen__abc_22171_n689) );
  OR2X2 OR2X2_1192 ( .A(u_sdrc_core_u_req_gen__abc_22171_n684), .B(u_sdrc_core_u_req_gen__abc_22171_n690), .Y(u_sdrc_core_u_req_gen_map_address_13_) );
  OR2X2 OR2X2_1193 ( .A(u_sdrc_core_u_req_gen__abc_22171_n681), .B(u_sdrc_core_u_req_gen_curr_sdr_addr_14_), .Y(u_sdrc_core_u_req_gen__abc_22171_n692) );
  OR2X2 OR2X2_1194 ( .A(u_sdrc_core_u_req_gen__abc_22171_n699), .B(u_sdrc_core_u_req_gen__abc_22171_n698), .Y(u_sdrc_core_u_req_gen__abc_22171_n700) );
  OR2X2 OR2X2_1195 ( .A(u_sdrc_core_u_req_gen__abc_22171_n700), .B(u_sdrc_core_u_req_gen__abc_22171_n697), .Y(u_sdrc_core_u_req_gen__abc_22171_n701) );
  OR2X2 OR2X2_1196 ( .A(u_sdrc_core_u_req_gen__abc_22171_n696), .B(u_sdrc_core_u_req_gen__abc_22171_n702), .Y(u_sdrc_core_u_req_gen_map_address_14_) );
  OR2X2 OR2X2_1197 ( .A(u_sdrc_core_u_req_gen__abc_22171_n705), .B(u_sdrc_core_u_req_gen__abc_22171_n706), .Y(u_sdrc_core_u_req_gen__abc_22171_n707) );
  OR2X2 OR2X2_1198 ( .A(u_sdrc_core_u_req_gen__abc_22171_n707), .B(u_sdrc_core_u_req_gen__abc_22171_n704), .Y(u_sdrc_core_u_req_gen__abc_22171_n708) );
  OR2X2 OR2X2_1199 ( .A(u_sdrc_core_u_req_gen__abc_22171_n693), .B(u_sdrc_core_u_req_gen_curr_sdr_addr_15_), .Y(u_sdrc_core_u_req_gen__abc_22171_n710) );
  OR2X2 OR2X2_12 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n237_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n234), .Y(u_sdrc_core_b2x_req) );
  OR2X2 OR2X2_120 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_len_0_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n488) );
  OR2X2 OR2X2_1200 ( .A(u_sdrc_core_u_req_gen__abc_22171_n717), .B(u_sdrc_core_u_req_gen__abc_22171_n709), .Y(u_sdrc_core_u_req_gen_map_address_15_) );
  OR2X2 OR2X2_1201 ( .A(u_sdrc_core_u_req_gen__abc_22171_n721), .B(u_sdrc_core_u_req_gen__abc_22171_n720), .Y(u_sdrc_core_u_req_gen__abc_22171_n722) );
  OR2X2 OR2X2_1202 ( .A(u_sdrc_core_u_req_gen__abc_22171_n722), .B(u_sdrc_core_u_req_gen__abc_22171_n719), .Y(u_sdrc_core_u_req_gen__abc_22171_n723) );
  OR2X2 OR2X2_1203 ( .A(u_sdrc_core_u_req_gen__abc_22171_n714), .B(u_sdrc_core_u_req_gen_curr_sdr_addr_16_), .Y(u_sdrc_core_u_req_gen__abc_22171_n727) );
  OR2X2 OR2X2_1204 ( .A(u_sdrc_core_u_req_gen__abc_22171_n729), .B(u_sdrc_core_u_req_gen__abc_22171_n724), .Y(u_sdrc_core_u_req_gen_map_address_16_) );
  OR2X2 OR2X2_1205 ( .A(u_sdrc_core_u_req_gen__abc_22171_n732), .B(u_sdrc_core_u_req_gen__abc_22171_n733), .Y(u_sdrc_core_u_req_gen__abc_22171_n734) );
  OR2X2 OR2X2_1206 ( .A(u_sdrc_core_u_req_gen__abc_22171_n734), .B(u_sdrc_core_u_req_gen__abc_22171_n731), .Y(u_sdrc_core_u_req_gen__abc_22171_n735) );
  OR2X2 OR2X2_1207 ( .A(u_sdrc_core_u_req_gen__abc_22171_n725), .B(u_sdrc_core_u_req_gen_curr_sdr_addr_17_), .Y(u_sdrc_core_u_req_gen__abc_22171_n740) );
  OR2X2 OR2X2_1208 ( .A(u_sdrc_core_u_req_gen__abc_22171_n742), .B(u_sdrc_core_u_req_gen__abc_22171_n736), .Y(u_sdrc_core_u_req_gen_map_address_17_) );
  OR2X2 OR2X2_1209 ( .A(u_sdrc_core_u_req_gen__abc_22171_n745), .B(u_sdrc_core_u_req_gen__abc_22171_n746), .Y(u_sdrc_core_u_req_gen__abc_22171_n747) );
  OR2X2 OR2X2_121 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n223_1_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_len_0_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n489) );
  OR2X2 OR2X2_1210 ( .A(u_sdrc_core_u_req_gen__abc_22171_n747), .B(u_sdrc_core_u_req_gen__abc_22171_n744), .Y(u_sdrc_core_u_req_gen__abc_22171_n748) );
  OR2X2 OR2X2_1211 ( .A(u_sdrc_core_u_req_gen__abc_22171_n750), .B(u_sdrc_core_u_req_gen__abc_22171_n752), .Y(u_sdrc_core_u_req_gen__abc_22171_n753) );
  OR2X2 OR2X2_1212 ( .A(u_sdrc_core_u_req_gen__abc_22171_n754), .B(u_sdrc_core_u_req_gen__abc_22171_n749), .Y(u_sdrc_core_u_req_gen_map_address_18_) );
  OR2X2 OR2X2_1213 ( .A(u_sdrc_core_u_req_gen__abc_22171_n757), .B(u_sdrc_core_u_req_gen_curr_sdr_addr_19_), .Y(u_sdrc_core_u_req_gen__abc_22171_n758) );
  OR2X2 OR2X2_1214 ( .A(u_sdrc_core_u_req_gen__abc_22171_n767), .B(u_sdrc_core_u_req_gen__abc_22171_n766), .Y(u_sdrc_core_u_req_gen__abc_22171_n768) );
  OR2X2 OR2X2_1215 ( .A(u_sdrc_core_u_req_gen__abc_22171_n768), .B(u_sdrc_core_u_req_gen__abc_22171_n765), .Y(u_sdrc_core_u_req_gen__abc_22171_n769) );
  OR2X2 OR2X2_1216 ( .A(u_sdrc_core_u_req_gen__abc_22171_n764), .B(u_sdrc_core_u_req_gen__abc_22171_n770), .Y(u_sdrc_core_u_req_gen_map_address_19_) );
  OR2X2 OR2X2_1217 ( .A(u_sdrc_core_u_req_gen__abc_22171_n773), .B(u_sdrc_core_u_req_gen__abc_22171_n774), .Y(u_sdrc_core_u_req_gen__abc_22171_n775) );
  OR2X2 OR2X2_1218 ( .A(u_sdrc_core_u_req_gen__abc_22171_n775), .B(u_sdrc_core_u_req_gen__abc_22171_n772), .Y(u_sdrc_core_u_req_gen__abc_22171_n776) );
  OR2X2 OR2X2_1219 ( .A(u_sdrc_core_u_req_gen__abc_22171_n761), .B(u_sdrc_core_u_req_gen_curr_sdr_addr_20_), .Y(u_sdrc_core_u_req_gen__abc_22171_n778) );
  OR2X2 OR2X2_122 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n490), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf3), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n491) );
  OR2X2 OR2X2_1220 ( .A(u_sdrc_core_u_req_gen__abc_22171_n783), .B(u_sdrc_core_u_req_gen__abc_22171_n777), .Y(u_sdrc_core_u_req_gen_map_address_20_) );
  OR2X2 OR2X2_1221 ( .A(u_sdrc_core_u_req_gen__abc_22171_n788), .B(u_sdrc_core_u_req_gen__abc_22171_n789), .Y(u_sdrc_core_u_req_gen__abc_22171_n790) );
  OR2X2 OR2X2_1222 ( .A(u_sdrc_core_u_req_gen__abc_22171_n780), .B(u_sdrc_core_u_req_gen_curr_sdr_addr_21_), .Y(u_sdrc_core_u_req_gen__abc_22171_n793) );
  OR2X2 OR2X2_1223 ( .A(u_sdrc_core_u_req_gen__abc_22171_n794), .B(u_sdrc_core_u_req_gen__abc_22171_n795), .Y(u_sdrc_core_u_req_gen__abc_22171_n796) );
  OR2X2 OR2X2_1224 ( .A(u_sdrc_core_u_req_gen__abc_22171_n797), .B(u_sdrc_core_u_req_gen__abc_22171_n792), .Y(u_sdrc_core_u_req_gen__abc_22171_n798) );
  OR2X2 OR2X2_1225 ( .A(u_sdrc_core_u_req_gen__abc_22171_n802), .B(u_sdrc_core_u_req_gen__abc_22171_n801), .Y(u_sdrc_core_u_req_gen__abc_22171_n803) );
  OR2X2 OR2X2_1226 ( .A(u_sdrc_core_u_req_gen__abc_22171_n803), .B(u_sdrc_core_u_req_gen__abc_22171_n800), .Y(u_sdrc_core_u_req_gen__abc_22171_n804) );
  OR2X2 OR2X2_1227 ( .A(u_sdrc_core_u_req_gen__abc_22171_n795), .B(u_sdrc_core_u_req_gen__abc_22171_n807), .Y(u_sdrc_core_u_req_gen__abc_22171_n810) );
  OR2X2 OR2X2_1228 ( .A(u_sdrc_core_u_req_gen__abc_22171_n812), .B(u_sdrc_core_u_req_gen__abc_22171_n806), .Y(u_sdrc_core_u_req_gen__abc_22171_n813) );
  OR2X2 OR2X2_1229 ( .A(u_sdrc_core_u_req_gen__abc_22171_n816), .B(u_sdrc_core_u_req_gen__abc_22171_n817), .Y(u_sdrc_core_u_req_gen__abc_22171_n818) );
  OR2X2 OR2X2_123 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n283_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_len_0_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n492) );
  OR2X2 OR2X2_1230 ( .A(u_sdrc_core_u_req_gen__abc_22171_n818), .B(u_sdrc_core_u_req_gen__abc_22171_n815), .Y(u_sdrc_core_u_req_gen__abc_22171_n819) );
  OR2X2 OR2X2_1231 ( .A(u_sdrc_core_u_req_gen__abc_22171_n828), .B(app_req_ack_bF_buf0), .Y(u_sdrc_core_u_req_gen__abc_22171_n829) );
  OR2X2 OR2X2_1232 ( .A(u_sdrc_core_u_req_gen__abc_22171_n829), .B(u_sdrc_core_u_req_gen__abc_22171_n827), .Y(u_sdrc_core_u_req_gen__abc_22171_n830) );
  OR2X2 OR2X2_1233 ( .A(u_sdrc_core_u_req_gen__abc_22171_n834), .B(u_sdrc_core_u_req_gen__abc_22171_n835), .Y(u_sdrc_core_u_req_gen__abc_22171_n836) );
  OR2X2 OR2X2_1234 ( .A(u_sdrc_core_u_req_gen__abc_22171_n836), .B(u_sdrc_core_u_req_gen__abc_22171_n833), .Y(u_sdrc_core_u_req_gen__abc_22171_n837) );
  OR2X2 OR2X2_1235 ( .A(u_sdrc_core_u_req_gen__abc_22171_n847), .B(app_req_ack_bF_buf5), .Y(u_sdrc_core_u_req_gen__abc_22171_n848) );
  OR2X2 OR2X2_1236 ( .A(u_sdrc_core_u_req_gen__abc_22171_n848), .B(u_sdrc_core_u_req_gen__abc_22171_n846), .Y(u_sdrc_core_u_req_gen__abc_22171_n849) );
  OR2X2 OR2X2_1237 ( .A(u_sdrc_core_u_req_gen__abc_22171_n853), .B(u_sdrc_core_u_req_gen__abc_22171_n854), .Y(u_sdrc_core_u_req_gen__abc_22171_n855) );
  OR2X2 OR2X2_1238 ( .A(u_sdrc_core_u_req_gen__abc_22171_n855), .B(u_sdrc_core_u_req_gen__abc_22171_n852), .Y(u_sdrc_core_u_req_gen__abc_22171_n856) );
  OR2X2 OR2X2_1239 ( .A(u_sdrc_core_u_req_gen__abc_22171_n863), .B(u_sdrc_core_u_req_gen__abc_22171_n859), .Y(u_sdrc_core_u_req_gen__abc_22171_n864) );
  OR2X2 OR2X2_124 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n494), .B(u_sdrc_core_u_bank_ctl__abc_21249_n487), .Y(u_sdrc_core_b2x_len_0_) );
  OR2X2 OR2X2_1240 ( .A(u_sdrc_core_u_req_gen__abc_22171_n865), .B(u_sdrc_core_u_req_gen_curr_sdr_addr_25_), .Y(u_sdrc_core_u_req_gen__abc_22171_n866) );
  OR2X2 OR2X2_1241 ( .A(u_sdrc_core_u_req_gen__abc_22171_n867), .B(app_req_ack_bF_buf3), .Y(u_sdrc_core_u_req_gen__abc_22171_n868) );
  OR2X2 OR2X2_1242 ( .A(u_sdrc_core_u_req_gen__abc_22171_n880), .B(u_sdrc_core_u_req_gen__abc_22171_n878), .Y(u_sdrc_core_u_req_gen__abc_22171_n881) );
  OR2X2 OR2X2_1243 ( .A(u_sdrc_core_u_req_gen__abc_22171_n881), .B(u_sdrc_core_u_req_gen__abc_22171_n875), .Y(u_sdrc_core_u_req_gen__abc_22171_n882) );
  OR2X2 OR2X2_1244 ( .A(u_sdrc_core_u_req_gen__abc_22171_n882), .B(u_sdrc_core_u_req_gen__abc_22171_n872), .Y(u_sdrc_core_u_req_gen_r2b_ba_0__FF_INPUT) );
  OR2X2 OR2X2_1245 ( .A(u_sdrc_core_u_req_gen__abc_22171_n889), .B(u_sdrc_core_u_req_gen__abc_22171_n877), .Y(u_sdrc_core_u_req_gen__abc_22171_n890) );
  OR2X2 OR2X2_1246 ( .A(u_sdrc_core_u_req_gen__abc_22171_n890), .B(u_sdrc_core_u_req_gen__abc_22171_n885), .Y(u_sdrc_core_u_req_gen__abc_22171_n891) );
  OR2X2 OR2X2_1247 ( .A(u_sdrc_core_u_req_gen__abc_22171_n891), .B(u_sdrc_core_u_req_gen__abc_22171_n884), .Y(u_sdrc_core_u_req_gen__abc_22171_n892) );
  OR2X2 OR2X2_1248 ( .A(u_sdrc_core_u_req_gen_map_address_9_), .B(u_sdrc_core_u_req_gen__abc_22171_n893_bF_buf3), .Y(u_sdrc_core_u_req_gen__abc_22171_n894) );
  OR2X2 OR2X2_1249 ( .A(u_sdrc_core_u_req_gen__abc_22171_n901), .B(u_sdrc_core_u_req_gen__abc_22171_n877), .Y(u_sdrc_core_u_req_gen__abc_22171_n902) );
  OR2X2 OR2X2_125 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_len_1_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n497) );
  OR2X2 OR2X2_1250 ( .A(u_sdrc_core_u_req_gen__abc_22171_n902), .B(u_sdrc_core_u_req_gen__abc_22171_n900), .Y(u_sdrc_core_u_req_gen__abc_22171_n903) );
  OR2X2 OR2X2_1251 ( .A(u_sdrc_core_u_req_gen__abc_22171_n903), .B(u_sdrc_core_u_req_gen__abc_22171_n899), .Y(u_sdrc_core_u_req_gen__abc_22171_n904) );
  OR2X2 OR2X2_1252 ( .A(u_sdrc_core_u_req_gen_map_address_10_), .B(u_sdrc_core_u_req_gen__abc_22171_n893_bF_buf1), .Y(u_sdrc_core_u_req_gen__abc_22171_n905) );
  OR2X2 OR2X2_1253 ( .A(u_sdrc_core_u_req_gen__abc_22171_n909), .B(u_sdrc_core_u_req_gen__abc_22171_n877), .Y(u_sdrc_core_u_req_gen__abc_22171_n910) );
  OR2X2 OR2X2_1254 ( .A(u_sdrc_core_u_req_gen__abc_22171_n910), .B(u_sdrc_core_u_req_gen__abc_22171_n908), .Y(u_sdrc_core_u_req_gen__abc_22171_n911) );
  OR2X2 OR2X2_1255 ( .A(u_sdrc_core_u_req_gen__abc_22171_n911), .B(u_sdrc_core_u_req_gen__abc_22171_n907), .Y(u_sdrc_core_u_req_gen__abc_22171_n912) );
  OR2X2 OR2X2_1256 ( .A(u_sdrc_core_u_req_gen_map_address_11_), .B(u_sdrc_core_u_req_gen__abc_22171_n893_bF_buf0), .Y(u_sdrc_core_u_req_gen__abc_22171_n913) );
  OR2X2 OR2X2_1257 ( .A(u_sdrc_core_u_req_gen__abc_22171_n917), .B(u_sdrc_core_u_req_gen__abc_22171_n877), .Y(u_sdrc_core_u_req_gen__abc_22171_n918) );
  OR2X2 OR2X2_1258 ( .A(u_sdrc_core_u_req_gen__abc_22171_n918), .B(u_sdrc_core_u_req_gen__abc_22171_n916), .Y(u_sdrc_core_u_req_gen__abc_22171_n919) );
  OR2X2 OR2X2_1259 ( .A(u_sdrc_core_u_req_gen__abc_22171_n919), .B(u_sdrc_core_u_req_gen__abc_22171_n915), .Y(u_sdrc_core_u_req_gen__abc_22171_n920) );
  OR2X2 OR2X2_126 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n223_1_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_len_1_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n498) );
  OR2X2 OR2X2_1260 ( .A(u_sdrc_core_u_req_gen_map_address_12_), .B(u_sdrc_core_u_req_gen__abc_22171_n893_bF_buf3), .Y(u_sdrc_core_u_req_gen__abc_22171_n921) );
  OR2X2 OR2X2_1261 ( .A(u_sdrc_core_u_req_gen__abc_22171_n926), .B(u_sdrc_core_u_req_gen__abc_22171_n925), .Y(u_sdrc_core_u_req_gen__abc_22171_n927) );
  OR2X2 OR2X2_1262 ( .A(u_sdrc_core_u_req_gen__abc_22171_n927), .B(u_sdrc_core_u_req_gen__abc_22171_n924), .Y(u_sdrc_core_u_req_gen__abc_22171_n928) );
  OR2X2 OR2X2_1263 ( .A(u_sdrc_core_u_req_gen__abc_22171_n928), .B(u_sdrc_core_u_req_gen__abc_22171_n923), .Y(u_sdrc_core_u_req_gen_r2b_raddr_3__FF_INPUT) );
  OR2X2 OR2X2_1264 ( .A(u_sdrc_core_u_req_gen__abc_22171_n932), .B(u_sdrc_core_u_req_gen__abc_22171_n877), .Y(u_sdrc_core_u_req_gen__abc_22171_n933) );
  OR2X2 OR2X2_1265 ( .A(u_sdrc_core_u_req_gen__abc_22171_n933), .B(u_sdrc_core_u_req_gen__abc_22171_n931), .Y(u_sdrc_core_u_req_gen__abc_22171_n934) );
  OR2X2 OR2X2_1266 ( .A(u_sdrc_core_u_req_gen__abc_22171_n934), .B(u_sdrc_core_u_req_gen__abc_22171_n930), .Y(u_sdrc_core_u_req_gen__abc_22171_n935) );
  OR2X2 OR2X2_1267 ( .A(u_sdrc_core_u_req_gen_map_address_14_), .B(u_sdrc_core_u_req_gen__abc_22171_n893_bF_buf2), .Y(u_sdrc_core_u_req_gen__abc_22171_n936) );
  OR2X2 OR2X2_1268 ( .A(u_sdrc_core_u_req_gen__abc_22171_n940), .B(u_sdrc_core_u_req_gen__abc_22171_n877), .Y(u_sdrc_core_u_req_gen__abc_22171_n941) );
  OR2X2 OR2X2_1269 ( .A(u_sdrc_core_u_req_gen__abc_22171_n941), .B(u_sdrc_core_u_req_gen__abc_22171_n939), .Y(u_sdrc_core_u_req_gen__abc_22171_n942) );
  OR2X2 OR2X2_127 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n499), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf2), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n500) );
  OR2X2 OR2X2_1270 ( .A(u_sdrc_core_u_req_gen__abc_22171_n942), .B(u_sdrc_core_u_req_gen__abc_22171_n938), .Y(u_sdrc_core_u_req_gen__abc_22171_n943) );
  OR2X2 OR2X2_1271 ( .A(u_sdrc_core_u_req_gen_map_address_15_), .B(u_sdrc_core_u_req_gen__abc_22171_n893_bF_buf1), .Y(u_sdrc_core_u_req_gen__abc_22171_n944) );
  OR2X2 OR2X2_1272 ( .A(u_sdrc_core_u_req_gen__abc_22171_n946), .B(u_sdrc_core_u_req_gen__abc_22171_n877), .Y(u_sdrc_core_u_req_gen__abc_22171_n947) );
  OR2X2 OR2X2_1273 ( .A(u_sdrc_core_u_req_gen__abc_22171_n948), .B(u_sdrc_core_u_req_gen__abc_22171_n949), .Y(u_sdrc_core_u_req_gen__abc_22171_n950) );
  OR2X2 OR2X2_1274 ( .A(u_sdrc_core_u_req_gen__abc_22171_n947), .B(u_sdrc_core_u_req_gen__abc_22171_n950), .Y(u_sdrc_core_u_req_gen__abc_22171_n951) );
  OR2X2 OR2X2_1275 ( .A(u_sdrc_core_u_req_gen_map_address_16_), .B(u_sdrc_core_u_req_gen__abc_22171_n893_bF_buf0), .Y(u_sdrc_core_u_req_gen__abc_22171_n952) );
  OR2X2 OR2X2_1276 ( .A(u_sdrc_core_u_req_gen__abc_22171_n956), .B(u_sdrc_core_u_req_gen__abc_22171_n877), .Y(u_sdrc_core_u_req_gen__abc_22171_n957) );
  OR2X2 OR2X2_1277 ( .A(u_sdrc_core_u_req_gen__abc_22171_n957), .B(u_sdrc_core_u_req_gen__abc_22171_n955), .Y(u_sdrc_core_u_req_gen__abc_22171_n958) );
  OR2X2 OR2X2_1278 ( .A(u_sdrc_core_u_req_gen__abc_22171_n958), .B(u_sdrc_core_u_req_gen__abc_22171_n954), .Y(u_sdrc_core_u_req_gen__abc_22171_n959) );
  OR2X2 OR2X2_1279 ( .A(u_sdrc_core_u_req_gen_map_address_17_), .B(u_sdrc_core_u_req_gen__abc_22171_n893_bF_buf3), .Y(u_sdrc_core_u_req_gen__abc_22171_n960) );
  OR2X2 OR2X2_128 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n283_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_len_1_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n501) );
  OR2X2 OR2X2_1280 ( .A(u_sdrc_core_u_req_gen__abc_22171_n964), .B(u_sdrc_core_u_req_gen__abc_22171_n877), .Y(u_sdrc_core_u_req_gen__abc_22171_n965) );
  OR2X2 OR2X2_1281 ( .A(u_sdrc_core_u_req_gen__abc_22171_n965), .B(u_sdrc_core_u_req_gen__abc_22171_n963), .Y(u_sdrc_core_u_req_gen__abc_22171_n966) );
  OR2X2 OR2X2_1282 ( .A(u_sdrc_core_u_req_gen__abc_22171_n966), .B(u_sdrc_core_u_req_gen__abc_22171_n962), .Y(u_sdrc_core_u_req_gen__abc_22171_n967) );
  OR2X2 OR2X2_1283 ( .A(u_sdrc_core_u_req_gen_map_address_18_), .B(u_sdrc_core_u_req_gen__abc_22171_n893_bF_buf2), .Y(u_sdrc_core_u_req_gen__abc_22171_n968) );
  OR2X2 OR2X2_1284 ( .A(u_sdrc_core_u_req_gen__abc_22171_n971), .B(u_sdrc_core_u_req_gen__abc_22171_n970), .Y(u_sdrc_core_u_req_gen__abc_22171_n972) );
  OR2X2 OR2X2_1285 ( .A(u_sdrc_core_u_req_gen__abc_22171_n973), .B(u_sdrc_core_u_req_gen__abc_22171_n974), .Y(u_sdrc_core_u_req_gen__abc_22171_n975) );
  OR2X2 OR2X2_1286 ( .A(u_sdrc_core_u_req_gen__abc_22171_n975), .B(u_sdrc_core_u_req_gen__abc_22171_n972), .Y(u_sdrc_core_u_req_gen_r2b_raddr_9__FF_INPUT) );
  OR2X2 OR2X2_1287 ( .A(u_sdrc_core_u_req_gen__abc_22171_n798), .B(u_sdrc_core_u_req_gen__abc_22171_n887), .Y(u_sdrc_core_u_req_gen__abc_22171_n977) );
  OR2X2 OR2X2_1288 ( .A(u_sdrc_core_u_req_gen__abc_22171_n813), .B(u_sdrc_core_u_req_gen__abc_22171_n886), .Y(u_sdrc_core_u_req_gen__abc_22171_n979) );
  OR2X2 OR2X2_1289 ( .A(u_sdrc_core_u_req_gen__abc_22171_n831), .B(u_sdrc_core_u_req_gen__abc_22171_n980), .Y(u_sdrc_core_u_req_gen__abc_22171_n981) );
  OR2X2 OR2X2_129 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n503), .B(u_sdrc_core_u_bank_ctl__abc_21249_n496), .Y(u_sdrc_core_b2x_len_1_) );
  OR2X2 OR2X2_1290 ( .A(u_sdrc_core_u_req_gen_map_address_20_), .B(u_sdrc_core_u_req_gen__abc_22171_n893_bF_buf0), .Y(u_sdrc_core_u_req_gen__abc_22171_n985) );
  OR2X2 OR2X2_1291 ( .A(u_sdrc_core_u_req_gen_map_address_21_), .B(u_sdrc_core_u_req_gen__abc_22171_n893_bF_buf3), .Y(u_sdrc_core_u_req_gen__abc_22171_n987) );
  OR2X2 OR2X2_1292 ( .A(u_sdrc_core_u_req_gen__abc_22171_n813), .B(u_sdrc_core_u_req_gen__abc_22171_n887), .Y(u_sdrc_core_u_req_gen__abc_22171_n988) );
  OR2X2 OR2X2_1293 ( .A(u_sdrc_core_u_req_gen__abc_22171_n831), .B(u_sdrc_core_u_req_gen__abc_22171_n886), .Y(u_sdrc_core_u_req_gen__abc_22171_n989) );
  OR2X2 OR2X2_1294 ( .A(u_sdrc_core_u_req_gen__abc_22171_n850), .B(u_sdrc_core_u_req_gen__abc_22171_n980), .Y(u_sdrc_core_u_req_gen__abc_22171_n991) );
  OR2X2 OR2X2_1295 ( .A(u_sdrc_core_u_req_gen__abc_22171_n869), .B(u_sdrc_core_u_req_gen__abc_22171_n980), .Y(u_sdrc_core_u_req_gen__abc_22171_n996) );
  OR2X2 OR2X2_1296 ( .A(u_sdrc_core_u_req_gen__abc_22171_n850), .B(u_sdrc_core_u_req_gen__abc_22171_n886), .Y(u_sdrc_core_u_req_gen__abc_22171_n998) );
  OR2X2 OR2X2_1297 ( .A(u_sdrc_core_u_req_gen__abc_22171_n831), .B(u_sdrc_core_u_req_gen__abc_22171_n887), .Y(u_sdrc_core_u_req_gen__abc_22171_n999) );
  OR2X2 OR2X2_1298 ( .A(u_sdrc_core_u_req_gen_map_address_22_), .B(u_sdrc_core_u_req_gen__abc_22171_n893_bF_buf0), .Y(u_sdrc_core_u_req_gen__abc_22171_n1003) );
  OR2X2 OR2X2_1299 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1007), .B(u_sdrc_core_u_req_gen_req_st_1_), .Y(u_sdrc_core_r2b_last) );
  OR2X2 OR2X2_13 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n241), .B(u_sdrc_core_u_bank_ctl__abc_21249_n239_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n242_1) );
  OR2X2 OR2X2_130 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_len_2_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n506) );
  OR2X2 OR2X2_1300 ( .A(u_sdrc_core_u_req_gen__abc_22171_n309), .B(u_sdrc_core_u_req_gen__abc_22171_n1009), .Y(u_sdrc_core_u_req_gen__abc_22171_n1012) );
  OR2X2 OR2X2_1301 ( .A(u_sdrc_core_u_req_gen__abc_22171_n391), .B(app_req_len_7_), .Y(u_sdrc_core_u_req_gen__abc_22171_n1014) );
  OR2X2 OR2X2_1302 ( .A(u_sdrc_core_u_req_gen__abc_22171_n241), .B(app_req_len_5_), .Y(u_sdrc_core_u_req_gen__abc_22171_n1015) );
  OR2X2 OR2X2_1303 ( .A(u_sdrc_core_u_req_gen__abc_22171_n416), .B(app_req_len_6_), .Y(u_sdrc_core_u_req_gen__abc_22171_n1016) );
  OR2X2 OR2X2_1304 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1024), .B(u_sdrc_core_u_req_gen__abc_22171_n1025), .Y(u_sdrc_core_u_req_gen__abc_22171_n1026) );
  OR2X2 OR2X2_1305 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1030), .B(u_sdrc_core_u_req_gen__abc_22171_n1031), .Y(u_sdrc_core_u_req_gen__abc_22171_n1032) );
  OR2X2 OR2X2_1306 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1032), .B(u_sdrc_core_u_req_gen__abc_22171_n1028), .Y(u_sdrc_core_u_req_gen__abc_22171_n1033) );
  OR2X2 OR2X2_1307 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1033), .B(u_sdrc_core_u_req_gen__abc_22171_n1027), .Y(u_sdrc_core_u_req_gen__abc_22171_n1034) );
  OR2X2 OR2X2_1308 ( .A(u_sdrc_core_u_req_gen__abc_22171_n278), .B(u_sdrc_core_u_req_gen__abc_22171_n1023), .Y(u_sdrc_core_u_req_gen__abc_22171_n1035) );
  OR2X2 OR2X2_1309 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1036), .B(u_sdrc_core_u_req_gen__abc_22171_n1037), .Y(u_sdrc_core_u_req_gen__abc_22171_n1038) );
  OR2X2 OR2X2_131 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n223_1_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_len_2_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n507) );
  OR2X2 OR2X2_1310 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1038), .B(u_sdrc_core_u_req_gen__abc_22171_n1034), .Y(u_sdrc_core_u_req_gen__abc_22171_n1039) );
  OR2X2 OR2X2_1311 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1039), .B(u_sdrc_core_u_req_gen__abc_22171_n1026), .Y(u_sdrc_core_u_req_gen__abc_22171_n1040) );
  OR2X2 OR2X2_1312 ( .A(u_sdrc_core_u_req_gen__abc_22171_n289), .B(u_sdrc_core_u_req_gen__abc_22171_n419), .Y(u_sdrc_core_u_req_gen__abc_22171_n1041) );
  OR2X2 OR2X2_1313 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1045), .B(u_sdrc_core_u_req_gen__abc_22171_n1031), .Y(u_sdrc_core_u_req_gen__abc_22171_n1046) );
  OR2X2 OR2X2_1314 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1047), .B(u_sdrc_core_u_req_gen__abc_22171_n1043), .Y(u_sdrc_core_u_req_gen__abc_22171_n1048) );
  OR2X2 OR2X2_1315 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1053), .B(u_sdrc_core_u_req_gen__abc_22171_n1051), .Y(u_sdrc_core_u_req_gen__abc_22171_n1054) );
  OR2X2 OR2X2_1316 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1050), .B(u_sdrc_core_u_req_gen__abc_22171_n1054), .Y(u_sdrc_core_u_req_gen__abc_22171_n1055) );
  OR2X2 OR2X2_1317 ( .A(u_sdrc_core_u_req_gen__abc_22171_n311), .B(u_sdrc_core_u_req_gen__abc_22171_n464_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n1056) );
  OR2X2 OR2X2_1318 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1052), .B(u_sdrc_core_u_req_gen__abc_22171_n442_1), .Y(u_sdrc_core_u_req_gen__abc_22171_n1057) );
  OR2X2 OR2X2_1319 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1059), .B(u_sdrc_core_u_req_gen__abc_22171_n1022), .Y(u_sdrc_core_u_req_gen__abc_22171_n1060) );
  OR2X2 OR2X2_132 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n508), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n509) );
  OR2X2 OR2X2_1320 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1068), .B(u_sdrc_core_u_req_gen__abc_22171_n1066), .Y(u_sdrc_core_u_req_gen__abc_22171_n1069) );
  OR2X2 OR2X2_1321 ( .A(u_sdrc_core_u_req_gen__abc_22171_n391), .B(app_req_len_8_), .Y(u_sdrc_core_u_req_gen__abc_22171_n1070) );
  OR2X2 OR2X2_1322 ( .A(u_sdrc_core_u_req_gen__abc_22171_n241), .B(app_req_len_6_), .Y(u_sdrc_core_u_req_gen__abc_22171_n1071) );
  OR2X2 OR2X2_1323 ( .A(u_sdrc_core_u_req_gen__abc_22171_n416), .B(app_req_len_7_), .Y(u_sdrc_core_u_req_gen__abc_22171_n1072) );
  OR2X2 OR2X2_1324 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1075), .B(u_sdrc_core_u_req_gen__abc_22171_n1063), .Y(u_sdrc_core_u_req_gen__abc_22171_n1076) );
  OR2X2 OR2X2_1325 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1061), .B(u_sdrc_core_u_req_gen__abc_22171_n1076), .Y(u_sdrc_core_u_req_gen__abc_22171_n1077) );
  OR2X2 OR2X2_1326 ( .A(u_sdrc_core_u_req_gen__abc_22171_n644), .B(u_sdrc_core_u_req_gen__abc_22171_n874), .Y(u_sdrc_core_u_req_gen__abc_22171_n1081) );
  OR2X2 OR2X2_1327 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1080), .B(u_sdrc_core_u_req_gen__abc_22171_n1081), .Y(u_sdrc_core_u_req_gen__abc_22171_n1084) );
  OR2X2 OR2X2_1328 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1085), .B(u_sdrc_core_u_req_gen__abc_22171_n876), .Y(u_sdrc_core_u_req_gen__abc_22171_n1086) );
  OR2X2 OR2X2_1329 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1097), .B(u_sdrc_core_u_req_gen__abc_22171_n1098), .Y(u_sdrc_core_u_req_gen__abc_22171_n1099) );
  OR2X2 OR2X2_133 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n283_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_len_2_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n510) );
  OR2X2 OR2X2_1330 ( .A(u_sdrc_core_u_req_gen__abc_22171_n1069), .B(u_sdrc_core_u_req_gen__abc_22171_n1074), .Y(u_sdrc_core_u_req_gen__abc_22171_n1100) );
  OR2X2 OR2X2_1331 ( .A(app_req_ack_bF_buf1), .B(u_sdrc_core_u_req_gen__abc_22171_n1105), .Y(u_sdrc_core_u_req_gen_r2b_start_FF_INPUT) );
  OR2X2 OR2X2_1332 ( .A(u_sdrc_core_u_xfr_ctl_tmr0_0_), .B(u_sdrc_core_u_xfr_ctl_tmr0_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n351_1) );
  OR2X2 OR2X2_1333 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n351_1), .B(u_sdrc_core_u_xfr_ctl_tmr0_2_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n352) );
  OR2X2 OR2X2_1334 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n352), .B(u_sdrc_core_u_xfr_ctl_tmr0_3_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n353_1) );
  OR2X2 OR2X2_1335 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n369_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n371), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n372_1) );
  OR2X2 OR2X2_1336 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n368), .B(\cfg_sdr_rfmax[1] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n373) );
  OR2X2 OR2X2_1337 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n366), .B(\cfg_sdr_rfmax[2] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n374_1) );
  OR2X2 OR2X2_1338 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n376), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n367_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n377_1) );
  OR2X2 OR2X2_1339 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n382_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n380_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n383) );
  OR2X2 OR2X2_134 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n512), .B(u_sdrc_core_u_bank_ctl__abc_21249_n505), .Y(u_sdrc_core_b2x_len_2_) );
  OR2X2 OR2X2_1340 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n383), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n365_1), .Y(u_sdrc_core_u_xfr_ctl__abc_16728_n35) );
  OR2X2 OR2X2_1341 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n401_1), .B(u_sdrc_core_u_xfr_ctl_mgmt_st_3_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n402_1) );
  OR2X2 OR2X2_1342 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n402_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n395), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n403_1) );
  OR2X2 OR2X2_1343 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n408_1), .B(u_sdrc_core_u_xfr_ctl_mgmt_st_2_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n409_1) );
  OR2X2 OR2X2_1344 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n407_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n411_1), .Y(u_sdrc_core_u_xfr_ctl__abc_16728_n43) );
  OR2X2 OR2X2_1345 ( .A(u_sdrc_core_u_xfr_ctl_mgmt_st_7_), .B(u_sdrc_core_u_xfr_ctl_mgmt_st_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n415) );
  OR2X2 OR2X2_1346 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n416_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n413_1), .Y(u_sdrc_core_u_xfr_ctl__abc_16728_n178) );
  OR2X2 OR2X2_1347 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n421), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n419), .Y(u_sdrc_core_u_xfr_ctl__abc_16728_n181) );
  OR2X2 OR2X2_1348 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n423), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n426), .Y(u_sdrc_core_u_xfr_ctl__abc_16728_n184) );
  OR2X2 OR2X2_1349 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n434_1), .B(u_sdrc_core_u_xfr_ctl_mgmt_st_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n435) );
  OR2X2 OR2X2_135 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_len_3_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n515) );
  OR2X2 OR2X2_1350 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n436_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n432_1), .Y(u_sdrc_core_u_xfr_ctl__abc_16728_n189) );
  OR2X2 OR2X2_1351 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n439), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n438_1), .Y(u_sdrc_core_u_xfr_ctl__abc_16728_n258) );
  OR2X2 OR2X2_1352 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n441), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n442_1), .Y(u_sdrc_core_u_xfr_ctl__abc_16728_n270) );
  OR2X2 OR2X2_1353 ( .A(u_sdrc_core_b2x_ba_1_), .B(u_sdrc_core_u_bank_ctl_xfr_bank_sel_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n466_1) );
  OR2X2 OR2X2_1354 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n475), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n476), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n477) );
  OR2X2 OR2X2_1355 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n480), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n465_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n481) );
  OR2X2 OR2X2_1356 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n482), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n486), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n487) );
  OR2X2 OR2X2_1357 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n488_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n446_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n489_1) );
  OR2X2 OR2X2_1358 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n496_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n386), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n497_1) );
  OR2X2 OR2X2_1359 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n499_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n502), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n503) );
  OR2X2 OR2X2_136 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n223_1_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_len_3_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n516) );
  OR2X2 OR2X2_1360 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n490_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n503), .Y(u_sdrc_core_u_bank_ctl_x2b_ack) );
  OR2X2 OR2X2_1361 ( .A(u_sdrc_core_u_bank_ctl_xfr_bank_sel_0_), .B(u_sdrc_core_b2x_ba_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n509) );
  OR2X2 OR2X2_1362 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n511_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n508), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n512_1) );
  OR2X2 OR2X2_1363 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n512_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n469_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n513_1) );
  OR2X2 OR2X2_1364 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n513_1), .B(u_sdrc_core_u_xfr_ctl_l_wrap), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n514) );
  OR2X2 OR2X2_1365 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n515), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n387_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n516_1) );
  OR2X2 OR2X2_1366 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n518_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n491_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n519) );
  OR2X2 OR2X2_1367 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n520_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n505_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n521_1) );
  OR2X2 OR2X2_1368 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n526_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_pre_ok), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n527) );
  OR2X2 OR2X2_1369 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n527), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n528), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n529_1) );
  OR2X2 OR2X2_137 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n517), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf0), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n518) );
  OR2X2 OR2X2_1370 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n530_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n532), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n533_1) );
  OR2X2 OR2X2_1371 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n429), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n396_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n535) );
  OR2X2 OR2X2_1372 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n405_1_bF_buf1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n536_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n537) );
  OR2X2 OR2X2_1373 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n538), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n539_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n540_1) );
  OR2X2 OR2X2_1374 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n534_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n540_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n541) );
  OR2X2 OR2X2_1375 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n399_1), .B(u_sdrc_core_u_xfr_ctl_mgmt_st_4_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n542_1) );
  OR2X2 OR2X2_1376 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n405_1_bF_buf0), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n542_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n543) );
  OR2X2 OR2X2_1377 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n551_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n546_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n552_1) );
  OR2X2 OR2X2_1378 ( .A(u_sdrc_core_u_xfr_ctl_l_rd_next_1_), .B(u_sdrc_core_u_xfr_ctl_l_rd_next_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n556) );
  OR2X2 OR2X2_1379 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n568), .B(u_sdrc_core_u_xfr_ctl_l_rd_next_4_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n569_1) );
  OR2X2 OR2X2_138 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n283_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_len_3_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n519) );
  OR2X2 OR2X2_1380 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n573), .B(u_sdrc_core_u_xfr_ctl_l_rd_next_2_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n574) );
  OR2X2 OR2X2_1381 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n570_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n574), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n575_1) );
  OR2X2 OR2X2_1382 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n576_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n556), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n577) );
  OR2X2 OR2X2_1383 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n581_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n580), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n582_1) );
  OR2X2 OR2X2_1384 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n578_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n582_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n583) );
  OR2X2 OR2X2_1385 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n584_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n552_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n585) );
  OR2X2 OR2X2_1386 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n491_1), .B(_auto_iopadmap_cc_313_execute_24701), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n587_1) );
  OR2X2 OR2X2_1387 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n589), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n446_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n590_1) );
  OR2X2 OR2X2_1388 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n591), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n592), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n593_1) );
  OR2X2 OR2X2_1389 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n593_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n588_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n594_1) );
  OR2X2 OR2X2_139 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n521), .B(u_sdrc_core_u_bank_ctl__abc_21249_n514), .Y(u_sdrc_core_b2x_len_3_) );
  OR2X2 OR2X2_1390 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n594_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n578_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n595) );
  OR2X2 OR2X2_1391 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n577), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n506_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n600_1) );
  OR2X2 OR2X2_1392 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n600_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n599_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n601) );
  OR2X2 OR2X2_1393 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n604_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n387_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n605) );
  OR2X2 OR2X2_1394 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n607), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n597), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n608) );
  OR2X2 OR2X2_1395 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n523_1_bF_buf2), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n461_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1) );
  OR2X2 OR2X2_1396 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n610_1), .B(u_sdrc_core_u_xfr_ctl_xfr_caddr_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n611) );
  OR2X2 OR2X2_1397 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n613), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n615), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n616) );
  OR2X2 OR2X2_1398 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n610_1), .B(u_sdrc_core_u_xfr_ctl_xfr_caddr_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n618_1) );
  OR2X2 OR2X2_1399 ( .A(u_sdrc_core_u_xfr_ctl_xfr_caddr_1_), .B(u_sdrc_core_u_xfr_ctl_xfr_caddr_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n620_1) );
  OR2X2 OR2X2_14 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n246_1), .B(u_sdrc_core_u_bank_ctl_rank_cnt_0_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n247_1) );
  OR2X2 OR2X2_140 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_len_4_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n524) );
  OR2X2 OR2X2_1400 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n607), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n621), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n622) );
  OR2X2 OR2X2_1401 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n624), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n625_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n626) );
  OR2X2 OR2X2_1402 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n610_1), .B(u_sdrc_core_u_xfr_ctl_xfr_caddr_2_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n628_1) );
  OR2X2 OR2X2_1403 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n492_1), .B(u_sdrc_core_u_xfr_ctl_xfr_caddr_2_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n631) );
  OR2X2 OR2X2_1404 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n607), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n632), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n633) );
  OR2X2 OR2X2_1405 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n635_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n636), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n637) );
  OR2X2 OR2X2_1406 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n610_1), .B(u_sdrc_core_u_xfr_ctl_xfr_caddr_3_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n639_1) );
  OR2X2 OR2X2_1407 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n629), .B(u_sdrc_core_u_xfr_ctl_xfr_caddr_3_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n642) );
  OR2X2 OR2X2_1408 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n607), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n643), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n644) );
  OR2X2 OR2X2_1409 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n646_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n647), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n648) );
  OR2X2 OR2X2_141 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n223_1_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_len_4_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n525) );
  OR2X2 OR2X2_1410 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n610_1), .B(u_sdrc_core_u_xfr_ctl_xfr_caddr_4_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n650) );
  OR2X2 OR2X2_1411 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n640), .B(u_sdrc_core_u_xfr_ctl_xfr_caddr_4_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n653_1) );
  OR2X2 OR2X2_1412 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n607), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n654), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n655) );
  OR2X2 OR2X2_1413 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n657_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n658), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n659) );
  OR2X2 OR2X2_1414 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n610_1), .B(u_sdrc_core_u_xfr_ctl_xfr_caddr_5_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n661) );
  OR2X2 OR2X2_1415 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n651), .B(u_sdrc_core_u_xfr_ctl_xfr_caddr_5_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n664) );
  OR2X2 OR2X2_1416 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n607), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n665), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n666) );
  OR2X2 OR2X2_1417 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n668), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n669), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n670) );
  OR2X2 OR2X2_1418 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n610_1), .B(u_sdrc_core_u_xfr_ctl_xfr_caddr_6_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n672_1) );
  OR2X2 OR2X2_1419 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n662), .B(u_sdrc_core_u_xfr_ctl_xfr_caddr_6_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n675) );
  OR2X2 OR2X2_142 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n526), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf4), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n527) );
  OR2X2 OR2X2_1420 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n607), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n676), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n677_1) );
  OR2X2 OR2X2_1421 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n679), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n680), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n681) );
  OR2X2 OR2X2_1422 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n610_1), .B(u_sdrc_core_u_xfr_ctl_xfr_caddr_7_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n683) );
  OR2X2 OR2X2_1423 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n673), .B(u_sdrc_core_u_xfr_ctl_xfr_caddr_7_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n686_1) );
  OR2X2 OR2X2_1424 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n607), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n687), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n688_1) );
  OR2X2 OR2X2_1425 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n690), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n691), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n692_1) );
  OR2X2 OR2X2_1426 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n610_1), .B(u_sdrc_core_u_xfr_ctl_xfr_caddr_8_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n694) );
  OR2X2 OR2X2_1427 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n684_1), .B(u_sdrc_core_u_xfr_ctl_xfr_caddr_8_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n697) );
  OR2X2 OR2X2_1428 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n607), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n698), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n699) );
  OR2X2 OR2X2_1429 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n701_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n702), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n703_1) );
  OR2X2 OR2X2_143 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n283_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_len_4_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n528) );
  OR2X2 OR2X2_1430 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n610_1), .B(u_sdrc_core_u_xfr_ctl_xfr_caddr_9_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n705) );
  OR2X2 OR2X2_1431 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n695_1), .B(u_sdrc_core_u_xfr_ctl_xfr_caddr_9_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n708_1) );
  OR2X2 OR2X2_1432 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n607), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n709), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n710_1) );
  OR2X2 OR2X2_1433 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n712), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n713), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n714) );
  OR2X2 OR2X2_1434 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n610_1), .B(u_sdrc_core_u_xfr_ctl_xfr_caddr_10_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n716_1) );
  OR2X2 OR2X2_1435 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n706), .B(u_sdrc_core_u_xfr_ctl_xfr_caddr_10_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n719_1) );
  OR2X2 OR2X2_1436 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n607), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n720), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n721) );
  OR2X2 OR2X2_1437 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n723_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n724), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n725_1) );
  OR2X2 OR2X2_1438 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n610_1), .B(u_sdrc_core_u_xfr_ctl_xfr_caddr_11_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n727) );
  OR2X2 OR2X2_1439 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n717), .B(u_sdrc_core_u_xfr_ctl_xfr_caddr_11_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n730) );
  OR2X2 OR2X2_144 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n530), .B(u_sdrc_core_u_bank_ctl__abc_21249_n523), .Y(u_sdrc_core_b2x_len_4_) );
  OR2X2 OR2X2_1440 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n607), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n731), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n732) );
  OR2X2 OR2X2_1441 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n734), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n735), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n736_1) );
  OR2X2 OR2X2_1442 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n610_1), .B(u_sdrc_core_u_xfr_ctl_xfr_caddr_12_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n738) );
  OR2X2 OR2X2_1443 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n728), .B(u_sdrc_core_u_xfr_ctl_xfr_caddr_12_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n739) );
  OR2X2 OR2X2_1444 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n607), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n742), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n743) );
  OR2X2 OR2X2_1445 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n745), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n746), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n747) );
  OR2X2 OR2X2_1446 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n765), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n766), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n767) );
  OR2X2 OR2X2_1447 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n769), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n770), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n771_1) );
  OR2X2 OR2X2_1448 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n614_bF_buf0), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n457), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n774) );
  OR2X2 OR2X2_1449 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n774), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n773), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n775_1) );
  OR2X2 OR2X2_145 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_len_5_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n533) );
  OR2X2 OR2X2_1450 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf4), .B(u_sdrc_core_b2x_len_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n776) );
  OR2X2 OR2X2_1451 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf3), .B(u_sdrc_core_b2x_len_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n779) );
  OR2X2 OR2X2_1452 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n780), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n781_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n782) );
  OR2X2 OR2X2_1453 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n614_bF_buf3), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n782), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n783) );
  OR2X2 OR2X2_1454 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n788_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n786), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n789_1) );
  OR2X2 OR2X2_1455 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n614_bF_buf2), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n789_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n790) );
  OR2X2 OR2X2_1456 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf2), .B(u_sdrc_core_b2x_len_2_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n791) );
  OR2X2 OR2X2_1457 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n796), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n794_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n797) );
  OR2X2 OR2X2_1458 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n798_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n799_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n800) );
  OR2X2 OR2X2_1459 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n804_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n802), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n805_1) );
  OR2X2 OR2X2_146 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n223_1_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_len_5_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n534) );
  OR2X2 OR2X2_1460 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n806_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n807_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n808_1) );
  OR2X2 OR2X2_1461 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n812_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n810_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n813_1) );
  OR2X2 OR2X2_1462 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n814_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n815_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n816_1) );
  OR2X2 OR2X2_1463 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n820_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n821_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n822_1) );
  OR2X2 OR2X2_1464 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n823_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n818_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n824_1) );
  OR2X2 OR2X2_1465 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n614_bF_buf1), .B(u_sdrc_core_u_xfr_ctl_l_last), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n843_1) );
  OR2X2 OR2X2_1466 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf2), .B(u_sdrc_core_b2x_last), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n844_1) );
  OR2X2 OR2X2_1467 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n848_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n849_1) );
  OR2X2 OR2X2_1468 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf0), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n854), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n855_1) );
  OR2X2 OR2X2_1469 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n609_1_bF_buf4), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n858), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n859_1) );
  OR2X2 OR2X2_147 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n535), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf3), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n536) );
  OR2X2 OR2X2_1470 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n458), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_pre_ok), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n869_1) );
  OR2X2 OR2X2_1471 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n875), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n877), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n878) );
  OR2X2 OR2X2_1472 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n433), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n878), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n879) );
  OR2X2 OR2X2_1473 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n874), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n879), .Y(u_sdrc_core_u_xfr_ctl_sdr_cke_FF_INPUT) );
  OR2X2 OR2X2_1474 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n882), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n538), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n883) );
  OR2X2 OR2X2_1475 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n883_bF_buf3), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n413_1), .Y(u_sdrc_core_u_xfr_ctl_sdr_cs_n_FF_INPUT) );
  OR2X2 OR2X2_1476 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n885), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n404_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n886) );
  OR2X2 OR2X2_1477 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n869_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n494_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n890) );
  OR2X2 OR2X2_1478 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n892), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n413_1), .Y(u_sdrc_core_u_xfr_ctl_sdr_cas_n_FF_INPUT) );
  OR2X2 OR2X2_1479 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n541), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n413_1), .Y(u_sdrc_core_u_xfr_ctl_sdr_we_n_FF_INPUT) );
  OR2X2 OR2X2_148 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n283_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_len_5_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n537) );
  OR2X2 OR2X2_1480 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n897), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n552_1), .Y(u_sdrc_core_u_bs_convert_x2a_wrnext) );
  OR2X2 OR2X2_1481 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n899), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n413_1), .Y(u_sdrc_core_u_xfr_ctl_sdr_dqm_0__FF_INPUT) );
  OR2X2 OR2X2_1482 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n901), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n413_1), .Y(u_sdrc_core_u_xfr_ctl_sdr_dqm_1__FF_INPUT) );
  OR2X2 OR2X2_1483 ( .A(u_sdrc_core_u_bank_ctl_x2b_ack_bF_buf3), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n905), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n906) );
  OR2X2 OR2X2_1484 ( .A(u_sdrc_core_u_bank_ctl_x2b_ack_bF_buf2), .B(u_sdrc_core_u_bank_ctl_xfr_bank_sel_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n907) );
  OR2X2 OR2X2_1485 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n523_1_bF_buf0), .B(u_sdrc_core_b2x_ba_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n908) );
  OR2X2 OR2X2_1486 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n914), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n910), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n915) );
  OR2X2 OR2X2_1487 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n915), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n904), .Y(u_sdrc_core_u_xfr_ctl_sdr_ba_0__FF_INPUT) );
  OR2X2 OR2X2_1488 ( .A(u_sdrc_core_u_bank_ctl_x2b_ack_bF_buf1), .B(u_sdrc_core_u_bank_ctl_xfr_bank_sel_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n918) );
  OR2X2 OR2X2_1489 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n523_1_bF_buf3), .B(u_sdrc_core_b2x_ba_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n919) );
  OR2X2 OR2X2_149 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n539), .B(u_sdrc_core_u_bank_ctl__abc_21249_n532), .Y(u_sdrc_core_b2x_len_5_) );
  OR2X2 OR2X2_1490 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n917), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n921), .Y(u_sdrc_core_u_xfr_ctl_sdr_ba_1__FF_INPUT) );
  OR2X2 OR2X2_1491 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n924), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n923), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n925) );
  OR2X2 OR2X2_1492 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n883_bF_buf3), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n927), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n928) );
  OR2X2 OR2X2_1493 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n928), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n926), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n929) );
  OR2X2 OR2X2_1494 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n911), .B(_auto_iopadmap_cc_313_execute_24675_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n930) );
  OR2X2 OR2X2_1495 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n932), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n933), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n934) );
  OR2X2 OR2X2_1496 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n883_bF_buf2), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n936), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n937) );
  OR2X2 OR2X2_1497 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n937), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n935), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n938) );
  OR2X2 OR2X2_1498 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n911), .B(_auto_iopadmap_cc_313_execute_24675_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n939) );
  OR2X2 OR2X2_1499 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n941), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n942), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n943) );
  OR2X2 OR2X2_15 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n245_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n217_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n248) );
  OR2X2 OR2X2_150 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_len_6_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n542) );
  OR2X2 OR2X2_1500 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n883_bF_buf1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n945), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n946) );
  OR2X2 OR2X2_1501 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n946), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n944), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n947) );
  OR2X2 OR2X2_1502 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n911), .B(_auto_iopadmap_cc_313_execute_24675_2_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n948) );
  OR2X2 OR2X2_1503 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n950), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n951), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n952) );
  OR2X2 OR2X2_1504 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n883_bF_buf0), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n954), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n955) );
  OR2X2 OR2X2_1505 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n955), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n953), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n956) );
  OR2X2 OR2X2_1506 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n911), .B(_auto_iopadmap_cc_313_execute_24675_3_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n957) );
  OR2X2 OR2X2_1507 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n959), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n960), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n961) );
  OR2X2 OR2X2_1508 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n883_bF_buf3), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n963), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n964) );
  OR2X2 OR2X2_1509 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n964), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n962), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n965) );
  OR2X2 OR2X2_151 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n223_1_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_len_6_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n543) );
  OR2X2 OR2X2_1510 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n911), .B(_auto_iopadmap_cc_313_execute_24675_4_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n966) );
  OR2X2 OR2X2_1511 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n968), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n969), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n970) );
  OR2X2 OR2X2_1512 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n883_bF_buf2), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n972), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n973) );
  OR2X2 OR2X2_1513 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n973), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n971), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n974) );
  OR2X2 OR2X2_1514 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n911), .B(_auto_iopadmap_cc_313_execute_24675_5_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n975) );
  OR2X2 OR2X2_1515 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n977), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n978), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n979) );
  OR2X2 OR2X2_1516 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n883_bF_buf1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n981), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n982) );
  OR2X2 OR2X2_1517 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n982), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n980), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n983) );
  OR2X2 OR2X2_1518 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n911), .B(_auto_iopadmap_cc_313_execute_24675_6_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n984) );
  OR2X2 OR2X2_1519 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n986), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n987), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n988) );
  OR2X2 OR2X2_152 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n544), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf2), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n545) );
  OR2X2 OR2X2_1520 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n883_bF_buf0), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n990), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n991) );
  OR2X2 OR2X2_1521 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n991), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n989), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n992) );
  OR2X2 OR2X2_1522 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n911), .B(_auto_iopadmap_cc_313_execute_24675_7_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n993) );
  OR2X2 OR2X2_1523 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n995), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n996), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n997) );
  OR2X2 OR2X2_1524 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n883_bF_buf3), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n999), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1000) );
  OR2X2 OR2X2_1525 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1000), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n998), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1001) );
  OR2X2 OR2X2_1526 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n911), .B(_auto_iopadmap_cc_313_execute_24675_8_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1002) );
  OR2X2 OR2X2_1527 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1004), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1005), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1006) );
  OR2X2 OR2X2_1528 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n883_bF_buf2), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1008), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1009) );
  OR2X2 OR2X2_1529 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1009), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1007), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1010) );
  OR2X2 OR2X2_153 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n283_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_len_6_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n546) );
  OR2X2 OR2X2_1530 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n911), .B(_auto_iopadmap_cc_313_execute_24675_9_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1011) );
  OR2X2 OR2X2_1531 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1013), .B(\cfg_sdr_mode_reg[10] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1014) );
  OR2X2 OR2X2_1532 ( .A(u_sdrc_core_u_bank_ctl_x2b_ack_bF_buf2), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n720), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1015) );
  OR2X2 OR2X2_1533 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n523_1_bF_buf0), .B(u_sdrc_core_b2x_addr_10_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1016) );
  OR2X2 OR2X2_1534 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1017), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n404_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1018) );
  OR2X2 OR2X2_1535 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1019), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n883_bF_buf1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1020) );
  OR2X2 OR2X2_1536 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n911), .B(_auto_iopadmap_cc_313_execute_24675_10_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1021) );
  OR2X2 OR2X2_1537 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n523_1_bF_buf3), .B(u_sdrc_core_b2x_addr_11_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1023) );
  OR2X2 OR2X2_1538 ( .A(u_sdrc_core_u_bank_ctl_x2b_ack_bF_buf1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n731), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1024) );
  OR2X2 OR2X2_1539 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n914), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1028), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1029) );
  OR2X2 OR2X2_154 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n548), .B(u_sdrc_core_u_bank_ctl__abc_21249_n541), .Y(u_sdrc_core_b2x_len_6_) );
  OR2X2 OR2X2_1540 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1029), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1027), .Y(u_sdrc_core_u_xfr_ctl_sdr_addr_11__FF_INPUT) );
  OR2X2 OR2X2_1541 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n742), .B(u_sdrc_core_u_bank_ctl_x2b_ack_bF_buf0), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1031) );
  OR2X2 OR2X2_1542 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n523_1_bF_buf2), .B(u_sdrc_core_b2x_addr_12_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1032) );
  OR2X2 OR2X2_1543 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n883_bF_buf3), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1035), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1036) );
  OR2X2 OR2X2_1544 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1036), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1034), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1037) );
  OR2X2 OR2X2_1545 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n911), .B(_auto_iopadmap_cc_313_execute_24675_12_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1038) );
  OR2X2 OR2X2_1546 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1046), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1048), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1049) );
  OR2X2 OR2X2_1547 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1049), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1044), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1050) );
  OR2X2 OR2X2_1548 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1055), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1051), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1056) );
  OR2X2 OR2X2_1549 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1058), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1059), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1060) );
  OR2X2 OR2X2_155 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_cmd_0_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n551) );
  OR2X2 OR2X2_1550 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1063), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1064), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1065) );
  OR2X2 OR2X2_1551 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1065), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1044), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1066) );
  OR2X2 OR2X2_1552 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1062), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1067), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1068) );
  OR2X2 OR2X2_1553 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1072), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1070), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1073) );
  OR2X2 OR2X2_1554 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1075), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1076), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1077) );
  OR2X2 OR2X2_1555 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1077), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1044), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1078) );
  OR2X2 OR2X2_1556 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1074), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1079), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1080) );
  OR2X2 OR2X2_1557 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1082), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1083), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1084) );
  OR2X2 OR2X2_1558 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1087), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1085), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1088) );
  OR2X2 OR2X2_1559 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1090), .B(u_sdrc_core_u_xfr_ctl_mgmt_st_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1091) );
  OR2X2 OR2X2_156 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n223_1_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_cmd_0_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n552) );
  OR2X2 OR2X2_1560 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1094), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1095), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1096) );
  OR2X2 OR2X2_1561 ( .A(u_sdrc_core_u_xfr_ctl_mgmt_st_1_), .B(u_sdrc_core_u_xfr_ctl_mgmt_st_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1098) );
  OR2X2 OR2X2_1562 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n402_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1098), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1099) );
  OR2X2 OR2X2_1563 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1099), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1100), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1101) );
  OR2X2 OR2X2_1564 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1102), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n413_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1103) );
  OR2X2 OR2X2_1565 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1097), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1103), .Y(u_sdrc_core_u_xfr_ctl_cntr1_0__FF_INPUT) );
  OR2X2 OR2X2_1566 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1106), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1107), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1108) );
  OR2X2 OR2X2_1567 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1099), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1110), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1111) );
  OR2X2 OR2X2_1568 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1112), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n413_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1113) );
  OR2X2 OR2X2_1569 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1109), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1113), .Y(u_sdrc_core_u_xfr_ctl_cntr1_1__FF_INPUT) );
  OR2X2 OR2X2_157 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n553), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n554) );
  OR2X2 OR2X2_1570 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1116), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1117), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1118) );
  OR2X2 OR2X2_1571 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1099), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1120), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1121) );
  OR2X2 OR2X2_1572 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1122), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n413_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1123) );
  OR2X2 OR2X2_1573 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1119), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1123), .Y(u_sdrc_core_u_xfr_ctl_cntr1_2__FF_INPUT) );
  OR2X2 OR2X2_1574 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1126), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1127), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1128) );
  OR2X2 OR2X2_1575 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1129), .B(u_sdrc_core_u_xfr_ctl_mgmt_st_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1130) );
  OR2X2 OR2X2_1576 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1133), .B(u_sdrc_core_u_xfr_ctl_rfsh_timer_5_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1134) );
  OR2X2 OR2X2_1577 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1135), .B(\cfg_sdr_rfsh[5] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1136) );
  OR2X2 OR2X2_1578 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1138), .B(u_sdrc_core_u_xfr_ctl_rfsh_timer_4_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1139) );
  OR2X2 OR2X2_1579 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1140), .B(\cfg_sdr_rfsh[4] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1141) );
  OR2X2 OR2X2_158 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n283_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_cmd_0_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n555) );
  OR2X2 OR2X2_1580 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1144), .B(u_sdrc_core_u_xfr_ctl_rfsh_timer_7_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1145) );
  OR2X2 OR2X2_1581 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1146), .B(\cfg_sdr_rfsh[7] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1147) );
  OR2X2 OR2X2_1582 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1150), .B(u_sdrc_core_u_xfr_ctl_rfsh_timer_11_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1151) );
  OR2X2 OR2X2_1583 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1152), .B(\cfg_sdr_rfsh[11] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1153) );
  OR2X2 OR2X2_1584 ( .A(\cfg_sdr_rfsh[9] ), .B(u_sdrc_core_u_xfr_ctl_rfsh_timer_9_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1155) );
  OR2X2 OR2X2_1585 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1163), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1160), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1164) );
  OR2X2 OR2X2_1586 ( .A(\cfg_sdr_rfsh[3] ), .B(u_sdrc_core_u_xfr_ctl_rfsh_timer_3_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1168) );
  OR2X2 OR2X2_1587 ( .A(\cfg_sdr_rfsh[1] ), .B(u_sdrc_core_u_xfr_ctl_rfsh_timer_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1173) );
  OR2X2 OR2X2_1588 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1180), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1178), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1181) );
  OR2X2 OR2X2_1589 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1184), .B(u_sdrc_core_u_xfr_ctl_rfsh_timer_2_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1185) );
  OR2X2 OR2X2_159 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n557), .B(u_sdrc_core_u_bank_ctl__abc_21249_n550), .Y(u_sdrc_core_b2x_cmd_0_) );
  OR2X2 OR2X2_1590 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1186), .B(\cfg_sdr_rfsh[2] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1187) );
  OR2X2 OR2X2_1591 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1192), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1189), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1193) );
  OR2X2 OR2X2_1592 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1197), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1194), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1198) );
  OR2X2 OR2X2_1593 ( .A(u_sdrc_core_u_xfr_ctl_rfsh_timer_0_), .B(u_sdrc_core_u_xfr_ctl_rfsh_timer_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1206) );
  OR2X2 OR2X2_1594 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1207), .B(u_sdrc_core_u_xfr_ctl_rfsh_timer_2_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1211) );
  OR2X2 OR2X2_1595 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1212), .B(u_sdrc_core_u_xfr_ctl_rfsh_timer_3_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1216) );
  OR2X2 OR2X2_1596 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1217), .B(u_sdrc_core_u_xfr_ctl_rfsh_timer_4_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1221) );
  OR2X2 OR2X2_1597 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1222), .B(u_sdrc_core_u_xfr_ctl_rfsh_timer_5_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1226) );
  OR2X2 OR2X2_1598 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1227), .B(u_sdrc_core_u_xfr_ctl_rfsh_timer_6_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1231) );
  OR2X2 OR2X2_1599 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1232), .B(u_sdrc_core_u_xfr_ctl_rfsh_timer_7_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1238) );
  OR2X2 OR2X2_16 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n252_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n257), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n258_1) );
  OR2X2 OR2X2_160 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n594), .B(u_sdrc_core_u_bank_ctl__abc_21249_n595), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n596) );
  OR2X2 OR2X2_1600 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1236), .B(u_sdrc_core_u_xfr_ctl_rfsh_timer_8_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1243) );
  OR2X2 OR2X2_1601 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1241), .B(u_sdrc_core_u_xfr_ctl_rfsh_timer_9_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1248) );
  OR2X2 OR2X2_1602 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1246), .B(u_sdrc_core_u_xfr_ctl_rfsh_timer_10_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1253) );
  OR2X2 OR2X2_1603 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1256), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1257), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1258) );
  OR2X2 OR2X2_1604 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1202), .B(u_sdrc_core_u_xfr_ctl_rfsh_row_cnt_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1262) );
  OR2X2 OR2X2_1605 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1260), .B(u_sdrc_core_u_xfr_ctl_rfsh_row_cnt_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1267) );
  OR2X2 OR2X2_1606 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1265), .B(u_sdrc_core_u_xfr_ctl_rfsh_row_cnt_2_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1272) );
  OR2X2 OR2X2_1607 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n567), .B(u_sdrc_core_u_xfr_ctl_l_rd_next_5_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1275) );
  OR2X2 OR2X2_1608 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n566_1), .B(u_sdrc_core_u_xfr_ctl_l_rd_next_6_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1276) );
  OR2X2 OR2X2_1609 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1277), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n562), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1278) );
  OR2X2 OR2X2_161 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n597), .B(u_sdrc_core_u_bank_ctl__abc_21249_n598), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n599) );
  OR2X2 OR2X2_1610 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n572_1), .B(u_sdrc_core_u_xfr_ctl_l_rd_next_3_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1279) );
  OR2X2 OR2X2_1611 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n563_1), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n564_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1280) );
  OR2X2 OR2X2_1612 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1280), .B(u_sdrc_core_u_xfr_ctl_l_rd_next_4_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1281) );
  OR2X2 OR2X2_1613 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1283), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n560_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1284) );
  OR2X2 OR2X2_1614 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n561), .B(u_sdrc_core_u_xfr_ctl_l_rd_next_2_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1285) );
  OR2X2 OR2X2_1615 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n567), .B(u_sdrc_core_u_xfr_ctl_l_rd_last_5_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1287) );
  OR2X2 OR2X2_1616 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n566_1), .B(u_sdrc_core_u_xfr_ctl_l_rd_last_6_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1288) );
  OR2X2 OR2X2_1617 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n571), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1291), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1292) );
  OR2X2 OR2X2_1618 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1290), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1292), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1293) );
  OR2X2 OR2X2_1619 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n572_1), .B(u_sdrc_core_u_xfr_ctl_l_rd_last_3_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1294) );
  OR2X2 OR2X2_162 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n599), .B(u_sdrc_core_u_bank_ctl__abc_21249_n596), .Y(u_sdrc_core_b2x_last) );
  OR2X2 OR2X2_1620 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1296), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1297), .Y(app_last_rd) );
  OR2X2 OR2X2_1621 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n602_bF_buf2), .B(u_sdrc_core_a2x_wrdt_0_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1311) );
  OR2X2 OR2X2_1622 ( .A(u_sdrc_core_u_bs_convert_x2a_wrnext_bF_buf2), .B(\sdr_dq[0] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1312) );
  OR2X2 OR2X2_1623 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n602_bF_buf1), .B(u_sdrc_core_a2x_wrdt_1_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1314) );
  OR2X2 OR2X2_1624 ( .A(u_sdrc_core_u_bs_convert_x2a_wrnext_bF_buf1), .B(\sdr_dq[1] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1315) );
  OR2X2 OR2X2_1625 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n602_bF_buf0), .B(u_sdrc_core_a2x_wrdt_2_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1317) );
  OR2X2 OR2X2_1626 ( .A(u_sdrc_core_u_bs_convert_x2a_wrnext_bF_buf0), .B(\sdr_dq[2] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1318) );
  OR2X2 OR2X2_1627 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n602_bF_buf3), .B(u_sdrc_core_a2x_wrdt_3_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1320) );
  OR2X2 OR2X2_1628 ( .A(u_sdrc_core_u_bs_convert_x2a_wrnext_bF_buf3), .B(\sdr_dq[3] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1321) );
  OR2X2 OR2X2_1629 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n602_bF_buf2), .B(u_sdrc_core_a2x_wrdt_4_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1323) );
  OR2X2 OR2X2_163 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n608), .B(u_sdrc_core_u_bank_ctl__abc_21249_n609), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n610) );
  OR2X2 OR2X2_1630 ( .A(u_sdrc_core_u_bs_convert_x2a_wrnext_bF_buf2), .B(\sdr_dq[4] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1324) );
  OR2X2 OR2X2_1631 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n602_bF_buf1), .B(u_sdrc_core_a2x_wrdt_5_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1326) );
  OR2X2 OR2X2_1632 ( .A(u_sdrc_core_u_bs_convert_x2a_wrnext_bF_buf1), .B(\sdr_dq[5] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1327) );
  OR2X2 OR2X2_1633 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n602_bF_buf0), .B(u_sdrc_core_a2x_wrdt_6_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1329) );
  OR2X2 OR2X2_1634 ( .A(u_sdrc_core_u_bs_convert_x2a_wrnext_bF_buf0), .B(\sdr_dq[6] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1330) );
  OR2X2 OR2X2_1635 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n602_bF_buf3), .B(u_sdrc_core_a2x_wrdt_7_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1332) );
  OR2X2 OR2X2_1636 ( .A(u_sdrc_core_u_bs_convert_x2a_wrnext_bF_buf3), .B(\sdr_dq[7] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1333) );
  OR2X2 OR2X2_1637 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n602_bF_buf2), .B(u_sdrc_core_a2x_wrdt_8_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1335) );
  OR2X2 OR2X2_1638 ( .A(u_sdrc_core_u_bs_convert_x2a_wrnext_bF_buf2), .B(\sdr_dq[8] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1336) );
  OR2X2 OR2X2_1639 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n602_bF_buf1), .B(u_sdrc_core_a2x_wrdt_9_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1338) );
  OR2X2 OR2X2_164 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n611), .B(u_sdrc_core_u_bank_ctl__abc_21249_n612), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n613) );
  OR2X2 OR2X2_1640 ( .A(u_sdrc_core_u_bs_convert_x2a_wrnext_bF_buf1), .B(\sdr_dq[9] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1339) );
  OR2X2 OR2X2_1641 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n602_bF_buf0), .B(u_sdrc_core_a2x_wrdt_10_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1341) );
  OR2X2 OR2X2_1642 ( .A(u_sdrc_core_u_bs_convert_x2a_wrnext_bF_buf0), .B(\sdr_dq[10] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1342) );
  OR2X2 OR2X2_1643 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n602_bF_buf3), .B(u_sdrc_core_a2x_wrdt_11_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1344) );
  OR2X2 OR2X2_1644 ( .A(u_sdrc_core_u_bs_convert_x2a_wrnext_bF_buf3), .B(\sdr_dq[11] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1345) );
  OR2X2 OR2X2_1645 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n602_bF_buf2), .B(u_sdrc_core_a2x_wrdt_12_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1347) );
  OR2X2 OR2X2_1646 ( .A(u_sdrc_core_u_bs_convert_x2a_wrnext_bF_buf2), .B(\sdr_dq[12] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1348) );
  OR2X2 OR2X2_1647 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n602_bF_buf1), .B(u_sdrc_core_a2x_wrdt_13_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1350) );
  OR2X2 OR2X2_1648 ( .A(u_sdrc_core_u_bs_convert_x2a_wrnext_bF_buf1), .B(\sdr_dq[13] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1351) );
  OR2X2 OR2X2_1649 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n602_bF_buf0), .B(u_sdrc_core_a2x_wrdt_14_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1353) );
  OR2X2 OR2X2_165 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n610), .B(u_sdrc_core_u_bank_ctl__abc_21249_n613), .Y(u_sdrc_core_b2x_wrap) );
  OR2X2 OR2X2_1650 ( .A(u_sdrc_core_u_bs_convert_x2a_wrnext_bF_buf0), .B(\sdr_dq[14] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1354) );
  OR2X2 OR2X2_1651 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n602_bF_buf3), .B(u_sdrc_core_a2x_wrdt_15_), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1356) );
  OR2X2 OR2X2_1652 ( .A(u_sdrc_core_u_bs_convert_x2a_wrnext_bF_buf3), .B(\sdr_dq[15] ), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1357) );
  OR2X2 OR2X2_1653 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n589), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n500_1), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1359) );
  OR2X2 OR2X2_1654 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n896), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1359), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1360) );
  OR2X2 OR2X2_1655 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n1364), .B(u_sdrc_core_u_xfr_ctl__abc_23098_n1363), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1365) );
  OR2X2 OR2X2_1656 ( .A(u_sdrc_core_u_xfr_ctl__abc_23098_n872), .B(_auto_iopadmap_cc_313_execute_24701), .Y(u_sdrc_core_u_xfr_ctl__abc_23098_n1370) );
  OR2X2 OR2X2_1657 ( .A(wb_we_i), .B(u_wb2sdrc_rddatafifo_empty), .Y(u_wb2sdrc__abc_24125_n35_1) );
  OR2X2 OR2X2_1658 ( .A(u_wb2sdrc__abc_24125_n34), .B(u_wb2sdrc__abc_24125_n35_1), .Y(u_wb2sdrc__abc_24125_n36_1) );
  OR2X2 OR2X2_1659 ( .A(u_wb2sdrc_rddatafifo_rd), .B(u_wb2sdrc_u_wrdatafifo_wr_en), .Y(_auto_iopadmap_cc_313_execute_24707) );
  OR2X2 OR2X2_166 ( .A(u_sdrc_core_u_bank_ctl_rank_cnt_1_), .B(\cfg_req_depth[1] ), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n617) );
  OR2X2 OR2X2_1660 ( .A(u_wb2sdrc_u_wrdatafifo_wr_en), .B(u_wb2sdrc__abc_24125_n41), .Y(u_wb2sdrc_cmdfifo_wr) );
  OR2X2 OR2X2_1661 ( .A(u_wb2sdrc__abc_24125_n47), .B(u_wb2sdrc__abc_24125_n41), .Y(u_wb2sdrc_pending_read_FF_INPUT) );
  OR2X2 OR2X2_1662 ( .A(u_wb2sdrc_u_cmdfifo_sync_rd_ptr_1_1_), .B(u_wb2sdrc_u_cmdfifo_sync_rd_ptr_2_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n399) );
  OR2X2 OR2X2_1663 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n407_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n409_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n410_1) );
  OR2X2 OR2X2_1664 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n404_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n413_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n414) );
  OR2X2 OR2X2_1665 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n411), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n414), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n415_1) );
  OR2X2 OR2X2_1666 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n419_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n420), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n421_1) );
  OR2X2 OR2X2_1667 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n425_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n423), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n426) );
  OR2X2 OR2X2_1668 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n430_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n429), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n431_1) );
  OR2X2 OR2X2_1669 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n411), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n432), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n433_1) );
  OR2X2 OR2X2_167 ( .A(u_sdrc_core_u_bank_ctl_rank_cnt_0_), .B(\cfg_req_depth[0] ), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n621) );
  OR2X2 OR2X2_1670 ( .A(u_wb2sdrc_u_cmdfifo_sync_wr_ptr_1_1_), .B(u_wb2sdrc_u_cmdfifo_sync_wr_ptr_2_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n437_1) );
  OR2X2 OR2X2_1671 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n445_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n438), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n446_1) );
  OR2X2 OR2X2_1672 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n447), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n449_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n450) );
  OR2X2 OR2X2_1673 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n450), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf7), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n451_1) );
  OR2X2 OR2X2_1674 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n452_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n441), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n453) );
  OR2X2 OR2X2_1675 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n455), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n441), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n456_1) );
  OR2X2 OR2X2_1676 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n444), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_2_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n457_1) );
  OR2X2 OR2X2_1677 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n458_1), .B(u_wb2sdrc_u_cmdfifo_sync_wr_ptr_2_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n459_1) );
  OR2X2 OR2X2_1678 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n440_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n448_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n463_1) );
  OR2X2 OR2X2_1679 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n446_1), .B(u_wb2sdrc_u_cmdfifo_sync_wr_ptr_1_0_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n464_1) );
  OR2X2 OR2X2_168 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n618), .B(u_sdrc_core_u_bank_ctl__abc_21249_n622), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n623) );
  OR2X2 OR2X2_1680 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n466_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n453), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n467_1) );
  OR2X2 OR2X2_1681 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n461_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n470_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n471_1) );
  OR2X2 OR2X2_1682 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n455), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n472_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n473_1) );
  OR2X2 OR2X2_1683 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n466_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n474_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n475_1) );
  OR2X2 OR2X2_1684 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_0__0_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n480_1) );
  OR2X2 OR2X2_1685 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf5), .B(\wb_addr_i[0] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n482_1) );
  OR2X2 OR2X2_1686 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_0__1_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n484_1) );
  OR2X2 OR2X2_1687 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf4), .B(\wb_addr_i[1] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n485_1) );
  OR2X2 OR2X2_1688 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_0__2_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n487_1) );
  OR2X2 OR2X2_1689 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf3), .B(\wb_addr_i[2] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n488_1) );
  OR2X2 OR2X2_169 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n254), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_12_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n255_1) );
  OR2X2 OR2X2_1690 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_0__3_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n490_1) );
  OR2X2 OR2X2_1691 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf2), .B(\wb_addr_i[3] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n491_1) );
  OR2X2 OR2X2_1692 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_0__4_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n493_1) );
  OR2X2 OR2X2_1693 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf1), .B(\wb_addr_i[4] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n494_1) );
  OR2X2 OR2X2_1694 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_0__5_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n496_1) );
  OR2X2 OR2X2_1695 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf0), .B(\wb_addr_i[5] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n497_1) );
  OR2X2 OR2X2_1696 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_0__6_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n499_1) );
  OR2X2 OR2X2_1697 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf5), .B(\wb_addr_i[6] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n500_1) );
  OR2X2 OR2X2_1698 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_0__7_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n502_1) );
  OR2X2 OR2X2_1699 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf4), .B(\wb_addr_i[7] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n503_1) );
  OR2X2 OR2X2_17 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n243), .B(u_sdrc_core_u_bank_ctl__abc_21249_n259_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n260_1) );
  OR2X2 OR2X2_170 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n256_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_11_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n257) );
  OR2X2 OR2X2_1700 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_0__8_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n505_1) );
  OR2X2 OR2X2_1701 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf3), .B(\wb_addr_i[8] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n506_1) );
  OR2X2 OR2X2_1702 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_0__9_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n508_1) );
  OR2X2 OR2X2_1703 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf2), .B(\wb_addr_i[9] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n509_1) );
  OR2X2 OR2X2_1704 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_0__10_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n511_1) );
  OR2X2 OR2X2_1705 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf1), .B(\wb_addr_i[10] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n512_1) );
  OR2X2 OR2X2_1706 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_0__11_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n514_1) );
  OR2X2 OR2X2_1707 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf0), .B(\wb_addr_i[11] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n515_1) );
  OR2X2 OR2X2_1708 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_0__12_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n517_1) );
  OR2X2 OR2X2_1709 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf5), .B(\wb_addr_i[12] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n518_1) );
  OR2X2 OR2X2_171 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n258_1), .B(u_sdrc_core_r2b_raddr_12_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n259_1) );
  OR2X2 OR2X2_1710 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_0__13_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n520_1) );
  OR2X2 OR2X2_1711 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf4), .B(\wb_addr_i[13] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n521_1) );
  OR2X2 OR2X2_1712 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_0__14_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n523_1) );
  OR2X2 OR2X2_1713 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf3), .B(\wb_addr_i[14] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n524_1) );
  OR2X2 OR2X2_1714 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_0__15_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n526_1) );
  OR2X2 OR2X2_1715 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf2), .B(\wb_addr_i[15] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n527_1) );
  OR2X2 OR2X2_1716 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_0__16_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n529) );
  OR2X2 OR2X2_1717 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf1), .B(\wb_addr_i[16] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n530_1) );
  OR2X2 OR2X2_1718 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_0__17_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n532_1) );
  OR2X2 OR2X2_1719 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf0), .B(\wb_addr_i[17] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n533_1) );
  OR2X2 OR2X2_172 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n262_1), .B(u_sdrc_core_r2b_raddr_11_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n263) );
  OR2X2 OR2X2_1720 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_0__18_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n535_1) );
  OR2X2 OR2X2_1721 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf5), .B(\wb_addr_i[18] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n536_1) );
  OR2X2 OR2X2_1722 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_0__19_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n538_1) );
  OR2X2 OR2X2_1723 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf4), .B(\wb_addr_i[19] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n539_1) );
  OR2X2 OR2X2_1724 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_0__20_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n541_1) );
  OR2X2 OR2X2_1725 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf3), .B(\wb_addr_i[20] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n542_1) );
  OR2X2 OR2X2_1726 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_0__21_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n544_1) );
  OR2X2 OR2X2_1727 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf2), .B(\wb_addr_i[21] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n545_1) );
  OR2X2 OR2X2_1728 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_0__22_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n547_1) );
  OR2X2 OR2X2_1729 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf1), .B(\wb_addr_i[22] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n548_1) );
  OR2X2 OR2X2_173 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n264_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_9_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n265_1) );
  OR2X2 OR2X2_1730 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_0__23_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n550_1) );
  OR2X2 OR2X2_1731 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf0), .B(\wb_addr_i[23] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n551_1) );
  OR2X2 OR2X2_1732 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_0__24_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n553_1) );
  OR2X2 OR2X2_1733 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf5), .B(\wb_addr_i[24] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n554_1) );
  OR2X2 OR2X2_1734 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_0__25_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n556_1) );
  OR2X2 OR2X2_1735 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf4), .B(\wb_addr_i[25] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n557_1) );
  OR2X2 OR2X2_1736 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_0__26_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n559_1) );
  OR2X2 OR2X2_1737 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_wr_data_26_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n560_1) );
  OR2X2 OR2X2_1738 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_0__27_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n562_1) );
  OR2X2 OR2X2_1739 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf2), .B(1'b1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n563_1) );
  OR2X2 OR2X2_174 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n267_1), .B(u_sdrc_core_r2b_raddr_9_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n268_1) );
  OR2X2 OR2X2_1740 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_0__28_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n565_1) );
  OR2X2 OR2X2_1741 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf1), .B(1'b0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n566) );
  OR2X2 OR2X2_1742 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_0__29_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n568) );
  OR2X2 OR2X2_1743 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf0), .B(1'b0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n569) );
  OR2X2 OR2X2_1744 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_0__30_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n571) );
  OR2X2 OR2X2_1745 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf5), .B(1'b0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n572) );
  OR2X2 OR2X2_1746 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_0__31_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n574) );
  OR2X2 OR2X2_1747 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf4), .B(1'b0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n575) );
  OR2X2 OR2X2_1748 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_0__32_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n577) );
  OR2X2 OR2X2_1749 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf3), .B(1'b0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n578) );
  OR2X2 OR2X2_175 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n269), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_7_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n270_1) );
  OR2X2 OR2X2_1750 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_0__33_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n580) );
  OR2X2 OR2X2_1751 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf2), .B(1'b0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n581) );
  OR2X2 OR2X2_1752 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_0__34_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n583) );
  OR2X2 OR2X2_1753 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf1), .B(1'b0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n584) );
  OR2X2 OR2X2_1754 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n479_1_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_0__35_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n586) );
  OR2X2 OR2X2_1755 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n481_1_bF_buf0), .B(1'b0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n587) );
  OR2X2 OR2X2_1756 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n589), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n591), .Y(u_wb2sdrc_u_cmdfifo_grey_rd_ptr_0__FF_INPUT) );
  OR2X2 OR2X2_1757 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n594), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n593), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n595) );
  OR2X2 OR2X2_1758 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n593), .B(u_wb2sdrc_u_cmdfifo_rd_ptr_2_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n598) );
  OR2X2 OR2X2_1759 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n605), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n602), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n606) );
  OR2X2 OR2X2_176 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n274_1), .B(u_sdrc_core_r2b_raddr_7_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n275) );
  OR2X2 OR2X2_1760 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n606), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n601), .Y(u_wb2sdrc_u_cmdfifo_grey_rd_ptr_1__FF_INPUT) );
  OR2X2 OR2X2_1761 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n600), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n608), .Y(u_wb2sdrc_u_cmdfifo_grey_rd_ptr_2__FF_INPUT) );
  OR2X2 OR2X2_1762 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n610), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n611), .Y(u_wb2sdrc_u_cmdfifo_rd_ptr_0__FF_INPUT) );
  OR2X2 OR2X2_1763 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n604), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n613), .Y(u_wb2sdrc_u_cmdfifo_rd_ptr_1__FF_INPUT) );
  OR2X2 OR2X2_1764 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n600), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n615), .Y(u_wb2sdrc_u_cmdfifo_rd_ptr_2__FF_INPUT) );
  OR2X2 OR2X2_1765 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n617), .B(u_wb2sdrc_cmdfifo_empty), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n618) );
  OR2X2 OR2X2_1766 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n621), .B(app_req_ack_bF_buf1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n622) );
  OR2X2 OR2X2_1767 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n478_1), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n625), .Y(u_wb2sdrc_u_cmdfifo_wr_ptr_0__FF_INPUT) );
  OR2X2 OR2X2_1768 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf5), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n628), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n631) );
  OR2X2 OR2X2_1769 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n631), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf5), .Y(u_wb2sdrc_u_cmdfifo_wr_ptr_1__FF_INPUT) );
  OR2X2 OR2X2_177 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n276_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_3_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n277_1) );
  OR2X2 OR2X2_1770 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n634), .B(u_wb2sdrc_u_cmdfifo_wr_ptr_2_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n637) );
  OR2X2 OR2X2_1771 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n639), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n633), .Y(u_wb2sdrc_u_cmdfifo_wr_ptr_2__FF_INPUT) );
  OR2X2 OR2X2_1772 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n629), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n641), .Y(u_wb2sdrc_u_cmdfifo_grey_wr_ptr_0__FF_INPUT) );
  OR2X2 OR2X2_1773 ( .A(u_wb2sdrc_cmdfifo_wr), .B(u_wb2sdrc_u_cmdfifo_grey_wr_ptr_1_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n643) );
  OR2X2 OR2X2_1774 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n645), .B(u_wb2sdrc_u_cmdfifo_wr_ptr_2_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n646) );
  OR2X2 OR2X2_1775 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n644), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n418_1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n647) );
  OR2X2 OR2X2_1776 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n648), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n624), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n649) );
  OR2X2 OR2X2_1777 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n639), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n651), .Y(u_wb2sdrc_u_cmdfifo_grey_wr_ptr_2__FF_INPUT) );
  OR2X2 OR2X2_1778 ( .A(u_wb2sdrc_u_cmdfifo_afull), .B(u_wb2sdrc_cmdfifo_full), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n653) );
  OR2X2 OR2X2_1779 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n654), .B(u_wb2sdrc_cmdfifo_wr), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n655) );
  OR2X2 OR2X2_178 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n279_1), .B(u_sdrc_core_r2b_raddr_6_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n280_1) );
  OR2X2 OR2X2_1780 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_0__0_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n657) );
  OR2X2 OR2X2_1781 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_1__0_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n658) );
  OR2X2 OR2X2_1782 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_3__0_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n661) );
  OR2X2 OR2X2_1783 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_2__0_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n662) );
  OR2X2 OR2X2_1784 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n660), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n664), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n349) );
  OR2X2 OR2X2_1785 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_0__1_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n666) );
  OR2X2 OR2X2_1786 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_1__1_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n667) );
  OR2X2 OR2X2_1787 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_3__1_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n670) );
  OR2X2 OR2X2_1788 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_2__1_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n671) );
  OR2X2 OR2X2_1789 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n669), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n673), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n351) );
  OR2X2 OR2X2_179 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n281), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_6_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n282_1) );
  OR2X2 OR2X2_1790 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf7), .B(u_wb2sdrc_u_cmdfifo_mem_0__2_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n675) );
  OR2X2 OR2X2_1791 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf7), .B(u_wb2sdrc_u_cmdfifo_mem_1__2_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n676) );
  OR2X2 OR2X2_1792 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf6), .B(u_wb2sdrc_u_cmdfifo_mem_3__2_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n679) );
  OR2X2 OR2X2_1793 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf6), .B(u_wb2sdrc_u_cmdfifo_mem_2__2_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n680) );
  OR2X2 OR2X2_1794 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n678), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n682), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n353) );
  OR2X2 OR2X2_1795 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_0__3_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n684) );
  OR2X2 OR2X2_1796 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_1__3_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n685) );
  OR2X2 OR2X2_1797 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_3__3_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n688) );
  OR2X2 OR2X2_1798 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_2__3_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n689) );
  OR2X2 OR2X2_1799 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n687), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n691), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n355) );
  OR2X2 OR2X2_18 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n261_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n251_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n262) );
  OR2X2 OR2X2_180 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n285), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_5_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n286_1) );
  OR2X2 OR2X2_1800 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_0__4_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n693) );
  OR2X2 OR2X2_1801 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_1__4_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n694) );
  OR2X2 OR2X2_1802 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_3__4_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n697) );
  OR2X2 OR2X2_1803 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_2__4_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n698) );
  OR2X2 OR2X2_1804 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n696), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n700), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n357) );
  OR2X2 OR2X2_1805 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_0__5_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n702) );
  OR2X2 OR2X2_1806 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_1__5_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n703) );
  OR2X2 OR2X2_1807 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_3__5_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n706) );
  OR2X2 OR2X2_1808 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_2__5_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n707) );
  OR2X2 OR2X2_1809 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n705), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n709), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n359) );
  OR2X2 OR2X2_181 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n287_1), .B(u_sdrc_core_r2b_raddr_1_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n288_1) );
  OR2X2 OR2X2_1810 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf7), .B(u_wb2sdrc_u_cmdfifo_mem_0__6_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n711) );
  OR2X2 OR2X2_1811 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf7), .B(u_wb2sdrc_u_cmdfifo_mem_1__6_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n712) );
  OR2X2 OR2X2_1812 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf6), .B(u_wb2sdrc_u_cmdfifo_mem_3__6_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n715) );
  OR2X2 OR2X2_1813 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf6), .B(u_wb2sdrc_u_cmdfifo_mem_2__6_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n716) );
  OR2X2 OR2X2_1814 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n714), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n718), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n361) );
  OR2X2 OR2X2_1815 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_0__7_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n720) );
  OR2X2 OR2X2_1816 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_1__7_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n721) );
  OR2X2 OR2X2_1817 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_3__7_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n724) );
  OR2X2 OR2X2_1818 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_2__7_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n725) );
  OR2X2 OR2X2_1819 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n723), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n727), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n363) );
  OR2X2 OR2X2_182 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n290_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_0_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n291_1) );
  OR2X2 OR2X2_1820 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_0__8_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n729) );
  OR2X2 OR2X2_1821 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_1__8_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n730) );
  OR2X2 OR2X2_1822 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_3__8_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n733) );
  OR2X2 OR2X2_1823 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_2__8_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n734) );
  OR2X2 OR2X2_1824 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n732), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n736), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n365) );
  OR2X2 OR2X2_1825 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_0__9_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n738) );
  OR2X2 OR2X2_1826 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_1__9_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n739) );
  OR2X2 OR2X2_1827 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_3__9_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n742) );
  OR2X2 OR2X2_1828 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_2__9_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n743) );
  OR2X2 OR2X2_1829 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n741), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n745), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n367) );
  OR2X2 OR2X2_183 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n292_1), .B(u_sdrc_core_r2b_raddr_0_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n293) );
  OR2X2 OR2X2_1830 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf7), .B(u_wb2sdrc_u_cmdfifo_mem_0__10_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n747) );
  OR2X2 OR2X2_1831 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf7), .B(u_wb2sdrc_u_cmdfifo_mem_1__10_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n748) );
  OR2X2 OR2X2_1832 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf6), .B(u_wb2sdrc_u_cmdfifo_mem_3__10_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n751) );
  OR2X2 OR2X2_1833 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf6), .B(u_wb2sdrc_u_cmdfifo_mem_2__10_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n752) );
  OR2X2 OR2X2_1834 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n750), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n754), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n369) );
  OR2X2 OR2X2_1835 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_0__11_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n756) );
  OR2X2 OR2X2_1836 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_1__11_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n757) );
  OR2X2 OR2X2_1837 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_3__11_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n760) );
  OR2X2 OR2X2_1838 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_2__11_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n761) );
  OR2X2 OR2X2_1839 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n759), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n763), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n371) );
  OR2X2 OR2X2_184 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n301), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n298_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n302_1) );
  OR2X2 OR2X2_1840 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_0__12_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n765) );
  OR2X2 OR2X2_1841 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_1__12_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n766) );
  OR2X2 OR2X2_1842 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_3__12_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n769) );
  OR2X2 OR2X2_1843 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_2__12_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n770) );
  OR2X2 OR2X2_1844 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n768), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n772), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n373) );
  OR2X2 OR2X2_1845 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_0__13_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n774) );
  OR2X2 OR2X2_1846 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_1__13_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n775) );
  OR2X2 OR2X2_1847 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_3__13_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n778) );
  OR2X2 OR2X2_1848 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_2__13_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n779) );
  OR2X2 OR2X2_1849 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n777), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n781), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n375) );
  OR2X2 OR2X2_185 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n306_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n303_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n307_1) );
  OR2X2 OR2X2_1850 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf7), .B(u_wb2sdrc_u_cmdfifo_mem_0__14_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n783) );
  OR2X2 OR2X2_1851 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf7), .B(u_wb2sdrc_u_cmdfifo_mem_1__14_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n784) );
  OR2X2 OR2X2_1852 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf6), .B(u_wb2sdrc_u_cmdfifo_mem_3__14_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n787) );
  OR2X2 OR2X2_1853 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf6), .B(u_wb2sdrc_u_cmdfifo_mem_2__14_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n788) );
  OR2X2 OR2X2_1854 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n786), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n790), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n377) );
  OR2X2 OR2X2_1855 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_0__15_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n792) );
  OR2X2 OR2X2_1856 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_1__15_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n793) );
  OR2X2 OR2X2_1857 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_3__15_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n796) );
  OR2X2 OR2X2_1858 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_2__15_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n797) );
  OR2X2 OR2X2_1859 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n795), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n799), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n379) );
  OR2X2 OR2X2_186 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n309), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_2_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n310_1) );
  OR2X2 OR2X2_1860 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_0__16_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n801) );
  OR2X2 OR2X2_1861 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_1__16_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n802) );
  OR2X2 OR2X2_1862 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_3__16_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n805) );
  OR2X2 OR2X2_1863 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_2__16_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n806) );
  OR2X2 OR2X2_1864 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n804), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n808), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n381) );
  OR2X2 OR2X2_1865 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_0__17_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n810) );
  OR2X2 OR2X2_1866 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_1__17_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n811) );
  OR2X2 OR2X2_1867 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_3__17_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n814) );
  OR2X2 OR2X2_1868 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_2__17_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n815) );
  OR2X2 OR2X2_1869 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n813), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n817), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n383) );
  OR2X2 OR2X2_187 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n311_1), .B(u_sdrc_core_r2b_raddr_3_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n312_1) );
  OR2X2 OR2X2_1870 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf7), .B(u_wb2sdrc_u_cmdfifo_mem_0__18_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n819) );
  OR2X2 OR2X2_1871 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf7), .B(u_wb2sdrc_u_cmdfifo_mem_1__18_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n820) );
  OR2X2 OR2X2_1872 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf6), .B(u_wb2sdrc_u_cmdfifo_mem_3__18_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n823) );
  OR2X2 OR2X2_1873 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf6), .B(u_wb2sdrc_u_cmdfifo_mem_2__18_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n824) );
  OR2X2 OR2X2_1874 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n822), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n826), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n385) );
  OR2X2 OR2X2_1875 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_0__19_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n828) );
  OR2X2 OR2X2_1876 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_1__19_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n829) );
  OR2X2 OR2X2_1877 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_3__19_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n832) );
  OR2X2 OR2X2_1878 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_2__19_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n833) );
  OR2X2 OR2X2_1879 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n831), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n835), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n387) );
  OR2X2 OR2X2_188 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n314_1), .B(u_sdrc_core_r2b_raddr_2_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n315_1) );
  OR2X2 OR2X2_1880 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_0__20_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n837) );
  OR2X2 OR2X2_1881 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_1__20_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n838) );
  OR2X2 OR2X2_1882 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_3__20_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n841) );
  OR2X2 OR2X2_1883 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_2__20_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n842) );
  OR2X2 OR2X2_1884 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n840), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n844), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n389) );
  OR2X2 OR2X2_1885 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_0__21_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n846) );
  OR2X2 OR2X2_1886 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_1__21_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n847) );
  OR2X2 OR2X2_1887 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_3__21_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n850) );
  OR2X2 OR2X2_1888 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_2__21_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n851) );
  OR2X2 OR2X2_1889 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n849), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n853), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n391) );
  OR2X2 OR2X2_189 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n316_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_1_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n317) );
  OR2X2 OR2X2_1890 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf7), .B(u_wb2sdrc_u_cmdfifo_mem_0__22_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n855) );
  OR2X2 OR2X2_1891 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf7), .B(u_wb2sdrc_u_cmdfifo_mem_1__22_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n856) );
  OR2X2 OR2X2_1892 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf6), .B(u_wb2sdrc_u_cmdfifo_mem_3__22_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n859) );
  OR2X2 OR2X2_1893 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf6), .B(u_wb2sdrc_u_cmdfifo_mem_2__22_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n860) );
  OR2X2 OR2X2_1894 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n858), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n862), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n393) );
  OR2X2 OR2X2_1895 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_0__23_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n864) );
  OR2X2 OR2X2_1896 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_1__23_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n865) );
  OR2X2 OR2X2_1897 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_3__23_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n868) );
  OR2X2 OR2X2_1898 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_2__23_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n869) );
  OR2X2 OR2X2_1899 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n867), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n871), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n395) );
  OR2X2 OR2X2_19 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n244_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n264), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n265_1) );
  OR2X2 OR2X2_190 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n320_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_4_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n321) );
  OR2X2 OR2X2_1900 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_0__24_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n873) );
  OR2X2 OR2X2_1901 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_1__24_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n874) );
  OR2X2 OR2X2_1902 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_3__24_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n877) );
  OR2X2 OR2X2_1903 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_2__24_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n878) );
  OR2X2 OR2X2_1904 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n876), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n880), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n397) );
  OR2X2 OR2X2_1905 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_0__25_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n882) );
  OR2X2 OR2X2_1906 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_1__25_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n883) );
  OR2X2 OR2X2_1907 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_3__25_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n886) );
  OR2X2 OR2X2_1908 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_2__25_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n887) );
  OR2X2 OR2X2_1909 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n885), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n889), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n399) );
  OR2X2 OR2X2_191 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n322_1), .B(u_sdrc_core_r2b_raddr_4_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n323_1) );
  OR2X2 OR2X2_1910 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf7), .B(u_wb2sdrc_u_cmdfifo_mem_0__26_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n891) );
  OR2X2 OR2X2_1911 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf7), .B(u_wb2sdrc_u_cmdfifo_mem_1__26_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n892) );
  OR2X2 OR2X2_1912 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf6), .B(u_wb2sdrc_u_cmdfifo_mem_3__26_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n895) );
  OR2X2 OR2X2_1913 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf6), .B(u_wb2sdrc_u_cmdfifo_mem_2__26_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n896) );
  OR2X2 OR2X2_1914 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n894), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n898), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n401) );
  OR2X2 OR2X2_1915 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_0__27_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n900) );
  OR2X2 OR2X2_1916 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_1__27_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n901) );
  OR2X2 OR2X2_1917 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_3__27_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n904) );
  OR2X2 OR2X2_1918 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_2__27_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n905) );
  OR2X2 OR2X2_1919 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n903), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n907), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n403) );
  OR2X2 OR2X2_192 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n325), .B(u_sdrc_core_r2b_raddr_5_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n326_1) );
  OR2X2 OR2X2_1920 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_0__28_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n909) );
  OR2X2 OR2X2_1921 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_1__28_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n910) );
  OR2X2 OR2X2_1922 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_3__28_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n913) );
  OR2X2 OR2X2_1923 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_2__28_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n914) );
  OR2X2 OR2X2_1924 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n912), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n916), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n405) );
  OR2X2 OR2X2_1925 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_0__29_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n918) );
  OR2X2 OR2X2_1926 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_1__29_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n919) );
  OR2X2 OR2X2_1927 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_3__29_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n922) );
  OR2X2 OR2X2_1928 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_2__29_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n923) );
  OR2X2 OR2X2_1929 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n921), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n925), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n407) );
  OR2X2 OR2X2_193 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n333), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n251), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_17422_n55) );
  OR2X2 OR2X2_1930 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf7), .B(u_wb2sdrc_u_cmdfifo_mem_0__30_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n927) );
  OR2X2 OR2X2_1931 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf7), .B(u_wb2sdrc_u_cmdfifo_mem_1__30_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n928) );
  OR2X2 OR2X2_1932 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf6), .B(u_wb2sdrc_u_cmdfifo_mem_3__30_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n931) );
  OR2X2 OR2X2_1933 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf6), .B(u_wb2sdrc_u_cmdfifo_mem_2__30_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n932) );
  OR2X2 OR2X2_1934 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n930), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n934), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n409) );
  OR2X2 OR2X2_1935 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_0__31_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n936) );
  OR2X2 OR2X2_1936 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_1__31_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n937) );
  OR2X2 OR2X2_1937 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_3__31_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n940) );
  OR2X2 OR2X2_1938 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_2__31_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n941) );
  OR2X2 OR2X2_1939 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n939), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n943), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n411) );
  OR2X2 OR2X2_194 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n340), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n335), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_17422_n61) );
  OR2X2 OR2X2_1940 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_0__32_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n945) );
  OR2X2 OR2X2_1941 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_1__32_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n946) );
  OR2X2 OR2X2_1942 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_3__32_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n949) );
  OR2X2 OR2X2_1943 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_2__32_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n950) );
  OR2X2 OR2X2_1944 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n948), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n952), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n413) );
  OR2X2 OR2X2_1945 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_0__33_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n954) );
  OR2X2 OR2X2_1946 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_1__33_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n955) );
  OR2X2 OR2X2_1947 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_3__33_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n958) );
  OR2X2 OR2X2_1948 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_2__33_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n959) );
  OR2X2 OR2X2_1949 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n957), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n961), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n415) );
  OR2X2 OR2X2_195 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n344_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n345), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n346) );
  OR2X2 OR2X2_1950 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf7), .B(u_wb2sdrc_u_cmdfifo_mem_0__34_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n963) );
  OR2X2 OR2X2_1951 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf7), .B(u_wb2sdrc_u_cmdfifo_mem_1__34_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n964) );
  OR2X2 OR2X2_1952 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf6), .B(u_wb2sdrc_u_cmdfifo_mem_3__34_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n967) );
  OR2X2 OR2X2_1953 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf6), .B(u_wb2sdrc_u_cmdfifo_mem_2__34_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n968) );
  OR2X2 OR2X2_1954 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n966), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n970), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n417) );
  OR2X2 OR2X2_1955 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_0__35_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n972) );
  OR2X2 OR2X2_1956 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_1__35_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n973) );
  OR2X2 OR2X2_1957 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n442_1_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_3__35_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n976) );
  OR2X2 OR2X2_1958 ( .A(u_wb2sdrc_u_cmdfifo_rd_ptr_0_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_2__35_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n977) );
  OR2X2 OR2X2_1959 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n975), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n979), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n419) );
  OR2X2 OR2X2_196 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n346), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n342), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_17422_n66) );
  OR2X2 OR2X2_1960 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n983), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n984), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n422) );
  OR2X2 OR2X2_1961 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n986), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n987), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n424) );
  OR2X2 OR2X2_1962 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n989), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n990), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n426) );
  OR2X2 OR2X2_1963 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n992), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n993), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n428) );
  OR2X2 OR2X2_1964 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n995), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n996), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n430) );
  OR2X2 OR2X2_1965 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n998), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n999), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n432) );
  OR2X2 OR2X2_1966 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1001), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1002), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n434) );
  OR2X2 OR2X2_1967 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1004), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1005), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n436) );
  OR2X2 OR2X2_1968 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1007), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1008), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n438) );
  OR2X2 OR2X2_1969 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1010), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1011), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n440) );
  OR2X2 OR2X2_197 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n349_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n348_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n350) );
  OR2X2 OR2X2_1970 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1013), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1014), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n442) );
  OR2X2 OR2X2_1971 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1016), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1017), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n444) );
  OR2X2 OR2X2_1972 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1019), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1020), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n446) );
  OR2X2 OR2X2_1973 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1022), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1023), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n448) );
  OR2X2 OR2X2_1974 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1025), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1026), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n450) );
  OR2X2 OR2X2_1975 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1028), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1029), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n452) );
  OR2X2 OR2X2_1976 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1031), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1032), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n454) );
  OR2X2 OR2X2_1977 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1034), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1035), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n456) );
  OR2X2 OR2X2_1978 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1037), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1038), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n458) );
  OR2X2 OR2X2_1979 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1040), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1041), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n460) );
  OR2X2 OR2X2_198 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n351), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n350), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_17422_n82) );
  OR2X2 OR2X2_1980 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1043), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1044), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n462) );
  OR2X2 OR2X2_1981 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1046), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1047), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n464) );
  OR2X2 OR2X2_1982 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1049), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1050), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n466) );
  OR2X2 OR2X2_1983 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1052), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1053), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n468) );
  OR2X2 OR2X2_1984 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1055), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1056), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n470) );
  OR2X2 OR2X2_1985 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1058), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1059), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n472) );
  OR2X2 OR2X2_1986 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1061), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1062), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n474) );
  OR2X2 OR2X2_1987 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1064), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1065), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n476) );
  OR2X2 OR2X2_1988 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1067), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1068), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n478) );
  OR2X2 OR2X2_1989 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1070), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1071), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n480) );
  OR2X2 OR2X2_199 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n359_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n361), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n362) );
  OR2X2 OR2X2_1990 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1073), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1074), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n482) );
  OR2X2 OR2X2_1991 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1076), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1077), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n484) );
  OR2X2 OR2X2_1992 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1079), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1080), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n486) );
  OR2X2 OR2X2_1993 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1082), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1083), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n488) );
  OR2X2 OR2X2_1994 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1085), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1086), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n490) );
  OR2X2 OR2X2_1995 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1088), .B(u_wb2sdrc_u_cmdfifo__abc_18561_n1089), .Y(u_wb2sdrc_u_cmdfifo__abc_14585_n492) );
  OR2X2 OR2X2_1996 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_1__0_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1091) );
  OR2X2 OR2X2_1997 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf5), .B(\wb_addr_i[0] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1093) );
  OR2X2 OR2X2_1998 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_1__1_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1095) );
  OR2X2 OR2X2_1999 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf4), .B(\wb_addr_i[1] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1096) );
  OR2X2 OR2X2_2 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2r_ack_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_b2r_ack_bF_buf4), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n208) );
  OR2X2 OR2X2_20 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n271), .B(u_sdrc_core_u_bank_ctl__abc_21249_n269), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n272_1) );
  OR2X2 OR2X2_200 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n362), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n354_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_17422_n90) );
  OR2X2 OR2X2_2000 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_1__2_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1098) );
  OR2X2 OR2X2_2001 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf3), .B(\wb_addr_i[2] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1099) );
  OR2X2 OR2X2_2002 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_1__3_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1101) );
  OR2X2 OR2X2_2003 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf2), .B(\wb_addr_i[3] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1102) );
  OR2X2 OR2X2_2004 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_1__4_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1104) );
  OR2X2 OR2X2_2005 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf1), .B(\wb_addr_i[4] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1105) );
  OR2X2 OR2X2_2006 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_1__5_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1107) );
  OR2X2 OR2X2_2007 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf0), .B(\wb_addr_i[5] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1108) );
  OR2X2 OR2X2_2008 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_1__6_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1110) );
  OR2X2 OR2X2_2009 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf5), .B(\wb_addr_i[6] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1111) );
  OR2X2 OR2X2_201 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n364_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_2_bF_buf1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n365) );
  OR2X2 OR2X2_2010 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_1__7_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1113) );
  OR2X2 OR2X2_2011 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf4), .B(\wb_addr_i[7] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1114) );
  OR2X2 OR2X2_2012 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_1__8_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1116) );
  OR2X2 OR2X2_2013 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf3), .B(\wb_addr_i[8] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1117) );
  OR2X2 OR2X2_2014 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_1__9_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1119) );
  OR2X2 OR2X2_2015 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf2), .B(\wb_addr_i[9] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1120) );
  OR2X2 OR2X2_2016 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_1__10_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1122) );
  OR2X2 OR2X2_2017 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf1), .B(\wb_addr_i[10] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1123) );
  OR2X2 OR2X2_2018 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_1__11_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1125) );
  OR2X2 OR2X2_2019 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf0), .B(\wb_addr_i[11] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1126) );
  OR2X2 OR2X2_202 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_3_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_prech_page_closed), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n368_1) );
  OR2X2 OR2X2_2020 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_1__12_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1128) );
  OR2X2 OR2X2_2021 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf5), .B(\wb_addr_i[12] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1129) );
  OR2X2 OR2X2_2022 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_1__13_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1131) );
  OR2X2 OR2X2_2023 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf4), .B(\wb_addr_i[13] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1132) );
  OR2X2 OR2X2_2024 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_1__14_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1134) );
  OR2X2 OR2X2_2025 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf3), .B(\wb_addr_i[14] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1135) );
  OR2X2 OR2X2_2026 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_1__15_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1137) );
  OR2X2 OR2X2_2027 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf2), .B(\wb_addr_i[15] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1138) );
  OR2X2 OR2X2_2028 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_1__16_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1140) );
  OR2X2 OR2X2_2029 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf1), .B(\wb_addr_i[16] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1141) );
  OR2X2 OR2X2_203 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n373_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n365), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n374_1) );
  OR2X2 OR2X2_2030 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_1__17_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1143) );
  OR2X2 OR2X2_2031 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf0), .B(\wb_addr_i[17] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1144) );
  OR2X2 OR2X2_2032 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_1__18_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1146) );
  OR2X2 OR2X2_2033 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf5), .B(\wb_addr_i[18] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1147) );
  OR2X2 OR2X2_2034 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_1__19_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1149) );
  OR2X2 OR2X2_2035 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf4), .B(\wb_addr_i[19] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1150) );
  OR2X2 OR2X2_2036 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_1__20_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1152) );
  OR2X2 OR2X2_2037 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf3), .B(\wb_addr_i[20] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1153) );
  OR2X2 OR2X2_2038 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_1__21_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1155) );
  OR2X2 OR2X2_2039 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf2), .B(\wb_addr_i[21] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1156) );
  OR2X2 OR2X2_204 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n377), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n337), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_cmd_r_1__FF_INPUT) );
  OR2X2 OR2X2_2040 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_1__22_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1158) );
  OR2X2 OR2X2_2041 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf1), .B(\wb_addr_i[22] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1159) );
  OR2X2 OR2X2_2042 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_1__23_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1161) );
  OR2X2 OR2X2_2043 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf0), .B(\wb_addr_i[23] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1162) );
  OR2X2 OR2X2_2044 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_1__24_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1164) );
  OR2X2 OR2X2_2045 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf5), .B(\wb_addr_i[24] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1165) );
  OR2X2 OR2X2_2046 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_1__25_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1167) );
  OR2X2 OR2X2_2047 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf4), .B(\wb_addr_i[25] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1168) );
  OR2X2 OR2X2_2048 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_1__26_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1170) );
  OR2X2 OR2X2_2049 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_wr_data_26_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1171) );
  OR2X2 OR2X2_205 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n249_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_cmd_1_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n380) );
  OR2X2 OR2X2_2050 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_1__27_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1173) );
  OR2X2 OR2X2_2051 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf2), .B(1'b1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1174) );
  OR2X2 OR2X2_2052 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_1__28_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1176) );
  OR2X2 OR2X2_2053 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf1), .B(1'b0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1177) );
  OR2X2 OR2X2_2054 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_1__29_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1179) );
  OR2X2 OR2X2_2055 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf0), .B(1'b0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1180) );
  OR2X2 OR2X2_2056 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_1__30_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1182) );
  OR2X2 OR2X2_2057 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf5), .B(1'b0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1183) );
  OR2X2 OR2X2_2058 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_1__31_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1185) );
  OR2X2 OR2X2_2059 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf4), .B(1'b0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1186) );
  OR2X2 OR2X2_206 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_tras_cntr_0_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_tras_cntr_1_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n384_1) );
  OR2X2 OR2X2_2060 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_1__32_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1188) );
  OR2X2 OR2X2_2061 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf3), .B(1'b0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1189) );
  OR2X2 OR2X2_2062 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_1__33_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1191) );
  OR2X2 OR2X2_2063 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf2), .B(1'b0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1192) );
  OR2X2 OR2X2_2064 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_1__34_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1194) );
  OR2X2 OR2X2_2065 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf1), .B(1'b0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1195) );
  OR2X2 OR2X2_2066 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n630_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_1__35_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1197) );
  OR2X2 OR2X2_2067 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1092_bF_buf0), .B(1'b0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1198) );
  OR2X2 OR2X2_2068 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_2__0_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1200) );
  OR2X2 OR2X2_2069 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf5), .B(\wb_addr_i[0] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1202) );
  OR2X2 OR2X2_207 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n384_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_tras_cntr_2_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n385) );
  OR2X2 OR2X2_2070 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_2__1_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1204) );
  OR2X2 OR2X2_2071 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf4), .B(\wb_addr_i[1] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1205) );
  OR2X2 OR2X2_2072 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_2__2_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1207) );
  OR2X2 OR2X2_2073 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf3), .B(\wb_addr_i[2] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1208) );
  OR2X2 OR2X2_2074 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_2__3_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1210) );
  OR2X2 OR2X2_2075 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf2), .B(\wb_addr_i[3] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1211) );
  OR2X2 OR2X2_2076 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_2__4_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1213) );
  OR2X2 OR2X2_2077 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf1), .B(\wb_addr_i[4] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1214) );
  OR2X2 OR2X2_2078 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_2__5_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1216) );
  OR2X2 OR2X2_2079 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf0), .B(\wb_addr_i[5] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1217) );
  OR2X2 OR2X2_208 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n385), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_tras_cntr_3_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n386_1) );
  OR2X2 OR2X2_2080 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_2__6_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1219) );
  OR2X2 OR2X2_2081 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf5), .B(\wb_addr_i[6] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1220) );
  OR2X2 OR2X2_2082 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_2__7_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1222) );
  OR2X2 OR2X2_2083 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf4), .B(\wb_addr_i[7] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1223) );
  OR2X2 OR2X2_2084 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_2__8_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1225) );
  OR2X2 OR2X2_2085 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf3), .B(\wb_addr_i[8] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1226) );
  OR2X2 OR2X2_2086 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_2__9_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1228) );
  OR2X2 OR2X2_2087 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf2), .B(\wb_addr_i[9] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1229) );
  OR2X2 OR2X2_2088 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_2__10_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1231) );
  OR2X2 OR2X2_2089 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf1), .B(\wb_addr_i[10] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1232) );
  OR2X2 OR2X2_209 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n388), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n389), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n390) );
  OR2X2 OR2X2_2090 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_2__11_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1234) );
  OR2X2 OR2X2_2091 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf0), .B(\wb_addr_i[11] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1235) );
  OR2X2 OR2X2_2092 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_2__12_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1237) );
  OR2X2 OR2X2_2093 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf5), .B(\wb_addr_i[12] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1238) );
  OR2X2 OR2X2_2094 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_2__13_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1240) );
  OR2X2 OR2X2_2095 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf4), .B(\wb_addr_i[13] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1241) );
  OR2X2 OR2X2_2096 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_2__14_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1243) );
  OR2X2 OR2X2_2097 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf3), .B(\wb_addr_i[14] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1244) );
  OR2X2 OR2X2_2098 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_2__15_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1246) );
  OR2X2 OR2X2_2099 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf2), .B(\wb_addr_i[15] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1247) );
  OR2X2 OR2X2_21 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n273_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n274_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n275_1) );
  OR2X2 OR2X2_210 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n393), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n394_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n395_1) );
  OR2X2 OR2X2_2100 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_2__16_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1249) );
  OR2X2 OR2X2_2101 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf1), .B(\wb_addr_i[16] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1250) );
  OR2X2 OR2X2_2102 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_2__17_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1252) );
  OR2X2 OR2X2_2103 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf0), .B(\wb_addr_i[17] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1253) );
  OR2X2 OR2X2_2104 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_2__18_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1255) );
  OR2X2 OR2X2_2105 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf5), .B(\wb_addr_i[18] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1256) );
  OR2X2 OR2X2_2106 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_2__19_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1258) );
  OR2X2 OR2X2_2107 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf4), .B(\wb_addr_i[19] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1259) );
  OR2X2 OR2X2_2108 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_2__20_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1261) );
  OR2X2 OR2X2_2109 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf3), .B(\wb_addr_i[20] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1262) );
  OR2X2 OR2X2_211 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n396_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n392_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n397_1) );
  OR2X2 OR2X2_2110 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_2__21_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1264) );
  OR2X2 OR2X2_2111 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf2), .B(\wb_addr_i[21] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1265) );
  OR2X2 OR2X2_2112 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_2__22_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1267) );
  OR2X2 OR2X2_2113 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf1), .B(\wb_addr_i[22] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1268) );
  OR2X2 OR2X2_2114 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_2__23_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1270) );
  OR2X2 OR2X2_2115 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf0), .B(\wb_addr_i[23] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1271) );
  OR2X2 OR2X2_2116 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_2__24_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1273) );
  OR2X2 OR2X2_2117 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf5), .B(\wb_addr_i[24] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1274) );
  OR2X2 OR2X2_2118 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_2__25_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1276) );
  OR2X2 OR2X2_2119 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf4), .B(\wb_addr_i[25] ), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1277) );
  OR2X2 OR2X2_212 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n400_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n401_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n402_1) );
  OR2X2 OR2X2_2120 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_2__26_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1279) );
  OR2X2 OR2X2_2121 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_wr_data_26_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1280) );
  OR2X2 OR2X2_2122 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_2__27_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1282) );
  OR2X2 OR2X2_2123 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf2), .B(1'b1), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1283) );
  OR2X2 OR2X2_2124 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_2__28_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1285) );
  OR2X2 OR2X2_2125 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf1), .B(1'b0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1286) );
  OR2X2 OR2X2_2126 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_2__29_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1288) );
  OR2X2 OR2X2_2127 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf0), .B(1'b0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1289) );
  OR2X2 OR2X2_2128 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf3), .B(u_wb2sdrc_u_cmdfifo_mem_2__30_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1291) );
  OR2X2 OR2X2_2129 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf5), .B(1'b0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1292) );
  OR2X2 OR2X2_213 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n403_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n399_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n404_1) );
  OR2X2 OR2X2_2130 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf2), .B(u_wb2sdrc_u_cmdfifo_mem_2__31_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1294) );
  OR2X2 OR2X2_2131 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf4), .B(1'b0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1295) );
  OR2X2 OR2X2_2132 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf1), .B(u_wb2sdrc_u_cmdfifo_mem_2__32_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1297) );
  OR2X2 OR2X2_2133 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf3), .B(1'b0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1298) );
  OR2X2 OR2X2_2134 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf0), .B(u_wb2sdrc_u_cmdfifo_mem_2__33_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1300) );
  OR2X2 OR2X2_2135 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf2), .B(1'b0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1301) );
  OR2X2 OR2X2_2136 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf5), .B(u_wb2sdrc_u_cmdfifo_mem_2__34_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1303) );
  OR2X2 OR2X2_2137 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf1), .B(1'b0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1304) );
  OR2X2 OR2X2_2138 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n627_bF_buf4), .B(u_wb2sdrc_u_cmdfifo_mem_2__35_), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1306) );
  OR2X2 OR2X2_2139 ( .A(u_wb2sdrc_u_cmdfifo__abc_18561_n1201_bF_buf0), .B(1'b0), .Y(u_wb2sdrc_u_cmdfifo__abc_18561_n1307) );
  OR2X2 OR2X2_214 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n406_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n382), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n407_1) );
  OR2X2 OR2X2_2140 ( .A(u_wb2sdrc_u_rddatafifo_sync_wr_ptr_1_1_), .B(u_wb2sdrc_u_rddatafifo_sync_wr_ptr_2_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n410) );
  OR2X2 OR2X2_2141 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n416_1), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n414), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n417) );
  OR2X2 OR2X2_2142 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n420_1), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n422), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n423_1) );
  OR2X2 OR2X2_2143 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n423_1), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n419_1_bF_buf5), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n424_1) );
  OR2X2 OR2X2_2144 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n426), .B(u_wb2sdrc_u_rddatafifo_rd_ptr_2_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n427_1) );
  OR2X2 OR2X2_2145 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n428_1), .B(u_wb2sdrc_u_rddatafifo_sync_wr_ptr_2_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n429) );
  OR2X2 OR2X2_2146 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n450_1), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n448), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n98) );
  OR2X2 OR2X2_2147 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n453_1), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n452_1), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n101) );
  OR2X2 OR2X2_2148 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n456_1), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n455_1), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n104) );
  OR2X2 OR2X2_2149 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n459_1), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n458_1), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n107) );
  OR2X2 OR2X2_215 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n383_1), .B(\cfg_sdr_tras_d[3] ), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n408_1) );
  OR2X2 OR2X2_2150 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n462_1), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n461_1), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n110) );
  OR2X2 OR2X2_2151 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n465_1), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n464_1), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n113) );
  OR2X2 OR2X2_2152 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n468_1), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n467_1), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n116) );
  OR2X2 OR2X2_2153 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n471_1), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n470_1), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n119) );
  OR2X2 OR2X2_2154 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n474_1), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n473_1), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n122) );
  OR2X2 OR2X2_2155 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n477_1), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n476_1), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n125) );
  OR2X2 OR2X2_2156 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n480_1), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n479_1), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n128) );
  OR2X2 OR2X2_2157 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n483_1), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n482_1), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n131) );
  OR2X2 OR2X2_2158 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n486_1), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n485), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n134) );
  OR2X2 OR2X2_2159 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n489_1), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n488), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n137) );
  OR2X2 OR2X2_216 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n380), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_cmd_0_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n411_1) );
  OR2X2 OR2X2_2160 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n492), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n491), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n140) );
  OR2X2 OR2X2_2161 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n495_1), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n494), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n143) );
  OR2X2 OR2X2_2162 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n498), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n497), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n146) );
  OR2X2 OR2X2_2163 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n501_1), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n500_1), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n149) );
  OR2X2 OR2X2_2164 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n504), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n503_1), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n152) );
  OR2X2 OR2X2_2165 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n507), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n506), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n155) );
  OR2X2 OR2X2_2166 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n510_1), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n509_1), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n158) );
  OR2X2 OR2X2_2167 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n513), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n512), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n161) );
  OR2X2 OR2X2_2168 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n516), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n515), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n164) );
  OR2X2 OR2X2_2169 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n519), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n518), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n167) );
  OR2X2 OR2X2_217 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_timer0_2_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_timer0_3_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n414_1) );
  OR2X2 OR2X2_2170 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n522_1), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n521_1), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n170) );
  OR2X2 OR2X2_2171 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n525), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n524_1), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n173) );
  OR2X2 OR2X2_2172 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n528), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n527_1), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n176) );
  OR2X2 OR2X2_2173 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n531), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n530), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n179) );
  OR2X2 OR2X2_2174 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n534), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n533), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n182) );
  OR2X2 OR2X2_2175 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n537), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n536), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n185) );
  OR2X2 OR2X2_2176 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n540), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n539), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n188) );
  OR2X2 OR2X2_2177 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n543), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n542), .Y(u_wb2sdrc_u_rddatafifo__abc_14216_n191) );
  OR2X2 OR2X2_2178 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_0__0_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n550) );
  OR2X2 OR2X2_2179 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf4), .B(app_rd_data_0_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n552) );
  OR2X2 OR2X2_218 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n414_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_timer0_1_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n415_1) );
  OR2X2 OR2X2_2180 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_0__1_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n554) );
  OR2X2 OR2X2_2181 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf3), .B(app_rd_data_1_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n555) );
  OR2X2 OR2X2_2182 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_0__2_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n557) );
  OR2X2 OR2X2_2183 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf2), .B(app_rd_data_2_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n558) );
  OR2X2 OR2X2_2184 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_0__3_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n560) );
  OR2X2 OR2X2_2185 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf1), .B(app_rd_data_3_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n561) );
  OR2X2 OR2X2_2186 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_0__4_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n563) );
  OR2X2 OR2X2_2187 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf0), .B(app_rd_data_4_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n564) );
  OR2X2 OR2X2_2188 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_0__5_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n566) );
  OR2X2 OR2X2_2189 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf4), .B(app_rd_data_5_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n567) );
  OR2X2 OR2X2_219 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n416), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n382), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n417_1) );
  OR2X2 OR2X2_2190 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_0__6_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n569) );
  OR2X2 OR2X2_2191 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf3), .B(app_rd_data_6_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n570) );
  OR2X2 OR2X2_2192 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_0__7_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n572) );
  OR2X2 OR2X2_2193 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf2), .B(app_rd_data_7_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n573) );
  OR2X2 OR2X2_2194 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_0__8_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n575) );
  OR2X2 OR2X2_2195 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf1), .B(app_rd_data_8_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n576) );
  OR2X2 OR2X2_2196 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_0__9_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n578) );
  OR2X2 OR2X2_2197 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf0), .B(app_rd_data_9_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n579) );
  OR2X2 OR2X2_2198 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_0__10_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n581) );
  OR2X2 OR2X2_2199 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf4), .B(app_rd_data_10_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n582) );
  OR2X2 OR2X2_22 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n275_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n267_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n276) );
  OR2X2 OR2X2_220 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n380), .B(\cfg_sdr_trcd_d[0] ), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n418) );
  OR2X2 OR2X2_2200 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_0__11_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n584) );
  OR2X2 OR2X2_2201 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf3), .B(app_rd_data_11_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n585) );
  OR2X2 OR2X2_2202 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_0__12_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n587) );
  OR2X2 OR2X2_2203 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf2), .B(app_rd_data_12_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n588) );
  OR2X2 OR2X2_2204 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_0__13_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n590) );
  OR2X2 OR2X2_2205 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf1), .B(app_rd_data_13_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n591) );
  OR2X2 OR2X2_2206 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_0__14_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n593) );
  OR2X2 OR2X2_2207 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf0), .B(app_rd_data_14_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n594) );
  OR2X2 OR2X2_2208 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_0__15_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n596) );
  OR2X2 OR2X2_2209 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf4), .B(app_rd_data_15_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n597) );
  OR2X2 OR2X2_221 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n419_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n412_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n420_1) );
  OR2X2 OR2X2_2210 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_0__16_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n599) );
  OR2X2 OR2X2_2211 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf3), .B(app_rd_data_16_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n600) );
  OR2X2 OR2X2_2212 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_0__17_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n602) );
  OR2X2 OR2X2_2213 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf2), .B(app_rd_data_17_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n603) );
  OR2X2 OR2X2_2214 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_0__18_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n605) );
  OR2X2 OR2X2_2215 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf1), .B(app_rd_data_18_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n606) );
  OR2X2 OR2X2_2216 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_0__19_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n608) );
  OR2X2 OR2X2_2217 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf0), .B(app_rd_data_19_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n609) );
  OR2X2 OR2X2_2218 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_0__20_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n611) );
  OR2X2 OR2X2_2219 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf4), .B(app_rd_data_20_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n612) );
  OR2X2 OR2X2_222 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n411_1), .B(\cfg_sdr_trp_d[0] ), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n421) );
  OR2X2 OR2X2_2220 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_0__21_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n614) );
  OR2X2 OR2X2_2221 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf3), .B(app_rd_data_21_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n615) );
  OR2X2 OR2X2_2222 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_0__22_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n617) );
  OR2X2 OR2X2_2223 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf2), .B(app_rd_data_22_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n618) );
  OR2X2 OR2X2_2224 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_0__23_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n620) );
  OR2X2 OR2X2_2225 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf1), .B(app_rd_data_23_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n621) );
  OR2X2 OR2X2_2226 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_0__24_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n623) );
  OR2X2 OR2X2_2227 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf0), .B(app_rd_data_24_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n624) );
  OR2X2 OR2X2_2228 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_0__25_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n626) );
  OR2X2 OR2X2_2229 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf4), .B(app_rd_data_25_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n627) );
  OR2X2 OR2X2_223 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_timer0_1_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_timer0_0_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n424) );
  OR2X2 OR2X2_2230 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_0__26_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n629) );
  OR2X2 OR2X2_2231 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf3), .B(app_rd_data_26_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n630) );
  OR2X2 OR2X2_2232 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_0__27_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n632) );
  OR2X2 OR2X2_2233 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf2), .B(app_rd_data_27_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n633) );
  OR2X2 OR2X2_2234 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_0__28_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n635) );
  OR2X2 OR2X2_2235 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf1), .B(app_rd_data_28_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n636) );
  OR2X2 OR2X2_2236 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_0__29_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n638) );
  OR2X2 OR2X2_2237 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf0), .B(app_rd_data_29_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n639) );
  OR2X2 OR2X2_2238 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_0__30_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n641) );
  OR2X2 OR2X2_2239 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf4), .B(app_rd_data_30_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n642) );
  OR2X2 OR2X2_224 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n425), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n426), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n427_1) );
  OR2X2 OR2X2_2240 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n549_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_0__31_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n644) );
  OR2X2 OR2X2_2241 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n551_bF_buf3), .B(app_rd_data_31_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n645) );
  OR2X2 OR2X2_2242 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_2__0_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n651) );
  OR2X2 OR2X2_2243 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf4), .B(app_rd_data_0_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n653) );
  OR2X2 OR2X2_2244 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_2__1_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n655) );
  OR2X2 OR2X2_2245 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf3), .B(app_rd_data_1_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n656) );
  OR2X2 OR2X2_2246 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_2__2_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n658) );
  OR2X2 OR2X2_2247 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf2), .B(app_rd_data_2_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n659) );
  OR2X2 OR2X2_2248 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_2__3_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n661) );
  OR2X2 OR2X2_2249 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf1), .B(app_rd_data_3_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n662) );
  OR2X2 OR2X2_225 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n414_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n424), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n428_1) );
  OR2X2 OR2X2_2250 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_2__4_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n664) );
  OR2X2 OR2X2_2251 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf0), .B(app_rd_data_4_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n665) );
  OR2X2 OR2X2_2252 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_2__5_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n667) );
  OR2X2 OR2X2_2253 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf4), .B(app_rd_data_5_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n668) );
  OR2X2 OR2X2_2254 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_2__6_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n670) );
  OR2X2 OR2X2_2255 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf3), .B(app_rd_data_6_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n671) );
  OR2X2 OR2X2_2256 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_2__7_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n673) );
  OR2X2 OR2X2_2257 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf2), .B(app_rd_data_7_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n674) );
  OR2X2 OR2X2_2258 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_2__8_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n676) );
  OR2X2 OR2X2_2259 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf1), .B(app_rd_data_8_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n677) );
  OR2X2 OR2X2_226 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n412_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n431_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n432) );
  OR2X2 OR2X2_2260 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_2__9_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n679) );
  OR2X2 OR2X2_2261 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf0), .B(app_rd_data_9_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n680) );
  OR2X2 OR2X2_2262 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_2__10_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n682) );
  OR2X2 OR2X2_2263 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf4), .B(app_rd_data_10_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n683) );
  OR2X2 OR2X2_2264 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_2__11_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n685) );
  OR2X2 OR2X2_2265 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf3), .B(app_rd_data_11_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n686) );
  OR2X2 OR2X2_2266 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_2__12_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n688) );
  OR2X2 OR2X2_2267 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf2), .B(app_rd_data_12_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n689) );
  OR2X2 OR2X2_2268 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_2__13_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n691) );
  OR2X2 OR2X2_2269 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf1), .B(app_rd_data_13_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n692) );
  OR2X2 OR2X2_227 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n430), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n432), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n433) );
  OR2X2 OR2X2_2270 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_2__14_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n694) );
  OR2X2 OR2X2_2271 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf0), .B(app_rd_data_14_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n695) );
  OR2X2 OR2X2_2272 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_2__15_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n697) );
  OR2X2 OR2X2_2273 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf4), .B(app_rd_data_15_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n698) );
  OR2X2 OR2X2_2274 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_2__16_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n700) );
  OR2X2 OR2X2_2275 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf3), .B(app_rd_data_16_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n701) );
  OR2X2 OR2X2_2276 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_2__17_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n703) );
  OR2X2 OR2X2_2277 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf2), .B(app_rd_data_17_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n704) );
  OR2X2 OR2X2_2278 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_2__18_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n706) );
  OR2X2 OR2X2_2279 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf1), .B(app_rd_data_18_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n707) );
  OR2X2 OR2X2_228 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n411_1), .B(\cfg_sdr_trp_d[1] ), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n434_1) );
  OR2X2 OR2X2_2280 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_2__19_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n709) );
  OR2X2 OR2X2_2281 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf0), .B(app_rd_data_19_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n710) );
  OR2X2 OR2X2_2282 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_2__20_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n712) );
  OR2X2 OR2X2_2283 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf4), .B(app_rd_data_20_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n713) );
  OR2X2 OR2X2_2284 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_2__21_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n715) );
  OR2X2 OR2X2_2285 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf3), .B(app_rd_data_21_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n716) );
  OR2X2 OR2X2_2286 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_2__22_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n718) );
  OR2X2 OR2X2_2287 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf2), .B(app_rd_data_22_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n719) );
  OR2X2 OR2X2_2288 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_2__23_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n721) );
  OR2X2 OR2X2_2289 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf1), .B(app_rd_data_23_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n722) );
  OR2X2 OR2X2_229 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n424), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_timer0_2_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n437_1) );
  OR2X2 OR2X2_2290 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_2__24_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n724) );
  OR2X2 OR2X2_2291 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf0), .B(app_rd_data_24_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n725) );
  OR2X2 OR2X2_2292 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_2__25_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n727) );
  OR2X2 OR2X2_2293 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf4), .B(app_rd_data_25_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n728) );
  OR2X2 OR2X2_2294 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_2__26_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n730) );
  OR2X2 OR2X2_2295 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf3), .B(app_rd_data_26_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n731) );
  OR2X2 OR2X2_2296 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_2__27_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n733) );
  OR2X2 OR2X2_2297 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf2), .B(app_rd_data_27_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n734) );
  OR2X2 OR2X2_2298 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_2__28_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n736) );
  OR2X2 OR2X2_2299 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf1), .B(app_rd_data_28_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n737) );
  OR2X2 OR2X2_23 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n285), .B(u_sdrc_core_u_bank_ctl__abc_21249_n287_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n288_1) );
  OR2X2 OR2X2_230 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n438_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n439_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n440_1) );
  OR2X2 OR2X2_2300 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_2__29_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n739) );
  OR2X2 OR2X2_2301 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf0), .B(app_rd_data_29_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n740) );
  OR2X2 OR2X2_2302 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_2__30_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n742) );
  OR2X2 OR2X2_2303 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf4), .B(app_rd_data_30_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n743) );
  OR2X2 OR2X2_2304 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n650_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_2__31_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n745) );
  OR2X2 OR2X2_2305 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n652_bF_buf3), .B(app_rd_data_31_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n746) );
  OR2X2 OR2X2_2306 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n751), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n752), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n753) );
  OR2X2 OR2X2_2307 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n758), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n756), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n759) );
  OR2X2 OR2X2_2308 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n754), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n759), .Y(_auto_iopadmap_cc_313_execute_24709_0_) );
  OR2X2 OR2X2_2309 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n761), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n762), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n763) );
  OR2X2 OR2X2_231 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n412_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n442), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n443) );
  OR2X2 OR2X2_2310 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n766), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n765), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n767) );
  OR2X2 OR2X2_2311 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n764), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n767), .Y(_auto_iopadmap_cc_313_execute_24709_1_) );
  OR2X2 OR2X2_2312 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n769), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n770), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n771) );
  OR2X2 OR2X2_2313 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n774), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n773), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n775) );
  OR2X2 OR2X2_2314 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n772), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n775), .Y(_auto_iopadmap_cc_313_execute_24709_2_) );
  OR2X2 OR2X2_2315 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n777), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n778), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n779) );
  OR2X2 OR2X2_2316 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n782), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n781), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n783) );
  OR2X2 OR2X2_2317 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n780), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n783), .Y(_auto_iopadmap_cc_313_execute_24709_3_) );
  OR2X2 OR2X2_2318 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n785), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n786), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n787) );
  OR2X2 OR2X2_2319 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n790), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n789), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n791) );
  OR2X2 OR2X2_232 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n441), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n443), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n444_1) );
  OR2X2 OR2X2_2320 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n788), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n791), .Y(_auto_iopadmap_cc_313_execute_24709_4_) );
  OR2X2 OR2X2_2321 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n793), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n794), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n795) );
  OR2X2 OR2X2_2322 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n798), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n797), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n799) );
  OR2X2 OR2X2_2323 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n796), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n799), .Y(_auto_iopadmap_cc_313_execute_24709_5_) );
  OR2X2 OR2X2_2324 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n801), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n802), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n803) );
  OR2X2 OR2X2_2325 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n806), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n805), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n807) );
  OR2X2 OR2X2_2326 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n804), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n807), .Y(_auto_iopadmap_cc_313_execute_24709_6_) );
  OR2X2 OR2X2_2327 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n809), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n810), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n811) );
  OR2X2 OR2X2_2328 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n814), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n813), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n815) );
  OR2X2 OR2X2_2329 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n812), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n815), .Y(_auto_iopadmap_cc_313_execute_24709_7_) );
  OR2X2 OR2X2_233 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n411_1), .B(\cfg_sdr_trp_d[2] ), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n445_1) );
  OR2X2 OR2X2_2330 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n817), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n818), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n819) );
  OR2X2 OR2X2_2331 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n822), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n821), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n823) );
  OR2X2 OR2X2_2332 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n820), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n823), .Y(_auto_iopadmap_cc_313_execute_24709_8_) );
  OR2X2 OR2X2_2333 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n825), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n826), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n827) );
  OR2X2 OR2X2_2334 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n830), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n829), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n831) );
  OR2X2 OR2X2_2335 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n828), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n831), .Y(_auto_iopadmap_cc_313_execute_24709_9_) );
  OR2X2 OR2X2_2336 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n833), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n834), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n835) );
  OR2X2 OR2X2_2337 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n838), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n837), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n839) );
  OR2X2 OR2X2_2338 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n836), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n839), .Y(_auto_iopadmap_cc_313_execute_24709_10_) );
  OR2X2 OR2X2_2339 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n841), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n842), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n843) );
  OR2X2 OR2X2_234 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n448_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n382), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n449_1) );
  OR2X2 OR2X2_2340 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n846), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n845), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n847) );
  OR2X2 OR2X2_2341 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n844), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n847), .Y(_auto_iopadmap_cc_313_execute_24709_11_) );
  OR2X2 OR2X2_2342 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n849), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n850), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n851) );
  OR2X2 OR2X2_2343 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n854), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n853), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n855) );
  OR2X2 OR2X2_2344 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n852), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n855), .Y(_auto_iopadmap_cc_313_execute_24709_12_) );
  OR2X2 OR2X2_2345 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n857), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n858), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n859) );
  OR2X2 OR2X2_2346 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n862), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n861), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n863) );
  OR2X2 OR2X2_2347 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n860), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n863), .Y(_auto_iopadmap_cc_313_execute_24709_13_) );
  OR2X2 OR2X2_2348 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n865), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n866), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n867) );
  OR2X2 OR2X2_2349 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n870), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n869), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n871) );
  OR2X2 OR2X2_235 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n380), .B(\cfg_sdr_trcd_d[3] ), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n450) );
  OR2X2 OR2X2_2350 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n868), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n871), .Y(_auto_iopadmap_cc_313_execute_24709_14_) );
  OR2X2 OR2X2_2351 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n873), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n874), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n875) );
  OR2X2 OR2X2_2352 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n878), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n877), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n879) );
  OR2X2 OR2X2_2353 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n876), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n879), .Y(_auto_iopadmap_cc_313_execute_24709_15_) );
  OR2X2 OR2X2_2354 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n881), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n882), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n883) );
  OR2X2 OR2X2_2355 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n886), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n885), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n887) );
  OR2X2 OR2X2_2356 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n884), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n887), .Y(_auto_iopadmap_cc_313_execute_24709_16_) );
  OR2X2 OR2X2_2357 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n889), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n890), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n891) );
  OR2X2 OR2X2_2358 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n894), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n893), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n895) );
  OR2X2 OR2X2_2359 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n892), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n895), .Y(_auto_iopadmap_cc_313_execute_24709_17_) );
  OR2X2 OR2X2_236 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n451), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n412_1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n452) );
  OR2X2 OR2X2_2360 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n897), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n898), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n899) );
  OR2X2 OR2X2_2361 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n902), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n901), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n903) );
  OR2X2 OR2X2_2362 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n900), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n903), .Y(_auto_iopadmap_cc_313_execute_24709_18_) );
  OR2X2 OR2X2_2363 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n905), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n906), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n907) );
  OR2X2 OR2X2_2364 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n910), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n909), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n911) );
  OR2X2 OR2X2_2365 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n908), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n911), .Y(_auto_iopadmap_cc_313_execute_24709_19_) );
  OR2X2 OR2X2_2366 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n913), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n914), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n915) );
  OR2X2 OR2X2_2367 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n918), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n917), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n919) );
  OR2X2 OR2X2_2368 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n916), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n919), .Y(_auto_iopadmap_cc_313_execute_24709_20_) );
  OR2X2 OR2X2_2369 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n921), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n922), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n923) );
  OR2X2 OR2X2_237 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n411_1), .B(\cfg_sdr_trp_d[3] ), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n453_1) );
  OR2X2 OR2X2_2370 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n926), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n925), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n927) );
  OR2X2 OR2X2_2371 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n924), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n927), .Y(_auto_iopadmap_cc_313_execute_24709_21_) );
  OR2X2 OR2X2_2372 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n929), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n930), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n931) );
  OR2X2 OR2X2_2373 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n934), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n933), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n935) );
  OR2X2 OR2X2_2374 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n932), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n935), .Y(_auto_iopadmap_cc_313_execute_24709_22_) );
  OR2X2 OR2X2_2375 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n937), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n938), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n939) );
  OR2X2 OR2X2_2376 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n942), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n941), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n943) );
  OR2X2 OR2X2_2377 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n940), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n943), .Y(_auto_iopadmap_cc_313_execute_24709_23_) );
  OR2X2 OR2X2_2378 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n945), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n946), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n947) );
  OR2X2 OR2X2_2379 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n950), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n949), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n951) );
  OR2X2 OR2X2_238 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n473), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n475), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_0__FF_INPUT) );
  OR2X2 OR2X2_2380 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n948), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n951), .Y(_auto_iopadmap_cc_313_execute_24709_24_) );
  OR2X2 OR2X2_2381 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n953), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n954), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n955) );
  OR2X2 OR2X2_2382 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n958), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n957), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n959) );
  OR2X2 OR2X2_2383 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n956), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n959), .Y(_auto_iopadmap_cc_313_execute_24709_25_) );
  OR2X2 OR2X2_2384 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n961), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n962), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n963) );
  OR2X2 OR2X2_2385 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n966), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n965), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n967) );
  OR2X2 OR2X2_2386 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n964), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n967), .Y(_auto_iopadmap_cc_313_execute_24709_26_) );
  OR2X2 OR2X2_2387 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n969), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n970), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n971) );
  OR2X2 OR2X2_2388 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n974), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n973), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n975) );
  OR2X2 OR2X2_2389 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n972), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n975), .Y(_auto_iopadmap_cc_313_execute_24709_27_) );
  OR2X2 OR2X2_239 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n477), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n479), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_1__FF_INPUT) );
  OR2X2 OR2X2_2390 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n977), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n978), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n979) );
  OR2X2 OR2X2_2391 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n982), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n981), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n983) );
  OR2X2 OR2X2_2392 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n980), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n983), .Y(_auto_iopadmap_cc_313_execute_24709_28_) );
  OR2X2 OR2X2_2393 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n985), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n986), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n987) );
  OR2X2 OR2X2_2394 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n990), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n989), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n991) );
  OR2X2 OR2X2_2395 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n988), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n991), .Y(_auto_iopadmap_cc_313_execute_24709_29_) );
  OR2X2 OR2X2_2396 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n993), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n994), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n995) );
  OR2X2 OR2X2_2397 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n998), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n997), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n999) );
  OR2X2 OR2X2_2398 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n996), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n999), .Y(_auto_iopadmap_cc_313_execute_24709_30_) );
  OR2X2 OR2X2_2399 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1001), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1002), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1003) );
  OR2X2 OR2X2_24 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n289_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n290), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n291_1) );
  OR2X2 OR2X2_240 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n481), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n483), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_2__FF_INPUT) );
  OR2X2 OR2X2_2400 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1006), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1005), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1007) );
  OR2X2 OR2X2_2401 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1004), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1007), .Y(_auto_iopadmap_cc_313_execute_24709_31_) );
  OR2X2 OR2X2_2402 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_1__0_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1019) );
  OR2X2 OR2X2_2403 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf4), .B(app_rd_data_0_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1021) );
  OR2X2 OR2X2_2404 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_1__1_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1023) );
  OR2X2 OR2X2_2405 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf3), .B(app_rd_data_1_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1024) );
  OR2X2 OR2X2_2406 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_1__2_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1026) );
  OR2X2 OR2X2_2407 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf2), .B(app_rd_data_2_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1027) );
  OR2X2 OR2X2_2408 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_1__3_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1029) );
  OR2X2 OR2X2_2409 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf1), .B(app_rd_data_3_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1030) );
  OR2X2 OR2X2_241 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n485), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n487), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_3__FF_INPUT) );
  OR2X2 OR2X2_2410 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_1__4_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1032) );
  OR2X2 OR2X2_2411 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf0), .B(app_rd_data_4_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1033) );
  OR2X2 OR2X2_2412 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_1__5_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1035) );
  OR2X2 OR2X2_2413 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf4), .B(app_rd_data_5_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1036) );
  OR2X2 OR2X2_2414 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_1__6_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1038) );
  OR2X2 OR2X2_2415 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf3), .B(app_rd_data_6_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1039) );
  OR2X2 OR2X2_2416 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_1__7_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1041) );
  OR2X2 OR2X2_2417 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf2), .B(app_rd_data_7_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1042) );
  OR2X2 OR2X2_2418 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_1__8_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1044) );
  OR2X2 OR2X2_2419 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf1), .B(app_rd_data_8_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1045) );
  OR2X2 OR2X2_242 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n489), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n491), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_4__FF_INPUT) );
  OR2X2 OR2X2_2420 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_1__9_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1047) );
  OR2X2 OR2X2_2421 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf0), .B(app_rd_data_9_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1048) );
  OR2X2 OR2X2_2422 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_1__10_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1050) );
  OR2X2 OR2X2_2423 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf4), .B(app_rd_data_10_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1051) );
  OR2X2 OR2X2_2424 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_1__11_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1053) );
  OR2X2 OR2X2_2425 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf3), .B(app_rd_data_11_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1054) );
  OR2X2 OR2X2_2426 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_1__12_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1056) );
  OR2X2 OR2X2_2427 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf2), .B(app_rd_data_12_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1057) );
  OR2X2 OR2X2_2428 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_1__13_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1059) );
  OR2X2 OR2X2_2429 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf1), .B(app_rd_data_13_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1060) );
  OR2X2 OR2X2_243 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n493), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n495), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_5__FF_INPUT) );
  OR2X2 OR2X2_2430 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_1__14_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1062) );
  OR2X2 OR2X2_2431 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf0), .B(app_rd_data_14_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1063) );
  OR2X2 OR2X2_2432 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_1__15_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1065) );
  OR2X2 OR2X2_2433 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf4), .B(app_rd_data_15_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1066) );
  OR2X2 OR2X2_2434 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_1__16_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1068) );
  OR2X2 OR2X2_2435 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf3), .B(app_rd_data_16_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1069) );
  OR2X2 OR2X2_2436 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_1__17_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1071) );
  OR2X2 OR2X2_2437 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf2), .B(app_rd_data_17_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1072) );
  OR2X2 OR2X2_2438 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_1__18_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1074) );
  OR2X2 OR2X2_2439 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf1), .B(app_rd_data_18_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1075) );
  OR2X2 OR2X2_244 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n497), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n499), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_6__FF_INPUT) );
  OR2X2 OR2X2_2440 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_1__19_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1077) );
  OR2X2 OR2X2_2441 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf0), .B(app_rd_data_19_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1078) );
  OR2X2 OR2X2_2442 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_1__20_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1080) );
  OR2X2 OR2X2_2443 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf4), .B(app_rd_data_20_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1081) );
  OR2X2 OR2X2_2444 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_1__21_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1083) );
  OR2X2 OR2X2_2445 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf3), .B(app_rd_data_21_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1084) );
  OR2X2 OR2X2_2446 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_1__22_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1086) );
  OR2X2 OR2X2_2447 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf2), .B(app_rd_data_22_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1087) );
  OR2X2 OR2X2_2448 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_1__23_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1089) );
  OR2X2 OR2X2_2449 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf1), .B(app_rd_data_23_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1090) );
  OR2X2 OR2X2_245 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n501), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n502), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n503) );
  OR2X2 OR2X2_2450 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_1__24_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1092) );
  OR2X2 OR2X2_2451 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf0), .B(app_rd_data_24_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1093) );
  OR2X2 OR2X2_2452 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_1__25_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1095) );
  OR2X2 OR2X2_2453 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf4), .B(app_rd_data_25_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1096) );
  OR2X2 OR2X2_2454 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_1__26_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1098) );
  OR2X2 OR2X2_2455 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf3), .B(app_rd_data_26_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1099) );
  OR2X2 OR2X2_2456 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf1), .B(u_wb2sdrc_u_rddatafifo_mem_1__27_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1101) );
  OR2X2 OR2X2_2457 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf2), .B(app_rd_data_27_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1102) );
  OR2X2 OR2X2_2458 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf0), .B(u_wb2sdrc_u_rddatafifo_mem_1__28_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1104) );
  OR2X2 OR2X2_2459 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf1), .B(app_rd_data_28_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1105) );
  OR2X2 OR2X2_246 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n505), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n506), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n507) );
  OR2X2 OR2X2_2460 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf4), .B(u_wb2sdrc_u_rddatafifo_mem_1__29_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1107) );
  OR2X2 OR2X2_2461 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf0), .B(app_rd_data_29_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1108) );
  OR2X2 OR2X2_2462 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf3), .B(u_wb2sdrc_u_rddatafifo_mem_1__30_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1110) );
  OR2X2 OR2X2_2463 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf4), .B(app_rd_data_30_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1111) );
  OR2X2 OR2X2_2464 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1018_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_mem_1__31_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1113) );
  OR2X2 OR2X2_2465 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1020_bF_buf3), .B(app_rd_data_31_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1114) );
  OR2X2 OR2X2_2466 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1120), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1121), .Y(u_wb2sdrc_u_rddatafifo_rd_ptr_0__FF_INPUT) );
  OR2X2 OR2X2_2467 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n757_bF_buf2), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1124), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1125) );
  OR2X2 OR2X2_2468 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1126), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1123), .Y(u_wb2sdrc_u_rddatafifo_rd_ptr_1__FF_INPUT) );
  OR2X2 OR2X2_2469 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n755_bF_buf2), .B(u_wb2sdrc_u_rddatafifo_rd_ptr_2_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1129) );
  OR2X2 OR2X2_247 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n509), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n510), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n511) );
  OR2X2 OR2X2_2470 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1133), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1128), .Y(u_wb2sdrc_u_rddatafifo_rd_ptr_2__FF_INPUT) );
  OR2X2 OR2X2_2471 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1017), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1152), .Y(u_wb2sdrc_u_rddatafifo_grey_wr_ptr_0__FF_INPUT) );
  OR2X2 OR2X2_2472 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1154), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n446), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1155) );
  OR2X2 OR2X2_2473 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n446), .B(u_wb2sdrc_u_rddatafifo_wr_ptr_2_), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1158) );
  OR2X2 OR2X2_2474 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1165), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1162), .Y(u_wb2sdrc_u_rddatafifo__abc_17752_n1166) );
  OR2X2 OR2X2_2475 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1166), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1161), .Y(u_wb2sdrc_u_rddatafifo_grey_wr_ptr_1__FF_INPUT) );
  OR2X2 OR2X2_2476 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1160), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1168), .Y(u_wb2sdrc_u_rddatafifo_grey_wr_ptr_2__FF_INPUT) );
  OR2X2 OR2X2_2477 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n548), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1170), .Y(u_wb2sdrc_u_rddatafifo_wr_ptr_0__FF_INPUT) );
  OR2X2 OR2X2_2478 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1164), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1172), .Y(u_wb2sdrc_u_rddatafifo_wr_ptr_1__FF_INPUT) );
  OR2X2 OR2X2_2479 ( .A(u_wb2sdrc_u_rddatafifo__abc_17752_n1160), .B(u_wb2sdrc_u_rddatafifo__abc_17752_n1174), .Y(u_wb2sdrc_u_rddatafifo_wr_ptr_2__FF_INPUT) );
  OR2X2 OR2X2_248 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n513), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n514), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n515) );
  OR2X2 OR2X2_2480 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n698), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n699_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n700) );
  OR2X2 OR2X2_2481 ( .A(u_wb2sdrc_u_wrdatafifo_sync_rd_ptr_1_2_), .B(u_wb2sdrc_u_wrdatafifo_sync_rd_ptr_1_3_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n703) );
  OR2X2 OR2X2_2482 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n705_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n702_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n706) );
  OR2X2 OR2X2_2483 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n700), .B(u_wb2sdrc_u_wrdatafifo_sync_rd_ptr_1_1_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n707) );
  OR2X2 OR2X2_2484 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n711_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n712), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n713) );
  OR2X2 OR2X2_2485 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n713), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n705_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n714_1) );
  OR2X2 OR2X2_2486 ( .A(u_wb2sdrc_u_wrdatafifo_sync_rd_ptr_1_0_), .B(u_wb2sdrc_u_wrdatafifo_sync_rd_ptr_1_1_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n715) );
  OR2X2 OR2X2_2487 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n700), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n717_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n718) );
  OR2X2 OR2X2_2488 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n719), .B(u_wb2sdrc_u_wrdatafifo_wr_ptr_0_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n720_1) );
  OR2X2 OR2X2_2489 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n708_1), .B(u_wb2sdrc_u_wrdatafifo_wr_ptr_1_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n721_1) );
  OR2X2 OR2X2_249 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n517), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n518), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n519) );
  OR2X2 OR2X2_2490 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n722), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n709_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n723_1) );
  OR2X2 OR2X2_2491 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n701), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n725), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n726_1) );
  OR2X2 OR2X2_2492 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n728_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n701), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n729_1) );
  OR2X2 OR2X2_2493 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n697_1), .B(u_wb2sdrc_u_wrdatafifo_wr_ptr_3_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n730) );
  OR2X2 OR2X2_2494 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n731), .B(u_wb2sdrc_u_wrdatafifo_sync_rd_ptr_1_3_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n732_1) );
  OR2X2 OR2X2_2495 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n729_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n734), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n735_1) );
  OR2X2 OR2X2_2496 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n739), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n740_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n741_1) );
  OR2X2 OR2X2_2497 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n744_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n745_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n746) );
  OR2X2 OR2X2_2498 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n742), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n747_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n748) );
  OR2X2 OR2X2_2499 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n749), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n726_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n750_1) );
  OR2X2 OR2X2_25 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n292_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n293), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n294_1) );
  OR2X2 OR2X2_250 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n521), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n522), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n523) );
  OR2X2 OR2X2_2500 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n751), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n733_1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n752_1) );
  OR2X2 OR2X2_2501 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n754), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n719), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n755) );
  OR2X2 OR2X2_2502 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n758), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n742), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n759_1) );
  OR2X2 OR2X2_2503 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n723_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n727), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n760) );
  OR2X2 OR2X2_2504 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_0__0_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n820_1) );
  OR2X2 OR2X2_2505 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf5), .B(\wb_dat_i[0] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n822_1) );
  OR2X2 OR2X2_2506 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_0__1_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n824_1) );
  OR2X2 OR2X2_2507 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf4), .B(\wb_dat_i[1] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n825_1) );
  OR2X2 OR2X2_2508 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_0__2_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n827_1) );
  OR2X2 OR2X2_2509 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf3), .B(\wb_dat_i[2] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n828_1) );
  OR2X2 OR2X2_251 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n525), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n526), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n527) );
  OR2X2 OR2X2_2510 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_0__3_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n830_1) );
  OR2X2 OR2X2_2511 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf2), .B(\wb_dat_i[3] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n831_1) );
  OR2X2 OR2X2_2512 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_0__4_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n833_1) );
  OR2X2 OR2X2_2513 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf1), .B(\wb_dat_i[4] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n834_1) );
  OR2X2 OR2X2_2514 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_0__5_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n836_1) );
  OR2X2 OR2X2_2515 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf0), .B(\wb_dat_i[5] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n837_1) );
  OR2X2 OR2X2_2516 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_0__6_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n839_1) );
  OR2X2 OR2X2_2517 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf5), .B(\wb_dat_i[6] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n840_1) );
  OR2X2 OR2X2_2518 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_0__7_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n842_1) );
  OR2X2 OR2X2_2519 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf4), .B(\wb_dat_i[7] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n843) );
  OR2X2 OR2X2_252 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n529), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n530), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n531) );
  OR2X2 OR2X2_2520 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_0__8_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n845_1) );
  OR2X2 OR2X2_2521 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf3), .B(\wb_dat_i[8] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n846_1) );
  OR2X2 OR2X2_2522 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_0__9_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n848_1) );
  OR2X2 OR2X2_2523 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf2), .B(\wb_dat_i[9] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n849_1) );
  OR2X2 OR2X2_2524 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_0__10_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n851_1) );
  OR2X2 OR2X2_2525 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf1), .B(\wb_dat_i[10] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n852_1) );
  OR2X2 OR2X2_2526 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_0__11_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n854_1) );
  OR2X2 OR2X2_2527 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf0), .B(\wb_dat_i[11] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n855_1) );
  OR2X2 OR2X2_2528 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_0__12_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n857_1) );
  OR2X2 OR2X2_2529 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf5), .B(\wb_dat_i[12] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n858_1) );
  OR2X2 OR2X2_253 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n533), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n534), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n535) );
  OR2X2 OR2X2_2530 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_0__13_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n860_1) );
  OR2X2 OR2X2_2531 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf4), .B(\wb_dat_i[13] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n861_1) );
  OR2X2 OR2X2_2532 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_0__14_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n863_1) );
  OR2X2 OR2X2_2533 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf3), .B(\wb_dat_i[14] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n864_1) );
  OR2X2 OR2X2_2534 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_0__15_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n866_1) );
  OR2X2 OR2X2_2535 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf2), .B(\wb_dat_i[15] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n867_1) );
  OR2X2 OR2X2_2536 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_0__16_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n869_1) );
  OR2X2 OR2X2_2537 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf1), .B(\wb_dat_i[16] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n870_1) );
  OR2X2 OR2X2_2538 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_0__17_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n872_1) );
  OR2X2 OR2X2_2539 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf0), .B(\wb_dat_i[17] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n873_1) );
  OR2X2 OR2X2_254 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n537), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n538), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n539) );
  OR2X2 OR2X2_2540 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_0__18_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n875_1) );
  OR2X2 OR2X2_2541 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf5), .B(\wb_dat_i[18] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n876_1) );
  OR2X2 OR2X2_2542 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_0__19_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n878_1) );
  OR2X2 OR2X2_2543 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf4), .B(\wb_dat_i[19] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n879_1) );
  OR2X2 OR2X2_2544 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_0__20_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n881_1) );
  OR2X2 OR2X2_2545 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf3), .B(\wb_dat_i[20] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n882_1) );
  OR2X2 OR2X2_2546 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_0__21_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n884_1) );
  OR2X2 OR2X2_2547 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf2), .B(\wb_dat_i[21] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n885_1) );
  OR2X2 OR2X2_2548 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_0__22_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n887_1) );
  OR2X2 OR2X2_2549 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf1), .B(\wb_dat_i[22] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n888_1) );
  OR2X2 OR2X2_255 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n541), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n542), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n543) );
  OR2X2 OR2X2_2550 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_0__23_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n890_1) );
  OR2X2 OR2X2_2551 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf0), .B(\wb_dat_i[23] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n891_1) );
  OR2X2 OR2X2_2552 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_0__24_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n893_1) );
  OR2X2 OR2X2_2553 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf5), .B(\wb_dat_i[24] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n894_1) );
  OR2X2 OR2X2_2554 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_0__25_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n896_1) );
  OR2X2 OR2X2_2555 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf4), .B(\wb_dat_i[25] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n897_1) );
  OR2X2 OR2X2_2556 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_0__26_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n899_1) );
  OR2X2 OR2X2_2557 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf3), .B(\wb_dat_i[26] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n900_1) );
  OR2X2 OR2X2_2558 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_0__27_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n902_1) );
  OR2X2 OR2X2_2559 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf2), .B(\wb_dat_i[27] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n903_1) );
  OR2X2 OR2X2_256 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n545), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n546), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n547) );
  OR2X2 OR2X2_2560 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_0__28_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n905_1) );
  OR2X2 OR2X2_2561 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf1), .B(\wb_dat_i[28] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n906_1) );
  OR2X2 OR2X2_2562 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_0__29_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n908_1) );
  OR2X2 OR2X2_2563 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf0), .B(\wb_dat_i[29] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n909_1) );
  OR2X2 OR2X2_2564 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_0__30_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n911_1) );
  OR2X2 OR2X2_2565 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf5), .B(\wb_dat_i[30] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n912_1) );
  OR2X2 OR2X2_2566 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_0__31_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n914_1) );
  OR2X2 OR2X2_2567 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf4), .B(\wb_dat_i[31] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n915_1) );
  OR2X2 OR2X2_2568 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_0__32_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n917) );
  OR2X2 OR2X2_2569 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_wr_data_32_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n918_1) );
  OR2X2 OR2X2_257 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n549), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n550), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n551) );
  OR2X2 OR2X2_2570 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_0__33_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n920_1) );
  OR2X2 OR2X2_2571 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_wr_data_33_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n921_1) );
  OR2X2 OR2X2_2572 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_0__34_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n923_1) );
  OR2X2 OR2X2_2573 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_wr_data_34_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n924_1) );
  OR2X2 OR2X2_2574 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n819_1_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_0__35_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n926_1) );
  OR2X2 OR2X2_2575 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n821_1_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_wr_data_35_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n927_1) );
  OR2X2 OR2X2_2576 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_4__0_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n931_1) );
  OR2X2 OR2X2_2577 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf5), .B(\wb_dat_i[0] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n933_1) );
  OR2X2 OR2X2_2578 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_4__1_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n935_1) );
  OR2X2 OR2X2_2579 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf4), .B(\wb_dat_i[1] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n936_1) );
  OR2X2 OR2X2_258 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n553), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n554), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n555) );
  OR2X2 OR2X2_2580 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_4__2_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n938_1) );
  OR2X2 OR2X2_2581 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf3), .B(\wb_dat_i[2] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n939_1) );
  OR2X2 OR2X2_2582 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_4__3_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n941_1) );
  OR2X2 OR2X2_2583 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf2), .B(\wb_dat_i[3] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n942_1) );
  OR2X2 OR2X2_2584 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_4__4_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n944_1) );
  OR2X2 OR2X2_2585 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf1), .B(\wb_dat_i[4] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n945_1) );
  OR2X2 OR2X2_2586 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_4__5_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n947_1) );
  OR2X2 OR2X2_2587 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf0), .B(\wb_dat_i[5] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n948_1) );
  OR2X2 OR2X2_2588 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_4__6_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n950_1) );
  OR2X2 OR2X2_2589 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf5), .B(\wb_dat_i[6] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n951_1) );
  OR2X2 OR2X2_259 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n557), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n558), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n559) );
  OR2X2 OR2X2_2590 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_4__7_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n953_1) );
  OR2X2 OR2X2_2591 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf4), .B(\wb_dat_i[7] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n954_1) );
  OR2X2 OR2X2_2592 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_4__8_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n956) );
  OR2X2 OR2X2_2593 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf3), .B(\wb_dat_i[8] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n957_1) );
  OR2X2 OR2X2_2594 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_4__9_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n959) );
  OR2X2 OR2X2_2595 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf2), .B(\wb_dat_i[9] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n960) );
  OR2X2 OR2X2_2596 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_4__10_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n962) );
  OR2X2 OR2X2_2597 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf1), .B(\wb_dat_i[10] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n963) );
  OR2X2 OR2X2_2598 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_4__11_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n965_1) );
  OR2X2 OR2X2_2599 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf0), .B(\wb_dat_i[11] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n966_1) );
  OR2X2 OR2X2_26 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n294_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n239_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n295_1) );
  OR2X2 OR2X2_260 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n561), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n562), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n563) );
  OR2X2 OR2X2_2600 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_4__12_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n968) );
  OR2X2 OR2X2_2601 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf5), .B(\wb_dat_i[12] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n969) );
  OR2X2 OR2X2_2602 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_4__13_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n971_1) );
  OR2X2 OR2X2_2603 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf4), .B(\wb_dat_i[13] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n972) );
  OR2X2 OR2X2_2604 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_4__14_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n974) );
  OR2X2 OR2X2_2605 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf3), .B(\wb_dat_i[14] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n975) );
  OR2X2 OR2X2_2606 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_4__15_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n977_1) );
  OR2X2 OR2X2_2607 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf2), .B(\wb_dat_i[15] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n978_1) );
  OR2X2 OR2X2_2608 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_4__16_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n980) );
  OR2X2 OR2X2_2609 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf1), .B(\wb_dat_i[16] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n981) );
  OR2X2 OR2X2_261 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n565), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n566), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n567) );
  OR2X2 OR2X2_2610 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_4__17_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n983) );
  OR2X2 OR2X2_2611 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf0), .B(\wb_dat_i[17] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n984_1) );
  OR2X2 OR2X2_2612 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_4__18_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n986) );
  OR2X2 OR2X2_2613 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf5), .B(\wb_dat_i[18] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n987) );
  OR2X2 OR2X2_2614 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_4__19_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n989_1) );
  OR2X2 OR2X2_2615 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf4), .B(\wb_dat_i[19] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n990) );
  OR2X2 OR2X2_2616 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_4__20_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n992) );
  OR2X2 OR2X2_2617 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf3), .B(\wb_dat_i[20] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n993_1) );
  OR2X2 OR2X2_2618 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_4__21_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n995) );
  OR2X2 OR2X2_2619 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf2), .B(\wb_dat_i[21] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n996) );
  OR2X2 OR2X2_262 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n569), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n570), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n571) );
  OR2X2 OR2X2_2620 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_4__22_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n998_1) );
  OR2X2 OR2X2_2621 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf1), .B(\wb_dat_i[22] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n999_1) );
  OR2X2 OR2X2_2622 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_4__23_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1001) );
  OR2X2 OR2X2_2623 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf0), .B(\wb_dat_i[23] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1002) );
  OR2X2 OR2X2_2624 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_4__24_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1004) );
  OR2X2 OR2X2_2625 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf5), .B(\wb_dat_i[24] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1005_1) );
  OR2X2 OR2X2_2626 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_4__25_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1007) );
  OR2X2 OR2X2_2627 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf4), .B(\wb_dat_i[25] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1008) );
  OR2X2 OR2X2_2628 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_4__26_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1010) );
  OR2X2 OR2X2_2629 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf3), .B(\wb_dat_i[26] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1011_1) );
  OR2X2 OR2X2_263 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n573), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n574), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n575) );
  OR2X2 OR2X2_2630 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_4__27_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1013_1) );
  OR2X2 OR2X2_2631 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf2), .B(\wb_dat_i[27] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1014) );
  OR2X2 OR2X2_2632 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_4__28_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1016) );
  OR2X2 OR2X2_2633 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf1), .B(\wb_dat_i[28] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1017) );
  OR2X2 OR2X2_2634 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_4__29_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1019) );
  OR2X2 OR2X2_2635 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf0), .B(\wb_dat_i[29] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1020) );
  OR2X2 OR2X2_2636 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_4__30_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1022_1) );
  OR2X2 OR2X2_2637 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf5), .B(\wb_dat_i[30] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1023_1) );
  OR2X2 OR2X2_2638 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_4__31_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1025) );
  OR2X2 OR2X2_2639 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf4), .B(\wb_dat_i[31] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1026) );
  OR2X2 OR2X2_264 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n577), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n578), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n579) );
  OR2X2 OR2X2_2640 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_4__32_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1028_1) );
  OR2X2 OR2X2_2641 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_wr_data_32_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1029) );
  OR2X2 OR2X2_2642 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_4__33_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1031_1) );
  OR2X2 OR2X2_2643 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_wr_data_33_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1032) );
  OR2X2 OR2X2_2644 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_4__34_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1034) );
  OR2X2 OR2X2_2645 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_wr_data_34_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1035_1) );
  OR2X2 OR2X2_2646 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n930_1_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_4__35_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1037_1) );
  OR2X2 OR2X2_2647 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n932_1_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_wr_data_35_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1038_1) );
  OR2X2 OR2X2_2648 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_3__0_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1043_1) );
  OR2X2 OR2X2_2649 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf5), .B(\wb_dat_i[0] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1045_1) );
  OR2X2 OR2X2_265 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n581), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n582), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n583) );
  OR2X2 OR2X2_2650 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_3__1_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1047_1) );
  OR2X2 OR2X2_2651 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf4), .B(\wb_dat_i[1] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1048_1) );
  OR2X2 OR2X2_2652 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_3__2_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1050_1) );
  OR2X2 OR2X2_2653 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf3), .B(\wb_dat_i[2] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1051_1) );
  OR2X2 OR2X2_2654 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_3__3_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1053_1) );
  OR2X2 OR2X2_2655 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf2), .B(\wb_dat_i[3] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1054_1) );
  OR2X2 OR2X2_2656 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_3__4_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1056_1) );
  OR2X2 OR2X2_2657 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf1), .B(\wb_dat_i[4] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1057_1) );
  OR2X2 OR2X2_2658 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_3__5_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1059_1) );
  OR2X2 OR2X2_2659 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf0), .B(\wb_dat_i[5] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1060_1) );
  OR2X2 OR2X2_266 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n585), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n586), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n587) );
  OR2X2 OR2X2_2660 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_3__6_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1062_1) );
  OR2X2 OR2X2_2661 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf5), .B(\wb_dat_i[6] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1063_1) );
  OR2X2 OR2X2_2662 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_3__7_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1065_1) );
  OR2X2 OR2X2_2663 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf4), .B(\wb_dat_i[7] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1066_1) );
  OR2X2 OR2X2_2664 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_3__8_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1068_1) );
  OR2X2 OR2X2_2665 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf3), .B(\wb_dat_i[8] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1069_1) );
  OR2X2 OR2X2_2666 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_3__9_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1071) );
  OR2X2 OR2X2_2667 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf2), .B(\wb_dat_i[9] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1072) );
  OR2X2 OR2X2_2668 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_3__10_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1074) );
  OR2X2 OR2X2_2669 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf1), .B(\wb_dat_i[10] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1075) );
  OR2X2 OR2X2_267 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n589), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n590), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n591) );
  OR2X2 OR2X2_2670 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_3__11_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1077) );
  OR2X2 OR2X2_2671 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf0), .B(\wb_dat_i[11] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1078) );
  OR2X2 OR2X2_2672 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_3__12_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1080) );
  OR2X2 OR2X2_2673 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf5), .B(\wb_dat_i[12] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1081) );
  OR2X2 OR2X2_2674 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_3__13_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1083) );
  OR2X2 OR2X2_2675 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf4), .B(\wb_dat_i[13] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1084) );
  OR2X2 OR2X2_2676 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_3__14_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1086) );
  OR2X2 OR2X2_2677 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf3), .B(\wb_dat_i[14] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1087) );
  OR2X2 OR2X2_2678 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_3__15_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1089) );
  OR2X2 OR2X2_2679 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf2), .B(\wb_dat_i[15] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1090) );
  OR2X2 OR2X2_268 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n593), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n594), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n595) );
  OR2X2 OR2X2_2680 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_3__16_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1092) );
  OR2X2 OR2X2_2681 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf1), .B(\wb_dat_i[16] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1093) );
  OR2X2 OR2X2_2682 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_3__17_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1095) );
  OR2X2 OR2X2_2683 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf0), .B(\wb_dat_i[17] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1096) );
  OR2X2 OR2X2_2684 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_3__18_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1098) );
  OR2X2 OR2X2_2685 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf5), .B(\wb_dat_i[18] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1099) );
  OR2X2 OR2X2_2686 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_3__19_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1101) );
  OR2X2 OR2X2_2687 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf4), .B(\wb_dat_i[19] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1102) );
  OR2X2 OR2X2_2688 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_3__20_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1104) );
  OR2X2 OR2X2_2689 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf3), .B(\wb_dat_i[20] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1105) );
  OR2X2 OR2X2_269 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n597), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n598), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n599) );
  OR2X2 OR2X2_2690 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_3__21_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1107) );
  OR2X2 OR2X2_2691 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf2), .B(\wb_dat_i[21] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1108) );
  OR2X2 OR2X2_2692 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_3__22_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1110) );
  OR2X2 OR2X2_2693 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf1), .B(\wb_dat_i[22] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1111) );
  OR2X2 OR2X2_2694 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_3__23_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1113) );
  OR2X2 OR2X2_2695 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf0), .B(\wb_dat_i[23] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1114) );
  OR2X2 OR2X2_2696 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_3__24_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1116) );
  OR2X2 OR2X2_2697 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf5), .B(\wb_dat_i[24] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1117) );
  OR2X2 OR2X2_2698 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_3__25_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1119) );
  OR2X2 OR2X2_2699 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf4), .B(\wb_dat_i[25] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1120) );
  OR2X2 OR2X2_27 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n295_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n281_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n296_1) );
  OR2X2 OR2X2_270 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n601), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n602), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n603) );
  OR2X2 OR2X2_2700 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_3__26_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1122) );
  OR2X2 OR2X2_2701 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf3), .B(\wb_dat_i[26] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1123) );
  OR2X2 OR2X2_2702 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_3__27_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1125) );
  OR2X2 OR2X2_2703 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf2), .B(\wb_dat_i[27] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1126) );
  OR2X2 OR2X2_2704 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_3__28_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1128) );
  OR2X2 OR2X2_2705 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf1), .B(\wb_dat_i[28] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1129) );
  OR2X2 OR2X2_2706 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_3__29_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1131) );
  OR2X2 OR2X2_2707 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf0), .B(\wb_dat_i[29] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1132) );
  OR2X2 OR2X2_2708 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_3__30_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1134) );
  OR2X2 OR2X2_2709 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf5), .B(\wb_dat_i[30] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1135) );
  OR2X2 OR2X2_271 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n368_1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n367), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n606) );
  OR2X2 OR2X2_2710 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_3__31_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1137) );
  OR2X2 OR2X2_2711 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf4), .B(\wb_dat_i[31] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1138) );
  OR2X2 OR2X2_2712 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_3__32_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1140) );
  OR2X2 OR2X2_2713 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_wr_data_32_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1141) );
  OR2X2 OR2X2_2714 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_3__33_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1143) );
  OR2X2 OR2X2_2715 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_wr_data_33_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1144) );
  OR2X2 OR2X2_2716 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_3__34_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1146) );
  OR2X2 OR2X2_2717 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_wr_data_34_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1147) );
  OR2X2 OR2X2_2718 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1042_1_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_3__35_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1149) );
  OR2X2 OR2X2_2719 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1044_1_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_wr_data_35_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1150) );
  OR2X2 OR2X2_272 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n607), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n605), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_0_) );
  OR2X2 OR2X2_2720 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1153), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1152), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1154) );
  OR2X2 OR2X2_2721 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1159), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf4), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1160) );
  OR2X2 OR2X2_2722 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1160), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1157), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1161) );
  OR2X2 OR2X2_2723 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1161), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1155), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1162) );
  OR2X2 OR2X2_2724 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1164), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1163), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1165) );
  OR2X2 OR2X2_2725 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1168), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf5), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1169) );
  OR2X2 OR2X2_2726 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1169), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1167), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1170) );
  OR2X2 OR2X2_2727 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1170), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1166), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1171) );
  OR2X2 OR2X2_2728 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1174), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1173), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1175) );
  OR2X2 OR2X2_2729 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1178), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf4), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1179) );
  OR2X2 OR2X2_273 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_0_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n609) );
  OR2X2 OR2X2_2730 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1179), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1177), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1180) );
  OR2X2 OR2X2_2731 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1180), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1176), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1181) );
  OR2X2 OR2X2_2732 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1183), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1182), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1184) );
  OR2X2 OR2X2_2733 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1187), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf3), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1188) );
  OR2X2 OR2X2_2734 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1188), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1186), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1189) );
  OR2X2 OR2X2_2735 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1189), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1185), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1190) );
  OR2X2 OR2X2_2736 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1193), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1192), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1194) );
  OR2X2 OR2X2_2737 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1197), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf2), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1198) );
  OR2X2 OR2X2_2738 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1198), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1196), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1199) );
  OR2X2 OR2X2_2739 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1199), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1195), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1200) );
  OR2X2 OR2X2_274 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_0_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_2_bF_buf3), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n610) );
  OR2X2 OR2X2_2740 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1202), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1201), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1203) );
  OR2X2 OR2X2_2741 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1206), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf3), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1207) );
  OR2X2 OR2X2_2742 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1207), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1205), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1208) );
  OR2X2 OR2X2_2743 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1208), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1204), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1209) );
  OR2X2 OR2X2_2744 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1212), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1211), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1213) );
  OR2X2 OR2X2_2745 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1216), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf2), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1217) );
  OR2X2 OR2X2_2746 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1217), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1215), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1218) );
  OR2X2 OR2X2_2747 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1218), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1214), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1219) );
  OR2X2 OR2X2_2748 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1221), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1220), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1222) );
  OR2X2 OR2X2_2749 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1225), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1226) );
  OR2X2 OR2X2_275 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n613), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n612), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_1_) );
  OR2X2 OR2X2_2750 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1226), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1224), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1227) );
  OR2X2 OR2X2_2751 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1227), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1223), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1228) );
  OR2X2 OR2X2_2752 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1231), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1230), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1232) );
  OR2X2 OR2X2_2753 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1235), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1236) );
  OR2X2 OR2X2_2754 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1236), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1234), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1237) );
  OR2X2 OR2X2_2755 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1237), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1233), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1238) );
  OR2X2 OR2X2_2756 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1240), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1239), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1241) );
  OR2X2 OR2X2_2757 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1244), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf0), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1245) );
  OR2X2 OR2X2_2758 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1245), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1243), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1246) );
  OR2X2 OR2X2_2759 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1246), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1242), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1247) );
  OR2X2 OR2X2_276 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_1_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n615) );
  OR2X2 OR2X2_2760 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1250), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1249), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1251) );
  OR2X2 OR2X2_2761 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1254), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf0), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1255) );
  OR2X2 OR2X2_2762 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1255), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1253), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1256) );
  OR2X2 OR2X2_2763 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1256), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1252), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1257) );
  OR2X2 OR2X2_2764 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1259), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1258), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1260) );
  OR2X2 OR2X2_2765 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1263), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf5), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1264) );
  OR2X2 OR2X2_2766 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1264), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1262), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1265) );
  OR2X2 OR2X2_2767 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1265), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1261), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1266) );
  OR2X2 OR2X2_2768 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1269), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1268), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1270) );
  OR2X2 OR2X2_2769 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1273), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf5), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1274) );
  OR2X2 OR2X2_277 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_1_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_2_bF_buf2), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n616) );
  OR2X2 OR2X2_2770 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1274), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1272), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1275) );
  OR2X2 OR2X2_2771 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1275), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1271), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1276) );
  OR2X2 OR2X2_2772 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1278), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1277), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1279) );
  OR2X2 OR2X2_2773 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1282), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf4), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1283) );
  OR2X2 OR2X2_2774 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1283), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1281), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1284) );
  OR2X2 OR2X2_2775 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1284), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1280), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1285) );
  OR2X2 OR2X2_2776 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1288), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1287), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1289) );
  OR2X2 OR2X2_2777 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1292), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf4), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1293) );
  OR2X2 OR2X2_2778 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1293), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1291), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1294) );
  OR2X2 OR2X2_2779 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1294), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1290), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1295) );
  OR2X2 OR2X2_278 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n619), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n618), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_2_) );
  OR2X2 OR2X2_2780 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1297), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1296), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1298) );
  OR2X2 OR2X2_2781 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1301), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf3), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1302) );
  OR2X2 OR2X2_2782 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1302), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1300), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1303) );
  OR2X2 OR2X2_2783 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1303), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1299), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1304) );
  OR2X2 OR2X2_2784 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1307), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1306), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1308) );
  OR2X2 OR2X2_2785 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1311), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf2), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1312) );
  OR2X2 OR2X2_2786 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1312), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1310), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1313) );
  OR2X2 OR2X2_2787 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1313), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1309), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1314) );
  OR2X2 OR2X2_2788 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1316), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1315), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1317) );
  OR2X2 OR2X2_2789 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1320), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf3), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1321) );
  OR2X2 OR2X2_279 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_2_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n621) );
  OR2X2 OR2X2_2790 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1321), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1319), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1322) );
  OR2X2 OR2X2_2791 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1322), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1318), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1323) );
  OR2X2 OR2X2_2792 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1326), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1325), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1327) );
  OR2X2 OR2X2_2793 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1330), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1331) );
  OR2X2 OR2X2_2794 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1331), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1329), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1332) );
  OR2X2 OR2X2_2795 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1332), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1328), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1333) );
  OR2X2 OR2X2_2796 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1335), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1334), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1336) );
  OR2X2 OR2X2_2797 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1339), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf2), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1340) );
  OR2X2 OR2X2_2798 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1340), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1338), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1341) );
  OR2X2 OR2X2_2799 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1341), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1337), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1342) );
  OR2X2 OR2X2_28 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n298_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n299_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n300) );
  OR2X2 OR2X2_280 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_2_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_2_bF_buf1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n622) );
  OR2X2 OR2X2_2800 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1345), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1344), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1346) );
  OR2X2 OR2X2_2801 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1349), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1350) );
  OR2X2 OR2X2_2802 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1350), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1348), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1351) );
  OR2X2 OR2X2_2803 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1351), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1347), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1352) );
  OR2X2 OR2X2_2804 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1354), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1353), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1355) );
  OR2X2 OR2X2_2805 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1358), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf0), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1359) );
  OR2X2 OR2X2_2806 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1359), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1357), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1360) );
  OR2X2 OR2X2_2807 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1360), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1356), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1361) );
  OR2X2 OR2X2_2808 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1364), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1363), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1365) );
  OR2X2 OR2X2_2809 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1367), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf0), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1368) );
  OR2X2 OR2X2_281 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n625), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n624), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_3_) );
  OR2X2 OR2X2_2810 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1368), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1369), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1370) );
  OR2X2 OR2X2_2811 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1370), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1366), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1371) );
  OR2X2 OR2X2_2812 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1373), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1372), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1374) );
  OR2X2 OR2X2_2813 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1377), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf5), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1378) );
  OR2X2 OR2X2_2814 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1378), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1376), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1379) );
  OR2X2 OR2X2_2815 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1379), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1375), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1380) );
  OR2X2 OR2X2_2816 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1383), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1382), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1384) );
  OR2X2 OR2X2_2817 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1387), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf4), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1388) );
  OR2X2 OR2X2_2818 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1388), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1386), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1389) );
  OR2X2 OR2X2_2819 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1389), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1385), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1390) );
  OR2X2 OR2X2_282 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_3_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n627) );
  OR2X2 OR2X2_2820 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1392), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1391), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1393) );
  OR2X2 OR2X2_2821 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1396), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf5), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1397) );
  OR2X2 OR2X2_2822 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1397), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1395), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1398) );
  OR2X2 OR2X2_2823 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1398), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1394), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1399) );
  OR2X2 OR2X2_2824 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1402), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1401), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1403) );
  OR2X2 OR2X2_2825 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1406), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf4), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1407) );
  OR2X2 OR2X2_2826 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1407), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1405), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1408) );
  OR2X2 OR2X2_2827 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1408), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1404), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1409) );
  OR2X2 OR2X2_2828 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1411), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1410), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1412) );
  OR2X2 OR2X2_2829 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1415), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf3), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1416) );
  OR2X2 OR2X2_283 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_3_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_2_bF_buf0), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n628) );
  OR2X2 OR2X2_2830 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1416), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1414), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1417) );
  OR2X2 OR2X2_2831 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1417), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1413), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1418) );
  OR2X2 OR2X2_2832 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1421), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1420), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1422) );
  OR2X2 OR2X2_2833 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1425), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf3), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1426) );
  OR2X2 OR2X2_2834 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1426), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1424), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1427) );
  OR2X2 OR2X2_2835 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1427), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1423), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1428) );
  OR2X2 OR2X2_2836 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1430), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1429), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1431) );
  OR2X2 OR2X2_2837 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1434), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf2), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1435) );
  OR2X2 OR2X2_2838 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1435), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1433), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1436) );
  OR2X2 OR2X2_2839 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1436), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1432), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1437) );
  OR2X2 OR2X2_284 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n631), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n630), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_4_) );
  OR2X2 OR2X2_2840 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1440), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1439), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1441) );
  OR2X2 OR2X2_2841 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1444), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1445) );
  OR2X2 OR2X2_2842 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1445), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1443), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1446) );
  OR2X2 OR2X2_2843 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1446), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1442), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1447) );
  OR2X2 OR2X2_2844 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1449), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1448), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1450) );
  OR2X2 OR2X2_2845 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1453), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf2), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1454) );
  OR2X2 OR2X2_2846 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1454), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1452), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1455) );
  OR2X2 OR2X2_2847 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1455), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1451), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1456) );
  OR2X2 OR2X2_2848 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1459), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1458), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1460) );
  OR2X2 OR2X2_2849 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1463), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf0), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1464) );
  OR2X2 OR2X2_285 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_4_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n633) );
  OR2X2 OR2X2_2850 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1464), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1462), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1465) );
  OR2X2 OR2X2_2851 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1465), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1461), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1466) );
  OR2X2 OR2X2_2852 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1468), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1467), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1469) );
  OR2X2 OR2X2_2853 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1472), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1473) );
  OR2X2 OR2X2_2854 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1473), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1471), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1474) );
  OR2X2 OR2X2_2855 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1474), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1470), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1475) );
  OR2X2 OR2X2_2856 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1478), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1477), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1479) );
  OR2X2 OR2X2_2857 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1482), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf0), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1483) );
  OR2X2 OR2X2_2858 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1483), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1481), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1484) );
  OR2X2 OR2X2_2859 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1484), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1480), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1485) );
  OR2X2 OR2X2_286 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_4_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_2_bF_buf3), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n634) );
  OR2X2 OR2X2_2860 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1487), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1486), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1488) );
  OR2X2 OR2X2_2861 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1491), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf5), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1492) );
  OR2X2 OR2X2_2862 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1492), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1490), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1493) );
  OR2X2 OR2X2_2863 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1493), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1489), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1494) );
  OR2X2 OR2X2_2864 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1497), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1496), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1498) );
  OR2X2 OR2X2_2865 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1501), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf4), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1502) );
  OR2X2 OR2X2_2866 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1502), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1500), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1503) );
  OR2X2 OR2X2_2867 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1503), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1499), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1504) );
  OR2X2 OR2X2_2868 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1506), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1505), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1507) );
  OR2X2 OR2X2_2869 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1510), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf5), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1511) );
  OR2X2 OR2X2_287 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n637), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n636), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_5_) );
  OR2X2 OR2X2_2870 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1511), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1509), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1512) );
  OR2X2 OR2X2_2871 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1512), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1508), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1513) );
  OR2X2 OR2X2_2872 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1516), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1515), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1517) );
  OR2X2 OR2X2_2873 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1520), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf3), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1521) );
  OR2X2 OR2X2_2874 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1521), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1519), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1522) );
  OR2X2 OR2X2_2875 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1522), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1518), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1523) );
  OR2X2 OR2X2_2876 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1525), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1524), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1526) );
  OR2X2 OR2X2_2877 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1529), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf4), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1530) );
  OR2X2 OR2X2_2878 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1530), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1528), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1531) );
  OR2X2 OR2X2_2879 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1531), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1527), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1532) );
  OR2X2 OR2X2_288 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_5_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n639) );
  OR2X2 OR2X2_2880 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1535), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1534), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1536) );
  OR2X2 OR2X2_2881 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1539), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf3), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1540) );
  OR2X2 OR2X2_2882 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1540), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1538), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1541) );
  OR2X2 OR2X2_2883 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1541), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1537), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1542) );
  OR2X2 OR2X2_2884 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1544), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1543), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1545) );
  OR2X2 OR2X2_2885 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1548), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf2), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1549) );
  OR2X2 OR2X2_2886 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1549), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1547), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1550) );
  OR2X2 OR2X2_2887 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1550), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1546), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1551) );
  OR2X2 OR2X2_2888 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1554), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1553), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1555) );
  OR2X2 OR2X2_2889 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1558), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1559) );
  OR2X2 OR2X2_289 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_5_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_2_bF_buf2), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n640) );
  OR2X2 OR2X2_2890 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1559), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1557), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1560) );
  OR2X2 OR2X2_2891 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1560), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1556), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1561) );
  OR2X2 OR2X2_2892 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1563), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1562), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1564) );
  OR2X2 OR2X2_2893 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1567), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf2), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1568) );
  OR2X2 OR2X2_2894 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1568), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1566), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1569) );
  OR2X2 OR2X2_2895 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1569), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1565), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1570) );
  OR2X2 OR2X2_2896 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1573), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1572), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1574) );
  OR2X2 OR2X2_2897 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1576), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf0), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1577) );
  OR2X2 OR2X2_2898 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1577), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1578), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1579) );
  OR2X2 OR2X2_2899 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1579), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1575), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1580) );
  OR2X2 OR2X2_29 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n303_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n278), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n304) );
  OR2X2 OR2X2_290 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n643), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n642), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_6_) );
  OR2X2 OR2X2_2900 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1582), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1581), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1583) );
  OR2X2 OR2X2_2901 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1586), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1587) );
  OR2X2 OR2X2_2902 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1587), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1585), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1588) );
  OR2X2 OR2X2_2903 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1588), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1584), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1589) );
  OR2X2 OR2X2_2904 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1592), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1591), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1593) );
  OR2X2 OR2X2_2905 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1596), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf0), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1597) );
  OR2X2 OR2X2_2906 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1597), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1595), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1598) );
  OR2X2 OR2X2_2907 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1598), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1594), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1599) );
  OR2X2 OR2X2_2908 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1601), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1600), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1602) );
  OR2X2 OR2X2_2909 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1605), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf5), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1606) );
  OR2X2 OR2X2_291 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_6_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n645) );
  OR2X2 OR2X2_2910 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1606), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1604), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1607) );
  OR2X2 OR2X2_2911 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1607), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1603), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1608) );
  OR2X2 OR2X2_2912 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1611), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1610), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1612) );
  OR2X2 OR2X2_2913 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1615), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf4), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1616) );
  OR2X2 OR2X2_2914 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1616), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1614), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1617) );
  OR2X2 OR2X2_2915 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1617), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1613), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1618) );
  OR2X2 OR2X2_2916 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1620), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1619), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1621) );
  OR2X2 OR2X2_2917 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1624), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf5), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1625) );
  OR2X2 OR2X2_2918 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1625), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1623), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1626) );
  OR2X2 OR2X2_2919 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1626), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1622), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1627) );
  OR2X2 OR2X2_292 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_6_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_2_bF_buf1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n646) );
  OR2X2 OR2X2_2920 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1630), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1629), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1631) );
  OR2X2 OR2X2_2921 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1634), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf4), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1635) );
  OR2X2 OR2X2_2922 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1635), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1633), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1636) );
  OR2X2 OR2X2_2923 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1636), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1632), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1637) );
  OR2X2 OR2X2_2924 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1639), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1638), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1640) );
  OR2X2 OR2X2_2925 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1643), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf3), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1644) );
  OR2X2 OR2X2_2926 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1644), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1642), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1645) );
  OR2X2 OR2X2_2927 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1645), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1641), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1646) );
  OR2X2 OR2X2_2928 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1649), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1648), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1650) );
  OR2X2 OR2X2_2929 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1653), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf3), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1654) );
  OR2X2 OR2X2_293 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n649), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n648), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_7_) );
  OR2X2 OR2X2_2930 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1654), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1652), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1655) );
  OR2X2 OR2X2_2931 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1655), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1651), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1656) );
  OR2X2 OR2X2_2932 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1658), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1657), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1659) );
  OR2X2 OR2X2_2933 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1662), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf2), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1663) );
  OR2X2 OR2X2_2934 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1663), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1661), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1664) );
  OR2X2 OR2X2_2935 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1664), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1660), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1665) );
  OR2X2 OR2X2_2936 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1668), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1667), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1669) );
  OR2X2 OR2X2_2937 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1672), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1673) );
  OR2X2 OR2X2_2938 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1673), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1671), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1674) );
  OR2X2 OR2X2_2939 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1674), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1670), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1675) );
  OR2X2 OR2X2_294 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_7_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n651) );
  OR2X2 OR2X2_2940 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1677), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1676), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1678) );
  OR2X2 OR2X2_2941 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1681), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf2), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1682) );
  OR2X2 OR2X2_2942 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1682), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1680), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1683) );
  OR2X2 OR2X2_2943 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1683), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1679), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1684) );
  OR2X2 OR2X2_2944 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1687), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1686), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1688) );
  OR2X2 OR2X2_2945 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1690), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf0), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1691) );
  OR2X2 OR2X2_2946 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1691), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1692), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1693) );
  OR2X2 OR2X2_2947 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1693), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1689), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1694) );
  OR2X2 OR2X2_2948 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1696), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1695), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1697) );
  OR2X2 OR2X2_2949 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1700), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1701) );
  OR2X2 OR2X2_295 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_7_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_2_bF_buf0), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n652) );
  OR2X2 OR2X2_2950 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1701), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1699), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1702) );
  OR2X2 OR2X2_2951 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1702), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1698), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1703) );
  OR2X2 OR2X2_2952 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1706), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1705), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1707) );
  OR2X2 OR2X2_2953 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1709), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf0), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1710) );
  OR2X2 OR2X2_2954 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1710), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1711), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1712) );
  OR2X2 OR2X2_2955 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1712), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1708), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1713) );
  OR2X2 OR2X2_2956 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1715), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1714), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1716) );
  OR2X2 OR2X2_2957 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1719), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf5), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1720) );
  OR2X2 OR2X2_2958 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1720), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1718), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1721) );
  OR2X2 OR2X2_2959 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1721), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1717), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1722) );
  OR2X2 OR2X2_296 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n655), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n654), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_8_) );
  OR2X2 OR2X2_2960 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1725), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1724), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1726) );
  OR2X2 OR2X2_2961 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1729), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf5), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1730) );
  OR2X2 OR2X2_2962 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1730), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1728), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1731) );
  OR2X2 OR2X2_2963 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1731), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1727), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1732) );
  OR2X2 OR2X2_2964 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1734), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1733), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1735) );
  OR2X2 OR2X2_2965 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1738), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf4), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1739) );
  OR2X2 OR2X2_2966 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1739), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1737), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1740) );
  OR2X2 OR2X2_2967 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1740), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1736), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1741) );
  OR2X2 OR2X2_2968 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1744), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1743), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1745) );
  OR2X2 OR2X2_2969 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1748), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf3), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1749) );
  OR2X2 OR2X2_297 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_8_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n657) );
  OR2X2 OR2X2_2970 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1749), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1747), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1750) );
  OR2X2 OR2X2_2971 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1750), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1746), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1751) );
  OR2X2 OR2X2_2972 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1753), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1752), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1754) );
  OR2X2 OR2X2_2973 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1757), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf4), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1758) );
  OR2X2 OR2X2_2974 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1758), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1756), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1759) );
  OR2X2 OR2X2_2975 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1759), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1755), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1760) );
  OR2X2 OR2X2_2976 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1763), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1762), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1764) );
  OR2X2 OR2X2_2977 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1767), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf3), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1768) );
  OR2X2 OR2X2_2978 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1768), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1766), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1769) );
  OR2X2 OR2X2_2979 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1769), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1765), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1770) );
  OR2X2 OR2X2_298 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_8_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_2_bF_buf3), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n658) );
  OR2X2 OR2X2_2980 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1772), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1771), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1773) );
  OR2X2 OR2X2_2981 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1776), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf2), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1777) );
  OR2X2 OR2X2_2982 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1777), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1775), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1778) );
  OR2X2 OR2X2_2983 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1778), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1774), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1779) );
  OR2X2 OR2X2_2984 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1782), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1781), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1783) );
  OR2X2 OR2X2_2985 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1786), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf2), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1787) );
  OR2X2 OR2X2_2986 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1787), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1785), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1788) );
  OR2X2 OR2X2_2987 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1788), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1784), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1789) );
  OR2X2 OR2X2_2988 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1791), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1790), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1792) );
  OR2X2 OR2X2_2989 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1795), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1796) );
  OR2X2 OR2X2_299 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n661), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n660), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_9_) );
  OR2X2 OR2X2_2990 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1796), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1794), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1797) );
  OR2X2 OR2X2_2991 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1797), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1793), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1798) );
  OR2X2 OR2X2_2992 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1801), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1800), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1802) );
  OR2X2 OR2X2_2993 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1805), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf0), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1806) );
  OR2X2 OR2X2_2994 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1806), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1804), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1807) );
  OR2X2 OR2X2_2995 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1807), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1803), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1808) );
  OR2X2 OR2X2_2996 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1810), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1809), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1811) );
  OR2X2 OR2X2_2997 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1814), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf1), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1815) );
  OR2X2 OR2X2_2998 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1815), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1813), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1816) );
  OR2X2 OR2X2_2999 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1816), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1812), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1817) );
  OR2X2 OR2X2_3 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n207_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n208), .Y(u_sdrc_core_b2r_ack) );
  OR2X2 OR2X2_30 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n301_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n305_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n306_1) );
  OR2X2 OR2X2_300 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_9_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n663) );
  OR2X2 OR2X2_3000 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1820), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1819), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1821) );
  OR2X2 OR2X2_3001 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1824), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf5), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1825) );
  OR2X2 OR2X2_3002 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1825), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1823), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1826) );
  OR2X2 OR2X2_3003 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1826), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1822), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1827) );
  OR2X2 OR2X2_3004 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1829), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1828), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1830) );
  OR2X2 OR2X2_3005 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1832), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n795_1_bF_buf0), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1833) );
  OR2X2 OR2X2_3006 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1833), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1834), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1835) );
  OR2X2 OR2X2_3007 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1835), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1831), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1836) );
  OR2X2 OR2X2_3008 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_6__0_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1840) );
  OR2X2 OR2X2_3009 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf5), .B(\wb_dat_i[0] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1842) );
  OR2X2 OR2X2_301 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_9_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_2_bF_buf2), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n664) );
  OR2X2 OR2X2_3010 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_6__1_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1844) );
  OR2X2 OR2X2_3011 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf4), .B(\wb_dat_i[1] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1845) );
  OR2X2 OR2X2_3012 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_6__2_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1847) );
  OR2X2 OR2X2_3013 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf3), .B(\wb_dat_i[2] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1848) );
  OR2X2 OR2X2_3014 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_6__3_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1850) );
  OR2X2 OR2X2_3015 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf2), .B(\wb_dat_i[3] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1851) );
  OR2X2 OR2X2_3016 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_6__4_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1853) );
  OR2X2 OR2X2_3017 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf1), .B(\wb_dat_i[4] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1854) );
  OR2X2 OR2X2_3018 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_6__5_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1856) );
  OR2X2 OR2X2_3019 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf0), .B(\wb_dat_i[5] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1857) );
  OR2X2 OR2X2_302 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n667), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n666), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_10_) );
  OR2X2 OR2X2_3020 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_6__6_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1859) );
  OR2X2 OR2X2_3021 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf5), .B(\wb_dat_i[6] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1860) );
  OR2X2 OR2X2_3022 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_6__7_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1862) );
  OR2X2 OR2X2_3023 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf4), .B(\wb_dat_i[7] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1863) );
  OR2X2 OR2X2_3024 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_6__8_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1865) );
  OR2X2 OR2X2_3025 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf3), .B(\wb_dat_i[8] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1866) );
  OR2X2 OR2X2_3026 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_6__9_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1868) );
  OR2X2 OR2X2_3027 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf2), .B(\wb_dat_i[9] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1869) );
  OR2X2 OR2X2_3028 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_6__10_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1871) );
  OR2X2 OR2X2_3029 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf1), .B(\wb_dat_i[10] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1872) );
  OR2X2 OR2X2_303 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_10_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n669) );
  OR2X2 OR2X2_3030 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_6__11_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1874) );
  OR2X2 OR2X2_3031 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf0), .B(\wb_dat_i[11] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1875) );
  OR2X2 OR2X2_3032 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_6__12_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1877) );
  OR2X2 OR2X2_3033 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf5), .B(\wb_dat_i[12] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1878) );
  OR2X2 OR2X2_3034 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_6__13_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1880) );
  OR2X2 OR2X2_3035 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf4), .B(\wb_dat_i[13] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1881) );
  OR2X2 OR2X2_3036 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_6__14_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1883) );
  OR2X2 OR2X2_3037 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf3), .B(\wb_dat_i[14] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1884) );
  OR2X2 OR2X2_3038 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_6__15_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1886) );
  OR2X2 OR2X2_3039 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf2), .B(\wb_dat_i[15] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1887) );
  OR2X2 OR2X2_304 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_10_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_2_bF_buf1), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n670) );
  OR2X2 OR2X2_3040 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_6__16_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1889) );
  OR2X2 OR2X2_3041 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf1), .B(\wb_dat_i[16] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1890) );
  OR2X2 OR2X2_3042 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_6__17_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1892) );
  OR2X2 OR2X2_3043 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf0), .B(\wb_dat_i[17] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1893) );
  OR2X2 OR2X2_3044 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_6__18_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1895) );
  OR2X2 OR2X2_3045 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf5), .B(\wb_dat_i[18] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1896) );
  OR2X2 OR2X2_3046 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_6__19_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1898) );
  OR2X2 OR2X2_3047 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf4), .B(\wb_dat_i[19] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1899) );
  OR2X2 OR2X2_3048 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_6__20_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1901) );
  OR2X2 OR2X2_3049 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf3), .B(\wb_dat_i[20] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1902) );
  OR2X2 OR2X2_305 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n673), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n672), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_11_) );
  OR2X2 OR2X2_3050 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_6__21_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1904) );
  OR2X2 OR2X2_3051 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf2), .B(\wb_dat_i[21] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1905) );
  OR2X2 OR2X2_3052 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_6__22_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1907) );
  OR2X2 OR2X2_3053 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf1), .B(\wb_dat_i[22] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1908) );
  OR2X2 OR2X2_3054 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_6__23_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1910) );
  OR2X2 OR2X2_3055 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf0), .B(\wb_dat_i[23] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1911) );
  OR2X2 OR2X2_3056 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_6__24_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1913) );
  OR2X2 OR2X2_3057 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf5), .B(\wb_dat_i[24] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1914) );
  OR2X2 OR2X2_3058 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_6__25_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1916) );
  OR2X2 OR2X2_3059 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf4), .B(\wb_dat_i[25] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1917) );
  OR2X2 OR2X2_306 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_11_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n675) );
  OR2X2 OR2X2_3060 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_6__26_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1919) );
  OR2X2 OR2X2_3061 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf3), .B(\wb_dat_i[26] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1920) );
  OR2X2 OR2X2_3062 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_6__27_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1922) );
  OR2X2 OR2X2_3063 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf2), .B(\wb_dat_i[27] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1923) );
  OR2X2 OR2X2_3064 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_6__28_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1925) );
  OR2X2 OR2X2_3065 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf1), .B(\wb_dat_i[28] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1926) );
  OR2X2 OR2X2_3066 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_6__29_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1928) );
  OR2X2 OR2X2_3067 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf0), .B(\wb_dat_i[29] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1929) );
  OR2X2 OR2X2_3068 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_6__30_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1931) );
  OR2X2 OR2X2_3069 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf5), .B(\wb_dat_i[30] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1932) );
  OR2X2 OR2X2_307 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_11_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_2_bF_buf0), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n676) );
  OR2X2 OR2X2_3070 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_6__31_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1934) );
  OR2X2 OR2X2_3071 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf4), .B(\wb_dat_i[31] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1935) );
  OR2X2 OR2X2_3072 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_6__32_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1937) );
  OR2X2 OR2X2_3073 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_wr_data_32_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1938) );
  OR2X2 OR2X2_3074 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_6__33_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1940) );
  OR2X2 OR2X2_3075 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_wr_data_33_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1941) );
  OR2X2 OR2X2_3076 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_6__34_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1943) );
  OR2X2 OR2X2_3077 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_wr_data_34_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1944) );
  OR2X2 OR2X2_3078 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1839_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_6__35_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1946) );
  OR2X2 OR2X2_3079 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1841_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_wr_data_35_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1947) );
  OR2X2 OR2X2_308 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n679), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n678), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_12_) );
  OR2X2 OR2X2_3080 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_1__0_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1950) );
  OR2X2 OR2X2_3081 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf5), .B(\wb_dat_i[0] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1952) );
  OR2X2 OR2X2_3082 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_1__1_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1954) );
  OR2X2 OR2X2_3083 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf4), .B(\wb_dat_i[1] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1955) );
  OR2X2 OR2X2_3084 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_1__2_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1957) );
  OR2X2 OR2X2_3085 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf3), .B(\wb_dat_i[2] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1958) );
  OR2X2 OR2X2_3086 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_1__3_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1960) );
  OR2X2 OR2X2_3087 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf2), .B(\wb_dat_i[3] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1961) );
  OR2X2 OR2X2_3088 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_1__4_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1963) );
  OR2X2 OR2X2_3089 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf1), .B(\wb_dat_i[4] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1964) );
  OR2X2 OR2X2_309 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_12_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n681) );
  OR2X2 OR2X2_3090 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_1__5_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1966) );
  OR2X2 OR2X2_3091 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf0), .B(\wb_dat_i[5] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1967) );
  OR2X2 OR2X2_3092 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_1__6_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1969) );
  OR2X2 OR2X2_3093 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf5), .B(\wb_dat_i[6] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1970) );
  OR2X2 OR2X2_3094 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_1__7_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1972) );
  OR2X2 OR2X2_3095 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf4), .B(\wb_dat_i[7] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1973) );
  OR2X2 OR2X2_3096 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_1__8_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1975) );
  OR2X2 OR2X2_3097 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf3), .B(\wb_dat_i[8] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1976) );
  OR2X2 OR2X2_3098 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_1__9_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1978) );
  OR2X2 OR2X2_3099 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf2), .B(\wb_dat_i[9] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1979) );
  OR2X2 OR2X2_31 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n308_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n309_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n310) );
  OR2X2 OR2X2_310 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_row_12_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_2_bF_buf3), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n682) );
  OR2X2 OR2X2_3100 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_1__10_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1981) );
  OR2X2 OR2X2_3101 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf1), .B(\wb_dat_i[10] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1982) );
  OR2X2 OR2X2_3102 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_1__11_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1984) );
  OR2X2 OR2X2_3103 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf0), .B(\wb_dat_i[11] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1985) );
  OR2X2 OR2X2_3104 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_1__12_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1987) );
  OR2X2 OR2X2_3105 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf5), .B(\wb_dat_i[12] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1988) );
  OR2X2 OR2X2_3106 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_1__13_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1990) );
  OR2X2 OR2X2_3107 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf4), .B(\wb_dat_i[13] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1991) );
  OR2X2 OR2X2_3108 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_1__14_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1993) );
  OR2X2 OR2X2_3109 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf3), .B(\wb_dat_i[14] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1994) );
  OR2X2 OR2X2_311 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_0_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_last), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n688) );
  OR2X2 OR2X2_3110 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_1__15_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1996) );
  OR2X2 OR2X2_3111 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf2), .B(\wb_dat_i[15] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1997) );
  OR2X2 OR2X2_3112 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_1__16_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n1999) );
  OR2X2 OR2X2_3113 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf1), .B(\wb_dat_i[16] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2000) );
  OR2X2 OR2X2_3114 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_1__17_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2002) );
  OR2X2 OR2X2_3115 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf0), .B(\wb_dat_i[17] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2003) );
  OR2X2 OR2X2_3116 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_1__18_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2005) );
  OR2X2 OR2X2_3117 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf5), .B(\wb_dat_i[18] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2006) );
  OR2X2 OR2X2_3118 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_1__19_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2008) );
  OR2X2 OR2X2_3119 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf4), .B(\wb_dat_i[19] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2009) );
  OR2X2 OR2X2_312 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n685), .B(u_sdrc_core_r2b_last), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n689) );
  OR2X2 OR2X2_3120 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_1__20_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2011) );
  OR2X2 OR2X2_3121 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf3), .B(\wb_dat_i[20] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2012) );
  OR2X2 OR2X2_3122 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_1__21_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2014) );
  OR2X2 OR2X2_3123 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf2), .B(\wb_dat_i[21] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2015) );
  OR2X2 OR2X2_3124 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_1__22_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2017) );
  OR2X2 OR2X2_3125 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf1), .B(\wb_dat_i[22] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2018) );
  OR2X2 OR2X2_3126 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_1__23_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2020) );
  OR2X2 OR2X2_3127 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf0), .B(\wb_dat_i[23] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2021) );
  OR2X2 OR2X2_3128 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_1__24_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2023) );
  OR2X2 OR2X2_3129 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf5), .B(\wb_dat_i[24] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2024) );
  OR2X2 OR2X2_313 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_0_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_0_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n703) );
  OR2X2 OR2X2_3130 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_1__25_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2026) );
  OR2X2 OR2X2_3131 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf4), .B(\wb_dat_i[25] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2027) );
  OR2X2 OR2X2_3132 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_1__26_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2029) );
  OR2X2 OR2X2_3133 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf3), .B(\wb_dat_i[26] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2030) );
  OR2X2 OR2X2_3134 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_1__27_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2032) );
  OR2X2 OR2X2_3135 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf2), .B(\wb_dat_i[27] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2033) );
  OR2X2 OR2X2_3136 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_1__28_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2035) );
  OR2X2 OR2X2_3137 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf1), .B(\wb_dat_i[28] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2036) );
  OR2X2 OR2X2_3138 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_1__29_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2038) );
  OR2X2 OR2X2_3139 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf0), .B(\wb_dat_i[29] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2039) );
  OR2X2 OR2X2_314 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n685), .B(u_sdrc_core_r2b_len_0_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n704) );
  OR2X2 OR2X2_3140 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_1__30_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2041) );
  OR2X2 OR2X2_3141 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf5), .B(\wb_dat_i[30] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2042) );
  OR2X2 OR2X2_3142 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_1__31_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2044) );
  OR2X2 OR2X2_3143 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf4), .B(\wb_dat_i[31] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2045) );
  OR2X2 OR2X2_3144 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_1__32_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2047) );
  OR2X2 OR2X2_3145 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_wr_data_32_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2048) );
  OR2X2 OR2X2_3146 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_1__33_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2050) );
  OR2X2 OR2X2_3147 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_wr_data_33_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2051) );
  OR2X2 OR2X2_3148 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_1__34_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2053) );
  OR2X2 OR2X2_3149 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_wr_data_34_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2054) );
  OR2X2 OR2X2_315 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_0_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_1_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n706) );
  OR2X2 OR2X2_3150 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1949_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_1__35_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2056) );
  OR2X2 OR2X2_3151 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1951_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_wr_data_35_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2057) );
  OR2X2 OR2X2_3152 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_2__0_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2060) );
  OR2X2 OR2X2_3153 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf5), .B(\wb_dat_i[0] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2062) );
  OR2X2 OR2X2_3154 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_2__1_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2064) );
  OR2X2 OR2X2_3155 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf4), .B(\wb_dat_i[1] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2065) );
  OR2X2 OR2X2_3156 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_2__2_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2067) );
  OR2X2 OR2X2_3157 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf3), .B(\wb_dat_i[2] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2068) );
  OR2X2 OR2X2_3158 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_2__3_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2070) );
  OR2X2 OR2X2_3159 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf2), .B(\wb_dat_i[3] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2071) );
  OR2X2 OR2X2_316 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n685), .B(u_sdrc_core_r2b_len_1_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n707) );
  OR2X2 OR2X2_3160 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_2__4_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2073) );
  OR2X2 OR2X2_3161 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf1), .B(\wb_dat_i[4] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2074) );
  OR2X2 OR2X2_3162 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_2__5_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2076) );
  OR2X2 OR2X2_3163 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf0), .B(\wb_dat_i[5] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2077) );
  OR2X2 OR2X2_3164 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_2__6_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2079) );
  OR2X2 OR2X2_3165 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf5), .B(\wb_dat_i[6] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2080) );
  OR2X2 OR2X2_3166 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_2__7_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2082) );
  OR2X2 OR2X2_3167 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf4), .B(\wb_dat_i[7] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2083) );
  OR2X2 OR2X2_3168 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_2__8_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2085) );
  OR2X2 OR2X2_3169 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf3), .B(\wb_dat_i[8] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2086) );
  OR2X2 OR2X2_317 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_0_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_2_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n709) );
  OR2X2 OR2X2_3170 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_2__9_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2088) );
  OR2X2 OR2X2_3171 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf2), .B(\wb_dat_i[9] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2089) );
  OR2X2 OR2X2_3172 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_2__10_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2091) );
  OR2X2 OR2X2_3173 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf1), .B(\wb_dat_i[10] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2092) );
  OR2X2 OR2X2_3174 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_2__11_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2094) );
  OR2X2 OR2X2_3175 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf0), .B(\wb_dat_i[11] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2095) );
  OR2X2 OR2X2_3176 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_2__12_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2097) );
  OR2X2 OR2X2_3177 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf5), .B(\wb_dat_i[12] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2098) );
  OR2X2 OR2X2_3178 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_2__13_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2100) );
  OR2X2 OR2X2_3179 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf4), .B(\wb_dat_i[13] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2101) );
  OR2X2 OR2X2_318 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n685), .B(u_sdrc_core_r2b_len_2_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n710) );
  OR2X2 OR2X2_3180 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_2__14_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2103) );
  OR2X2 OR2X2_3181 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf3), .B(\wb_dat_i[14] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2104) );
  OR2X2 OR2X2_3182 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_2__15_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2106) );
  OR2X2 OR2X2_3183 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf2), .B(\wb_dat_i[15] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2107) );
  OR2X2 OR2X2_3184 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_2__16_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2109) );
  OR2X2 OR2X2_3185 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf1), .B(\wb_dat_i[16] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2110) );
  OR2X2 OR2X2_3186 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_2__17_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2112) );
  OR2X2 OR2X2_3187 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf0), .B(\wb_dat_i[17] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2113) );
  OR2X2 OR2X2_3188 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_2__18_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2115) );
  OR2X2 OR2X2_3189 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf5), .B(\wb_dat_i[18] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2116) );
  OR2X2 OR2X2_319 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_0_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_3_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n712) );
  OR2X2 OR2X2_3190 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_2__19_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2118) );
  OR2X2 OR2X2_3191 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf4), .B(\wb_dat_i[19] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2119) );
  OR2X2 OR2X2_3192 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_2__20_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2121) );
  OR2X2 OR2X2_3193 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf3), .B(\wb_dat_i[20] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2122) );
  OR2X2 OR2X2_3194 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_2__21_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2124) );
  OR2X2 OR2X2_3195 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf2), .B(\wb_dat_i[21] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2125) );
  OR2X2 OR2X2_3196 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_2__22_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2127) );
  OR2X2 OR2X2_3197 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf1), .B(\wb_dat_i[22] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2128) );
  OR2X2 OR2X2_3198 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_2__23_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2130) );
  OR2X2 OR2X2_3199 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf0), .B(\wb_dat_i[23] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2131) );
  OR2X2 OR2X2_32 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n311_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n312), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n313_1) );
  OR2X2 OR2X2_320 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n685), .B(u_sdrc_core_r2b_len_3_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n713) );
  OR2X2 OR2X2_3200 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_2__24_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2133) );
  OR2X2 OR2X2_3201 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf5), .B(\wb_dat_i[24] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2134) );
  OR2X2 OR2X2_3202 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_2__25_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2136) );
  OR2X2 OR2X2_3203 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf4), .B(\wb_dat_i[25] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2137) );
  OR2X2 OR2X2_3204 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_2__26_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2139) );
  OR2X2 OR2X2_3205 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf3), .B(\wb_dat_i[26] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2140) );
  OR2X2 OR2X2_3206 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_2__27_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2142) );
  OR2X2 OR2X2_3207 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf2), .B(\wb_dat_i[27] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2143) );
  OR2X2 OR2X2_3208 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_2__28_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2145) );
  OR2X2 OR2X2_3209 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf1), .B(\wb_dat_i[28] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2146) );
  OR2X2 OR2X2_321 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_0_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_4_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n715) );
  OR2X2 OR2X2_3210 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_2__29_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2148) );
  OR2X2 OR2X2_3211 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf0), .B(\wb_dat_i[29] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2149) );
  OR2X2 OR2X2_3212 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_2__30_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2151) );
  OR2X2 OR2X2_3213 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf5), .B(\wb_dat_i[30] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2152) );
  OR2X2 OR2X2_3214 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_2__31_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2154) );
  OR2X2 OR2X2_3215 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf4), .B(\wb_dat_i[31] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2155) );
  OR2X2 OR2X2_3216 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_2__32_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2157) );
  OR2X2 OR2X2_3217 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_wr_data_32_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2158) );
  OR2X2 OR2X2_3218 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_2__33_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2160) );
  OR2X2 OR2X2_3219 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_wr_data_33_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2161) );
  OR2X2 OR2X2_322 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n685), .B(u_sdrc_core_r2b_len_4_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n716) );
  OR2X2 OR2X2_3220 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_2__34_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2163) );
  OR2X2 OR2X2_3221 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_wr_data_34_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2164) );
  OR2X2 OR2X2_3222 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2059_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_2__35_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2166) );
  OR2X2 OR2X2_3223 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2061_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_wr_data_35_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2167) );
  OR2X2 OR2X2_3224 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_5__0_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2170) );
  OR2X2 OR2X2_3225 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf5), .B(\wb_dat_i[0] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2172) );
  OR2X2 OR2X2_3226 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_5__1_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2174) );
  OR2X2 OR2X2_3227 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf4), .B(\wb_dat_i[1] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2175) );
  OR2X2 OR2X2_3228 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_5__2_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2177) );
  OR2X2 OR2X2_3229 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf3), .B(\wb_dat_i[2] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2178) );
  OR2X2 OR2X2_323 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_0_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_5_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n718) );
  OR2X2 OR2X2_3230 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_5__3_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2180) );
  OR2X2 OR2X2_3231 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf2), .B(\wb_dat_i[3] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2181) );
  OR2X2 OR2X2_3232 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_5__4_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2183) );
  OR2X2 OR2X2_3233 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf1), .B(\wb_dat_i[4] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2184) );
  OR2X2 OR2X2_3234 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_5__5_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2186) );
  OR2X2 OR2X2_3235 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf0), .B(\wb_dat_i[5] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2187) );
  OR2X2 OR2X2_3236 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_5__6_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2189) );
  OR2X2 OR2X2_3237 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf5), .B(\wb_dat_i[6] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2190) );
  OR2X2 OR2X2_3238 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_5__7_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2192) );
  OR2X2 OR2X2_3239 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf4), .B(\wb_dat_i[7] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2193) );
  OR2X2 OR2X2_324 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n685), .B(u_sdrc_core_r2b_len_5_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n719) );
  OR2X2 OR2X2_3240 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_5__8_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2195) );
  OR2X2 OR2X2_3241 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf3), .B(\wb_dat_i[8] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2196) );
  OR2X2 OR2X2_3242 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_5__9_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2198) );
  OR2X2 OR2X2_3243 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf2), .B(\wb_dat_i[9] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2199) );
  OR2X2 OR2X2_3244 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_5__10_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2201) );
  OR2X2 OR2X2_3245 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf1), .B(\wb_dat_i[10] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2202) );
  OR2X2 OR2X2_3246 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_5__11_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2204) );
  OR2X2 OR2X2_3247 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf0), .B(\wb_dat_i[11] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2205) );
  OR2X2 OR2X2_3248 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_5__12_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2207) );
  OR2X2 OR2X2_3249 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf5), .B(\wb_dat_i[12] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2208) );
  OR2X2 OR2X2_325 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_0_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_len_6_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n721) );
  OR2X2 OR2X2_3250 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_5__13_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2210) );
  OR2X2 OR2X2_3251 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf4), .B(\wb_dat_i[13] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2211) );
  OR2X2 OR2X2_3252 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_5__14_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2213) );
  OR2X2 OR2X2_3253 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf3), .B(\wb_dat_i[14] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2214) );
  OR2X2 OR2X2_3254 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_5__15_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2216) );
  OR2X2 OR2X2_3255 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf2), .B(\wb_dat_i[15] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2217) );
  OR2X2 OR2X2_3256 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_5__16_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2219) );
  OR2X2 OR2X2_3257 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf1), .B(\wb_dat_i[16] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2220) );
  OR2X2 OR2X2_3258 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_5__17_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2222) );
  OR2X2 OR2X2_3259 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf0), .B(\wb_dat_i[17] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2223) );
  OR2X2 OR2X2_326 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n685), .B(u_sdrc_core_r2b_len_6_), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n722) );
  OR2X2 OR2X2_3260 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_5__18_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2225) );
  OR2X2 OR2X2_3261 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf5), .B(\wb_dat_i[18] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2226) );
  OR2X2 OR2X2_3262 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_5__19_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2228) );
  OR2X2 OR2X2_3263 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf4), .B(\wb_dat_i[19] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2229) );
  OR2X2 OR2X2_3264 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_5__20_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2231) );
  OR2X2 OR2X2_3265 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf3), .B(\wb_dat_i[20] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2232) );
  OR2X2 OR2X2_3266 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_5__21_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2234) );
  OR2X2 OR2X2_3267 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf2), .B(\wb_dat_i[21] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2235) );
  OR2X2 OR2X2_3268 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_5__22_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2237) );
  OR2X2 OR2X2_3269 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf1), .B(\wb_dat_i[22] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2238) );
  OR2X2 OR2X2_327 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_st_0_), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_l_wrap), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n724) );
  OR2X2 OR2X2_3270 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_5__23_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2240) );
  OR2X2 OR2X2_3271 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf0), .B(\wb_dat_i[23] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2241) );
  OR2X2 OR2X2_3272 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_5__24_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2243) );
  OR2X2 OR2X2_3273 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf5), .B(\wb_dat_i[24] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2244) );
  OR2X2 OR2X2_3274 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_5__25_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2246) );
  OR2X2 OR2X2_3275 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf4), .B(\wb_dat_i[25] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2247) );
  OR2X2 OR2X2_3276 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_5__26_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2249) );
  OR2X2 OR2X2_3277 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf3), .B(\wb_dat_i[26] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2250) );
  OR2X2 OR2X2_3278 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_5__27_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2252) );
  OR2X2 OR2X2_3279 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf2), .B(\wb_dat_i[27] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2253) );
  OR2X2 OR2X2_328 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n685), .B(u_sdrc_core_r2b_wrap), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n725) );
  OR2X2 OR2X2_3280 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_5__28_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2255) );
  OR2X2 OR2X2_3281 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf1), .B(\wb_dat_i[28] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2256) );
  OR2X2 OR2X2_3282 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_5__29_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2258) );
  OR2X2 OR2X2_3283 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf0), .B(\wb_dat_i[29] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2259) );
  OR2X2 OR2X2_3284 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf4), .B(u_wb2sdrc_u_wrdatafifo_mem_5__30_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2261) );
  OR2X2 OR2X2_3285 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf5), .B(\wb_dat_i[30] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2262) );
  OR2X2 OR2X2_3286 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_mem_5__31_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2264) );
  OR2X2 OR2X2_3287 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf4), .B(\wb_dat_i[31] ), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2265) );
  OR2X2 OR2X2_3288 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_mem_5__32_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2267) );
  OR2X2 OR2X2_3289 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf3), .B(u_wb2sdrc_u_wrdatafifo_wr_data_32_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2268) );
  OR2X2 OR2X2_329 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n730), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_wrok_r), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n731) );
  OR2X2 OR2X2_3290 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_mem_5__33_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2270) );
  OR2X2 OR2X2_3291 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf2), .B(u_wb2sdrc_u_wrdatafifo_wr_data_33_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2271) );
  OR2X2 OR2X2_3292 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_mem_5__34_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2273) );
  OR2X2 OR2X2_3293 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf1), .B(u_wb2sdrc_u_wrdatafifo_wr_data_34_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2274) );
  OR2X2 OR2X2_3294 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2169_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_mem_5__35_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2276) );
  OR2X2 OR2X2_3295 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2171_bF_buf0), .B(u_wb2sdrc_u_wrdatafifo_wr_data_35_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2277) );
  OR2X2 OR2X2_3296 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2280), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2281), .Y(u_wb2sdrc_u_wrdatafifo_rd_ptr_0__FF_INPUT) );
  OR2X2 OR2X2_3297 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2284), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf7), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2285) );
  OR2X2 OR2X2_3298 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2285), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2279), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2286) );
  OR2X2 OR2X2_3299 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2287), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2283), .Y(u_wb2sdrc_u_wrdatafifo_rd_ptr_1__FF_INPUT) );
  OR2X2 OR2X2_33 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n295_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n316), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n317_1) );
  OR2X2 OR2X2_330 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm_l_write), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_x2b_rdok_r), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n732) );
  OR2X2 OR2X2_3300 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n1156_bF_buf5), .B(u_wb2sdrc_u_wrdatafifo_rd_ptr_2_bF_buf2), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2292) );
  OR2X2 OR2X2_3301 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2294), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2289), .Y(u_wb2sdrc_u_wrdatafifo_rd_ptr_2__FF_INPUT) );
  OR2X2 OR2X2_3302 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2297), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2298), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2299) );
  OR2X2 OR2X2_3303 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2300), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2296), .Y(u_wb2sdrc_u_wrdatafifo_rd_ptr_3__FF_INPUT) );
  OR2X2 OR2X2_3304 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2302), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2303), .Y(u_wb2sdrc_u_wrdatafifo_grey_rd_ptr_0__FF_INPUT) );
  OR2X2 OR2X2_3305 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2307), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2306), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2308) );
  OR2X2 OR2X2_3306 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2308), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2305), .Y(u_wb2sdrc_u_wrdatafifo_grey_rd_ptr_1__FF_INPUT) );
  OR2X2 OR2X2_3307 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2313), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2312), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2314) );
  OR2X2 OR2X2_3308 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2314), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2311), .Y(u_wb2sdrc_u_wrdatafifo_grey_rd_ptr_2__FF_INPUT) );
  OR2X2 OR2X2_3309 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2300), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2316), .Y(u_wb2sdrc_u_wrdatafifo_grey_rd_ptr_3__FF_INPUT) );
  OR2X2 OR2X2_331 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n735), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n729), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n736) );
  OR2X2 OR2X2_3310 ( .A(u_wb2sdrc_u_wrdatafifo_afull), .B(u_wb2sdrc_u_wrdatafifo_full), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2318) );
  OR2X2 OR2X2_3311 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2319), .B(u_wb2sdrc_u_wrdatafifo_wr_en), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2320) );
  OR2X2 OR2X2_3312 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2326), .B(u_wb2sdrc_u_wrdatafifo_wr_ptr_2_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2327) );
  OR2X2 OR2X2_3313 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2332), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2326), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2333) );
  OR2X2 OR2X2_3314 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2333), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2323), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2334) );
  OR2X2 OR2X2_3315 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2328), .B(u_wb2sdrc_u_wrdatafifo_wr_ptr_3_), .Y(u_wb2sdrc_u_wrdatafifo__abc_19472_n2344) );
  OR2X2 OR2X2_3316 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n817_1), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2354), .Y(u_wb2sdrc_u_wrdatafifo_wr_ptr_0__FF_INPUT) );
  OR2X2 OR2X2_3317 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2335), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2356), .Y(u_wb2sdrc_u_wrdatafifo_wr_ptr_1__FF_INPUT) );
  OR2X2 OR2X2_3318 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2331), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2358), .Y(u_wb2sdrc_u_wrdatafifo_wr_ptr_2__FF_INPUT) );
  OR2X2 OR2X2_3319 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2346), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2360), .Y(u_wb2sdrc_u_wrdatafifo_wr_ptr_3__FF_INPUT) );
  OR2X2 OR2X2_332 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n737), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n728), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_req) );
  OR2X2 OR2X2_3320 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2364), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2365), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1070) );
  OR2X2 OR2X2_3321 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2367), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2368), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1071) );
  OR2X2 OR2X2_3322 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2370), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2371), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1072) );
  OR2X2 OR2X2_3323 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2373), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2374), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1073) );
  OR2X2 OR2X2_3324 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2376), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2377), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1074) );
  OR2X2 OR2X2_3325 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2379), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2380), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1075) );
  OR2X2 OR2X2_3326 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2382), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2383), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1076) );
  OR2X2 OR2X2_3327 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2385), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2386), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1077) );
  OR2X2 OR2X2_3328 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2388), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2389), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1078) );
  OR2X2 OR2X2_3329 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2391), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2392), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1079) );
  OR2X2 OR2X2_333 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n382), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_bank_valid), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n749) );
  OR2X2 OR2X2_3330 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2394), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2395), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1080) );
  OR2X2 OR2X2_3331 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2397), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2398), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1081) );
  OR2X2 OR2X2_3332 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2400), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2401), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1082) );
  OR2X2 OR2X2_3333 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2403), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2404), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1083) );
  OR2X2 OR2X2_3334 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2406), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2407), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1084) );
  OR2X2 OR2X2_3335 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2409), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2410), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1085) );
  OR2X2 OR2X2_3336 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2412), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2413), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1086) );
  OR2X2 OR2X2_3337 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2415), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2416), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1087) );
  OR2X2 OR2X2_3338 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2418), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2419), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1088) );
  OR2X2 OR2X2_3339 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2421), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2422), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1089) );
  OR2X2 OR2X2_334 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n756), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n757), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n758) );
  OR2X2 OR2X2_3340 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2424), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2425), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1090) );
  OR2X2 OR2X2_3341 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2427), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2428), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1091) );
  OR2X2 OR2X2_3342 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2430), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2431), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1092) );
  OR2X2 OR2X2_3343 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2433), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2434), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1093) );
  OR2X2 OR2X2_3344 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2436), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2437), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1094) );
  OR2X2 OR2X2_3345 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2439), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2440), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1095) );
  OR2X2 OR2X2_3346 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2442), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2443), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1096) );
  OR2X2 OR2X2_3347 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2445), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2446), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1097) );
  OR2X2 OR2X2_3348 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2448), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2449), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1098) );
  OR2X2 OR2X2_3349 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2451), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2452), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1099) );
  OR2X2 OR2X2_335 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n760), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n761), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n762) );
  OR2X2 OR2X2_3350 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2454), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2455), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1100) );
  OR2X2 OR2X2_3351 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2457), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2458), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1101) );
  OR2X2 OR2X2_3352 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2460), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2461), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1102) );
  OR2X2 OR2X2_3353 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2463), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2464), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1103) );
  OR2X2 OR2X2_3354 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2466), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2467), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1104) );
  OR2X2 OR2X2_3355 ( .A(u_wb2sdrc_u_wrdatafifo__abc_19472_n2469), .B(u_wb2sdrc_u_wrdatafifo__abc_19472_n2470), .Y(u_wb2sdrc_u_wrdatafifo__abc_14975_n1105) );
  OR2X2 OR2X2_336 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n764), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n765), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n766) );
  OR2X2 OR2X2_337 ( .A(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n768), .B(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n769), .Y(u_sdrc_core_u_bank_ctl_bank0_fsm__abc_24150_n770) );
  OR2X2 OR2X2_338 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n254), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_12_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n255_1) );
  OR2X2 OR2X2_339 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n256_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_11_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n257) );
  OR2X2 OR2X2_34 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n242_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n281_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n318) );
  OR2X2 OR2X2_340 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n258_1), .B(u_sdrc_core_r2b_raddr_12_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n259_1) );
  OR2X2 OR2X2_341 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n262_1), .B(u_sdrc_core_r2b_raddr_11_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n263) );
  OR2X2 OR2X2_342 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n264_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_9_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n265_1) );
  OR2X2 OR2X2_343 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n267_1), .B(u_sdrc_core_r2b_raddr_9_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n268_1) );
  OR2X2 OR2X2_344 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n269), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_7_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n270_1) );
  OR2X2 OR2X2_345 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n274_1), .B(u_sdrc_core_r2b_raddr_7_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n275) );
  OR2X2 OR2X2_346 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n276_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_3_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n277_1) );
  OR2X2 OR2X2_347 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n279_1), .B(u_sdrc_core_r2b_raddr_6_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n280_1) );
  OR2X2 OR2X2_348 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n281), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_6_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n282_1) );
  OR2X2 OR2X2_349 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n285), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_5_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n286_1) );
  OR2X2 OR2X2_35 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n321), .B(u_sdrc_core_u_bank_ctl__abc_21249_n322_1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n323) );
  OR2X2 OR2X2_350 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n287_1), .B(u_sdrc_core_r2b_raddr_1_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n288_1) );
  OR2X2 OR2X2_351 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n290_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_0_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n291_1) );
  OR2X2 OR2X2_352 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n292_1), .B(u_sdrc_core_r2b_raddr_0_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n293) );
  OR2X2 OR2X2_353 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n301), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n298_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n302_1) );
  OR2X2 OR2X2_354 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n306_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n303_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n307_1) );
  OR2X2 OR2X2_355 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n309), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_2_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n310_1) );
  OR2X2 OR2X2_356 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n311_1), .B(u_sdrc_core_r2b_raddr_3_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n312_1) );
  OR2X2 OR2X2_357 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n314_1), .B(u_sdrc_core_r2b_raddr_2_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n315_1) );
  OR2X2 OR2X2_358 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n316_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_1_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n317) );
  OR2X2 OR2X2_359 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n320_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_4_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n321) );
  OR2X2 OR2X2_36 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n320_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n323), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n324_1) );
  OR2X2 OR2X2_360 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n322_1), .B(u_sdrc_core_r2b_raddr_4_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n323_1) );
  OR2X2 OR2X2_361 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n325), .B(u_sdrc_core_r2b_raddr_5_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n326_1) );
  OR2X2 OR2X2_362 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n333), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n251), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_17422_n55) );
  OR2X2 OR2X2_363 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n340), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n335), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_17422_n61) );
  OR2X2 OR2X2_364 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n344_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n345), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n346) );
  OR2X2 OR2X2_365 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n346), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n342), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_17422_n66) );
  OR2X2 OR2X2_366 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n349_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n348_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n350) );
  OR2X2 OR2X2_367 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n351), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n350), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_17422_n82) );
  OR2X2 OR2X2_368 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n359_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n361), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n362) );
  OR2X2 OR2X2_369 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n362), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n354_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_17422_n90) );
  OR2X2 OR2X2_37 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n319), .B(u_sdrc_core_r2b_ba_0_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n325_1) );
  OR2X2 OR2X2_370 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n364_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_2_bF_buf1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n365) );
  OR2X2 OR2X2_371 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_3_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_prech_page_closed), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n368_1) );
  OR2X2 OR2X2_372 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n373_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n365), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n374_1) );
  OR2X2 OR2X2_373 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n377), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n337), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_cmd_r_1__FF_INPUT) );
  OR2X2 OR2X2_374 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n249_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_cmd_1_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n380) );
  OR2X2 OR2X2_375 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_tras_cntr_0_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_tras_cntr_1_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n384_1) );
  OR2X2 OR2X2_376 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n384_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_tras_cntr_2_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n385) );
  OR2X2 OR2X2_377 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n385), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_tras_cntr_3_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n386_1) );
  OR2X2 OR2X2_378 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n388), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n389), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n390) );
  OR2X2 OR2X2_379 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n393), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n394_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n395_1) );
  OR2X2 OR2X2_38 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n328_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n329), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n330) );
  OR2X2 OR2X2_380 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n396_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n392_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n397_1) );
  OR2X2 OR2X2_381 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n400_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n401_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n402_1) );
  OR2X2 OR2X2_382 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n403_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n399_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n404_1) );
  OR2X2 OR2X2_383 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n406_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n382), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n407_1) );
  OR2X2 OR2X2_384 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n383_1), .B(\cfg_sdr_tras_d[3] ), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n408_1) );
  OR2X2 OR2X2_385 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n380), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_cmd_0_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n411_1) );
  OR2X2 OR2X2_386 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_timer0_2_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_timer0_3_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n414_1) );
  OR2X2 OR2X2_387 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n414_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_timer0_1_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n415_1) );
  OR2X2 OR2X2_388 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n416), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n382), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n417_1) );
  OR2X2 OR2X2_389 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n380), .B(\cfg_sdr_trcd_d[0] ), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n418) );
  OR2X2 OR2X2_39 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n320_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n330), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n331) );
  OR2X2 OR2X2_390 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n419_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n412_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n420_1) );
  OR2X2 OR2X2_391 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n411_1), .B(\cfg_sdr_trp_d[0] ), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n421) );
  OR2X2 OR2X2_392 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_timer0_1_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_timer0_0_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n424) );
  OR2X2 OR2X2_393 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n425), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n426), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n427_1) );
  OR2X2 OR2X2_394 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n414_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n424), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n428_1) );
  OR2X2 OR2X2_395 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n412_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n431_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n432) );
  OR2X2 OR2X2_396 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n430), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n432), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n433) );
  OR2X2 OR2X2_397 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n411_1), .B(\cfg_sdr_trp_d[1] ), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n434_1) );
  OR2X2 OR2X2_398 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n424), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_timer0_2_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n437_1) );
  OR2X2 OR2X2_399 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n438_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n439_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n440_1) );
  OR2X2 OR2X2_4 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_cmd_1_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n222) );
  OR2X2 OR2X2_40 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n319), .B(u_sdrc_core_r2b_ba_1_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n332) );
  OR2X2 OR2X2_400 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n412_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n442), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n443) );
  OR2X2 OR2X2_401 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n441), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n443), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n444_1) );
  OR2X2 OR2X2_402 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n411_1), .B(\cfg_sdr_trp_d[2] ), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n445_1) );
  OR2X2 OR2X2_403 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n448_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n382), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n449_1) );
  OR2X2 OR2X2_404 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n380), .B(\cfg_sdr_trcd_d[3] ), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n450) );
  OR2X2 OR2X2_405 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n451), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n412_1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n452) );
  OR2X2 OR2X2_406 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n411_1), .B(\cfg_sdr_trp_d[3] ), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n453_1) );
  OR2X2 OR2X2_407 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n473), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n475), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_0__FF_INPUT) );
  OR2X2 OR2X2_408 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n477), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n479), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_1__FF_INPUT) );
  OR2X2 OR2X2_409 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n481), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n483), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_2__FF_INPUT) );
  OR2X2 OR2X2_41 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n295_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n335), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n336) );
  OR2X2 OR2X2_410 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n485), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n487), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_3__FF_INPUT) );
  OR2X2 OR2X2_411 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n489), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n491), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_4__FF_INPUT) );
  OR2X2 OR2X2_412 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n493), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n495), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_5__FF_INPUT) );
  OR2X2 OR2X2_413 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n497), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n499), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_6__FF_INPUT) );
  OR2X2 OR2X2_414 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n501), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n502), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n503) );
  OR2X2 OR2X2_415 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n505), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n506), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n507) );
  OR2X2 OR2X2_416 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n509), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n510), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n511) );
  OR2X2 OR2X2_417 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n513), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n514), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n515) );
  OR2X2 OR2X2_418 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n517), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n518), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n519) );
  OR2X2 OR2X2_419 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n521), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n522), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n523) );
  OR2X2 OR2X2_42 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n242_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n316), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n337) );
  OR2X2 OR2X2_420 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n525), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n526), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n527) );
  OR2X2 OR2X2_421 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n529), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n530), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n531) );
  OR2X2 OR2X2_422 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n533), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n534), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n535) );
  OR2X2 OR2X2_423 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n537), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n538), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n539) );
  OR2X2 OR2X2_424 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n541), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n542), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n543) );
  OR2X2 OR2X2_425 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n545), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n546), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n547) );
  OR2X2 OR2X2_426 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n549), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n550), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n551) );
  OR2X2 OR2X2_427 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n553), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n554), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n555) );
  OR2X2 OR2X2_428 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n557), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n558), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n559) );
  OR2X2 OR2X2_429 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n561), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n562), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n563) );
  OR2X2 OR2X2_43 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n340), .B(u_sdrc_core_u_bank_ctl__abc_21249_n341), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n342) );
  OR2X2 OR2X2_430 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n565), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n566), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n567) );
  OR2X2 OR2X2_431 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n569), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n570), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n571) );
  OR2X2 OR2X2_432 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n573), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n574), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n575) );
  OR2X2 OR2X2_433 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n577), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n578), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n579) );
  OR2X2 OR2X2_434 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n581), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n582), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n583) );
  OR2X2 OR2X2_435 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n585), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n586), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n587) );
  OR2X2 OR2X2_436 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n589), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n590), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n591) );
  OR2X2 OR2X2_437 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n593), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n594), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n595) );
  OR2X2 OR2X2_438 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n597), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n598), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n599) );
  OR2X2 OR2X2_439 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n601), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n602), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n603) );
  OR2X2 OR2X2_44 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n339), .B(u_sdrc_core_u_bank_ctl__abc_21249_n342), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n343) );
  OR2X2 OR2X2_440 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n368_1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n367), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n606) );
  OR2X2 OR2X2_441 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n607), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n605), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_0_) );
  OR2X2 OR2X2_442 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_0_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n609) );
  OR2X2 OR2X2_443 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_0_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_2_bF_buf3), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n610) );
  OR2X2 OR2X2_444 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n613), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n612), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_1_) );
  OR2X2 OR2X2_445 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_1_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n615) );
  OR2X2 OR2X2_446 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_1_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_2_bF_buf2), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n616) );
  OR2X2 OR2X2_447 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n619), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n618), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_2_) );
  OR2X2 OR2X2_448 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_2_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n621) );
  OR2X2 OR2X2_449 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_2_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_2_bF_buf1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n622) );
  OR2X2 OR2X2_45 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n338), .B(u_sdrc_core_r2b_ba_0_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n344) );
  OR2X2 OR2X2_450 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n625), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n624), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_3_) );
  OR2X2 OR2X2_451 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_3_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n627) );
  OR2X2 OR2X2_452 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_3_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_2_bF_buf0), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n628) );
  OR2X2 OR2X2_453 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n631), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n630), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_4_) );
  OR2X2 OR2X2_454 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_4_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n633) );
  OR2X2 OR2X2_455 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_4_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_2_bF_buf3), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n634) );
  OR2X2 OR2X2_456 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n637), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n636), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_5_) );
  OR2X2 OR2X2_457 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_5_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n639) );
  OR2X2 OR2X2_458 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_5_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_2_bF_buf2), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n640) );
  OR2X2 OR2X2_459 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n643), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n642), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_6_) );
  OR2X2 OR2X2_46 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n347), .B(u_sdrc_core_u_bank_ctl__abc_21249_n348), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n349) );
  OR2X2 OR2X2_460 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_6_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n645) );
  OR2X2 OR2X2_461 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_6_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_2_bF_buf1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n646) );
  OR2X2 OR2X2_462 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n649), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n648), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_7_) );
  OR2X2 OR2X2_463 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_7_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n651) );
  OR2X2 OR2X2_464 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_7_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_2_bF_buf0), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n652) );
  OR2X2 OR2X2_465 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n655), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n654), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_8_) );
  OR2X2 OR2X2_466 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_8_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n657) );
  OR2X2 OR2X2_467 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_8_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_2_bF_buf3), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n658) );
  OR2X2 OR2X2_468 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n661), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n660), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_9_) );
  OR2X2 OR2X2_469 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_9_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n663) );
  OR2X2 OR2X2_47 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n339), .B(u_sdrc_core_u_bank_ctl__abc_21249_n349), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n350) );
  OR2X2 OR2X2_470 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_9_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_2_bF_buf2), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n664) );
  OR2X2 OR2X2_471 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n667), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n666), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_10_) );
  OR2X2 OR2X2_472 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_10_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n669) );
  OR2X2 OR2X2_473 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_10_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_2_bF_buf1), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n670) );
  OR2X2 OR2X2_474 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n673), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n672), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_11_) );
  OR2X2 OR2X2_475 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_11_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n675) );
  OR2X2 OR2X2_476 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_11_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_2_bF_buf0), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n676) );
  OR2X2 OR2X2_477 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n679), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n678), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_12_) );
  OR2X2 OR2X2_478 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_12_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n681) );
  OR2X2 OR2X2_479 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_row_12_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_2_bF_buf3), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n682) );
  OR2X2 OR2X2_48 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n338), .B(u_sdrc_core_r2b_ba_1_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n351) );
  OR2X2 OR2X2_480 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_0_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_last), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n688) );
  OR2X2 OR2X2_481 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n685), .B(u_sdrc_core_r2b_last), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n689) );
  OR2X2 OR2X2_482 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_0_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_0_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n703) );
  OR2X2 OR2X2_483 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n685), .B(u_sdrc_core_r2b_len_0_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n704) );
  OR2X2 OR2X2_484 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_0_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_1_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n706) );
  OR2X2 OR2X2_485 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n685), .B(u_sdrc_core_r2b_len_1_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n707) );
  OR2X2 OR2X2_486 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_0_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_2_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n709) );
  OR2X2 OR2X2_487 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n685), .B(u_sdrc_core_r2b_len_2_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n710) );
  OR2X2 OR2X2_488 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_0_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_3_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n712) );
  OR2X2 OR2X2_489 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n685), .B(u_sdrc_core_r2b_len_3_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n713) );
  OR2X2 OR2X2_49 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n242_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n335), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n354) );
  OR2X2 OR2X2_490 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_0_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_4_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n715) );
  OR2X2 OR2X2_491 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n685), .B(u_sdrc_core_r2b_len_4_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n716) );
  OR2X2 OR2X2_492 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_0_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_5_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n718) );
  OR2X2 OR2X2_493 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n685), .B(u_sdrc_core_r2b_len_5_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n719) );
  OR2X2 OR2X2_494 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_0_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_len_6_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n721) );
  OR2X2 OR2X2_495 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n685), .B(u_sdrc_core_r2b_len_6_), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n722) );
  OR2X2 OR2X2_496 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_st_0_), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_l_wrap), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n724) );
  OR2X2 OR2X2_497 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n685), .B(u_sdrc_core_r2b_wrap), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n725) );
  OR2X2 OR2X2_498 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n730), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_x2b_wrok_r), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n731) );
  OR2X2 OR2X2_499 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_l_write), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_x2b_rdok_r), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n732) );
  OR2X2 OR2X2_5 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n211_1), .B(u_sdrc_core_b2x_ba_1_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n223_1) );
  OR2X2 OR2X2_50 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n295_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n356), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n357) );
  OR2X2 OR2X2_500 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n735), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n729), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n736) );
  OR2X2 OR2X2_501 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n737), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n728), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_req) );
  OR2X2 OR2X2_502 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n382), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_bank_valid), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n749) );
  OR2X2 OR2X2_503 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n756), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n757), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n758) );
  OR2X2 OR2X2_504 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n760), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n761), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n762) );
  OR2X2 OR2X2_505 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n764), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n765), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n766) );
  OR2X2 OR2X2_506 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n768), .B(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n769), .Y(u_sdrc_core_u_bank_ctl_bank1_fsm__abc_24150_n770) );
  OR2X2 OR2X2_507 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n254), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_12_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n255_1) );
  OR2X2 OR2X2_508 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n256_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_11_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n257) );
  OR2X2 OR2X2_509 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n258_1), .B(u_sdrc_core_r2b_raddr_12_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n259_1) );
  OR2X2 OR2X2_51 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n359), .B(u_sdrc_core_u_bank_ctl__abc_21249_n360), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n361) );
  OR2X2 OR2X2_510 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n262_1), .B(u_sdrc_core_r2b_raddr_11_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n263) );
  OR2X2 OR2X2_511 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n264_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_9_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n265_1) );
  OR2X2 OR2X2_512 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n267_1), .B(u_sdrc_core_r2b_raddr_9_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n268_1) );
  OR2X2 OR2X2_513 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n269), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_7_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n270_1) );
  OR2X2 OR2X2_514 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n274_1), .B(u_sdrc_core_r2b_raddr_7_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n275) );
  OR2X2 OR2X2_515 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n276_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_3_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n277_1) );
  OR2X2 OR2X2_516 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n279_1), .B(u_sdrc_core_r2b_raddr_6_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n280_1) );
  OR2X2 OR2X2_517 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n281), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_6_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n282_1) );
  OR2X2 OR2X2_518 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n285), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_5_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n286_1) );
  OR2X2 OR2X2_519 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n287_1), .B(u_sdrc_core_r2b_raddr_1_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n288_1) );
  OR2X2 OR2X2_52 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n358), .B(u_sdrc_core_r2b_ba_0_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n362) );
  OR2X2 OR2X2_520 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n290_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_0_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n291_1) );
  OR2X2 OR2X2_521 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n292_1), .B(u_sdrc_core_r2b_raddr_0_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n293) );
  OR2X2 OR2X2_522 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n301), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n298_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n302_1) );
  OR2X2 OR2X2_523 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n306_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n303_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n307_1) );
  OR2X2 OR2X2_524 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n309), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_2_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n310_1) );
  OR2X2 OR2X2_525 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n311_1), .B(u_sdrc_core_r2b_raddr_3_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n312_1) );
  OR2X2 OR2X2_526 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n314_1), .B(u_sdrc_core_r2b_raddr_2_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n315_1) );
  OR2X2 OR2X2_527 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n316_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_1_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n317) );
  OR2X2 OR2X2_528 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n320_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_4_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n321) );
  OR2X2 OR2X2_529 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n322_1), .B(u_sdrc_core_r2b_raddr_4_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n323_1) );
  OR2X2 OR2X2_53 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n359), .B(u_sdrc_core_u_bank_ctl__abc_21249_n365), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n366) );
  OR2X2 OR2X2_530 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n325), .B(u_sdrc_core_r2b_raddr_5_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n326_1) );
  OR2X2 OR2X2_531 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n333), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n251), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_17422_n55) );
  OR2X2 OR2X2_532 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n340), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n335), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_17422_n61) );
  OR2X2 OR2X2_533 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n344_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n345), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n346) );
  OR2X2 OR2X2_534 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n346), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n342), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_17422_n66) );
  OR2X2 OR2X2_535 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n349_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n348_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n350) );
  OR2X2 OR2X2_536 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n351), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n350), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_17422_n82) );
  OR2X2 OR2X2_537 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n359_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n361), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n362) );
  OR2X2 OR2X2_538 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n362), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n354_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_17422_n90) );
  OR2X2 OR2X2_539 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n364_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_2_bF_buf1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n365) );
  OR2X2 OR2X2_54 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n358), .B(u_sdrc_core_r2b_ba_1_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n367) );
  OR2X2 OR2X2_540 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_3_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_prech_page_closed), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n368_1) );
  OR2X2 OR2X2_541 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n373_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n365), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n374_1) );
  OR2X2 OR2X2_542 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n377), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n337), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_cmd_r_1__FF_INPUT) );
  OR2X2 OR2X2_543 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n249_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_cmd_1_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n380) );
  OR2X2 OR2X2_544 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_tras_cntr_0_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_tras_cntr_1_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n384_1) );
  OR2X2 OR2X2_545 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n384_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_tras_cntr_2_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n385) );
  OR2X2 OR2X2_546 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n385), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_tras_cntr_3_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n386_1) );
  OR2X2 OR2X2_547 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n388), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n389), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n390) );
  OR2X2 OR2X2_548 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n393), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n394_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n395_1) );
  OR2X2 OR2X2_549 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n396_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n392_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n397_1) );
  OR2X2 OR2X2_55 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_0_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n371) );
  OR2X2 OR2X2_550 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n400_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n401_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n402_1) );
  OR2X2 OR2X2_551 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n403_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n399_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n404_1) );
  OR2X2 OR2X2_552 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n406_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n382), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n407_1) );
  OR2X2 OR2X2_553 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n383_1), .B(\cfg_sdr_tras_d[3] ), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n408_1) );
  OR2X2 OR2X2_554 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n380), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_cmd_0_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n411_1) );
  OR2X2 OR2X2_555 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_timer0_2_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_timer0_3_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n414_1) );
  OR2X2 OR2X2_556 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n414_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_timer0_1_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n415_1) );
  OR2X2 OR2X2_557 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n416), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n382), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n417_1) );
  OR2X2 OR2X2_558 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n380), .B(\cfg_sdr_trcd_d[0] ), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n418) );
  OR2X2 OR2X2_559 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n419_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n412_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n420_1) );
  OR2X2 OR2X2_56 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n223_1_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_0_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n372) );
  OR2X2 OR2X2_560 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n411_1), .B(\cfg_sdr_trp_d[0] ), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n421) );
  OR2X2 OR2X2_561 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_timer0_1_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_timer0_0_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n424) );
  OR2X2 OR2X2_562 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n425), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n426), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n427_1) );
  OR2X2 OR2X2_563 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n414_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n424), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n428_1) );
  OR2X2 OR2X2_564 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n412_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n431_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n432) );
  OR2X2 OR2X2_565 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n430), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n432), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n433) );
  OR2X2 OR2X2_566 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n411_1), .B(\cfg_sdr_trp_d[1] ), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n434_1) );
  OR2X2 OR2X2_567 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n424), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_timer0_2_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n437_1) );
  OR2X2 OR2X2_568 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n438_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n439_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n440_1) );
  OR2X2 OR2X2_569 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n412_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n442), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n443) );
  OR2X2 OR2X2_57 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n373), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n374) );
  OR2X2 OR2X2_570 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n441), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n443), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n444_1) );
  OR2X2 OR2X2_571 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n411_1), .B(\cfg_sdr_trp_d[2] ), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n445_1) );
  OR2X2 OR2X2_572 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n448_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n382), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n449_1) );
  OR2X2 OR2X2_573 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n380), .B(\cfg_sdr_trcd_d[3] ), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n450) );
  OR2X2 OR2X2_574 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n451), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n412_1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n452) );
  OR2X2 OR2X2_575 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n411_1), .B(\cfg_sdr_trp_d[3] ), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n453_1) );
  OR2X2 OR2X2_576 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n473), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n475), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_0__FF_INPUT) );
  OR2X2 OR2X2_577 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n477), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n479), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_1__FF_INPUT) );
  OR2X2 OR2X2_578 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n481), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n483), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_2__FF_INPUT) );
  OR2X2 OR2X2_579 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n485), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n487), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_3__FF_INPUT) );
  OR2X2 OR2X2_58 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n283_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_0_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n375) );
  OR2X2 OR2X2_580 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n489), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n491), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_4__FF_INPUT) );
  OR2X2 OR2X2_581 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n493), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n495), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_5__FF_INPUT) );
  OR2X2 OR2X2_582 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n497), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n499), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_6__FF_INPUT) );
  OR2X2 OR2X2_583 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n501), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n502), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n503) );
  OR2X2 OR2X2_584 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n505), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n506), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n507) );
  OR2X2 OR2X2_585 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n509), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n510), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n511) );
  OR2X2 OR2X2_586 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n513), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n514), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n515) );
  OR2X2 OR2X2_587 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n517), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n518), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n519) );
  OR2X2 OR2X2_588 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n521), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n522), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n523) );
  OR2X2 OR2X2_589 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n525), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n526), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n527) );
  OR2X2 OR2X2_59 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n377), .B(u_sdrc_core_u_bank_ctl__abc_21249_n370), .Y(u_sdrc_core_b2x_addr_0_) );
  OR2X2 OR2X2_590 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n529), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n530), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n531) );
  OR2X2 OR2X2_591 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n533), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n534), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n535) );
  OR2X2 OR2X2_592 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n537), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n538), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n539) );
  OR2X2 OR2X2_593 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n541), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n542), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n543) );
  OR2X2 OR2X2_594 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n545), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n546), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n547) );
  OR2X2 OR2X2_595 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n549), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n550), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n551) );
  OR2X2 OR2X2_596 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n553), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n554), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n555) );
  OR2X2 OR2X2_597 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n557), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n558), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n559) );
  OR2X2 OR2X2_598 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n561), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n562), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n563) );
  OR2X2 OR2X2_599 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n565), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n566), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n567) );
  OR2X2 OR2X2_6 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n223_1_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_cmd_1_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n224_1) );
  OR2X2 OR2X2_60 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_1_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n380) );
  OR2X2 OR2X2_600 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n569), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n570), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n571) );
  OR2X2 OR2X2_601 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n573), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n574), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n575) );
  OR2X2 OR2X2_602 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n577), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n578), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n579) );
  OR2X2 OR2X2_603 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n581), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n582), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n583) );
  OR2X2 OR2X2_604 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n585), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n586), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n587) );
  OR2X2 OR2X2_605 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n589), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n590), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n591) );
  OR2X2 OR2X2_606 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n593), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n594), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n595) );
  OR2X2 OR2X2_607 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n597), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n598), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n599) );
  OR2X2 OR2X2_608 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n601), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n602), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n603) );
  OR2X2 OR2X2_609 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n368_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n367), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n606) );
  OR2X2 OR2X2_61 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n223_1_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_1_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n381) );
  OR2X2 OR2X2_610 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n607), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n605), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_0_) );
  OR2X2 OR2X2_611 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_0_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n609) );
  OR2X2 OR2X2_612 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_0_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_2_bF_buf3), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n610) );
  OR2X2 OR2X2_613 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n613), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n612), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_1_) );
  OR2X2 OR2X2_614 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_1_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n615) );
  OR2X2 OR2X2_615 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_1_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_2_bF_buf2), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n616) );
  OR2X2 OR2X2_616 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n619), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n618), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_2_) );
  OR2X2 OR2X2_617 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_2_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n621) );
  OR2X2 OR2X2_618 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_2_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_2_bF_buf1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n622) );
  OR2X2 OR2X2_619 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n625), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n624), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_3_) );
  OR2X2 OR2X2_62 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n382), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf0), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n383) );
  OR2X2 OR2X2_620 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_3_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n627) );
  OR2X2 OR2X2_621 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_3_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_2_bF_buf0), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n628) );
  OR2X2 OR2X2_622 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n631), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n630), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_4_) );
  OR2X2 OR2X2_623 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_4_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n633) );
  OR2X2 OR2X2_624 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_4_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_2_bF_buf3), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n634) );
  OR2X2 OR2X2_625 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n637), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n636), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_5_) );
  OR2X2 OR2X2_626 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_5_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n639) );
  OR2X2 OR2X2_627 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_5_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_2_bF_buf2), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n640) );
  OR2X2 OR2X2_628 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n643), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n642), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_6_) );
  OR2X2 OR2X2_629 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_6_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n645) );
  OR2X2 OR2X2_63 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n283_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_1_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n384) );
  OR2X2 OR2X2_630 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_6_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_2_bF_buf1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n646) );
  OR2X2 OR2X2_631 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n649), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n648), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_7_) );
  OR2X2 OR2X2_632 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_7_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n651) );
  OR2X2 OR2X2_633 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_7_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_2_bF_buf0), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n652) );
  OR2X2 OR2X2_634 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n655), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n654), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_8_) );
  OR2X2 OR2X2_635 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_8_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n657) );
  OR2X2 OR2X2_636 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_8_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_2_bF_buf3), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n658) );
  OR2X2 OR2X2_637 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n661), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n660), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_9_) );
  OR2X2 OR2X2_638 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_9_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n663) );
  OR2X2 OR2X2_639 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_9_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_2_bF_buf2), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n664) );
  OR2X2 OR2X2_64 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n386), .B(u_sdrc_core_u_bank_ctl__abc_21249_n379), .Y(u_sdrc_core_b2x_addr_1_) );
  OR2X2 OR2X2_640 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n667), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n666), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_10_) );
  OR2X2 OR2X2_641 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_10_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n669) );
  OR2X2 OR2X2_642 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_10_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_2_bF_buf1), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n670) );
  OR2X2 OR2X2_643 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n673), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n672), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_11_) );
  OR2X2 OR2X2_644 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_11_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n675) );
  OR2X2 OR2X2_645 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_11_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_2_bF_buf0), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n676) );
  OR2X2 OR2X2_646 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n679), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n678), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_12_) );
  OR2X2 OR2X2_647 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_12_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n681) );
  OR2X2 OR2X2_648 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_row_12_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_2_bF_buf3), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n682) );
  OR2X2 OR2X2_649 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_0_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_last), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n688) );
  OR2X2 OR2X2_65 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_2_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n389) );
  OR2X2 OR2X2_650 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n685), .B(u_sdrc_core_r2b_last), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n689) );
  OR2X2 OR2X2_651 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_0_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_0_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n703) );
  OR2X2 OR2X2_652 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n685), .B(u_sdrc_core_r2b_len_0_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n704) );
  OR2X2 OR2X2_653 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_0_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_1_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n706) );
  OR2X2 OR2X2_654 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n685), .B(u_sdrc_core_r2b_len_1_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n707) );
  OR2X2 OR2X2_655 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_0_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_2_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n709) );
  OR2X2 OR2X2_656 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n685), .B(u_sdrc_core_r2b_len_2_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n710) );
  OR2X2 OR2X2_657 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_0_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_3_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n712) );
  OR2X2 OR2X2_658 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n685), .B(u_sdrc_core_r2b_len_3_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n713) );
  OR2X2 OR2X2_659 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_0_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_4_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n715) );
  OR2X2 OR2X2_66 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n223_1_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_2_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n390) );
  OR2X2 OR2X2_660 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n685), .B(u_sdrc_core_r2b_len_4_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n716) );
  OR2X2 OR2X2_661 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_0_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_5_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n718) );
  OR2X2 OR2X2_662 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n685), .B(u_sdrc_core_r2b_len_5_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n719) );
  OR2X2 OR2X2_663 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_0_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_len_6_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n721) );
  OR2X2 OR2X2_664 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n685), .B(u_sdrc_core_r2b_len_6_), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n722) );
  OR2X2 OR2X2_665 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_st_0_), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_l_wrap), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n724) );
  OR2X2 OR2X2_666 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n685), .B(u_sdrc_core_r2b_wrap), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n725) );
  OR2X2 OR2X2_667 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n730), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_x2b_wrok_r), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n731) );
  OR2X2 OR2X2_668 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm_l_write), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_x2b_rdok_r), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n732) );
  OR2X2 OR2X2_669 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n735), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n729), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n736) );
  OR2X2 OR2X2_67 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n391), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf4), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n392) );
  OR2X2 OR2X2_670 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n737), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n728), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_req) );
  OR2X2 OR2X2_671 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n382), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_bank_valid), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n749) );
  OR2X2 OR2X2_672 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n756), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n757), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n758) );
  OR2X2 OR2X2_673 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n760), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n761), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n762) );
  OR2X2 OR2X2_674 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n764), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n765), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n766) );
  OR2X2 OR2X2_675 ( .A(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n768), .B(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n769), .Y(u_sdrc_core_u_bank_ctl_bank2_fsm__abc_24150_n770) );
  OR2X2 OR2X2_676 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n254), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_12_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n255_1) );
  OR2X2 OR2X2_677 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n256_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_11_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n257) );
  OR2X2 OR2X2_678 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n258_1), .B(u_sdrc_core_r2b_raddr_12_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n259_1) );
  OR2X2 OR2X2_679 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n262_1), .B(u_sdrc_core_r2b_raddr_11_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n263) );
  OR2X2 OR2X2_68 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n283_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_2_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n393) );
  OR2X2 OR2X2_680 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n264_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_9_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n265_1) );
  OR2X2 OR2X2_681 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n267_1), .B(u_sdrc_core_r2b_raddr_9_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n268_1) );
  OR2X2 OR2X2_682 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n269), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_7_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n270_1) );
  OR2X2 OR2X2_683 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n274_1), .B(u_sdrc_core_r2b_raddr_7_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n275) );
  OR2X2 OR2X2_684 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n276_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_3_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n277_1) );
  OR2X2 OR2X2_685 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n279_1), .B(u_sdrc_core_r2b_raddr_6_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n280_1) );
  OR2X2 OR2X2_686 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n281), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_6_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n282_1) );
  OR2X2 OR2X2_687 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n285), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_5_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n286_1) );
  OR2X2 OR2X2_688 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n287_1), .B(u_sdrc_core_r2b_raddr_1_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n288_1) );
  OR2X2 OR2X2_689 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n290_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_0_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n291_1) );
  OR2X2 OR2X2_69 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n395), .B(u_sdrc_core_u_bank_ctl__abc_21249_n388), .Y(u_sdrc_core_b2x_addr_2_) );
  OR2X2 OR2X2_690 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n292_1), .B(u_sdrc_core_r2b_raddr_0_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n293) );
  OR2X2 OR2X2_691 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n301), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n298_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n302_1) );
  OR2X2 OR2X2_692 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n306_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n303_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n307_1) );
  OR2X2 OR2X2_693 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n309), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_2_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n310_1) );
  OR2X2 OR2X2_694 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n311_1), .B(u_sdrc_core_r2b_raddr_3_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n312_1) );
  OR2X2 OR2X2_695 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n314_1), .B(u_sdrc_core_r2b_raddr_2_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n315_1) );
  OR2X2 OR2X2_696 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n316_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_1_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n317) );
  OR2X2 OR2X2_697 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n320_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_4_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n321) );
  OR2X2 OR2X2_698 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n322_1), .B(u_sdrc_core_r2b_raddr_4_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n323_1) );
  OR2X2 OR2X2_699 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n325), .B(u_sdrc_core_r2b_raddr_5_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n326_1) );
  OR2X2 OR2X2_7 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n225_1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf4), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n226_1) );
  OR2X2 OR2X2_70 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_3_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n398) );
  OR2X2 OR2X2_700 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n333), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n251), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_17422_n55) );
  OR2X2 OR2X2_701 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n340), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n335), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_17422_n61) );
  OR2X2 OR2X2_702 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n344_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n345), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n346) );
  OR2X2 OR2X2_703 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n346), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n342), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_17422_n66) );
  OR2X2 OR2X2_704 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n349_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n348_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n350) );
  OR2X2 OR2X2_705 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n351), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n350), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_17422_n82) );
  OR2X2 OR2X2_706 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n359_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n361), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n362) );
  OR2X2 OR2X2_707 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n362), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n354_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_17422_n90) );
  OR2X2 OR2X2_708 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n364_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_2_bF_buf1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n365) );
  OR2X2 OR2X2_709 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_3_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_prech_page_closed), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n368_1) );
  OR2X2 OR2X2_71 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n223_1_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_3_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n399) );
  OR2X2 OR2X2_710 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n373_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n365), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n374_1) );
  OR2X2 OR2X2_711 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n377), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n337), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_cmd_r_1__FF_INPUT) );
  OR2X2 OR2X2_712 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n249_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_cmd_1_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n380) );
  OR2X2 OR2X2_713 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_tras_cntr_0_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_tras_cntr_1_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n384_1) );
  OR2X2 OR2X2_714 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n384_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_tras_cntr_2_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n385) );
  OR2X2 OR2X2_715 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n385), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_tras_cntr_3_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n386_1) );
  OR2X2 OR2X2_716 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n388), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n389), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n390) );
  OR2X2 OR2X2_717 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n393), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n394_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n395_1) );
  OR2X2 OR2X2_718 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n396_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n392_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n397_1) );
  OR2X2 OR2X2_719 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n400_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n401_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n402_1) );
  OR2X2 OR2X2_72 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n400), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf3), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n401) );
  OR2X2 OR2X2_720 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n403_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n399_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n404_1) );
  OR2X2 OR2X2_721 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n406_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n382), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n407_1) );
  OR2X2 OR2X2_722 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n383_1), .B(\cfg_sdr_tras_d[3] ), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n408_1) );
  OR2X2 OR2X2_723 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n380), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_cmd_0_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n411_1) );
  OR2X2 OR2X2_724 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_timer0_2_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_timer0_3_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n414_1) );
  OR2X2 OR2X2_725 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n414_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_timer0_1_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n415_1) );
  OR2X2 OR2X2_726 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n416), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n382), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n417_1) );
  OR2X2 OR2X2_727 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n380), .B(\cfg_sdr_trcd_d[0] ), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n418) );
  OR2X2 OR2X2_728 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n419_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n412_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n420_1) );
  OR2X2 OR2X2_729 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n411_1), .B(\cfg_sdr_trp_d[0] ), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n421) );
  OR2X2 OR2X2_73 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n283_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_3_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n402) );
  OR2X2 OR2X2_730 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_timer0_1_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_timer0_0_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n424) );
  OR2X2 OR2X2_731 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n425), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n426), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n427_1) );
  OR2X2 OR2X2_732 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n414_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n424), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n428_1) );
  OR2X2 OR2X2_733 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n412_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n431_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n432) );
  OR2X2 OR2X2_734 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n430), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n432), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n433) );
  OR2X2 OR2X2_735 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n411_1), .B(\cfg_sdr_trp_d[1] ), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n434_1) );
  OR2X2 OR2X2_736 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n424), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_timer0_2_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n437_1) );
  OR2X2 OR2X2_737 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n438_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n439_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n440_1) );
  OR2X2 OR2X2_738 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n412_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n442), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n443) );
  OR2X2 OR2X2_739 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n441), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n443), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n444_1) );
  OR2X2 OR2X2_74 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n404), .B(u_sdrc_core_u_bank_ctl__abc_21249_n397), .Y(u_sdrc_core_b2x_addr_3_) );
  OR2X2 OR2X2_740 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n411_1), .B(\cfg_sdr_trp_d[2] ), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n445_1) );
  OR2X2 OR2X2_741 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n448_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n382), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n449_1) );
  OR2X2 OR2X2_742 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n380), .B(\cfg_sdr_trcd_d[3] ), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n450) );
  OR2X2 OR2X2_743 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n451), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n412_1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n452) );
  OR2X2 OR2X2_744 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n411_1), .B(\cfg_sdr_trp_d[3] ), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n453_1) );
  OR2X2 OR2X2_745 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n473), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n475), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_0__FF_INPUT) );
  OR2X2 OR2X2_746 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n477), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n479), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_1__FF_INPUT) );
  OR2X2 OR2X2_747 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n481), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n483), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_2__FF_INPUT) );
  OR2X2 OR2X2_748 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n485), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n487), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_3__FF_INPUT) );
  OR2X2 OR2X2_749 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n489), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n491), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_4__FF_INPUT) );
  OR2X2 OR2X2_75 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_4_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n407) );
  OR2X2 OR2X2_750 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n493), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n495), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_5__FF_INPUT) );
  OR2X2 OR2X2_751 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n497), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n499), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_6__FF_INPUT) );
  OR2X2 OR2X2_752 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n501), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n502), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n503) );
  OR2X2 OR2X2_753 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n505), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n506), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n507) );
  OR2X2 OR2X2_754 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n509), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n510), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n511) );
  OR2X2 OR2X2_755 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n513), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n514), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n515) );
  OR2X2 OR2X2_756 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n517), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n518), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n519) );
  OR2X2 OR2X2_757 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n521), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n522), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n523) );
  OR2X2 OR2X2_758 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n525), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n526), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n527) );
  OR2X2 OR2X2_759 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n529), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n530), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n531) );
  OR2X2 OR2X2_76 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n223_1_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_4_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n408) );
  OR2X2 OR2X2_760 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n533), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n534), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n535) );
  OR2X2 OR2X2_761 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n537), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n538), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n539) );
  OR2X2 OR2X2_762 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n541), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n542), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n543) );
  OR2X2 OR2X2_763 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n545), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n546), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n547) );
  OR2X2 OR2X2_764 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n549), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n550), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n551) );
  OR2X2 OR2X2_765 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n553), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n554), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n555) );
  OR2X2 OR2X2_766 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n557), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n558), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n559) );
  OR2X2 OR2X2_767 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n561), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n562), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n563) );
  OR2X2 OR2X2_768 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n565), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n566), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n567) );
  OR2X2 OR2X2_769 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n569), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n570), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n571) );
  OR2X2 OR2X2_77 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n409), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf2), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n410) );
  OR2X2 OR2X2_770 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n573), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n574), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n575) );
  OR2X2 OR2X2_771 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n577), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n578), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n579) );
  OR2X2 OR2X2_772 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n581), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n582), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n583) );
  OR2X2 OR2X2_773 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n585), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n586), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n587) );
  OR2X2 OR2X2_774 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n589), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n590), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n591) );
  OR2X2 OR2X2_775 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n593), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n594), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n595) );
  OR2X2 OR2X2_776 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n597), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n598), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n599) );
  OR2X2 OR2X2_777 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n601), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n602), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n603) );
  OR2X2 OR2X2_778 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n368_1), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n367), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n606) );
  OR2X2 OR2X2_779 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n607), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n605), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_0_) );
  OR2X2 OR2X2_78 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n283_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_4_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n411) );
  OR2X2 OR2X2_780 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_0_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n609) );
  OR2X2 OR2X2_781 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_0_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_2_bF_buf3), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n610) );
  OR2X2 OR2X2_782 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n613), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n612), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_1_) );
  OR2X2 OR2X2_783 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_1_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n615) );
  OR2X2 OR2X2_784 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_1_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_2_bF_buf2), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n616) );
  OR2X2 OR2X2_785 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n619), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n618), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_2_) );
  OR2X2 OR2X2_786 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_2_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n621) );
  OR2X2 OR2X2_787 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_2_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_2_bF_buf1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n622) );
  OR2X2 OR2X2_788 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n625), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n624), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_3_) );
  OR2X2 OR2X2_789 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_3_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n627) );
  OR2X2 OR2X2_79 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n413), .B(u_sdrc_core_u_bank_ctl__abc_21249_n406), .Y(u_sdrc_core_b2x_addr_4_) );
  OR2X2 OR2X2_790 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_3_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_2_bF_buf0), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n628) );
  OR2X2 OR2X2_791 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n631), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n630), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_4_) );
  OR2X2 OR2X2_792 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_4_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n633) );
  OR2X2 OR2X2_793 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_4_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_2_bF_buf3), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n634) );
  OR2X2 OR2X2_794 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n637), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n636), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_5_) );
  OR2X2 OR2X2_795 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_5_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n639) );
  OR2X2 OR2X2_796 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_5_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_2_bF_buf2), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n640) );
  OR2X2 OR2X2_797 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n643), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n642), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_6_) );
  OR2X2 OR2X2_798 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_6_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n645) );
  OR2X2 OR2X2_799 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_6_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_2_bF_buf1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n646) );
  OR2X2 OR2X2_8 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n213), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_cmd_1_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n228_1) );
  OR2X2 OR2X2_80 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_5_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n416) );
  OR2X2 OR2X2_800 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n649), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n648), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_7_) );
  OR2X2 OR2X2_801 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_7_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n651) );
  OR2X2 OR2X2_802 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_7_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_2_bF_buf0), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n652) );
  OR2X2 OR2X2_803 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n655), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n654), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_8_) );
  OR2X2 OR2X2_804 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_8_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n657) );
  OR2X2 OR2X2_805 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_8_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_2_bF_buf3), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n658) );
  OR2X2 OR2X2_806 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n661), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n660), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_9_) );
  OR2X2 OR2X2_807 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_9_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n663) );
  OR2X2 OR2X2_808 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_9_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_2_bF_buf2), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n664) );
  OR2X2 OR2X2_809 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n667), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n666), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_10_) );
  OR2X2 OR2X2_81 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n223_1_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_5_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n417) );
  OR2X2 OR2X2_810 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_10_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n669) );
  OR2X2 OR2X2_811 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_10_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_2_bF_buf1), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n670) );
  OR2X2 OR2X2_812 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n673), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n672), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_11_) );
  OR2X2 OR2X2_813 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_11_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n675) );
  OR2X2 OR2X2_814 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_11_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_2_bF_buf0), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n676) );
  OR2X2 OR2X2_815 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n679), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n678), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_12_) );
  OR2X2 OR2X2_816 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_addr_12_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n366), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n681) );
  OR2X2 OR2X2_817 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_row_12_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_2_bF_buf3), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n682) );
  OR2X2 OR2X2_818 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_0_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_last), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n688) );
  OR2X2 OR2X2_819 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n685), .B(u_sdrc_core_r2b_last), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n689) );
  OR2X2 OR2X2_82 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n418), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf1), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n419) );
  OR2X2 OR2X2_820 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_0_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_0_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n703) );
  OR2X2 OR2X2_821 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n685), .B(u_sdrc_core_r2b_len_0_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n704) );
  OR2X2 OR2X2_822 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_0_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_1_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n706) );
  OR2X2 OR2X2_823 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n685), .B(u_sdrc_core_r2b_len_1_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n707) );
  OR2X2 OR2X2_824 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_0_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_2_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n709) );
  OR2X2 OR2X2_825 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n685), .B(u_sdrc_core_r2b_len_2_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n710) );
  OR2X2 OR2X2_826 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_0_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_3_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n712) );
  OR2X2 OR2X2_827 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n685), .B(u_sdrc_core_r2b_len_3_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n713) );
  OR2X2 OR2X2_828 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_0_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_4_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n715) );
  OR2X2 OR2X2_829 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n685), .B(u_sdrc_core_r2b_len_4_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n716) );
  OR2X2 OR2X2_83 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n283_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_5_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n420) );
  OR2X2 OR2X2_830 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_0_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_5_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n718) );
  OR2X2 OR2X2_831 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n685), .B(u_sdrc_core_r2b_len_5_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n719) );
  OR2X2 OR2X2_832 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_0_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_len_6_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n721) );
  OR2X2 OR2X2_833 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n685), .B(u_sdrc_core_r2b_len_6_), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n722) );
  OR2X2 OR2X2_834 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_st_0_), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_l_wrap), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n724) );
  OR2X2 OR2X2_835 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n685), .B(u_sdrc_core_r2b_wrap), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n725) );
  OR2X2 OR2X2_836 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n730), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_x2b_wrok_r), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n731) );
  OR2X2 OR2X2_837 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm_l_write), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_x2b_rdok_r), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n732) );
  OR2X2 OR2X2_838 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n735), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n729), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n736) );
  OR2X2 OR2X2_839 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n737), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n728), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm_b2x_req) );
  OR2X2 OR2X2_84 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n422), .B(u_sdrc_core_u_bank_ctl__abc_21249_n415), .Y(u_sdrc_core_b2x_addr_5_) );
  OR2X2 OR2X2_840 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n382), .B(u_sdrc_core_u_bank_ctl_bank3_fsm_bank_valid), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n749) );
  OR2X2 OR2X2_841 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n756), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n757), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n758) );
  OR2X2 OR2X2_842 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n760), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n761), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n762) );
  OR2X2 OR2X2_843 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n764), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n765), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n766) );
  OR2X2 OR2X2_844 ( .A(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n768), .B(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n769), .Y(u_sdrc_core_u_bank_ctl_bank3_fsm__abc_24150_n770) );
  OR2X2 OR2X2_845 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n171_1_bF_buf3), .B(app_wr_data_0_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n172_1) );
  OR2X2 OR2X2_846 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n173_1), .B(u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf4), .Y(u_sdrc_core_u_bs_convert__abc_21684_n174_1) );
  OR2X2 OR2X2_847 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n175_1), .B(u_sdrc_core_u_bs_convert_wr_xfr_count_1_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n176_1) );
  OR2X2 OR2X2_848 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n179_1), .B(u_sdrc_core_u_bs_convert_wr_xfr_count_1_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n180_1) );
  OR2X2 OR2X2_849 ( .A(app_wr_data_16_), .B(u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n181_1) );
  OR2X2 OR2X2_85 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_6_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n425) );
  OR2X2 OR2X2_850 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n178_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n182_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n183_1) );
  OR2X2 OR2X2_851 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n175_1), .B(app_wr_data_16_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n192_1) );
  OR2X2 OR2X2_852 ( .A(app_wr_data_0_), .B(u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf4), .Y(u_sdrc_core_u_bs_convert__abc_21684_n193_1) );
  OR2X2 OR2X2_853 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n195_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n170_1_bF_buf2), .Y(u_sdrc_core_u_bs_convert__abc_21684_n196) );
  OR2X2 OR2X2_854 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n191_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n196), .Y(u_sdrc_core_u_bs_convert__abc_21684_n197_1) );
  OR2X2 OR2X2_855 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n200_1), .B(u_sdrc_core_u_bs_convert_wr_xfr_count_1_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n201_1) );
  OR2X2 OR2X2_856 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf2), .B(app_wr_data_17_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n202) );
  OR2X2 OR2X2_857 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n199), .B(u_sdrc_core_u_bs_convert__abc_21684_n203_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n204_1) );
  OR2X2 OR2X2_858 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n210_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n170_1_bF_buf1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n211) );
  OR2X2 OR2X2_859 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n212_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n214), .Y(u_sdrc_core_u_bs_convert__abc_21684_n215_1) );
  OR2X2 OR2X2_86 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n223_1_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_6_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n426) );
  OR2X2 OR2X2_860 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n209_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n215_1), .Y(u_sdrc_core_a2x_wrdt_1_) );
  OR2X2 OR2X2_861 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_1_), .B(app_wr_data_10_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n218_1) );
  OR2X2 OR2X2_862 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n219), .B(u_sdrc_core_u_bs_convert__abc_21684_n220_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n221) );
  OR2X2 OR2X2_863 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n217), .B(u_sdrc_core_u_bs_convert__abc_21684_n221), .Y(u_sdrc_core_u_bs_convert__abc_21684_n222_1) );
  OR2X2 OR2X2_864 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n228_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n230_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n231) );
  OR2X2 OR2X2_865 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n227), .B(u_sdrc_core_u_bs_convert__abc_21684_n231), .Y(u_sdrc_core_a2x_wrdt_2_) );
  OR2X2 OR2X2_866 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_1_), .B(app_wr_data_11_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n234_1) );
  OR2X2 OR2X2_867 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n235_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n236_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n237) );
  OR2X2 OR2X2_868 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n233), .B(u_sdrc_core_u_bs_convert__abc_21684_n237), .Y(u_sdrc_core_u_bs_convert__abc_21684_n238_1) );
  OR2X2 OR2X2_869 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n244_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n246_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n247) );
  OR2X2 OR2X2_87 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n427), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf0), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n428) );
  OR2X2 OR2X2_870 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n243), .B(u_sdrc_core_u_bs_convert__abc_21684_n247), .Y(u_sdrc_core_a2x_wrdt_3_) );
  OR2X2 OR2X2_871 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n187_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n252), .Y(u_sdrc_core_u_bs_convert__abc_21684_n253_1) );
  OR2X2 OR2X2_872 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n251_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n253_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n254) );
  OR2X2 OR2X2_873 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n249), .B(u_sdrc_core_u_bs_convert__abc_21684_n254), .Y(u_sdrc_core_u_bs_convert__abc_21684_n255_1) );
  OR2X2 OR2X2_874 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n175_1), .B(app_wr_data_20_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n262) );
  OR2X2 OR2X2_875 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf0), .B(app_wr_data_4_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n263) );
  OR2X2 OR2X2_876 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n265), .B(u_sdrc_core_u_bs_convert__abc_21684_n261), .Y(u_sdrc_core_u_bs_convert__abc_21684_n266) );
  OR2X2 OR2X2_877 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n260), .B(u_sdrc_core_u_bs_convert__abc_21684_n266), .Y(u_sdrc_core_a2x_wrdt_4_) );
  OR2X2 OR2X2_878 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n187_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n270_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n271) );
  OR2X2 OR2X2_879 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n269), .B(u_sdrc_core_u_bs_convert__abc_21684_n271), .Y(u_sdrc_core_u_bs_convert__abc_21684_n272) );
  OR2X2 OR2X2_88 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n283_bF_buf0), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_6_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n429) );
  OR2X2 OR2X2_880 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n268), .B(u_sdrc_core_u_bs_convert__abc_21684_n272), .Y(u_sdrc_core_u_bs_convert__abc_21684_n273) );
  OR2X2 OR2X2_881 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n175_1), .B(app_wr_data_21_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n279_1) );
  OR2X2 OR2X2_882 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf4), .B(app_wr_data_5_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n280) );
  OR2X2 OR2X2_883 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n282), .B(u_sdrc_core_u_bs_convert__abc_21684_n170_1_bF_buf3), .Y(u_sdrc_core_u_bs_convert__abc_21684_n283) );
  OR2X2 OR2X2_884 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n278), .B(u_sdrc_core_u_bs_convert__abc_21684_n283), .Y(u_sdrc_core_u_bs_convert__abc_21684_n284) );
  OR2X2 OR2X2_885 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n171_1_bF_buf2), .B(app_wr_data_5_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n285) );
  OR2X2 OR2X2_886 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n187_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n289), .Y(u_sdrc_core_u_bs_convert__abc_21684_n290) );
  OR2X2 OR2X2_887 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n288_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n290), .Y(u_sdrc_core_u_bs_convert__abc_21684_n291) );
  OR2X2 OR2X2_888 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n287), .B(u_sdrc_core_u_bs_convert__abc_21684_n291), .Y(u_sdrc_core_u_bs_convert__abc_21684_n292) );
  OR2X2 OR2X2_889 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n298), .B(u_sdrc_core_u_bs_convert__abc_21684_n300), .Y(u_sdrc_core_u_bs_convert__abc_21684_n301) );
  OR2X2 OR2X2_89 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n431), .B(u_sdrc_core_u_bank_ctl__abc_21249_n424), .Y(u_sdrc_core_b2x_addr_6_) );
  OR2X2 OR2X2_890 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n297_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n301), .Y(u_sdrc_core_a2x_wrdt_6_) );
  OR2X2 OR2X2_891 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n187_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n305), .Y(u_sdrc_core_u_bs_convert__abc_21684_n306_1) );
  OR2X2 OR2X2_892 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n304), .B(u_sdrc_core_u_bs_convert__abc_21684_n306_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n307) );
  OR2X2 OR2X2_893 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n303), .B(u_sdrc_core_u_bs_convert__abc_21684_n307), .Y(u_sdrc_core_u_bs_convert__abc_21684_n308) );
  OR2X2 OR2X2_894 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n175_1), .B(app_wr_data_23_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n314) );
  OR2X2 OR2X2_895 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf2), .B(app_wr_data_7_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n315_1) );
  OR2X2 OR2X2_896 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n317), .B(u_sdrc_core_u_bs_convert__abc_21684_n170_1_bF_buf2), .Y(u_sdrc_core_u_bs_convert__abc_21684_n318) );
  OR2X2 OR2X2_897 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n313), .B(u_sdrc_core_u_bs_convert__abc_21684_n318), .Y(u_sdrc_core_u_bs_convert__abc_21684_n319) );
  OR2X2 OR2X2_898 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n171_1_bF_buf1), .B(app_wr_data_7_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n320) );
  OR2X2 OR2X2_899 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n322), .B(u_sdrc_core_u_bs_convert__abc_21684_n324_1), .Y(u_sdrc_core_a2x_wrdt_8_) );
  OR2X2 OR2X2_9 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n230_1), .B(u_sdrc_core_u_bank_ctl__abc_21249_n221_1), .Y(u_sdrc_core_b2x_cmd_1_) );
  OR2X2 OR2X2_90 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf4), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_7_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n434) );
  OR2X2 OR2X2_900 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n326), .B(u_sdrc_core_u_bs_convert__abc_21684_n328), .Y(u_sdrc_core_a2x_wrdt_9_) );
  OR2X2 OR2X2_901 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n330), .B(u_sdrc_core_u_bs_convert__abc_21684_n332), .Y(u_sdrc_core_a2x_wrdt_10_) );
  OR2X2 OR2X2_902 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n334), .B(u_sdrc_core_u_bs_convert__abc_21684_n336), .Y(u_sdrc_core_a2x_wrdt_11_) );
  OR2X2 OR2X2_903 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n338), .B(u_sdrc_core_u_bs_convert__abc_21684_n340), .Y(u_sdrc_core_a2x_wrdt_12_) );
  OR2X2 OR2X2_904 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n342), .B(u_sdrc_core_u_bs_convert__abc_21684_n344), .Y(u_sdrc_core_a2x_wrdt_13_) );
  OR2X2 OR2X2_905 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n346), .B(u_sdrc_core_u_bs_convert__abc_21684_n348), .Y(u_sdrc_core_a2x_wrdt_14_) );
  OR2X2 OR2X2_906 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n350), .B(u_sdrc_core_u_bs_convert__abc_21684_n352), .Y(u_sdrc_core_a2x_wrdt_15_) );
  OR2X2 OR2X2_907 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n187_1), .B(u_sdrc_core_u_bs_convert__abc_21684_n356), .Y(u_sdrc_core_u_bs_convert__abc_21684_n357_1) );
  OR2X2 OR2X2_908 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n355), .B(u_sdrc_core_u_bs_convert__abc_21684_n357_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n358) );
  OR2X2 OR2X2_909 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n354), .B(u_sdrc_core_u_bs_convert__abc_21684_n358), .Y(u_sdrc_core_u_bs_convert__abc_21684_n359) );
  OR2X2 OR2X2_91 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n223_1_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_7_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n435) );
  OR2X2 OR2X2_910 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n175_1), .B(app_wr_en_n_2_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n365_1) );
  OR2X2 OR2X2_911 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf3), .B(app_wr_en_n_0_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n366) );
  OR2X2 OR2X2_912 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n368), .B(u_sdrc_core_u_bs_convert__abc_21684_n170_1_bF_buf1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n369) );
  OR2X2 OR2X2_913 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n364), .B(u_sdrc_core_u_bs_convert__abc_21684_n369), .Y(u_sdrc_core_u_bs_convert__abc_21684_n370) );
  OR2X2 OR2X2_914 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n171_1_bF_buf0), .B(app_wr_en_n_0_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n371_1) );
  OR2X2 OR2X2_915 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n373), .B(u_sdrc_core_u_bs_convert__abc_21684_n375), .Y(u_sdrc_core_a2x_wren_n_1_) );
  OR2X2 OR2X2_916 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n168_1), .B(u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n377) );
  OR2X2 OR2X2_917 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n378), .B(u_sdrc_core_u_bs_convert__abc_21684_n187_1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n379) );
  OR2X2 OR2X2_918 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n170_1_bF_buf0), .B(u_sdrc_core_u_bs_convert_saved_rd_data_0_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n381_1) );
  OR2X2 OR2X2_919 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n171_1_bF_buf3), .B(u_sdrc_core_pad_sdr_din2_0_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n382) );
  OR2X2 OR2X2_92 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n436), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf4), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n437) );
  OR2X2 OR2X2_920 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n170_1_bF_buf3), .B(u_sdrc_core_u_bs_convert_saved_rd_data_1_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n384) );
  OR2X2 OR2X2_921 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n171_1_bF_buf2), .B(u_sdrc_core_pad_sdr_din2_1_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n385) );
  OR2X2 OR2X2_922 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n170_1_bF_buf2), .B(u_sdrc_core_u_bs_convert_saved_rd_data_2_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n387) );
  OR2X2 OR2X2_923 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n171_1_bF_buf1), .B(u_sdrc_core_pad_sdr_din2_2_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n388) );
  OR2X2 OR2X2_924 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n170_1_bF_buf1), .B(u_sdrc_core_u_bs_convert_saved_rd_data_3_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n390) );
  OR2X2 OR2X2_925 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n171_1_bF_buf0), .B(u_sdrc_core_pad_sdr_din2_3_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n391_1) );
  OR2X2 OR2X2_926 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n170_1_bF_buf0), .B(u_sdrc_core_u_bs_convert_saved_rd_data_4_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n393) );
  OR2X2 OR2X2_927 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n171_1_bF_buf3), .B(u_sdrc_core_pad_sdr_din2_4_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n394) );
  OR2X2 OR2X2_928 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n170_1_bF_buf3), .B(u_sdrc_core_u_bs_convert_saved_rd_data_5_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n396_1) );
  OR2X2 OR2X2_929 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n171_1_bF_buf2), .B(u_sdrc_core_pad_sdr_din2_5_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n397) );
  OR2X2 OR2X2_93 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n283_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_7_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n438) );
  OR2X2 OR2X2_930 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n170_1_bF_buf2), .B(u_sdrc_core_u_bs_convert_saved_rd_data_6_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n399) );
  OR2X2 OR2X2_931 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n171_1_bF_buf1), .B(u_sdrc_core_pad_sdr_din2_6_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n400) );
  OR2X2 OR2X2_932 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n170_1_bF_buf1), .B(u_sdrc_core_u_bs_convert_saved_rd_data_7_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n402) );
  OR2X2 OR2X2_933 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n171_1_bF_buf0), .B(u_sdrc_core_pad_sdr_din2_7_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n403) );
  OR2X2 OR2X2_934 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n170_1_bF_buf0), .B(u_sdrc_core_u_bs_convert_saved_rd_data_8_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n405) );
  OR2X2 OR2X2_935 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n171_1_bF_buf3), .B(u_sdrc_core_pad_sdr_din2_8_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n406_1) );
  OR2X2 OR2X2_936 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n170_1_bF_buf3), .B(u_sdrc_core_u_bs_convert_saved_rd_data_9_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n408) );
  OR2X2 OR2X2_937 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n171_1_bF_buf2), .B(u_sdrc_core_pad_sdr_din2_9_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n409) );
  OR2X2 OR2X2_938 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n170_1_bF_buf2), .B(u_sdrc_core_u_bs_convert_saved_rd_data_10_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n411) );
  OR2X2 OR2X2_939 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n171_1_bF_buf1), .B(u_sdrc_core_pad_sdr_din2_10_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n412) );
  OR2X2 OR2X2_94 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n440), .B(u_sdrc_core_u_bank_ctl__abc_21249_n433), .Y(u_sdrc_core_b2x_addr_7_) );
  OR2X2 OR2X2_940 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n170_1_bF_buf1), .B(u_sdrc_core_u_bs_convert_saved_rd_data_11_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n414) );
  OR2X2 OR2X2_941 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n171_1_bF_buf0), .B(u_sdrc_core_pad_sdr_din2_11_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n415) );
  OR2X2 OR2X2_942 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n170_1_bF_buf0), .B(u_sdrc_core_u_bs_convert_saved_rd_data_12_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n417) );
  OR2X2 OR2X2_943 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n171_1_bF_buf3), .B(u_sdrc_core_pad_sdr_din2_12_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n418) );
  OR2X2 OR2X2_944 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n170_1_bF_buf3), .B(u_sdrc_core_u_bs_convert_saved_rd_data_13_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n420) );
  OR2X2 OR2X2_945 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n171_1_bF_buf2), .B(u_sdrc_core_pad_sdr_din2_13_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n421) );
  OR2X2 OR2X2_946 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n170_1_bF_buf2), .B(u_sdrc_core_u_bs_convert_saved_rd_data_14_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n423) );
  OR2X2 OR2X2_947 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n171_1_bF_buf1), .B(u_sdrc_core_pad_sdr_din2_14_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n424) );
  OR2X2 OR2X2_948 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n170_1_bF_buf1), .B(u_sdrc_core_u_bs_convert_saved_rd_data_15_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n426) );
  OR2X2 OR2X2_949 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n171_1_bF_buf0), .B(u_sdrc_core_pad_sdr_din2_15_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n427) );
  OR2X2 OR2X2_95 ( .A(u_sdrc_core_u_bank_ctl_bank1_fsm_xfr_ok_bF_buf3), .B(u_sdrc_core_u_bank_ctl_bank0_fsm_b2x_addr_8_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n443) );
  OR2X2 OR2X2_950 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n429), .B(u_sdrc_core_u_bs_convert__abc_21684_n430), .Y(app_rd_data_16_) );
  OR2X2 OR2X2_951 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n432), .B(u_sdrc_core_u_bs_convert__abc_21684_n433), .Y(app_rd_data_17_) );
  OR2X2 OR2X2_952 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n435), .B(u_sdrc_core_u_bs_convert__abc_21684_n436), .Y(app_rd_data_18_) );
  OR2X2 OR2X2_953 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n438), .B(u_sdrc_core_u_bs_convert__abc_21684_n439), .Y(app_rd_data_19_) );
  OR2X2 OR2X2_954 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n441), .B(u_sdrc_core_u_bs_convert__abc_21684_n442), .Y(app_rd_data_20_) );
  OR2X2 OR2X2_955 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n444), .B(u_sdrc_core_u_bs_convert__abc_21684_n445), .Y(app_rd_data_21_) );
  OR2X2 OR2X2_956 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n447), .B(u_sdrc_core_u_bs_convert__abc_21684_n448), .Y(app_rd_data_22_) );
  OR2X2 OR2X2_957 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n450), .B(u_sdrc_core_u_bs_convert__abc_21684_n451), .Y(app_rd_data_23_) );
  OR2X2 OR2X2_958 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n453), .B(u_sdrc_core_u_bs_convert__abc_21684_n454), .Y(app_rd_data_24_) );
  OR2X2 OR2X2_959 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n456), .B(u_sdrc_core_u_bs_convert__abc_21684_n457), .Y(app_rd_data_25_) );
  OR2X2 OR2X2_96 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n223_1_bF_buf1), .B(u_sdrc_core_u_bank_ctl_bank1_fsm_b2x_addr_8_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n444) );
  OR2X2 OR2X2_960 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n459), .B(u_sdrc_core_u_bs_convert__abc_21684_n460), .Y(app_rd_data_26_) );
  OR2X2 OR2X2_961 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n462), .B(u_sdrc_core_u_bs_convert__abc_21684_n463), .Y(app_rd_data_27_) );
  OR2X2 OR2X2_962 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n465), .B(u_sdrc_core_u_bs_convert__abc_21684_n466), .Y(app_rd_data_28_) );
  OR2X2 OR2X2_963 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n468), .B(u_sdrc_core_u_bs_convert__abc_21684_n469), .Y(app_rd_data_29_) );
  OR2X2 OR2X2_964 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n471), .B(u_sdrc_core_u_bs_convert__abc_21684_n472), .Y(app_rd_data_30_) );
  OR2X2 OR2X2_965 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n474), .B(u_sdrc_core_u_bs_convert__abc_21684_n475), .Y(app_rd_data_31_) );
  OR2X2 OR2X2_966 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n170_1_bF_buf0), .B(u_sdrc_core_u_bs_convert_rd_xfr_count_0_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n477) );
  OR2X2 OR2X2_967 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n169_1), .B(u_sdrc_core_u_bs_convert_rd_xfr_count_1_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n478) );
  OR2X2 OR2X2_968 ( .A(u_sdrc_core_u_bs_convert_wr_xfr_count_0_bF_buf4), .B(u_sdrc_core_u_bs_convert_x2a_wrnext_bF_buf1), .Y(u_sdrc_core_u_bs_convert__abc_21684_n485) );
  OR2X2 OR2X2_969 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n483), .B(u_sdrc_core_u_bs_convert_wr_xfr_count_1_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n490) );
  OR2X2 OR2X2_97 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n445), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_xfr_ok_bF_buf3), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n446) );
  OR2X2 OR2X2_970 ( .A(u_sdrc_core_u_bs_convert_x2a_rdok), .B(u_sdrc_core_u_bs_convert_rd_xfr_count_0_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n497) );
  OR2X2 OR2X2_971 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n495), .B(u_sdrc_core_u_bs_convert_rd_xfr_count_1_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n502) );
  OR2X2 OR2X2_972 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n511), .B(u_sdrc_core_u_bs_convert__abc_21684_n509), .Y(u_sdrc_core_u_bs_convert__abc_21684_n512) );
  OR2X2 OR2X2_973 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n515), .B(u_sdrc_core_u_bs_convert__abc_21684_n514), .Y(u_sdrc_core_u_bs_convert__abc_21684_n516) );
  OR2X2 OR2X2_974 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n519), .B(u_sdrc_core_u_bs_convert__abc_21684_n518), .Y(u_sdrc_core_u_bs_convert__abc_21684_n520) );
  OR2X2 OR2X2_975 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n523), .B(u_sdrc_core_u_bs_convert__abc_21684_n522), .Y(u_sdrc_core_u_bs_convert__abc_21684_n524) );
  OR2X2 OR2X2_976 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n527), .B(u_sdrc_core_u_bs_convert__abc_21684_n526), .Y(u_sdrc_core_u_bs_convert__abc_21684_n528) );
  OR2X2 OR2X2_977 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n531), .B(u_sdrc_core_u_bs_convert__abc_21684_n530), .Y(u_sdrc_core_u_bs_convert__abc_21684_n532) );
  OR2X2 OR2X2_978 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n535), .B(u_sdrc_core_u_bs_convert__abc_21684_n534), .Y(u_sdrc_core_u_bs_convert__abc_21684_n536) );
  OR2X2 OR2X2_979 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n539), .B(u_sdrc_core_u_bs_convert__abc_21684_n538), .Y(u_sdrc_core_u_bs_convert__abc_21684_n540) );
  OR2X2 OR2X2_98 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n283_bF_buf2), .B(u_sdrc_core_u_bank_ctl_bank2_fsm_b2x_addr_8_), .Y(u_sdrc_core_u_bank_ctl__abc_21249_n447) );
  OR2X2 OR2X2_980 ( .A(u_sdrc_core_u_bs_convert_rd_xfr_count_0_), .B(u_sdrc_core_u_bs_convert_rd_xfr_count_1_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n543) );
  OR2X2 OR2X2_981 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n544), .B(u_sdrc_core_u_bs_convert__abc_21684_n542), .Y(u_sdrc_core_u_bs_convert__abc_21684_n545) );
  OR2X2 OR2X2_982 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n546), .B(u_sdrc_core_u_bs_convert_saved_rd_data_0_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n547) );
  OR2X2 OR2X2_983 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n545), .B(u_sdrc_core_pad_sdr_din2_0_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n548) );
  OR2X2 OR2X2_984 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n546), .B(u_sdrc_core_u_bs_convert_saved_rd_data_1_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n551) );
  OR2X2 OR2X2_985 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n545), .B(u_sdrc_core_pad_sdr_din2_1_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n552) );
  OR2X2 OR2X2_986 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n546), .B(u_sdrc_core_u_bs_convert_saved_rd_data_2_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n555) );
  OR2X2 OR2X2_987 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n545), .B(u_sdrc_core_pad_sdr_din2_2_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n556) );
  OR2X2 OR2X2_988 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n546), .B(u_sdrc_core_u_bs_convert_saved_rd_data_3_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n559) );
  OR2X2 OR2X2_989 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n545), .B(u_sdrc_core_pad_sdr_din2_3_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n560) );
  OR2X2 OR2X2_99 ( .A(u_sdrc_core_u_bank_ctl__abc_21249_n449), .B(u_sdrc_core_u_bank_ctl__abc_21249_n442), .Y(u_sdrc_core_b2x_addr_8_) );
  OR2X2 OR2X2_990 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n546), .B(u_sdrc_core_u_bs_convert_saved_rd_data_4_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n563) );
  OR2X2 OR2X2_991 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n545), .B(u_sdrc_core_pad_sdr_din2_4_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n564) );
  OR2X2 OR2X2_992 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n546), .B(u_sdrc_core_u_bs_convert_saved_rd_data_5_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n567) );
  OR2X2 OR2X2_993 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n545), .B(u_sdrc_core_pad_sdr_din2_5_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n568) );
  OR2X2 OR2X2_994 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n546), .B(u_sdrc_core_u_bs_convert_saved_rd_data_6_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n571) );
  OR2X2 OR2X2_995 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n545), .B(u_sdrc_core_pad_sdr_din2_6_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n572) );
  OR2X2 OR2X2_996 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n546), .B(u_sdrc_core_u_bs_convert_saved_rd_data_7_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n575) );
  OR2X2 OR2X2_997 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n545), .B(u_sdrc_core_pad_sdr_din2_7_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n576) );
  OR2X2 OR2X2_998 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n505), .B(u_sdrc_core_u_bs_convert_rd_xfr_count_1_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n579) );
  OR2X2 OR2X2_999 ( .A(u_sdrc_core_u_bs_convert__abc_21684_n580), .B(u_sdrc_core_u_bs_convert_saved_rd_data_8_), .Y(u_sdrc_core_u_bs_convert__abc_21684_n581) );
endmodule
