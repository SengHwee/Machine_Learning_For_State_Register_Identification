module b08_reset(clock, RESET_G, nRESET_G, START, I_7_, I_6_, I_5_, I_4_, I_3_, I_2_, I_1_, I_0_, O_REG_3_, O_REG_2_, O_REG_1_, O_REG_0_);
  wire IN_R_REG_0_;
  wire IN_R_REG_1_;
  wire IN_R_REG_2_;
  wire IN_R_REG_3_;
  wire IN_R_REG_4_;
  wire IN_R_REG_5_;
  wire IN_R_REG_6_;
  wire IN_R_REG_7_;
  input I_0_;
  input I_1_;
  input I_2_;
  input I_3_;
  input I_4_;
  input I_5_;
  input I_6_;
  input I_7_;
  wire MAR_REG_0_;
  wire MAR_REG_1_;
  wire MAR_REG_2_;
  wire OUT_R_REG_0_;
  wire OUT_R_REG_1_;
  wire OUT_R_REG_2_;
  wire OUT_R_REG_3_;
  output O_REG_0_;
  output O_REG_1_;
  output O_REG_2_;
  output O_REG_3_;
  input RESET_G;
  input START;
  wire STATO_REG_0_;
  wire STATO_REG_1_;
  wire _abc_1014_n100_1;
  wire _abc_1014_n101;
  wire _abc_1014_n102;
  wire _abc_1014_n103;
  wire _abc_1014_n104_1;
  wire _abc_1014_n105;
  wire _abc_1014_n106;
  wire _abc_1014_n107;
  wire _abc_1014_n108;
  wire _abc_1014_n109;
  wire _abc_1014_n110;
  wire _abc_1014_n111;
  wire _abc_1014_n112;
  wire _abc_1014_n113;
  wire _abc_1014_n114_1;
  wire _abc_1014_n115;
  wire _abc_1014_n116_1;
  wire _abc_1014_n117;
  wire _abc_1014_n118_1;
  wire _abc_1014_n119;
  wire _abc_1014_n120_1;
  wire _abc_1014_n121;
  wire _abc_1014_n122;
  wire _abc_1014_n123_1;
  wire _abc_1014_n124_1;
  wire _abc_1014_n125;
  wire _abc_1014_n126;
  wire _abc_1014_n127_1;
  wire _abc_1014_n128_1;
  wire _abc_1014_n129;
  wire _abc_1014_n130_1;
  wire _abc_1014_n131;
  wire _abc_1014_n132;
  wire _abc_1014_n133_1;
  wire _abc_1014_n134_1;
  wire _abc_1014_n135;
  wire _abc_1014_n136;
  wire _abc_1014_n137;
  wire _abc_1014_n138;
  wire _abc_1014_n139_1;
  wire _abc_1014_n140;
  wire _abc_1014_n141_1;
  wire _abc_1014_n142;
  wire _abc_1014_n143;
  wire _abc_1014_n144;
  wire _abc_1014_n145;
  wire _abc_1014_n146_1;
  wire _abc_1014_n147;
  wire _abc_1014_n148_1;
  wire _abc_1014_n149_1;
  wire _abc_1014_n150;
  wire _abc_1014_n151;
  wire _abc_1014_n152_1;
  wire _abc_1014_n153_1;
  wire _abc_1014_n154;
  wire _abc_1014_n155;
  wire _abc_1014_n156_1;
  wire _abc_1014_n157_1;
  wire _abc_1014_n158;
  wire _abc_1014_n159;
  wire _abc_1014_n160_1;
  wire _abc_1014_n161_1;
  wire _abc_1014_n163;
  wire _abc_1014_n164_1;
  wire _abc_1014_n165_1;
  wire _abc_1014_n166;
  wire _abc_1014_n167;
  wire _abc_1014_n169_1;
  wire _abc_1014_n170;
  wire _abc_1014_n171;
  wire _abc_1014_n172_1;
  wire _abc_1014_n174;
  wire _abc_1014_n175;
  wire _abc_1014_n176;
  wire _abc_1014_n177;
  wire _abc_1014_n179;
  wire _abc_1014_n180;
  wire _abc_1014_n181;
  wire _abc_1014_n183;
  wire _abc_1014_n184;
  wire _abc_1014_n185;
  wire _abc_1014_n186;
  wire _abc_1014_n188;
  wire _abc_1014_n189;
  wire _abc_1014_n190;
  wire _abc_1014_n192;
  wire _abc_1014_n193;
  wire _abc_1014_n194;
  wire _abc_1014_n195;
  wire _abc_1014_n196;
  wire _abc_1014_n197;
  wire _abc_1014_n199;
  wire _abc_1014_n200;
  wire _abc_1014_n201;
  wire _abc_1014_n203;
  wire _abc_1014_n204;
  wire _abc_1014_n205;
  wire _abc_1014_n207;
  wire _abc_1014_n208;
  wire _abc_1014_n209;
  wire _abc_1014_n211;
  wire _abc_1014_n212;
  wire _abc_1014_n213;
  wire _abc_1014_n215;
  wire _abc_1014_n216;
  wire _abc_1014_n217;
  wire _abc_1014_n219;
  wire _abc_1014_n220;
  wire _abc_1014_n221;
  wire _abc_1014_n223;
  wire _abc_1014_n224;
  wire _abc_1014_n225;
  wire _abc_1014_n53;
  wire _abc_1014_n54;
  wire _abc_1014_n55;
  wire _abc_1014_n56;
  wire _abc_1014_n57;
  wire _abc_1014_n57_bF_buf0;
  wire _abc_1014_n57_bF_buf1;
  wire _abc_1014_n57_bF_buf2;
  wire _abc_1014_n57_bF_buf3;
  wire _abc_1014_n58;
  wire _abc_1014_n59;
  wire _abc_1014_n61;
  wire _abc_1014_n62;
  wire _abc_1014_n63;
  wire _abc_1014_n65;
  wire _abc_1014_n66;
  wire _abc_1014_n67;
  wire _abc_1014_n68;
  wire _abc_1014_n69;
  wire _abc_1014_n70;
  wire _abc_1014_n71_1;
  wire _abc_1014_n72;
  wire _abc_1014_n73;
  wire _abc_1014_n74;
  wire _abc_1014_n76;
  wire _abc_1014_n77;
  wire _abc_1014_n78_1;
  wire _abc_1014_n80;
  wire _abc_1014_n81;
  wire _abc_1014_n82;
  wire _abc_1014_n84;
  wire _abc_1014_n85;
  wire _abc_1014_n86;
  wire _abc_1014_n88;
  wire _abc_1014_n89;
  wire _abc_1014_n90;
  wire _abc_1014_n91;
  wire _abc_1014_n92;
  wire _abc_1014_n93;
  wire _abc_1014_n94;
  wire _abc_1014_n95;
  wire _abc_1014_n96;
  wire _abc_1014_n97;
  wire _abc_1014_n98;
  wire _abc_1014_n99;
  input clock;
  wire clock_bF_buf0;
  wire clock_bF_buf1;
  wire clock_bF_buf2;
  wire clock_bF_buf3;
  wire n101;
  wire n106;
  wire n111;
  wire n116;
  wire n121;
  wire n125;
  wire n129;
  wire n32;
  wire n36;
  wire n41;
  wire n46;
  wire n51;
  wire n56;
  wire n61;
  wire n66;
  wire n71;
  wire n76;
  wire n81;
  wire n86;
  wire n91;
  wire n96;
  input nRESET_G;
  AND2X2 AND2X2_1 ( .A(_abc_1014_n55), .B(I_1_), .Y(_abc_1014_n56) );
  AND2X2 AND2X2_10 ( .A(_abc_1014_n71_1), .B(O_REG_3_), .Y(_abc_1014_n72) );
  AND2X2 AND2X2_11 ( .A(_abc_1014_n70), .B(OUT_R_REG_3_), .Y(_abc_1014_n73) );
  AND2X2 AND2X2_12 ( .A(_abc_1014_n71_1), .B(O_REG_2_), .Y(_abc_1014_n76) );
  AND2X2 AND2X2_13 ( .A(_abc_1014_n70), .B(OUT_R_REG_2_), .Y(_abc_1014_n77) );
  AND2X2 AND2X2_14 ( .A(_abc_1014_n71_1), .B(O_REG_1_), .Y(_abc_1014_n80) );
  AND2X2 AND2X2_15 ( .A(_abc_1014_n70), .B(OUT_R_REG_1_), .Y(_abc_1014_n81) );
  AND2X2 AND2X2_16 ( .A(_abc_1014_n71_1), .B(O_REG_0_), .Y(_abc_1014_n84) );
  AND2X2 AND2X2_17 ( .A(_abc_1014_n70), .B(OUT_R_REG_0_), .Y(_abc_1014_n85) );
  AND2X2 AND2X2_18 ( .A(_abc_1014_n54), .B(OUT_R_REG_0_), .Y(_abc_1014_n88) );
  AND2X2 AND2X2_19 ( .A(_abc_1014_n92), .B(_abc_1014_n93), .Y(_abc_1014_n94) );
  AND2X2 AND2X2_2 ( .A(_abc_1014_n54), .B(IN_R_REG_1_), .Y(_abc_1014_n58) );
  AND2X2 AND2X2_20 ( .A(_abc_1014_n94), .B(_abc_1014_n89), .Y(_abc_1014_n95) );
  AND2X2 AND2X2_21 ( .A(_abc_1014_n93), .B(MAR_REG_2_), .Y(_abc_1014_n96) );
  AND2X2 AND2X2_22 ( .A(_abc_1014_n96), .B(MAR_REG_1_), .Y(_abc_1014_n97) );
  AND2X2 AND2X2_23 ( .A(MAR_REG_1_), .B(MAR_REG_0_), .Y(_abc_1014_n99) );
  AND2X2 AND2X2_24 ( .A(_abc_1014_n99), .B(_abc_1014_n92), .Y(_abc_1014_n100_1) );
  AND2X2 AND2X2_25 ( .A(_abc_1014_n89), .B(MAR_REG_2_), .Y(_abc_1014_n101) );
  AND2X2 AND2X2_26 ( .A(_abc_1014_n90), .B(_abc_1014_n105), .Y(_abc_1014_n106) );
  AND2X2 AND2X2_27 ( .A(_abc_1014_n103), .B(_abc_1014_n107), .Y(_abc_1014_n108) );
  AND2X2 AND2X2_28 ( .A(_abc_1014_n92), .B(MAR_REG_0_), .Y(_abc_1014_n112) );
  AND2X2 AND2X2_29 ( .A(_abc_1014_n112), .B(_abc_1014_n89), .Y(_abc_1014_n113) );
  AND2X2 AND2X2_3 ( .A(_abc_1014_n55), .B(I_0_), .Y(_abc_1014_n61) );
  AND2X2 AND2X2_30 ( .A(_abc_1014_n115), .B(_abc_1014_n105), .Y(_abc_1014_n116_1) );
  AND2X2 AND2X2_31 ( .A(_abc_1014_n117), .B(_abc_1014_n111), .Y(_abc_1014_n118_1) );
  AND2X2 AND2X2_32 ( .A(_abc_1014_n109), .B(_abc_1014_n118_1), .Y(_abc_1014_n119) );
  AND2X2 AND2X2_33 ( .A(_abc_1014_n122), .B(_abc_1014_n121), .Y(_abc_1014_n123_1) );
  AND2X2 AND2X2_34 ( .A(_abc_1014_n127_1), .B(_abc_1014_n125), .Y(_abc_1014_n128_1) );
  AND2X2 AND2X2_35 ( .A(_abc_1014_n124_1), .B(_abc_1014_n128_1), .Y(_abc_1014_n129) );
  AND2X2 AND2X2_36 ( .A(_abc_1014_n122), .B(_abc_1014_n105), .Y(_abc_1014_n133_1) );
  AND2X2 AND2X2_37 ( .A(_abc_1014_n132), .B(_abc_1014_n134_1), .Y(_abc_1014_n135) );
  AND2X2 AND2X2_38 ( .A(_abc_1014_n130_1), .B(_abc_1014_n135), .Y(_abc_1014_n136) );
  AND2X2 AND2X2_39 ( .A(_abc_1014_n126), .B(MAR_REG_1_), .Y(_abc_1014_n137) );
  AND2X2 AND2X2_4 ( .A(_abc_1014_n54), .B(IN_R_REG_0_), .Y(_abc_1014_n62) );
  AND2X2 AND2X2_40 ( .A(_abc_1014_n140), .B(_abc_1014_n141_1), .Y(_abc_1014_n142) );
  AND2X2 AND2X2_41 ( .A(_abc_1014_n148_1), .B(_abc_1014_n150), .Y(_abc_1014_n151) );
  AND2X2 AND2X2_42 ( .A(_abc_1014_n53), .B(STATO_REG_1_), .Y(_abc_1014_n152_1) );
  AND2X2 AND2X2_43 ( .A(_abc_1014_n153_1), .B(_abc_1014_n152_1), .Y(_abc_1014_n154) );
  AND2X2 AND2X2_44 ( .A(_abc_1014_n151), .B(_abc_1014_n154), .Y(_abc_1014_n155) );
  AND2X2 AND2X2_45 ( .A(_abc_1014_n155), .B(_abc_1014_n146_1), .Y(_abc_1014_n156_1) );
  AND2X2 AND2X2_46 ( .A(_abc_1014_n143), .B(_abc_1014_n156_1), .Y(_abc_1014_n157_1) );
  AND2X2 AND2X2_47 ( .A(_abc_1014_n136), .B(_abc_1014_n157_1), .Y(_abc_1014_n158) );
  AND2X2 AND2X2_48 ( .A(_abc_1014_n120_1), .B(_abc_1014_n158), .Y(_abc_1014_n159) );
  AND2X2 AND2X2_49 ( .A(_abc_1014_n159), .B(_abc_1014_n91), .Y(_abc_1014_n160_1) );
  AND2X2 AND2X2_5 ( .A(MAR_REG_2_), .B(MAR_REG_0_), .Y(_abc_1014_n66) );
  AND2X2 AND2X2_50 ( .A(_abc_1014_n90), .B(_abc_1014_n163), .Y(_abc_1014_n164_1) );
  AND2X2 AND2X2_51 ( .A(_abc_1014_n159), .B(_abc_1014_n164_1), .Y(_abc_1014_n165_1) );
  AND2X2 AND2X2_52 ( .A(_abc_1014_n54), .B(OUT_R_REG_1_), .Y(_abc_1014_n166) );
  AND2X2 AND2X2_53 ( .A(_abc_1014_n138), .B(_abc_1014_n115), .Y(_abc_1014_n169_1) );
  AND2X2 AND2X2_54 ( .A(_abc_1014_n159), .B(_abc_1014_n169_1), .Y(_abc_1014_n170) );
  AND2X2 AND2X2_55 ( .A(_abc_1014_n54), .B(OUT_R_REG_2_), .Y(_abc_1014_n171) );
  AND2X2 AND2X2_56 ( .A(_abc_1014_n54), .B(OUT_R_REG_3_), .Y(_abc_1014_n174) );
  AND2X2 AND2X2_57 ( .A(_abc_1014_n159), .B(_abc_1014_n175), .Y(_abc_1014_n176) );
  AND2X2 AND2X2_58 ( .A(_abc_1014_n100_1), .B(_abc_1014_n69), .Y(_abc_1014_n179) );
  AND2X2 AND2X2_59 ( .A(_abc_1014_n54), .B(MAR_REG_2_), .Y(_abc_1014_n180) );
  AND2X2 AND2X2_6 ( .A(_abc_1014_n66), .B(MAR_REG_1_), .Y(_abc_1014_n67) );
  AND2X2 AND2X2_60 ( .A(_abc_1014_n184), .B(_abc_1014_n54), .Y(_abc_1014_n185) );
  AND2X2 AND2X2_61 ( .A(_abc_1014_n185), .B(START), .Y(_abc_1014_n186) );
  AND2X2 AND2X2_62 ( .A(_abc_1014_n188), .B(STATO_REG_0_), .Y(_abc_1014_n189) );
  AND2X2 AND2X2_63 ( .A(_abc_1014_n54), .B(MAR_REG_1_), .Y(_abc_1014_n193) );
  AND2X2 AND2X2_64 ( .A(_abc_1014_n192), .B(_abc_1014_n193), .Y(_abc_1014_n194) );
  AND2X2 AND2X2_65 ( .A(_abc_1014_n89), .B(MAR_REG_0_), .Y(_abc_1014_n195) );
  AND2X2 AND2X2_66 ( .A(_abc_1014_n195), .B(_abc_1014_n69), .Y(_abc_1014_n196) );
  AND2X2 AND2X2_67 ( .A(_abc_1014_n185), .B(MAR_REG_0_), .Y(_abc_1014_n199) );
  AND2X2 AND2X2_68 ( .A(_abc_1014_n69), .B(_abc_1014_n93), .Y(_abc_1014_n200) );
  AND2X2 AND2X2_69 ( .A(_abc_1014_n55), .B(I_7_), .Y(_abc_1014_n203) );
  AND2X2 AND2X2_7 ( .A(_abc_1014_n67), .B(_abc_1014_n65), .Y(_abc_1014_n68) );
  AND2X2 AND2X2_70 ( .A(_abc_1014_n54), .B(IN_R_REG_7_), .Y(_abc_1014_n204) );
  AND2X2 AND2X2_71 ( .A(_abc_1014_n55), .B(I_6_), .Y(_abc_1014_n207) );
  AND2X2 AND2X2_72 ( .A(_abc_1014_n54), .B(IN_R_REG_6_), .Y(_abc_1014_n208) );
  AND2X2 AND2X2_73 ( .A(_abc_1014_n55), .B(I_5_), .Y(_abc_1014_n211) );
  AND2X2 AND2X2_74 ( .A(_abc_1014_n54), .B(IN_R_REG_5_), .Y(_abc_1014_n212) );
  AND2X2 AND2X2_75 ( .A(_abc_1014_n55), .B(I_4_), .Y(_abc_1014_n215) );
  AND2X2 AND2X2_76 ( .A(_abc_1014_n54), .B(IN_R_REG_4_), .Y(_abc_1014_n216) );
  AND2X2 AND2X2_77 ( .A(_abc_1014_n55), .B(I_3_), .Y(_abc_1014_n219) );
  AND2X2 AND2X2_78 ( .A(_abc_1014_n54), .B(IN_R_REG_3_), .Y(_abc_1014_n220) );
  AND2X2 AND2X2_79 ( .A(_abc_1014_n55), .B(I_2_), .Y(_abc_1014_n223) );
  AND2X2 AND2X2_8 ( .A(STATO_REG_0_), .B(STATO_REG_1_), .Y(_abc_1014_n69) );
  AND2X2 AND2X2_80 ( .A(_abc_1014_n54), .B(IN_R_REG_2_), .Y(_abc_1014_n224) );
  AND2X2 AND2X2_9 ( .A(_abc_1014_n68), .B(_abc_1014_n69), .Y(_abc_1014_n70) );
  DFFPOSX1 DFFPOSX1_1 ( .CLK(clock), .D(n121), .Q(O_REG_3_) );
  DFFPOSX1 DFFPOSX1_10 ( .CLK(clock), .D(n61), .Q(IN_R_REG_7_) );
  DFFPOSX1 DFFPOSX1_11 ( .CLK(clock), .D(n66), .Q(IN_R_REG_6_) );
  DFFPOSX1 DFFPOSX1_12 ( .CLK(clock), .D(n71), .Q(IN_R_REG_5_) );
  DFFPOSX1 DFFPOSX1_13 ( .CLK(clock), .D(n76), .Q(IN_R_REG_4_) );
  DFFPOSX1 DFFPOSX1_14 ( .CLK(clock), .D(n81), .Q(IN_R_REG_3_) );
  DFFPOSX1 DFFPOSX1_15 ( .CLK(clock), .D(n86), .Q(IN_R_REG_2_) );
  DFFPOSX1 DFFPOSX1_16 ( .CLK(clock), .D(n91), .Q(IN_R_REG_1_) );
  DFFPOSX1 DFFPOSX1_17 ( .CLK(clock), .D(n96), .Q(IN_R_REG_0_) );
  DFFPOSX1 DFFPOSX1_18 ( .CLK(clock), .D(n101), .Q(OUT_R_REG_3_) );
  DFFPOSX1 DFFPOSX1_19 ( .CLK(clock), .D(n106), .Q(OUT_R_REG_2_) );
  DFFPOSX1 DFFPOSX1_2 ( .CLK(clock), .D(n125), .Q(O_REG_2_) );
  DFFPOSX1 DFFPOSX1_20 ( .CLK(clock), .D(n111), .Q(OUT_R_REG_1_) );
  DFFPOSX1 DFFPOSX1_21 ( .CLK(clock), .D(n116), .Q(OUT_R_REG_0_) );
  DFFPOSX1 DFFPOSX1_3 ( .CLK(clock), .D(n129), .Q(O_REG_1_) );
  DFFPOSX1 DFFPOSX1_4 ( .CLK(clock), .D(n32), .Q(O_REG_0_) );
  DFFPOSX1 DFFPOSX1_5 ( .CLK(clock), .D(n36), .Q(STATO_REG_1_) );
  DFFPOSX1 DFFPOSX1_6 ( .CLK(clock), .D(n41), .Q(STATO_REG_0_) );
  DFFPOSX1 DFFPOSX1_7 ( .CLK(clock), .D(n46), .Q(MAR_REG_2_) );
  DFFPOSX1 DFFPOSX1_8 ( .CLK(clock), .D(n51), .Q(MAR_REG_1_) );
  DFFPOSX1 DFFPOSX1_9 ( .CLK(clock), .D(n56), .Q(MAR_REG_0_) );
  INVX1 INVX1_1 ( .A(STATO_REG_0_), .Y(_abc_1014_n53) );
  INVX1 INVX1_10 ( .A(IN_R_REG_4_), .Y(_abc_1014_n121) );
  INVX1 INVX1_11 ( .A(_abc_1014_n96), .Y(_abc_1014_n122) );
  INVX1 INVX1_12 ( .A(IN_R_REG_5_), .Y(_abc_1014_n131) );
  INVX1 INVX1_13 ( .A(IN_R_REG_7_), .Y(_abc_1014_n144) );
  INVX1 INVX1_14 ( .A(IN_R_REG_0_), .Y(_abc_1014_n147) );
  INVX1 INVX1_15 ( .A(_abc_1014_n66), .Y(_abc_1014_n163) );
  INVX1 INVX1_16 ( .A(_abc_1014_n68), .Y(_abc_1014_n188) );
  INVX1 INVX1_2 ( .A(START), .Y(_abc_1014_n65) );
  INVX1 INVX1_3 ( .A(_abc_1014_n70), .Y(_abc_1014_n71_1) );
  INVX1 INVX1_4 ( .A(_abc_1014_n90), .Y(_abc_1014_n91) );
  INVX1 INVX1_5 ( .A(MAR_REG_2_), .Y(_abc_1014_n92) );
  INVX1 INVX1_6 ( .A(IN_R_REG_6_), .Y(_abc_1014_n98) );
  INVX1 INVX1_7 ( .A(IN_R_REG_1_), .Y(_abc_1014_n104_1) );
  INVX1 INVX1_8 ( .A(IN_R_REG_2_), .Y(_abc_1014_n110) );
  INVX1 INVX1_9 ( .A(_abc_1014_n97), .Y(_abc_1014_n115) );
  INVX2 INVX2_1 ( .A(_abc_1014_n54), .Y(_abc_1014_n55) );
  INVX2 INVX2_2 ( .A(MAR_REG_1_), .Y(_abc_1014_n89) );
  INVX2 INVX2_3 ( .A(MAR_REG_0_), .Y(_abc_1014_n93) );
  INVX8 INVX8_1 ( .A(nRESET_G), .Y(_abc_1014_n57) );
  OR2X2 OR2X2_1 ( .A(_abc_1014_n53), .B(STATO_REG_1_), .Y(_abc_1014_n54) );
  OR2X2 OR2X2_10 ( .A(_abc_1014_n81), .B(_abc_1014_n57), .Y(_abc_1014_n82) );
  OR2X2 OR2X2_11 ( .A(_abc_1014_n82), .B(_abc_1014_n80), .Y(n129) );
  OR2X2 OR2X2_12 ( .A(_abc_1014_n85), .B(_abc_1014_n57), .Y(_abc_1014_n86) );
  OR2X2 OR2X2_13 ( .A(_abc_1014_n86), .B(_abc_1014_n84), .Y(n32) );
  OR2X2 OR2X2_14 ( .A(_abc_1014_n89), .B(MAR_REG_0_), .Y(_abc_1014_n90) );
  OR2X2 OR2X2_15 ( .A(_abc_1014_n100_1), .B(_abc_1014_n101), .Y(_abc_1014_n102) );
  OR2X2 OR2X2_16 ( .A(_abc_1014_n102), .B(_abc_1014_n98), .Y(_abc_1014_n103) );
  OR2X2 OR2X2_17 ( .A(MAR_REG_1_), .B(MAR_REG_2_), .Y(_abc_1014_n105) );
  OR2X2 OR2X2_18 ( .A(_abc_1014_n106), .B(_abc_1014_n104_1), .Y(_abc_1014_n107) );
  OR2X2 OR2X2_19 ( .A(_abc_1014_n108), .B(_abc_1014_n97), .Y(_abc_1014_n109) );
  OR2X2 OR2X2_2 ( .A(_abc_1014_n58), .B(_abc_1014_n57), .Y(_abc_1014_n59) );
  OR2X2 OR2X2_20 ( .A(_abc_1014_n106), .B(_abc_1014_n110), .Y(_abc_1014_n111) );
  OR2X2 OR2X2_21 ( .A(_abc_1014_n113), .B(IN_R_REG_1_), .Y(_abc_1014_n114_1) );
  OR2X2 OR2X2_22 ( .A(_abc_1014_n116_1), .B(_abc_1014_n114_1), .Y(_abc_1014_n117) );
  OR2X2 OR2X2_23 ( .A(_abc_1014_n119), .B(_abc_1014_n95), .Y(_abc_1014_n120_1) );
  OR2X2 OR2X2_24 ( .A(_abc_1014_n123_1), .B(IN_R_REG_7_), .Y(_abc_1014_n124_1) );
  OR2X2 OR2X2_25 ( .A(_abc_1014_n112), .B(_abc_1014_n121), .Y(_abc_1014_n125) );
  OR2X2 OR2X2_26 ( .A(_abc_1014_n93), .B(MAR_REG_2_), .Y(_abc_1014_n126) );
  OR2X2 OR2X2_27 ( .A(_abc_1014_n126), .B(IN_R_REG_4_), .Y(_abc_1014_n127_1) );
  OR2X2 OR2X2_28 ( .A(_abc_1014_n129), .B(_abc_1014_n89), .Y(_abc_1014_n130_1) );
  OR2X2 OR2X2_29 ( .A(_abc_1014_n115), .B(_abc_1014_n131), .Y(_abc_1014_n132) );
  OR2X2 OR2X2_3 ( .A(_abc_1014_n59), .B(_abc_1014_n56), .Y(n91) );
  OR2X2 OR2X2_30 ( .A(_abc_1014_n133_1), .B(IN_R_REG_3_), .Y(_abc_1014_n134_1) );
  OR2X2 OR2X2_31 ( .A(_abc_1014_n137), .B(_abc_1014_n96), .Y(_abc_1014_n138) );
  OR2X2 OR2X2_32 ( .A(_abc_1014_n138), .B(_abc_1014_n113), .Y(_abc_1014_n139_1) );
  OR2X2 OR2X2_33 ( .A(_abc_1014_n95), .B(IN_R_REG_2_), .Y(_abc_1014_n140) );
  OR2X2 OR2X2_34 ( .A(_abc_1014_n100_1), .B(IN_R_REG_6_), .Y(_abc_1014_n141_1) );
  OR2X2 OR2X2_35 ( .A(_abc_1014_n139_1), .B(_abc_1014_n142), .Y(_abc_1014_n143) );
  OR2X2 OR2X2_36 ( .A(_abc_1014_n91), .B(_abc_1014_n144), .Y(_abc_1014_n145) );
  OR2X2 OR2X2_37 ( .A(_abc_1014_n145), .B(_abc_1014_n102), .Y(_abc_1014_n146_1) );
  OR2X2 OR2X2_38 ( .A(_abc_1014_n90), .B(_abc_1014_n147), .Y(_abc_1014_n148_1) );
  OR2X2 OR2X2_39 ( .A(IN_R_REG_0_), .B(MAR_REG_1_), .Y(_abc_1014_n149_1) );
  OR2X2 OR2X2_4 ( .A(_abc_1014_n62), .B(_abc_1014_n57), .Y(_abc_1014_n63) );
  OR2X2 OR2X2_40 ( .A(_abc_1014_n94), .B(_abc_1014_n149_1), .Y(_abc_1014_n150) );
  OR2X2 OR2X2_41 ( .A(_abc_1014_n105), .B(IN_R_REG_5_), .Y(_abc_1014_n153_1) );
  OR2X2 OR2X2_42 ( .A(_abc_1014_n160_1), .B(_abc_1014_n57), .Y(_abc_1014_n161_1) );
  OR2X2 OR2X2_43 ( .A(_abc_1014_n161_1), .B(_abc_1014_n88), .Y(n116) );
  OR2X2 OR2X2_44 ( .A(_abc_1014_n165_1), .B(_abc_1014_n166), .Y(_abc_1014_n167) );
  OR2X2 OR2X2_45 ( .A(_abc_1014_n161_1), .B(_abc_1014_n167), .Y(n111) );
  OR2X2 OR2X2_46 ( .A(_abc_1014_n171), .B(_abc_1014_n57), .Y(_abc_1014_n172_1) );
  OR2X2 OR2X2_47 ( .A(_abc_1014_n170), .B(_abc_1014_n172_1), .Y(n106) );
  OR2X2 OR2X2_48 ( .A(_abc_1014_n102), .B(_abc_1014_n95), .Y(_abc_1014_n175) );
  OR2X2 OR2X2_49 ( .A(_abc_1014_n176), .B(_abc_1014_n174), .Y(_abc_1014_n177) );
  OR2X2 OR2X2_5 ( .A(_abc_1014_n63), .B(_abc_1014_n61), .Y(n96) );
  OR2X2 OR2X2_50 ( .A(_abc_1014_n161_1), .B(_abc_1014_n177), .Y(n101) );
  OR2X2 OR2X2_51 ( .A(_abc_1014_n180), .B(_abc_1014_n57), .Y(_abc_1014_n181) );
  OR2X2 OR2X2_52 ( .A(_abc_1014_n181), .B(_abc_1014_n179), .Y(n46) );
  OR2X2 OR2X2_53 ( .A(_abc_1014_n152_1), .B(_abc_1014_n57), .Y(_abc_1014_n183) );
  OR2X2 OR2X2_54 ( .A(_abc_1014_n67), .B(_abc_1014_n53), .Y(_abc_1014_n184) );
  OR2X2 OR2X2_55 ( .A(_abc_1014_n186), .B(_abc_1014_n183), .Y(n41) );
  OR2X2 OR2X2_56 ( .A(_abc_1014_n183), .B(_abc_1014_n55), .Y(_abc_1014_n190) );
  OR2X2 OR2X2_57 ( .A(_abc_1014_n189), .B(_abc_1014_n190), .Y(n36) );
  OR2X2 OR2X2_58 ( .A(_abc_1014_n184), .B(_abc_1014_n93), .Y(_abc_1014_n192) );
  OR2X2 OR2X2_59 ( .A(_abc_1014_n196), .B(_abc_1014_n57), .Y(_abc_1014_n197) );
  OR2X2 OR2X2_6 ( .A(_abc_1014_n73), .B(_abc_1014_n57), .Y(_abc_1014_n74) );
  OR2X2 OR2X2_60 ( .A(_abc_1014_n194), .B(_abc_1014_n197), .Y(n51) );
  OR2X2 OR2X2_61 ( .A(_abc_1014_n200), .B(_abc_1014_n57), .Y(_abc_1014_n201) );
  OR2X2 OR2X2_62 ( .A(_abc_1014_n199), .B(_abc_1014_n201), .Y(n56) );
  OR2X2 OR2X2_63 ( .A(_abc_1014_n204), .B(_abc_1014_n57), .Y(_abc_1014_n205) );
  OR2X2 OR2X2_64 ( .A(_abc_1014_n205), .B(_abc_1014_n203), .Y(n61) );
  OR2X2 OR2X2_65 ( .A(_abc_1014_n208), .B(_abc_1014_n57), .Y(_abc_1014_n209) );
  OR2X2 OR2X2_66 ( .A(_abc_1014_n209), .B(_abc_1014_n207), .Y(n66) );
  OR2X2 OR2X2_67 ( .A(_abc_1014_n212), .B(_abc_1014_n57), .Y(_abc_1014_n213) );
  OR2X2 OR2X2_68 ( .A(_abc_1014_n213), .B(_abc_1014_n211), .Y(n71) );
  OR2X2 OR2X2_69 ( .A(_abc_1014_n216), .B(_abc_1014_n57), .Y(_abc_1014_n217) );
  OR2X2 OR2X2_7 ( .A(_abc_1014_n74), .B(_abc_1014_n72), .Y(n121) );
  OR2X2 OR2X2_70 ( .A(_abc_1014_n217), .B(_abc_1014_n215), .Y(n76) );
  OR2X2 OR2X2_71 ( .A(_abc_1014_n220), .B(_abc_1014_n57), .Y(_abc_1014_n221) );
  OR2X2 OR2X2_72 ( .A(_abc_1014_n221), .B(_abc_1014_n219), .Y(n81) );
  OR2X2 OR2X2_73 ( .A(_abc_1014_n224), .B(_abc_1014_n57), .Y(_abc_1014_n225) );
  OR2X2 OR2X2_74 ( .A(_abc_1014_n225), .B(_abc_1014_n223), .Y(n86) );
  OR2X2 OR2X2_8 ( .A(_abc_1014_n77), .B(_abc_1014_n57), .Y(_abc_1014_n78_1) );
  OR2X2 OR2X2_9 ( .A(_abc_1014_n78_1), .B(_abc_1014_n76), .Y(n125) );
endmodule