module b02_reset(clock, RESET_G, nRESET_G, LINEA, U_REG);

input LINEA;
input RESET_G;
wire STATO_REG_0_; 
wire STATO_REG_1_; 
wire STATO_REG_2_; 
output U_REG;
wire _abc_181_new_n10_; 
wire _abc_181_new_n11_; 
wire _abc_181_new_n13_; 
wire _abc_181_new_n14_; 
wire _abc_181_new_n15_; 
wire _abc_181_new_n16_; 
wire _abc_181_new_n17_; 
wire _abc_181_new_n18_; 
wire _abc_181_new_n20_; 
wire _abc_181_new_n21_; 
wire _abc_181_new_n22_; 
wire _abc_181_new_n23_; 
wire _abc_181_new_n24_; 
wire _abc_181_new_n25_; 
wire _abc_181_new_n27_; 
wire _abc_181_new_n28_; 
wire _auto_iopadmap_cc_368_execute_202; 
input clock;
wire n10; 
wire n14; 
wire n19; 
wire n24; 
input nRESET_G;
AOI21X1 AOI21X1_1 ( .A(_abc_181_new_n14_), .B(LINEA), .C(_abc_181_new_n13_), .Y(_abc_181_new_n15_));
AOI21X1 AOI21X1_2 ( .A(_abc_181_new_n17_), .B(_abc_181_new_n13_), .C(_abc_181_new_n16_), .Y(_abc_181_new_n18_));
BUFX2 BUFX2_1 ( .A(_auto_iopadmap_cc_368_execute_202), .Y(U_REG));
DFFPOSX1 DFFPOSX1_1 ( .CLK(clock), .D(n24), .Q(STATO_REG_0_));
DFFPOSX1 DFFPOSX1_2 ( .CLK(clock), .D(n19), .Q(STATO_REG_1_));
DFFPOSX1 DFFPOSX1_3 ( .CLK(clock), .D(n10), .Q(_auto_iopadmap_cc_368_execute_202));
DFFPOSX1 DFFPOSX1_4 ( .CLK(clock), .D(n14), .Q(STATO_REG_2_));
INVX1 INVX1_1 ( .A(STATO_REG_1_), .Y(_abc_181_new_n10_));
INVX1 INVX1_2 ( .A(STATO_REG_2_), .Y(_abc_181_new_n14_));
INVX1 INVX1_3 ( .A(nRESET_G), .Y(_abc_181_new_n16_));
INVX1 INVX1_4 ( .A(LINEA), .Y(_abc_181_new_n20_));
INVX2 INVX2_1 ( .A(STATO_REG_0_), .Y(_abc_181_new_n13_));
NAND2X1 NAND2X1_1 ( .A(_abc_181_new_n10_), .B(_abc_181_new_n23_), .Y(_abc_181_new_n24_));
NAND2X1 NAND2X1_2 ( .A(nRESET_G), .B(_abc_181_new_n25_), .Y(n14));
NAND3X1 NAND3X1_1 ( .A(nRESET_G), .B(STATO_REG_2_), .C(_abc_181_new_n10_), .Y(_abc_181_new_n11_));
NAND3X1 NAND3X1_2 ( .A(STATO_REG_1_), .B(_abc_181_new_n13_), .C(_abc_181_new_n14_), .Y(_abc_181_new_n28_));
NAND3X1 NAND3X1_3 ( .A(nRESET_G), .B(_abc_181_new_n28_), .C(_abc_181_new_n27_), .Y(n19));
NOR2X1 NOR2X1_1 ( .A(STATO_REG_0_), .B(_abc_181_new_n11_), .Y(n10));
NOR2X1 NOR2X1_2 ( .A(STATO_REG_2_), .B(LINEA), .Y(_abc_181_new_n17_));
NOR2X1 NOR2X1_3 ( .A(STATO_REG_2_), .B(_abc_181_new_n20_), .Y(_abc_181_new_n21_));
OAI21X1 OAI21X1_1 ( .A(STATO_REG_1_), .B(_abc_181_new_n15_), .C(_abc_181_new_n18_), .Y(n24));
OAI21X1 OAI21X1_2 ( .A(LINEA), .B(_abc_181_new_n14_), .C(_abc_181_new_n13_), .Y(_abc_181_new_n22_));
OAI21X1 OAI21X1_3 ( .A(STATO_REG_2_), .B(LINEA), .C(STATO_REG_0_), .Y(_abc_181_new_n23_));
OAI21X1 OAI21X1_4 ( .A(_abc_181_new_n21_), .B(_abc_181_new_n22_), .C(_abc_181_new_n24_), .Y(_abc_181_new_n25_));
OAI21X1 OAI21X1_5 ( .A(_abc_181_new_n10_), .B(STATO_REG_2_), .C(_abc_181_new_n15_), .Y(_abc_181_new_n27_));


endmodule